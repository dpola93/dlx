
module SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_16 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net338260, net338262, net338263, net338266;
  assign net338260 = CLK;
  assign ENCLK = net338262;
  assign net338263 = EN;

  DLL_X1 latch ( .D(net338263), .GN(net338260), .Q(net338266) );
  AND2_X1 main_gate ( .A1(net338266), .A2(net338260), .ZN(net338262) );
endmodule


module SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_15 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net338260, net338262, net338263, net338266;
  assign net338260 = CLK;
  assign ENCLK = net338262;
  assign net338263 = EN;

  DLL_X1 latch ( .D(net338263), .GN(net338260), .Q(net338266) );
  AND2_X1 main_gate ( .A1(net338266), .A2(net338260), .ZN(net338262) );
endmodule


module SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_14 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net338260, net338262, net338263, net338266;
  assign net338260 = CLK;
  assign ENCLK = net338262;
  assign net338263 = EN;

  DLL_X1 latch ( .D(net338263), .GN(net338260), .Q(net338266) );
  AND2_X1 main_gate ( .A1(net338266), .A2(net338260), .ZN(net338262) );
endmodule


module SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_13 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net338260, net338262, net338263, net338266;
  assign net338260 = CLK;
  assign ENCLK = net338262;
  assign net338263 = EN;

  DLL_X1 latch ( .D(net338263), .GN(net338260), .Q(net338266) );
  AND2_X1 main_gate ( .A1(net338266), .A2(net338260), .ZN(net338262) );
endmodule


module SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_12 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net338260, net338262, net338263, net338266;
  assign net338260 = CLK;
  assign ENCLK = net338262;
  assign net338263 = EN;

  DLL_X1 latch ( .D(net338263), .GN(net338260), .Q(net338266) );
  AND2_X1 main_gate ( .A1(net338266), .A2(net338260), .ZN(net338262) );
endmodule


module SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_11 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net338260, net338262, net338263, net338266;
  assign net338260 = CLK;
  assign ENCLK = net338262;
  assign net338263 = EN;

  DLL_X1 latch ( .D(net338263), .GN(net338260), .Q(net338266) );
  AND2_X1 main_gate ( .A1(net338266), .A2(net338260), .ZN(net338262) );
endmodule


module SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_10 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net338260, net338262, net338263, net338266;
  assign net338260 = CLK;
  assign ENCLK = net338262;
  assign net338263 = EN;

  DLL_X1 latch ( .D(net338263), .GN(net338260), .Q(net338266) );
  AND2_X1 main_gate ( .A1(net338266), .A2(net338260), .ZN(net338262) );
endmodule


module SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_9 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net338260, net338262, net338263, net338266;
  assign net338260 = CLK;
  assign ENCLK = net338262;
  assign net338263 = EN;

  DLL_X1 latch ( .D(net338263), .GN(net338260), .Q(net338266) );
  AND2_X1 main_gate ( .A1(net338266), .A2(net338260), .ZN(net338262) );
endmodule


module SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_8 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net338260, net338262, net338263, net338266;
  assign net338260 = CLK;
  assign ENCLK = net338262;
  assign net338263 = EN;

  DLL_X1 latch ( .D(net338263), .GN(net338260), .Q(net338266) );
  AND2_X1 main_gate ( .A1(net338266), .A2(net338260), .ZN(net338262) );
endmodule


module SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_7 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net338260, net338262, net338263, net338266;
  assign net338260 = CLK;
  assign ENCLK = net338262;
  assign net338263 = EN;

  DLL_X1 latch ( .D(net338263), .GN(net338260), .Q(net338266) );
  AND2_X1 main_gate ( .A1(net338266), .A2(net338260), .ZN(net338262) );
endmodule


module SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_6 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net338260, net338262, net338263, net338266;
  assign net338260 = CLK;
  assign ENCLK = net338262;
  assign net338263 = EN;

  DLL_X1 latch ( .D(net338263), .GN(net338260), .Q(net338266) );
  AND2_X1 main_gate ( .A1(net338266), .A2(net338260), .ZN(net338262) );
endmodule


module SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_5 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net338260, net338262, net338263, net338266;
  assign net338260 = CLK;
  assign ENCLK = net338262;
  assign net338263 = EN;

  DLL_X1 latch ( .D(net338263), .GN(net338260), .Q(net338266) );
  AND2_X1 main_gate ( .A1(net338266), .A2(net338260), .ZN(net338262) );
endmodule


module SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_4 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net338260, net338262, net338263, net338266;
  assign net338260 = CLK;
  assign ENCLK = net338262;
  assign net338263 = EN;

  DLL_X1 latch ( .D(net338263), .GN(net338260), .Q(net338266) );
  AND2_X1 main_gate ( .A1(net338266), .A2(net338260), .ZN(net338262) );
endmodule


module SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_3 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net338260, net338262, net338263, net338266;
  assign net338260 = CLK;
  assign ENCLK = net338262;
  assign net338263 = EN;

  DLL_X1 latch ( .D(net338263), .GN(net338260), .Q(net338266) );
  AND2_X1 main_gate ( .A1(net338266), .A2(net338260), .ZN(net338262) );
endmodule


module SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_2 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net338260, net338262, net338263, net338266;
  assign net338260 = CLK;
  assign ENCLK = net338262;
  assign net338263 = EN;

  DLL_X1 latch ( .D(net338263), .GN(net338260), .Q(net338266) );
  AND2_X1 main_gate ( .A1(net338266), .A2(net338260), .ZN(net338262) );
endmodule


module SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_1 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net338260, net338262, net338263, net338266;
  assign net338260 = CLK;
  assign ENCLK = net338262;
  assign net338263 = EN;

  DLL_X1 latch ( .D(net338263), .GN(net338260), .Q(net338266) );
  AND2_X1 main_gate ( .A1(net338266), .A2(net338260), .ZN(net338262) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ff32_en_1 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net338245, net338247, net338248, net338251;
  assign net338245 = CLK;
  assign ENCLK = net338247;
  assign net338248 = EN;

  DLL_X1 latch ( .D(net338248), .GN(net338245), .Q(net338251) );
  AND2_X1 main_gate ( .A1(net338251), .A2(net338245), .ZN(net338247) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dlx_regfile_33 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net338030, net338032, net338033, net338036;
  assign net338030 = CLK;
  assign ENCLK = net338032;
  assign net338033 = EN;

  DLL_X1 latch ( .D(net338033), .GN(net338030), .Q(net338036) );
  AND2_X1 main_gate ( .A1(net338036), .A2(net338030), .ZN(net338032) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dlx_regfile_32 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net338030, net338032, net338033, net338036;
  assign net338030 = CLK;
  assign ENCLK = net338032;
  assign net338033 = EN;

  DLL_X1 latch ( .D(net338033), .GN(net338030), .Q(net338036) );
  AND2_X1 main_gate ( .A1(net338036), .A2(net338030), .ZN(net338032) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dlx_regfile_31 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net338030, net338032, net338033, net338036;
  assign net338030 = CLK;
  assign ENCLK = net338032;
  assign net338033 = EN;

  DLL_X1 latch ( .D(net338033), .GN(net338030), .Q(net338036) );
  AND2_X1 main_gate ( .A1(net338036), .A2(net338030), .ZN(net338032) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dlx_regfile_30 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net338030, net338032, net338033, net338036;
  assign net338030 = CLK;
  assign ENCLK = net338032;
  assign net338033 = EN;

  DLL_X1 latch ( .D(net338033), .GN(net338030), .Q(net338036) );
  AND2_X1 main_gate ( .A1(net338036), .A2(net338030), .ZN(net338032) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dlx_regfile_29 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net338030, net338032, net338033, net338036;
  assign net338030 = CLK;
  assign ENCLK = net338032;
  assign net338033 = EN;

  DLL_X1 latch ( .D(net338033), .GN(net338030), .Q(net338036) );
  AND2_X1 main_gate ( .A1(net338036), .A2(net338030), .ZN(net338032) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dlx_regfile_28 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net338030, net338032, net338033, net338036;
  assign net338030 = CLK;
  assign ENCLK = net338032;
  assign net338033 = EN;

  DLL_X1 latch ( .D(net338033), .GN(net338030), .Q(net338036) );
  AND2_X1 main_gate ( .A1(net338036), .A2(net338030), .ZN(net338032) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dlx_regfile_27 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net338030, net338032, net338033, net338036;
  assign net338030 = CLK;
  assign ENCLK = net338032;
  assign net338033 = EN;

  DLL_X1 latch ( .D(net338033), .GN(net338030), .Q(net338036) );
  AND2_X1 main_gate ( .A1(net338036), .A2(net338030), .ZN(net338032) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dlx_regfile_26 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net338030, net338032, net338033, net338036;
  assign net338030 = CLK;
  assign ENCLK = net338032;
  assign net338033 = EN;

  DLL_X1 latch ( .D(net338033), .GN(net338030), .Q(net338036) );
  AND2_X1 main_gate ( .A1(net338036), .A2(net338030), .ZN(net338032) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dlx_regfile_25 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net338030, net338032, net338033, net338036;
  assign net338030 = CLK;
  assign ENCLK = net338032;
  assign net338033 = EN;

  DLL_X1 latch ( .D(net338033), .GN(net338030), .Q(net338036) );
  AND2_X1 main_gate ( .A1(net338036), .A2(net338030), .ZN(net338032) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dlx_regfile_24 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net338030, net338032, net338033, net338036;
  assign net338030 = CLK;
  assign ENCLK = net338032;
  assign net338033 = EN;

  DLL_X1 latch ( .D(net338033), .GN(net338030), .Q(net338036) );
  AND2_X1 main_gate ( .A1(net338036), .A2(net338030), .ZN(net338032) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dlx_regfile_23 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net338030, net338032, net338033, net338036;
  assign net338030 = CLK;
  assign ENCLK = net338032;
  assign net338033 = EN;

  DLL_X1 latch ( .D(net338033), .GN(net338030), .Q(net338036) );
  AND2_X1 main_gate ( .A1(net338036), .A2(net338030), .ZN(net338032) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dlx_regfile_22 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net338030, net338032, net338033, net338036;
  assign net338030 = CLK;
  assign ENCLK = net338032;
  assign net338033 = EN;

  DLL_X1 latch ( .D(net338033), .GN(net338030), .Q(net338036) );
  AND2_X1 main_gate ( .A1(net338036), .A2(net338030), .ZN(net338032) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dlx_regfile_21 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net338030, net338032, net338033, net338036;
  assign net338030 = CLK;
  assign ENCLK = net338032;
  assign net338033 = EN;

  DLL_X1 latch ( .D(net338033), .GN(net338030), .Q(net338036) );
  AND2_X1 main_gate ( .A1(net338036), .A2(net338030), .ZN(net338032) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dlx_regfile_20 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net338030, net338032, net338033, net338036;
  assign net338030 = CLK;
  assign ENCLK = net338032;
  assign net338033 = EN;

  DLL_X1 latch ( .D(net338033), .GN(net338030), .Q(net338036) );
  AND2_X1 main_gate ( .A1(net338036), .A2(net338030), .ZN(net338032) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dlx_regfile_19 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net338030, net338032, net338033, net338036;
  assign net338030 = CLK;
  assign ENCLK = net338032;
  assign net338033 = EN;

  DLL_X1 latch ( .D(net338033), .GN(net338030), .Q(net338036) );
  AND2_X1 main_gate ( .A1(net338036), .A2(net338030), .ZN(net338032) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dlx_regfile_18 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net338030, net338032, net338033, net338036;
  assign net338030 = CLK;
  assign ENCLK = net338032;
  assign net338033 = EN;

  DLL_X1 latch ( .D(net338033), .GN(net338030), .Q(net338036) );
  AND2_X1 main_gate ( .A1(net338036), .A2(net338030), .ZN(net338032) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dlx_regfile_17 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net338030, net338032, net338033, net338036;
  assign net338030 = CLK;
  assign ENCLK = net338032;
  assign net338033 = EN;

  DLL_X1 latch ( .D(net338033), .GN(net338030), .Q(net338036) );
  AND2_X1 main_gate ( .A1(net338036), .A2(net338030), .ZN(net338032) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dlx_regfile_16 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net338030, net338032, net338033, net338036;
  assign net338030 = CLK;
  assign ENCLK = net338032;
  assign net338033 = EN;

  DLL_X1 latch ( .D(net338033), .GN(net338030), .Q(net338036) );
  AND2_X1 main_gate ( .A1(net338036), .A2(net338030), .ZN(net338032) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dlx_regfile_15 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net338030, net338032, net338033, net338036;
  assign net338030 = CLK;
  assign ENCLK = net338032;
  assign net338033 = EN;

  DLL_X1 latch ( .D(net338033), .GN(net338030), .Q(net338036) );
  AND2_X1 main_gate ( .A1(net338036), .A2(net338030), .ZN(net338032) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dlx_regfile_14 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net338030, net338032, net338033, net338036;
  assign net338030 = CLK;
  assign ENCLK = net338032;
  assign net338033 = EN;

  DLL_X1 latch ( .D(net338033), .GN(net338030), .Q(net338036) );
  AND2_X1 main_gate ( .A1(net338036), .A2(net338030), .ZN(net338032) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dlx_regfile_13 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net338030, net338032, net338033, net338036;
  assign net338030 = CLK;
  assign ENCLK = net338032;
  assign net338033 = EN;

  DLL_X1 latch ( .D(net338033), .GN(net338030), .Q(net338036) );
  AND2_X1 main_gate ( .A1(net338036), .A2(net338030), .ZN(net338032) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dlx_regfile_12 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net338030, net338032, net338033, net338036;
  assign net338030 = CLK;
  assign ENCLK = net338032;
  assign net338033 = EN;

  DLL_X1 latch ( .D(net338033), .GN(net338030), .Q(net338036) );
  AND2_X1 main_gate ( .A1(net338036), .A2(net338030), .ZN(net338032) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dlx_regfile_11 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net338030, net338032, net338033, net338036;
  assign net338030 = CLK;
  assign ENCLK = net338032;
  assign net338033 = EN;

  DLL_X1 latch ( .D(net338033), .GN(net338030), .Q(net338036) );
  AND2_X1 main_gate ( .A1(net338036), .A2(net338030), .ZN(net338032) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dlx_regfile_10 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net338030, net338032, net338033, net338036;
  assign net338030 = CLK;
  assign ENCLK = net338032;
  assign net338033 = EN;

  DLL_X1 latch ( .D(net338033), .GN(net338030), .Q(net338036) );
  AND2_X1 main_gate ( .A1(net338036), .A2(net338030), .ZN(net338032) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dlx_regfile_9 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net338030, net338032, net338033, net338036;
  assign net338030 = CLK;
  assign ENCLK = net338032;
  assign net338033 = EN;

  DLL_X1 latch ( .D(net338033), .GN(net338030), .Q(net338036) );
  AND2_X1 main_gate ( .A1(net338036), .A2(net338030), .ZN(net338032) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dlx_regfile_8 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net338030, net338032, net338033, net338036;
  assign net338030 = CLK;
  assign ENCLK = net338032;
  assign net338033 = EN;

  DLL_X1 latch ( .D(net338033), .GN(net338030), .Q(net338036) );
  AND2_X1 main_gate ( .A1(net338036), .A2(net338030), .ZN(net338032) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dlx_regfile_7 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net338030, net338032, net338033, net338036;
  assign net338030 = CLK;
  assign ENCLK = net338032;
  assign net338033 = EN;

  DLL_X1 latch ( .D(net338033), .GN(net338030), .Q(net338036) );
  AND2_X1 main_gate ( .A1(net338036), .A2(net338030), .ZN(net338032) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dlx_regfile_6 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net338030, net338032, net338033, net338036;
  assign net338030 = CLK;
  assign ENCLK = net338032;
  assign net338033 = EN;

  DLL_X1 latch ( .D(net338033), .GN(net338030), .Q(net338036) );
  AND2_X1 main_gate ( .A1(net338036), .A2(net338030), .ZN(net338032) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dlx_regfile_5 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net338030, net338032, net338033, net338036;
  assign net338030 = CLK;
  assign ENCLK = net338032;
  assign net338033 = EN;

  DLL_X1 latch ( .D(net338033), .GN(net338030), .Q(net338036) );
  AND2_X1 main_gate ( .A1(net338036), .A2(net338030), .ZN(net338032) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dlx_regfile_4 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net338030, net338032, net338033, net338036;
  assign net338030 = CLK;
  assign ENCLK = net338032;
  assign net338033 = EN;

  DLL_X1 latch ( .D(net338033), .GN(net338030), .Q(net338036) );
  AND2_X1 main_gate ( .A1(net338036), .A2(net338030), .ZN(net338032) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dlx_regfile_3 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net338030, net338032, net338033, net338036;
  assign net338030 = CLK;
  assign ENCLK = net338032;
  assign net338033 = EN;

  DLL_X1 latch ( .D(net338033), .GN(net338030), .Q(net338036) );
  AND2_X1 main_gate ( .A1(net338036), .A2(net338030), .ZN(net338032) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dlx_regfile_2 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net338030, net338032, net338033, net338036;
  assign net338030 = CLK;
  assign ENCLK = net338032;
  assign net338033 = EN;

  DLL_X1 latch ( .D(net338033), .GN(net338030), .Q(net338036) );
  AND2_X1 main_gate ( .A1(net338036), .A2(net338030), .ZN(net338032) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dlx_regfile_1 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net338030, net338032, net338033, net338036;
  assign net338030 = CLK;
  assign ENCLK = net338032;
  assign net338033 = EN;

  DLL_X1 latch ( .D(net338033), .GN(net338030), .Q(net338036) );
  AND2_X1 main_gate ( .A1(net338036), .A2(net338030), .ZN(net338032) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ff32_en_SIZE5_3 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net338000, net338002, net338003, net338006;
  assign net338000 = CLK;
  assign ENCLK = net338002;
  assign net338003 = EN;

  DLL_X1 latch ( .D(net338003), .GN(net338000), .Q(net338006) );
  AND2_X1 main_gate ( .A1(net338006), .A2(net338000), .ZN(net338002) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ff32_en_SIZE5_2 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net338000, net338002, net338003, net338006;
  assign net338000 = CLK;
  assign ENCLK = net338002;
  assign net338003 = EN;

  DLL_X1 latch ( .D(net338003), .GN(net338000), .Q(net338006) );
  AND2_X1 main_gate ( .A1(net338006), .A2(net338000), .ZN(net338002) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ff32_en_SIZE32_5 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net337985, net337987, net337988, net337991;
  assign net337985 = CLK;
  assign ENCLK = net337987;
  assign net337988 = EN;

  DLL_X1 latch ( .D(net337988), .GN(net337985), .Q(net337991) );
  AND2_X1 main_gate ( .A1(net337991), .A2(net337985), .ZN(net337987) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ff32_en_SIZE32_4 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net337985, net337987, net337988, net337991;
  assign net337985 = CLK;
  assign ENCLK = net337987;
  assign net337988 = EN;

  DLL_X1 latch ( .D(net337988), .GN(net337985), .Q(net337991) );
  AND2_X1 main_gate ( .A1(net337991), .A2(net337985), .ZN(net337987) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ff32_en_SIZE32_1 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net337985, net337987, net337988, net337991;
  assign net337985 = CLK;
  assign ENCLK = net337987;
  assign net337988 = EN;

  DLL_X1 latch ( .D(net337988), .GN(net337985), .Q(net337991) );
  AND2_X1 main_gate ( .A1(net337991), .A2(net337985), .ZN(net337987) );
endmodule


module FA_127 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6;

  OAI21_X1 U5 ( .B1(Ci), .B2(B), .A(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(B), .A2(Ci), .ZN(n4) );
  NAND2_X1 U3 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n6) );
  XNOR2_X1 U1 ( .A(n6), .B(B), .ZN(S) );
endmodule


module FA_126 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6;

  OAI21_X1 U5 ( .B1(Ci), .B2(B), .A(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(B), .A2(Ci), .ZN(n4) );
  NAND2_X1 U3 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n6) );
  XNOR2_X1 U1 ( .A(n6), .B(B), .ZN(S) );
endmodule


module FA_125 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2;

  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n2) );
  XNOR2_X1 U1 ( .A(n2), .B(B), .ZN(S) );
endmodule


module FA_120 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(S) );
  AND2_X1 U2 ( .A1(B), .A2(A), .ZN(Co) );
endmodule


module FA_119 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6;

  OAI21_X1 U5 ( .B1(Ci), .B2(B), .A(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(B), .A2(Ci), .ZN(n4) );
  NAND2_X1 U3 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n6) );
  XNOR2_X1 U1 ( .A(n6), .B(B), .ZN(S) );
endmodule


module FA_118 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6;

  OAI21_X1 U5 ( .B1(Ci), .B2(B), .A(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(B), .A2(Ci), .ZN(n4) );
  NAND2_X1 U3 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n6) );
  XNOR2_X1 U1 ( .A(n6), .B(B), .ZN(S) );
endmodule


module FA_117 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2;

  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n2) );
  XNOR2_X1 U1 ( .A(n2), .B(B), .ZN(S) );
endmodule


module FA_116 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(S) );
  OR2_X1 U2 ( .A1(A), .A2(B), .ZN(Co) );
endmodule


module FA_115 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6;

  OAI21_X1 U5 ( .B1(Ci), .B2(B), .A(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(B), .A2(Ci), .ZN(n4) );
  NAND2_X1 U3 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n6) );
  XNOR2_X1 U1 ( .A(n6), .B(B), .ZN(S) );
endmodule


module FA_114 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6;

  OAI21_X1 U5 ( .B1(Ci), .B2(B), .A(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(B), .A2(Ci), .ZN(n4) );
  NAND2_X1 U3 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n6) );
  XNOR2_X1 U1 ( .A(n6), .B(B), .ZN(S) );
endmodule


module FA_113 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2;

  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n2) );
  XNOR2_X1 U1 ( .A(n2), .B(B), .ZN(S) );
endmodule


module FA_112 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(S) );
  AND2_X1 U2 ( .A1(B), .A2(A), .ZN(Co) );
endmodule


module FA_111 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6;

  OAI21_X1 U5 ( .B1(Ci), .B2(B), .A(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(B), .A2(Ci), .ZN(n4) );
  NAND2_X1 U3 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n6) );
  XNOR2_X1 U1 ( .A(n6), .B(B), .ZN(S) );
endmodule


module FA_110 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6;

  OAI21_X1 U5 ( .B1(Ci), .B2(B), .A(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(B), .A2(Ci), .ZN(n4) );
  NAND2_X1 U3 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n6) );
  XNOR2_X1 U1 ( .A(n6), .B(B), .ZN(S) );
endmodule


module FA_109 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2;

  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n2) );
  XNOR2_X1 U1 ( .A(n2), .B(B), .ZN(S) );
endmodule


module FA_108 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(S) );
endmodule


module FA_107 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6;

  OAI21_X1 U5 ( .B1(Ci), .B2(B), .A(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(B), .A2(Ci), .ZN(n4) );
  NAND2_X1 U3 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n6) );
  XNOR2_X1 U1 ( .A(n6), .B(B), .ZN(S) );
endmodule


module FA_106 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6;

  OAI21_X1 U5 ( .B1(Ci), .B2(B), .A(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(B), .A2(Ci), .ZN(n4) );
  NAND2_X1 U3 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n6) );
  XNOR2_X1 U1 ( .A(n6), .B(B), .ZN(S) );
endmodule


module FA_105 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2;

  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n2) );
  XNOR2_X1 U1 ( .A(n2), .B(B), .ZN(S) );
endmodule


module FA_104 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(S) );
  AND2_X1 U2 ( .A1(B), .A2(A), .ZN(Co) );
endmodule


module FA_103 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6;

  OAI21_X1 U5 ( .B1(Ci), .B2(B), .A(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(B), .A2(Ci), .ZN(n4) );
  NAND2_X1 U3 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n6) );
  XNOR2_X1 U1 ( .A(n6), .B(B), .ZN(S) );
endmodule


module FA_102 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6;

  OAI21_X1 U5 ( .B1(Ci), .B2(B), .A(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(B), .A2(Ci), .ZN(n4) );
  NAND2_X1 U3 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n6) );
  XNOR2_X1 U1 ( .A(n6), .B(B), .ZN(S) );
endmodule


module FA_101 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2;

  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n2) );
  XNOR2_X1 U1 ( .A(n2), .B(B), .ZN(S) );
endmodule


module FA_100 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(S) );
  OR2_X1 U2 ( .A1(A), .A2(B), .ZN(Co) );
endmodule


module FA_99 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6;

  OAI21_X1 U5 ( .B1(Ci), .B2(B), .A(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(B), .A2(Ci), .ZN(n4) );
  NAND2_X1 U3 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n6) );
  XNOR2_X1 U1 ( .A(n6), .B(B), .ZN(S) );
endmodule


module FA_98 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6;

  OAI21_X1 U5 ( .B1(Ci), .B2(B), .A(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(B), .A2(Ci), .ZN(n4) );
  NAND2_X1 U3 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n6) );
  XNOR2_X1 U1 ( .A(n6), .B(B), .ZN(S) );
endmodule


module FA_97 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2;

  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n2) );
  XNOR2_X1 U1 ( .A(n2), .B(B), .ZN(S) );
endmodule


module FA_96 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(S) );
  AND2_X1 U2 ( .A1(B), .A2(A), .ZN(Co) );
endmodule


module FA_95 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6;

  OAI21_X1 U5 ( .B1(Ci), .B2(B), .A(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(B), .A2(Ci), .ZN(n4) );
  NAND2_X1 U3 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n6) );
  XNOR2_X1 U1 ( .A(n6), .B(B), .ZN(S) );
endmodule


module FA_94 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6;

  OAI21_X1 U5 ( .B1(Ci), .B2(B), .A(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(B), .A2(Ci), .ZN(n4) );
  NAND2_X1 U3 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n6) );
  XNOR2_X1 U1 ( .A(n6), .B(B), .ZN(S) );
endmodule


module FA_93 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2;

  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n2) );
  XNOR2_X1 U1 ( .A(n2), .B(B), .ZN(S) );
endmodule


module FA_92 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  NAND2_X1 U3 ( .A1(n3), .A2(n1), .ZN(Co) );
  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(S) );
  INV_X1 U2 ( .A(B), .ZN(n1) );
  INV_X1 U4 ( .A(A), .ZN(n3) );
endmodule


module FA_91 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6;

  OAI21_X1 U5 ( .B1(Ci), .B2(B), .A(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(B), .A2(Ci), .ZN(n4) );
  NAND2_X1 U3 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n6) );
  XNOR2_X1 U1 ( .A(n6), .B(B), .ZN(S) );
endmodule


module FA_90 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6;

  OAI21_X1 U5 ( .B1(Ci), .B2(B), .A(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(B), .A2(Ci), .ZN(n4) );
  NAND2_X1 U3 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n6) );
  XNOR2_X1 U1 ( .A(n6), .B(B), .ZN(S) );
endmodule


module FA_89 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2;

  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n2) );
  XNOR2_X1 U1 ( .A(n2), .B(B), .ZN(S) );
endmodule


module FA_88 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(S) );
  AND2_X1 U2 ( .A1(B), .A2(A), .ZN(Co) );
endmodule


module FA_87 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6;

  OAI21_X1 U5 ( .B1(Ci), .B2(B), .A(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(B), .A2(Ci), .ZN(n4) );
  NAND2_X1 U3 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n6) );
  XNOR2_X1 U1 ( .A(n6), .B(B), .ZN(S) );
endmodule


module FA_86 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6;

  OAI21_X1 U5 ( .B1(Ci), .B2(B), .A(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(B), .A2(Ci), .ZN(n4) );
  NAND2_X1 U3 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n6) );
  XNOR2_X1 U1 ( .A(n6), .B(B), .ZN(S) );
endmodule


module FA_85 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2;

  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n2) );
  XNOR2_X1 U1 ( .A(n2), .B(B), .ZN(S) );
endmodule


module FA_84 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Co) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(S) );
endmodule


module FA_83 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6;

  OAI21_X1 U5 ( .B1(Ci), .B2(B), .A(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(B), .A2(Ci), .ZN(n4) );
  NAND2_X1 U3 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n6) );
  XNOR2_X1 U1 ( .A(n6), .B(B), .ZN(S) );
endmodule


module FA_82 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6;

  OAI21_X1 U5 ( .B1(Ci), .B2(B), .A(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(B), .A2(Ci), .ZN(n4) );
  NAND2_X1 U3 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n6) );
  XNOR2_X1 U1 ( .A(n6), .B(B), .ZN(S) );
endmodule


module FA_81 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2;

  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n2) );
  XNOR2_X1 U1 ( .A(n2), .B(B), .ZN(S) );
endmodule


module FA_80 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(S) );
  AND2_X1 U2 ( .A1(B), .A2(A), .ZN(Co) );
endmodule


module FA_79 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6;

  OAI21_X1 U5 ( .B1(Ci), .B2(B), .A(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(B), .A2(Ci), .ZN(n4) );
  NAND2_X1 U3 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n6) );
  XNOR2_X1 U1 ( .A(n6), .B(B), .ZN(S) );
endmodule


module FA_78 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6;

  OAI21_X1 U5 ( .B1(Ci), .B2(B), .A(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(B), .A2(Ci), .ZN(n4) );
  NAND2_X1 U3 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n6) );
  XNOR2_X1 U1 ( .A(n6), .B(B), .ZN(S) );
endmodule


module FA_77 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2;

  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n2) );
  XNOR2_X1 U1 ( .A(n2), .B(B), .ZN(S) );
endmodule


module FA_76 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(S) );
endmodule


module FA_75 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6;

  OAI21_X1 U5 ( .B1(Ci), .B2(B), .A(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(B), .A2(Ci), .ZN(n4) );
  NAND2_X1 U3 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n6) );
  XNOR2_X1 U1 ( .A(n6), .B(B), .ZN(S) );
endmodule


module FA_74 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6;

  OAI21_X1 U5 ( .B1(Ci), .B2(B), .A(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(B), .A2(Ci), .ZN(n4) );
  NAND2_X1 U3 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n6) );
  XNOR2_X1 U1 ( .A(n6), .B(B), .ZN(S) );
endmodule


module FA_73 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2;

  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n2) );
  XNOR2_X1 U1 ( .A(n2), .B(B), .ZN(S) );
endmodule


module FA_72 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(S) );
  AND2_X1 U2 ( .A1(B), .A2(A), .ZN(Co) );
endmodule


module FA_71 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6;

  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n6) );
  XNOR2_X1 U1 ( .A(n6), .B(B), .ZN(S) );
  OAI21_X1 U5 ( .B1(Ci), .B2(B), .A(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(B), .A2(Ci), .ZN(n4) );
  NAND2_X1 U3 ( .A1(n5), .A2(n4), .ZN(Co) );
endmodule


module FA_70 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6;

  OAI21_X1 U5 ( .B1(Ci), .B2(B), .A(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(B), .A2(Ci), .ZN(n4) );
  NAND2_X1 U3 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n6) );
  XNOR2_X1 U1 ( .A(n6), .B(B), .ZN(S) );
endmodule


module FA_69 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2;

  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n2) );
  XNOR2_X1 U1 ( .A(n2), .B(B), .ZN(S) );
endmodule


module FA_68 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Co) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(S) );
endmodule


module FA_67 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6;

  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n6) );
  XNOR2_X1 U1 ( .A(n6), .B(B), .ZN(S) );
  OAI21_X1 U5 ( .B1(Ci), .B2(B), .A(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(B), .A2(Ci), .ZN(n4) );
  NAND2_X1 U3 ( .A1(n5), .A2(n4), .ZN(Co) );
endmodule


module FA_66 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6;

  OAI21_X1 U5 ( .B1(Ci), .B2(B), .A(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(B), .A2(Ci), .ZN(n4) );
  NAND2_X1 U3 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n6) );
  XNOR2_X1 U1 ( .A(n6), .B(B), .ZN(S) );
endmodule


module FA_65 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2;

  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n2) );
  XNOR2_X1 U1 ( .A(n2), .B(B), .ZN(S) );
endmodule


module FA_64 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(S) );
  AND2_X1 U2 ( .A1(B), .A2(A), .ZN(Co) );
endmodule


module FA_63 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6;

  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n6) );
  XNOR2_X1 U1 ( .A(n6), .B(B), .ZN(S) );
  OAI21_X1 U5 ( .B1(Ci), .B2(B), .A(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(B), .A2(Ci), .ZN(n4) );
  NAND2_X1 U3 ( .A1(n5), .A2(n4), .ZN(Co) );
endmodule


module FA_62 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6;

  OAI21_X1 U5 ( .B1(Ci), .B2(B), .A(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(B), .A2(Ci), .ZN(n4) );
  NAND2_X1 U3 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n6) );
  XNOR2_X1 U1 ( .A(n6), .B(B), .ZN(S) );
endmodule


module FA_61 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2;

  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n2) );
  XNOR2_X1 U1 ( .A(n2), .B(B), .ZN(S) );
endmodule


module FA_60 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Co) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(S) );
endmodule


module FA_59 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6;

  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n6) );
  XNOR2_X1 U1 ( .A(n6), .B(B), .ZN(S) );
  OAI21_X1 U5 ( .B1(Ci), .B2(B), .A(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(B), .A2(Ci), .ZN(n4) );
  NAND2_X1 U3 ( .A1(n5), .A2(n4), .ZN(Co) );
endmodule


module FA_58 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6;

  OAI21_X1 U5 ( .B1(Ci), .B2(B), .A(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(B), .A2(Ci), .ZN(n4) );
  NAND2_X1 U3 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n6) );
  XNOR2_X1 U1 ( .A(n6), .B(B), .ZN(S) );
endmodule


module FA_57 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2;

  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n2) );
  XNOR2_X1 U1 ( .A(n2), .B(B), .ZN(S) );
endmodule


module FA_56 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(S) );
  AND2_X1 U2 ( .A1(B), .A2(A), .ZN(Co) );
endmodule


module FA_55 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6;

  OAI21_X1 U5 ( .B1(Ci), .B2(B), .A(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(B), .A2(Ci), .ZN(n4) );
  NAND2_X1 U3 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n6) );
  XNOR2_X1 U1 ( .A(n6), .B(B), .ZN(S) );
endmodule


module FA_54 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6;

  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n6) );
  XNOR2_X1 U1 ( .A(n6), .B(B), .ZN(S) );
  OAI21_X1 U5 ( .B1(Ci), .B2(B), .A(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(B), .A2(Ci), .ZN(n4) );
  NAND2_X1 U3 ( .A1(n5), .A2(n4), .ZN(Co) );
endmodule


module FA_53 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2;

  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n2) );
  XNOR2_X1 U1 ( .A(n2), .B(B), .ZN(S) );
endmodule


module FA_52 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Co) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(S) );
endmodule


module FA_51 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6;

  OAI21_X1 U5 ( .B1(Ci), .B2(B), .A(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(B), .A2(Ci), .ZN(n4) );
  NAND2_X1 U3 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n6) );
  XNOR2_X1 U1 ( .A(n6), .B(B), .ZN(S) );
endmodule


module FA_50 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6;

  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n6) );
  XNOR2_X1 U1 ( .A(n6), .B(B), .ZN(S) );
  OAI21_X1 U5 ( .B1(Ci), .B2(B), .A(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(B), .A2(Ci), .ZN(n4) );
  NAND2_X1 U3 ( .A1(n5), .A2(n4), .ZN(Co) );
endmodule


module FA_49 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2;

  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n2) );
  XNOR2_X1 U1 ( .A(n2), .B(B), .ZN(S) );
endmodule


module FA_48 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(S) );
  AND2_X1 U2 ( .A1(B), .A2(A), .ZN(Co) );
endmodule


module FA_47 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6;

  OAI21_X1 U5 ( .B1(Ci), .B2(B), .A(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(B), .A2(Ci), .ZN(n4) );
  NAND2_X1 U3 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n6) );
  XNOR2_X1 U1 ( .A(n6), .B(B), .ZN(S) );
endmodule


module FA_46 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6;

  OAI21_X1 U5 ( .B1(Ci), .B2(B), .A(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(B), .A2(Ci), .ZN(n4) );
  NAND2_X1 U3 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n6) );
  XNOR2_X1 U1 ( .A(n6), .B(B), .ZN(S) );
endmodule


module FA_45 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2;

  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n2) );
  XNOR2_X1 U1 ( .A(n2), .B(B), .ZN(S) );
endmodule


module FA_44 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(S) );
endmodule


module FA_43 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6;

  OAI21_X1 U5 ( .B1(Ci), .B2(B), .A(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(B), .A2(Ci), .ZN(n4) );
  NAND2_X1 U3 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n6) );
  XNOR2_X1 U1 ( .A(n6), .B(B), .ZN(S) );
endmodule


module FA_42 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6;

  OAI21_X1 U5 ( .B1(Ci), .B2(B), .A(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(B), .A2(Ci), .ZN(n4) );
  NAND2_X1 U3 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n6) );
  XNOR2_X1 U1 ( .A(n6), .B(B), .ZN(S) );
endmodule


module FA_41 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2;

  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n2) );
  XNOR2_X1 U1 ( .A(n2), .B(B), .ZN(S) );
endmodule


module FA_40 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(S) );
  AND2_X1 U2 ( .A1(B), .A2(A), .ZN(Co) );
endmodule


module FA_39 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6;

  OAI21_X1 U5 ( .B1(Ci), .B2(B), .A(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(B), .A2(Ci), .ZN(n4) );
  NAND2_X1 U3 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n6) );
  XNOR2_X1 U1 ( .A(n6), .B(B), .ZN(S) );
endmodule


module FA_38 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6;

  OAI21_X1 U5 ( .B1(Ci), .B2(B), .A(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(B), .A2(Ci), .ZN(n4) );
  NAND2_X1 U3 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n6) );
  XNOR2_X1 U1 ( .A(n6), .B(B), .ZN(S) );
endmodule


module FA_37 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2;

  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n2) );
  XNOR2_X1 U1 ( .A(n2), .B(B), .ZN(S) );
endmodule


module FA_36 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n3;

  NAND2_X1 U3 ( .A1(n3), .A2(n1), .ZN(Co) );
  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(S) );
  INV_X1 U2 ( .A(B), .ZN(n1) );
  INV_X1 U4 ( .A(A), .ZN(n3) );
endmodule


module FA_35 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6;

  OAI21_X1 U5 ( .B1(Ci), .B2(B), .A(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(B), .A2(Ci), .ZN(n4) );
  NAND2_X1 U3 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n6) );
  XNOR2_X1 U1 ( .A(n6), .B(B), .ZN(S) );
endmodule


module FA_34 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6;

  OAI21_X1 U5 ( .B1(Ci), .B2(B), .A(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(B), .A2(Ci), .ZN(n4) );
  NAND2_X1 U3 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n6) );
  XNOR2_X1 U1 ( .A(n6), .B(B), .ZN(S) );
endmodule


module FA_33 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2;

  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n2) );
  XNOR2_X1 U1 ( .A(n2), .B(B), .ZN(S) );
endmodule


module FA_32 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(S) );
  AND2_X1 U2 ( .A1(B), .A2(A), .ZN(Co) );
endmodule


module FA_31 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6;

  OAI21_X1 U5 ( .B1(Ci), .B2(B), .A(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(B), .A2(Ci), .ZN(n4) );
  NAND2_X1 U3 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n6) );
  XNOR2_X1 U1 ( .A(n6), .B(B), .ZN(S) );
endmodule


module FA_30 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6;

  OAI21_X1 U5 ( .B1(Ci), .B2(B), .A(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(B), .A2(Ci), .ZN(n4) );
  NAND2_X1 U3 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n6) );
  XNOR2_X1 U1 ( .A(n6), .B(B), .ZN(S) );
endmodule


module FA_29 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2;

  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n2) );
  XNOR2_X1 U1 ( .A(n2), .B(B), .ZN(S) );
endmodule


module FA_28 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(S) );
endmodule


module FA_27 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6;

  OAI21_X1 U5 ( .B1(Ci), .B2(B), .A(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(B), .A2(Ci), .ZN(n4) );
  NAND2_X1 U3 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n6) );
  XNOR2_X1 U1 ( .A(n6), .B(B), .ZN(S) );
endmodule


module FA_26 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6;

  OAI21_X1 U5 ( .B1(Ci), .B2(B), .A(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(B), .A2(Ci), .ZN(n4) );
  NAND2_X1 U3 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n6) );
  XNOR2_X1 U1 ( .A(n6), .B(B), .ZN(S) );
endmodule


module FA_25 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2;

  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n2) );
  XNOR2_X1 U1 ( .A(n2), .B(B), .ZN(S) );
endmodule


module FA_24 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(S) );
  AND2_X1 U2 ( .A1(B), .A2(A), .ZN(Co) );
endmodule


module FA_23 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6;

  OAI21_X1 U5 ( .B1(Ci), .B2(B), .A(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(B), .A2(Ci), .ZN(n4) );
  NAND2_X1 U3 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n6) );
  XNOR2_X1 U1 ( .A(n6), .B(B), .ZN(S) );
endmodule


module FA_22 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6;

  OAI21_X1 U5 ( .B1(Ci), .B2(B), .A(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(B), .A2(Ci), .ZN(n4) );
  NAND2_X1 U3 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n6) );
  XNOR2_X1 U1 ( .A(n6), .B(B), .ZN(S) );
endmodule


module FA_21 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2;

  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n2) );
  XNOR2_X1 U1 ( .A(n2), .B(B), .ZN(S) );
endmodule


module FA_20 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(S) );
endmodule


module FA_19 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6;

  OAI21_X1 U5 ( .B1(Ci), .B2(B), .A(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(B), .A2(Ci), .ZN(n4) );
  NAND2_X1 U3 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n6) );
  XNOR2_X1 U1 ( .A(n6), .B(B), .ZN(S) );
endmodule


module FA_18 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6;

  OAI21_X1 U5 ( .B1(Ci), .B2(B), .A(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(B), .A2(Ci), .ZN(n4) );
  NAND2_X1 U3 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n6) );
  XNOR2_X1 U1 ( .A(n6), .B(B), .ZN(S) );
endmodule


module FA_17 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2;

  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n2) );
  XNOR2_X1 U1 ( .A(n2), .B(B), .ZN(S) );
endmodule


module FA_16 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(S) );
  AND2_X1 U2 ( .A1(B), .A2(A), .ZN(Co) );
endmodule


module FA_15 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6;

  OAI21_X1 U5 ( .B1(Ci), .B2(B), .A(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(B), .A2(Ci), .ZN(n4) );
  NAND2_X1 U3 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n6) );
  XNOR2_X1 U1 ( .A(n6), .B(B), .ZN(S) );
endmodule


module FA_14 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6;

  OAI21_X1 U5 ( .B1(Ci), .B2(B), .A(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(B), .A2(Ci), .ZN(n4) );
  NAND2_X1 U3 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n6) );
  XNOR2_X1 U1 ( .A(n6), .B(B), .ZN(S) );
endmodule


module FA_13 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2;

  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n2) );
  XNOR2_X1 U1 ( .A(n2), .B(B), .ZN(S) );
endmodule


module FA_12 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(S) );
endmodule


module FA_11 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6;

  OAI21_X1 U5 ( .B1(Ci), .B2(B), .A(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(B), .A2(Ci), .ZN(n4) );
  NAND2_X1 U3 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n6) );
  XNOR2_X1 U1 ( .A(n6), .B(B), .ZN(S) );
endmodule


module FA_10 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6;

  OAI21_X1 U5 ( .B1(Ci), .B2(B), .A(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(B), .A2(Ci), .ZN(n4) );
  NAND2_X1 U3 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n6) );
  XNOR2_X1 U1 ( .A(n6), .B(B), .ZN(S) );
endmodule


module FA_9 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2;

  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n2) );
  XNOR2_X1 U1 ( .A(n2), .B(B), .ZN(S) );
endmodule


module FA_8 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(S) );
  AND2_X1 U2 ( .A1(B), .A2(A), .ZN(Co) );
endmodule


module FA_7 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6;

  OAI21_X1 U5 ( .B1(Ci), .B2(B), .A(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(B), .A2(Ci), .ZN(n4) );
  NAND2_X1 U3 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n6) );
  XNOR2_X1 U1 ( .A(n6), .B(B), .ZN(S) );
endmodule


module FA_6 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6;

  OAI21_X1 U5 ( .B1(Ci), .B2(B), .A(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(B), .A2(Ci), .ZN(n4) );
  NAND2_X1 U3 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n6) );
  XNOR2_X1 U1 ( .A(n6), .B(B), .ZN(S) );
endmodule


module FA_5 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2;

  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n2) );
  XNOR2_X1 U1 ( .A(n2), .B(B), .ZN(S) );
endmodule


module FA_4 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(S) );
endmodule


module FA_3 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6;

  OAI21_X1 U5 ( .B1(Ci), .B2(B), .A(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(B), .A2(Ci), .ZN(n4) );
  NAND2_X1 U3 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n6) );
  XNOR2_X1 U1 ( .A(n6), .B(B), .ZN(S) );
endmodule


module FA_2 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5, n6;

  OAI21_X1 U5 ( .B1(Ci), .B2(B), .A(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(B), .A2(Ci), .ZN(n4) );
  NAND2_X1 U3 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n6) );
  XNOR2_X1 U1 ( .A(n6), .B(B), .ZN(S) );
endmodule


module FA_1 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2;

  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n2) );
  XNOR2_X1 U1 ( .A(n2), .B(B), .ZN(S) );
endmodule


module mux21_SIZE4_15 ( IN0, IN1, CTRL, OUT1 );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] OUT1;
  input CTRL;


  MUX2_X1 U1 ( .A(IN0[3]), .B(IN1[3]), .S(CTRL), .Z(OUT1[3]) );
  MUX2_X1 U2 ( .A(IN0[2]), .B(IN1[2]), .S(CTRL), .Z(OUT1[2]) );
  MUX2_X1 U3 ( .A(IN0[1]), .B(IN1[1]), .S(CTRL), .Z(OUT1[1]) );
  MUX2_X1 U4 ( .A(IN0[0]), .B(IN1[0]), .S(CTRL), .Z(OUT1[0]) );
endmodule


module mux21_SIZE4_14 ( IN0, IN1, CTRL, OUT1 );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] OUT1;
  input CTRL;


  MUX2_X1 U1 ( .A(IN0[3]), .B(IN1[3]), .S(CTRL), .Z(OUT1[3]) );
  MUX2_X1 U2 ( .A(IN0[2]), .B(IN1[2]), .S(CTRL), .Z(OUT1[2]) );
  MUX2_X1 U3 ( .A(IN0[1]), .B(IN1[1]), .S(CTRL), .Z(OUT1[1]) );
  MUX2_X1 U4 ( .A(IN0[0]), .B(IN1[0]), .S(CTRL), .Z(OUT1[0]) );
endmodule


module mux21_SIZE4_13 ( IN0, IN1, CTRL, OUT1 );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] OUT1;
  input CTRL;


  MUX2_X1 U1 ( .A(IN0[3]), .B(IN1[3]), .S(CTRL), .Z(OUT1[3]) );
  MUX2_X1 U2 ( .A(IN0[2]), .B(IN1[2]), .S(CTRL), .Z(OUT1[2]) );
  MUX2_X1 U3 ( .A(IN0[1]), .B(IN1[1]), .S(CTRL), .Z(OUT1[1]) );
  MUX2_X1 U4 ( .A(IN0[0]), .B(IN1[0]), .S(CTRL), .Z(OUT1[0]) );
endmodule


module mux21_SIZE4_12 ( IN0, IN1, CTRL, OUT1 );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] OUT1;
  input CTRL;


  MUX2_X1 U1 ( .A(IN0[3]), .B(IN1[3]), .S(CTRL), .Z(OUT1[3]) );
  MUX2_X1 U2 ( .A(IN0[2]), .B(IN1[2]), .S(CTRL), .Z(OUT1[2]) );
  MUX2_X1 U3 ( .A(IN0[1]), .B(IN1[1]), .S(CTRL), .Z(OUT1[1]) );
  MUX2_X1 U4 ( .A(IN0[0]), .B(IN1[0]), .S(CTRL), .Z(OUT1[0]) );
endmodule


module mux21_SIZE4_11 ( IN0, IN1, CTRL, OUT1 );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] OUT1;
  input CTRL;


  MUX2_X1 U1 ( .A(IN0[3]), .B(IN1[3]), .S(CTRL), .Z(OUT1[3]) );
  MUX2_X1 U2 ( .A(IN0[2]), .B(IN1[2]), .S(CTRL), .Z(OUT1[2]) );
  MUX2_X1 U3 ( .A(IN0[1]), .B(IN1[1]), .S(CTRL), .Z(OUT1[1]) );
  MUX2_X1 U4 ( .A(IN0[0]), .B(IN1[0]), .S(CTRL), .Z(OUT1[0]) );
endmodule


module mux21_SIZE4_10 ( IN0, IN1, CTRL, OUT1 );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] OUT1;
  input CTRL;


  MUX2_X1 U1 ( .A(IN0[3]), .B(IN1[3]), .S(CTRL), .Z(OUT1[3]) );
  MUX2_X1 U2 ( .A(IN0[2]), .B(IN1[2]), .S(CTRL), .Z(OUT1[2]) );
  MUX2_X1 U3 ( .A(IN0[1]), .B(IN1[1]), .S(CTRL), .Z(OUT1[1]) );
  MUX2_X1 U4 ( .A(IN0[0]), .B(IN1[0]), .S(CTRL), .Z(OUT1[0]) );
endmodule


module mux21_SIZE4_9 ( IN0, IN1, CTRL, OUT1 );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] OUT1;
  input CTRL;


  MUX2_X1 U1 ( .A(IN0[3]), .B(IN1[3]), .S(CTRL), .Z(OUT1[3]) );
  MUX2_X1 U2 ( .A(IN0[2]), .B(IN1[2]), .S(CTRL), .Z(OUT1[2]) );
  MUX2_X1 U3 ( .A(IN0[1]), .B(IN1[1]), .S(CTRL), .Z(OUT1[1]) );
  MUX2_X1 U4 ( .A(IN0[0]), .B(IN1[0]), .S(CTRL), .Z(OUT1[0]) );
endmodule


module mux21_SIZE4_8 ( IN0, IN1, CTRL, OUT1 );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] OUT1;
  input CTRL;


  MUX2_X1 U1 ( .A(IN0[3]), .B(IN1[3]), .S(CTRL), .Z(OUT1[3]) );
  MUX2_X1 U2 ( .A(IN0[2]), .B(IN1[2]), .S(CTRL), .Z(OUT1[2]) );
  MUX2_X1 U3 ( .A(IN0[1]), .B(IN1[1]), .S(CTRL), .Z(OUT1[1]) );
  MUX2_X1 U4 ( .A(IN0[0]), .B(IN1[0]), .S(CTRL), .Z(OUT1[0]) );
endmodule


module mux21_SIZE4_7 ( IN0, IN1, CTRL, OUT1 );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] OUT1;
  input CTRL;


  MUX2_X1 U1 ( .A(IN0[3]), .B(IN1[3]), .S(CTRL), .Z(OUT1[3]) );
  MUX2_X1 U2 ( .A(IN0[2]), .B(IN1[2]), .S(CTRL), .Z(OUT1[2]) );
  MUX2_X1 U3 ( .A(IN0[1]), .B(IN1[1]), .S(CTRL), .Z(OUT1[1]) );
  MUX2_X1 U4 ( .A(IN0[0]), .B(IN1[0]), .S(CTRL), .Z(OUT1[0]) );
endmodule


module mux21_SIZE4_6 ( IN0, IN1, CTRL, OUT1 );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] OUT1;
  input CTRL;


  MUX2_X1 U1 ( .A(IN0[3]), .B(IN1[3]), .S(CTRL), .Z(OUT1[3]) );
  MUX2_X1 U2 ( .A(IN0[2]), .B(IN1[2]), .S(CTRL), .Z(OUT1[2]) );
  MUX2_X1 U3 ( .A(IN0[1]), .B(IN1[1]), .S(CTRL), .Z(OUT1[1]) );
  MUX2_X1 U4 ( .A(IN0[0]), .B(IN1[0]), .S(CTRL), .Z(OUT1[0]) );
endmodule


module mux21_SIZE4_5 ( IN0, IN1, CTRL, OUT1 );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] OUT1;
  input CTRL;


  MUX2_X1 U1 ( .A(IN0[3]), .B(IN1[3]), .S(CTRL), .Z(OUT1[3]) );
  MUX2_X1 U2 ( .A(IN0[2]), .B(IN1[2]), .S(CTRL), .Z(OUT1[2]) );
  MUX2_X1 U3 ( .A(IN0[1]), .B(IN1[1]), .S(CTRL), .Z(OUT1[1]) );
  MUX2_X1 U4 ( .A(IN0[0]), .B(IN1[0]), .S(CTRL), .Z(OUT1[0]) );
endmodule


module mux21_SIZE4_4 ( IN0, IN1, CTRL, OUT1 );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] OUT1;
  input CTRL;


  MUX2_X1 U1 ( .A(IN0[3]), .B(IN1[3]), .S(CTRL), .Z(OUT1[3]) );
  MUX2_X1 U2 ( .A(IN0[2]), .B(IN1[2]), .S(CTRL), .Z(OUT1[2]) );
  MUX2_X1 U3 ( .A(IN0[1]), .B(IN1[1]), .S(CTRL), .Z(OUT1[1]) );
  MUX2_X1 U4 ( .A(IN0[0]), .B(IN1[0]), .S(CTRL), .Z(OUT1[0]) );
endmodule


module mux21_SIZE4_3 ( IN0, IN1, CTRL, OUT1 );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] OUT1;
  input CTRL;


  MUX2_X1 U1 ( .A(IN0[3]), .B(IN1[3]), .S(CTRL), .Z(OUT1[3]) );
  MUX2_X1 U2 ( .A(IN0[2]), .B(IN1[2]), .S(CTRL), .Z(OUT1[2]) );
  MUX2_X1 U3 ( .A(IN0[1]), .B(IN1[1]), .S(CTRL), .Z(OUT1[1]) );
  MUX2_X1 U4 ( .A(IN0[0]), .B(IN1[0]), .S(CTRL), .Z(OUT1[0]) );
endmodule


module mux21_SIZE4_2 ( IN0, IN1, CTRL, OUT1 );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] OUT1;
  input CTRL;


  MUX2_X1 U1 ( .A(IN0[3]), .B(IN1[3]), .S(CTRL), .Z(OUT1[3]) );
  MUX2_X1 U2 ( .A(IN0[2]), .B(IN1[2]), .S(CTRL), .Z(OUT1[2]) );
  MUX2_X1 U3 ( .A(IN0[1]), .B(IN1[1]), .S(CTRL), .Z(OUT1[1]) );
  MUX2_X1 U4 ( .A(IN0[0]), .B(IN1[0]), .S(CTRL), .Z(OUT1[0]) );
endmodule


module mux21_SIZE4_1 ( IN0, IN1, CTRL, OUT1 );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] OUT1;
  input CTRL;


  MUX2_X1 U1 ( .A(IN0[3]), .B(IN1[3]), .S(CTRL), .Z(OUT1[3]) );
  MUX2_X1 U2 ( .A(IN0[2]), .B(IN1[2]), .S(CTRL), .Z(OUT1[2]) );
  MUX2_X1 U3 ( .A(IN0[1]), .B(IN1[1]), .S(CTRL), .Z(OUT1[1]) );
  MUX2_X1 U4 ( .A(IN0[0]), .B(IN1[0]), .S(CTRL), .Z(OUT1[0]) );
endmodule


module RCA_N4_30 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_120 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(1'b0), .S(S[0]), .Co(CTMP[1]) );
  FA_119 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_118 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_117 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module RCA_N4_29 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_116 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(1'b1), .S(S[0]), .Co(CTMP[1]) );
  FA_115 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_114 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_113 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module RCA_N4_28 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_112 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(1'b0), .S(S[0]), .Co(CTMP[1]) );
  FA_111 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_110 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_109 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module RCA_N4_27 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_108 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(1'b1), .S(S[0]), .Co(CTMP[1]) );
  FA_107 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_106 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_105 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module RCA_N4_26 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_104 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(1'b0), .S(S[0]), .Co(CTMP[1]) );
  FA_103 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_102 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_101 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module RCA_N4_25 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_100 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(1'b1), .S(S[0]), .Co(CTMP[1]) );
  FA_99 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_98 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_97 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module RCA_N4_24 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_96 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(1'b0), .S(S[0]), .Co(CTMP[1]) );
  FA_95 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_94 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_93 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module RCA_N4_23 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_92 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(1'b1), .S(S[0]), .Co(CTMP[1]) );
  FA_91 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_90 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_89 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module RCA_N4_22 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_88 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(1'b0), .S(S[0]), .Co(CTMP[1]) );
  FA_87 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_86 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_85 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module RCA_N4_21 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_84 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(1'b1), .S(S[0]), .Co(CTMP[1]) );
  FA_83 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_82 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_81 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module RCA_N4_20 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_80 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(1'b0), .S(S[0]), .Co(CTMP[1]) );
  FA_79 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_78 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_77 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module RCA_N4_19 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_76 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(1'b1), .S(S[0]), .Co(CTMP[1]) );
  FA_75 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_74 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_73 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module RCA_N4_18 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_72 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(1'b0), .S(S[0]), .Co(CTMP[1]) );
  FA_71 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_70 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_69 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module RCA_N4_17 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_68 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(1'b1), .S(S[0]), .Co(CTMP[1]) );
  FA_67 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_66 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_65 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module RCA_N4_16 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_64 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(1'b0), .S(S[0]), .Co(CTMP[1]) );
  FA_63 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_62 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_61 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module RCA_N4_15 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_60 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(1'b1), .S(S[0]), .Co(CTMP[1]) );
  FA_59 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_58 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_57 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module RCA_N4_14 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_56 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(1'b0), .S(S[0]), .Co(CTMP[1]) );
  FA_55 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_54 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_53 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module RCA_N4_13 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_52 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(1'b1), .S(S[0]), .Co(CTMP[1]) );
  FA_51 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_50 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_49 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module RCA_N4_12 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_48 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(1'b0), .S(S[0]), .Co(CTMP[1]) );
  FA_47 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_46 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_45 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module RCA_N4_11 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_44 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(1'b1), .S(S[0]), .Co(CTMP[1]) );
  FA_43 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_42 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_41 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module RCA_N4_10 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_40 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(1'b0), .S(S[0]), .Co(CTMP[1]) );
  FA_39 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_38 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_37 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module RCA_N4_9 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_36 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(1'b1), .S(S[0]), .Co(CTMP[1]) );
  FA_35 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_34 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_33 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module RCA_N4_8 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_32 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(1'b0), .S(S[0]), .Co(CTMP[1]) );
  FA_31 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_30 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_29 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module RCA_N4_7 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_28 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(1'b1), .S(S[0]), .Co(CTMP[1]) );
  FA_27 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_26 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_25 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module RCA_N4_6 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_24 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(1'b0), .S(S[0]), .Co(CTMP[1]) );
  FA_23 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_22 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_21 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module RCA_N4_5 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_20 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(1'b1), .S(S[0]), .Co(CTMP[1]) );
  FA_19 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_18 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_17 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module RCA_N4_4 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_16 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(1'b0), .S(S[0]), .Co(CTMP[1]) );
  FA_15 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_14 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_13 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module RCA_N4_3 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_12 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(1'b1), .S(S[0]), .Co(CTMP[1]) );
  FA_11 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_10 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_9 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module RCA_N4_2 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_8 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(1'b0), .S(S[0]), .Co(CTMP[1]) );
  FA_7 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_6 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_5 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module RCA_N4_1 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_4 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(1'b1), .S(S[0]), .Co(CTMP[1]) );
  FA_3 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_2 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module shift_N9_2 ( Clock, ALOAD, D, SO );
  input [8:0] D;
  input Clock, ALOAD;
  output SO;
  wire   N11;
  wire   [8:1] tmp;

  DFF_X1 \tmp_reg[8]  ( .D(N11), .CK(Clock), .Q(tmp[8]) );
  SDFF_X1 \tmp_reg[7]  ( .D(tmp[8]), .SI(D[7]), .SE(ALOAD), .CK(Clock), .Q(
        tmp[7]) );
  SDFF_X1 \tmp_reg[6]  ( .D(tmp[7]), .SI(D[6]), .SE(ALOAD), .CK(Clock), .Q(
        tmp[6]) );
  SDFF_X1 \tmp_reg[5]  ( .D(tmp[6]), .SI(D[5]), .SE(ALOAD), .CK(Clock), .Q(
        tmp[5]) );
  SDFF_X1 \tmp_reg[4]  ( .D(tmp[5]), .SI(D[4]), .SE(ALOAD), .CK(Clock), .Q(
        tmp[4]) );
  SDFF_X1 \tmp_reg[3]  ( .D(tmp[4]), .SI(D[3]), .SE(ALOAD), .CK(Clock), .Q(
        tmp[3]) );
  SDFF_X1 \tmp_reg[2]  ( .D(tmp[3]), .SI(D[2]), .SE(ALOAD), .CK(Clock), .Q(
        tmp[2]) );
  SDFF_X1 \tmp_reg[1]  ( .D(tmp[2]), .SI(D[1]), .SE(ALOAD), .CK(Clock), .Q(
        tmp[1]) );
  SDFF_X1 \tmp_reg[0]  ( .D(tmp[1]), .SI(D[0]), .SE(ALOAD), .CK(Clock), .Q(SO)
         );
  AND2_X1 U3 ( .A1(ALOAD), .A2(D[8]), .ZN(N11) );
endmodule


module shift_N9_1 ( Clock, ALOAD, D, SO );
  input [8:0] D;
  input Clock, ALOAD;
  output SO;
  wire   N11;
  wire   [8:1] tmp;

  DFF_X1 \tmp_reg[8]  ( .D(N11), .CK(Clock), .Q(tmp[8]) );
  SDFF_X1 \tmp_reg[7]  ( .D(tmp[8]), .SI(D[7]), .SE(ALOAD), .CK(Clock), .Q(
        tmp[7]) );
  SDFF_X1 \tmp_reg[6]  ( .D(tmp[7]), .SI(D[6]), .SE(ALOAD), .CK(Clock), .Q(
        tmp[6]) );
  SDFF_X1 \tmp_reg[5]  ( .D(tmp[6]), .SI(D[5]), .SE(ALOAD), .CK(Clock), .Q(
        tmp[5]) );
  SDFF_X1 \tmp_reg[4]  ( .D(tmp[5]), .SI(D[4]), .SE(ALOAD), .CK(Clock), .Q(
        tmp[4]) );
  SDFF_X1 \tmp_reg[3]  ( .D(tmp[4]), .SI(D[3]), .SE(ALOAD), .CK(Clock), .Q(
        tmp[3]) );
  SDFF_X1 \tmp_reg[2]  ( .D(tmp[3]), .SI(D[2]), .SE(ALOAD), .CK(Clock), .Q(
        tmp[2]) );
  SDFF_X1 \tmp_reg[1]  ( .D(tmp[2]), .SI(D[1]), .SE(ALOAD), .CK(Clock), .Q(
        tmp[1]) );
  SDFF_X1 \tmp_reg[0]  ( .D(tmp[1]), .SI(D[0]), .SE(ALOAD), .CK(Clock), .Q(SO)
         );
  AND2_X1 U3 ( .A1(ALOAD), .A2(D[8]), .ZN(N11) );
endmodule


module booth_encoder_8 ( B_in, A_out );
  input [2:0] B_in;
  output [2:0] A_out;
  wire   N53, N55, N57, n1, n5, n6, n7;
  assign A_out[0] = N53;
  assign A_out[1] = N55;
  assign A_out[2] = N57;

  OAI33_X1 U6 ( .A1(B_in[0]), .A2(B_in[1]), .A3(n1), .B1(n7), .B2(n6), .B3(
        B_in[2]), .ZN(N53) );
  NAND2_X1 U4 ( .A1(B_in[2]), .A2(n7), .ZN(n5) );
  OAI221_X1 U3 ( .B1(B_in[1]), .B2(n7), .C1(n6), .C2(B_in[2]), .A(n5), .ZN(N57) );
  AOI21_X1 U5 ( .B1(B_in[0]), .B2(B_in[1]), .A(n1), .ZN(N55) );
  INV_X1 U8 ( .A(B_in[0]), .ZN(n7) );
  INV_X1 U7 ( .A(B_in[1]), .ZN(n6) );
  INV_X1 U9 ( .A(B_in[2]), .ZN(n1) );
endmodule


module booth_encoder_7 ( B_in, A_out );
  input [2:0] B_in;
  output [2:0] A_out;
  wire   N53, N55, N57, n1, n5, n6, n7;
  assign A_out[0] = N53;
  assign A_out[1] = N55;
  assign A_out[2] = N57;

  OAI33_X1 U6 ( .A1(B_in[0]), .A2(B_in[1]), .A3(n1), .B1(n7), .B2(n6), .B3(
        B_in[2]), .ZN(N53) );
  NAND2_X1 U4 ( .A1(B_in[2]), .A2(n7), .ZN(n5) );
  OAI221_X1 U3 ( .B1(B_in[1]), .B2(n7), .C1(n6), .C2(B_in[2]), .A(n5), .ZN(N57) );
  AOI21_X1 U5 ( .B1(B_in[0]), .B2(B_in[1]), .A(n1), .ZN(N55) );
  INV_X1 U8 ( .A(B_in[0]), .ZN(n7) );
  INV_X1 U7 ( .A(B_in[1]), .ZN(n6) );
  INV_X1 U9 ( .A(B_in[2]), .ZN(n1) );
endmodule


module booth_encoder_6 ( B_in, A_out );
  input [2:0] B_in;
  output [2:0] A_out;
  wire   N53, N55, N57, n1, n5, n6, n7;
  assign A_out[0] = N53;
  assign A_out[1] = N55;
  assign A_out[2] = N57;

  OAI33_X1 U6 ( .A1(B_in[0]), .A2(B_in[1]), .A3(n1), .B1(n7), .B2(n6), .B3(
        B_in[2]), .ZN(N53) );
  NAND2_X1 U4 ( .A1(B_in[2]), .A2(n7), .ZN(n5) );
  OAI221_X1 U3 ( .B1(B_in[1]), .B2(n7), .C1(n6), .C2(B_in[2]), .A(n5), .ZN(N57) );
  AOI21_X1 U5 ( .B1(B_in[0]), .B2(B_in[1]), .A(n1), .ZN(N55) );
  INV_X1 U8 ( .A(B_in[0]), .ZN(n7) );
  INV_X1 U7 ( .A(B_in[1]), .ZN(n6) );
  INV_X1 U9 ( .A(B_in[2]), .ZN(n1) );
endmodule


module booth_encoder_5 ( B_in, A_out );
  input [2:0] B_in;
  output [2:0] A_out;
  wire   N53, N55, N57, n1, n5, n6, n7;
  assign A_out[0] = N53;
  assign A_out[1] = N55;
  assign A_out[2] = N57;

  OAI33_X1 U6 ( .A1(B_in[0]), .A2(B_in[1]), .A3(n1), .B1(n7), .B2(n6), .B3(
        B_in[2]), .ZN(N53) );
  NAND2_X1 U4 ( .A1(B_in[2]), .A2(n7), .ZN(n5) );
  OAI221_X1 U3 ( .B1(B_in[1]), .B2(n7), .C1(n6), .C2(B_in[2]), .A(n5), .ZN(N57) );
  AOI21_X1 U5 ( .B1(B_in[0]), .B2(B_in[1]), .A(n1), .ZN(N55) );
  INV_X1 U8 ( .A(B_in[0]), .ZN(n7) );
  INV_X1 U7 ( .A(B_in[1]), .ZN(n6) );
  INV_X1 U9 ( .A(B_in[2]), .ZN(n1) );
endmodule


module booth_encoder_4 ( B_in, A_out );
  input [2:0] B_in;
  output [2:0] A_out;
  wire   N53, N55, N57, n1, n5, n6, n7;
  assign A_out[0] = N53;
  assign A_out[1] = N55;
  assign A_out[2] = N57;

  OAI33_X1 U6 ( .A1(B_in[0]), .A2(B_in[1]), .A3(n1), .B1(n7), .B2(n6), .B3(
        B_in[2]), .ZN(N53) );
  NAND2_X1 U4 ( .A1(B_in[2]), .A2(n7), .ZN(n5) );
  OAI221_X1 U3 ( .B1(B_in[1]), .B2(n7), .C1(n6), .C2(B_in[2]), .A(n5), .ZN(N57) );
  AOI21_X1 U5 ( .B1(B_in[0]), .B2(B_in[1]), .A(n1), .ZN(N55) );
  INV_X1 U8 ( .A(B_in[0]), .ZN(n7) );
  INV_X1 U7 ( .A(B_in[1]), .ZN(n6) );
  INV_X1 U9 ( .A(B_in[2]), .ZN(n1) );
endmodule


module booth_encoder_3 ( B_in, A_out );
  input [2:0] B_in;
  output [2:0] A_out;
  wire   N53, N55, N57, n1, n5, n6, n7;
  assign A_out[0] = N53;
  assign A_out[1] = N55;
  assign A_out[2] = N57;

  OAI33_X1 U6 ( .A1(B_in[0]), .A2(B_in[1]), .A3(n1), .B1(n7), .B2(n6), .B3(
        B_in[2]), .ZN(N53) );
  NAND2_X1 U4 ( .A1(B_in[2]), .A2(n7), .ZN(n5) );
  OAI221_X1 U3 ( .B1(B_in[1]), .B2(n7), .C1(n6), .C2(B_in[2]), .A(n5), .ZN(N57) );
  AOI21_X1 U5 ( .B1(B_in[0]), .B2(B_in[1]), .A(n1), .ZN(N55) );
  INV_X1 U8 ( .A(B_in[0]), .ZN(n7) );
  INV_X1 U7 ( .A(B_in[1]), .ZN(n6) );
  INV_X1 U9 ( .A(B_in[2]), .ZN(n1) );
endmodule


module booth_encoder_2 ( B_in, A_out );
  input [2:0] B_in;
  output [2:0] A_out;
  wire   N53, N55, N57, n1, n5, n6, n7;
  assign A_out[0] = N53;
  assign A_out[1] = N55;
  assign A_out[2] = N57;

  OAI33_X1 U6 ( .A1(B_in[0]), .A2(B_in[1]), .A3(n1), .B1(n7), .B2(n6), .B3(
        B_in[2]), .ZN(N53) );
  NAND2_X1 U4 ( .A1(B_in[2]), .A2(n7), .ZN(n5) );
  OAI221_X1 U3 ( .B1(B_in[1]), .B2(n7), .C1(n6), .C2(B_in[2]), .A(n5), .ZN(N57) );
  AOI21_X1 U5 ( .B1(B_in[0]), .B2(B_in[1]), .A(n1), .ZN(N55) );
  INV_X1 U8 ( .A(B_in[0]), .ZN(n7) );
  INV_X1 U7 ( .A(B_in[1]), .ZN(n6) );
  INV_X1 U9 ( .A(B_in[2]), .ZN(n1) );
endmodule


module booth_encoder_1 ( B_in, A_out );
  input [2:0] B_in;
  output [2:0] A_out;
  wire   N53, N55, N57, n1, n4, n5;
  assign A_out[0] = N53;
  assign A_out[1] = N55;
  assign A_out[2] = N57;

  OAI33_X1 U6 ( .A1(B_in[0]), .A2(B_in[1]), .A3(n4), .B1(n5), .B2(n4), .B3(
        B_in[2]), .ZN(N53) );
  AOI21_X1 U5 ( .B1(B_in[0]), .B2(B_in[1]), .A(n4), .ZN(N55) );
  NAND2_X1 U4 ( .A1(B_in[2]), .A2(n5), .ZN(n1) );
  OAI221_X1 U3 ( .B1(B_in[1]), .B2(n5), .C1(n4), .C2(B_in[2]), .A(n1), .ZN(N57) );
  INV_X1 U8 ( .A(B_in[0]), .ZN(n5) );
  INV_X1 U7 ( .A(B_in[1]), .ZN(n4) );
endmodule


module carry_sel_gen_N4_15 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:0] nocarry_sum_to_mux;
  wire   [3:0] carry_sum_to_mux;

  RCA_N4_30 rca_nocarry ( .A(A), .B(B), .Ci(1'b0), .S(nocarry_sum_to_mux) );
  RCA_N4_29 rca_carry ( .A(A), .B(B), .Ci(1'b1), .S(carry_sum_to_mux) );
  mux21_SIZE4_15 outmux ( .IN0(nocarry_sum_to_mux), .IN1(carry_sum_to_mux), 
        .CTRL(Ci), .OUT1(S) );
endmodule


module carry_sel_gen_N4_14 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:0] nocarry_sum_to_mux;
  wire   [3:0] carry_sum_to_mux;

  RCA_N4_28 rca_nocarry ( .A(A), .B(B), .Ci(1'b0), .S(nocarry_sum_to_mux) );
  RCA_N4_27 rca_carry ( .A(A), .B(B), .Ci(1'b1), .S(carry_sum_to_mux) );
  mux21_SIZE4_14 outmux ( .IN0(nocarry_sum_to_mux), .IN1(carry_sum_to_mux), 
        .CTRL(Ci), .OUT1(S) );
endmodule


module carry_sel_gen_N4_13 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:0] nocarry_sum_to_mux;
  wire   [3:0] carry_sum_to_mux;

  RCA_N4_26 rca_nocarry ( .A(A), .B(B), .Ci(1'b0), .S(nocarry_sum_to_mux) );
  RCA_N4_25 rca_carry ( .A(A), .B(B), .Ci(1'b1), .S(carry_sum_to_mux) );
  mux21_SIZE4_13 outmux ( .IN0(nocarry_sum_to_mux), .IN1(carry_sum_to_mux), 
        .CTRL(Ci), .OUT1(S) );
endmodule


module carry_sel_gen_N4_12 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:0] nocarry_sum_to_mux;
  wire   [3:0] carry_sum_to_mux;

  RCA_N4_24 rca_nocarry ( .A(A), .B(B), .Ci(1'b0), .S(nocarry_sum_to_mux) );
  RCA_N4_23 rca_carry ( .A(A), .B(B), .Ci(1'b1), .S(carry_sum_to_mux) );
  mux21_SIZE4_12 outmux ( .IN0(nocarry_sum_to_mux), .IN1(carry_sum_to_mux), 
        .CTRL(Ci), .OUT1(S) );
endmodule


module carry_sel_gen_N4_11 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:0] nocarry_sum_to_mux;
  wire   [3:0] carry_sum_to_mux;

  RCA_N4_22 rca_nocarry ( .A(A), .B(B), .Ci(1'b0), .S(nocarry_sum_to_mux) );
  RCA_N4_21 rca_carry ( .A(A), .B(B), .Ci(1'b1), .S(carry_sum_to_mux) );
  mux21_SIZE4_11 outmux ( .IN0(nocarry_sum_to_mux), .IN1(carry_sum_to_mux), 
        .CTRL(Ci), .OUT1(S) );
endmodule


module carry_sel_gen_N4_10 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:0] nocarry_sum_to_mux;
  wire   [3:0] carry_sum_to_mux;

  RCA_N4_20 rca_nocarry ( .A(A), .B(B), .Ci(1'b0), .S(nocarry_sum_to_mux) );
  RCA_N4_19 rca_carry ( .A(A), .B(B), .Ci(1'b1), .S(carry_sum_to_mux) );
  mux21_SIZE4_10 outmux ( .IN0(nocarry_sum_to_mux), .IN1(carry_sum_to_mux), 
        .CTRL(Ci), .OUT1(S) );
endmodule


module carry_sel_gen_N4_9 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:0] nocarry_sum_to_mux;
  wire   [3:0] carry_sum_to_mux;

  RCA_N4_18 rca_nocarry ( .A(A), .B(B), .Ci(1'b0), .S(nocarry_sum_to_mux) );
  RCA_N4_17 rca_carry ( .A(A), .B(B), .Ci(1'b1), .S(carry_sum_to_mux) );
  mux21_SIZE4_9 outmux ( .IN0(nocarry_sum_to_mux), .IN1(carry_sum_to_mux), 
        .CTRL(Ci), .OUT1(S) );
endmodule


module carry_sel_gen_N4_8 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:0] nocarry_sum_to_mux;
  wire   [3:0] carry_sum_to_mux;

  RCA_N4_16 rca_nocarry ( .A(A), .B(B), .Ci(1'b0), .S(nocarry_sum_to_mux) );
  RCA_N4_15 rca_carry ( .A(A), .B(B), .Ci(1'b1), .S(carry_sum_to_mux) );
  mux21_SIZE4_8 outmux ( .IN0(nocarry_sum_to_mux), .IN1(carry_sum_to_mux), 
        .CTRL(Ci), .OUT1(S) );
endmodule


module carry_sel_gen_N4_7 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:0] nocarry_sum_to_mux;
  wire   [3:0] carry_sum_to_mux;

  RCA_N4_14 rca_nocarry ( .A(A), .B(B), .Ci(1'b0), .S(nocarry_sum_to_mux) );
  RCA_N4_13 rca_carry ( .A(A), .B(B), .Ci(1'b1), .S(carry_sum_to_mux) );
  mux21_SIZE4_7 outmux ( .IN0(nocarry_sum_to_mux), .IN1(carry_sum_to_mux), 
        .CTRL(Ci), .OUT1(S) );
endmodule


module carry_sel_gen_N4_6 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:0] nocarry_sum_to_mux;
  wire   [3:0] carry_sum_to_mux;

  RCA_N4_12 rca_nocarry ( .A(A), .B(B), .Ci(1'b0), .S(nocarry_sum_to_mux) );
  RCA_N4_11 rca_carry ( .A(A), .B(B), .Ci(1'b1), .S(carry_sum_to_mux) );
  mux21_SIZE4_6 outmux ( .IN0(nocarry_sum_to_mux), .IN1(carry_sum_to_mux), 
        .CTRL(Ci), .OUT1(S) );
endmodule


module carry_sel_gen_N4_5 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:0] nocarry_sum_to_mux;
  wire   [3:0] carry_sum_to_mux;

  RCA_N4_10 rca_nocarry ( .A(A), .B(B), .Ci(1'b0), .S(nocarry_sum_to_mux) );
  RCA_N4_9 rca_carry ( .A(A), .B(B), .Ci(1'b1), .S(carry_sum_to_mux) );
  mux21_SIZE4_5 outmux ( .IN0(nocarry_sum_to_mux), .IN1(carry_sum_to_mux), 
        .CTRL(Ci), .OUT1(S) );
endmodule


module carry_sel_gen_N4_4 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:0] nocarry_sum_to_mux;
  wire   [3:0] carry_sum_to_mux;

  RCA_N4_8 rca_nocarry ( .A(A), .B(B), .Ci(1'b0), .S(nocarry_sum_to_mux) );
  RCA_N4_7 rca_carry ( .A(A), .B(B), .Ci(1'b1), .S(carry_sum_to_mux) );
  mux21_SIZE4_4 outmux ( .IN0(nocarry_sum_to_mux), .IN1(carry_sum_to_mux), 
        .CTRL(Ci), .OUT1(S) );
endmodule


module carry_sel_gen_N4_3 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:0] nocarry_sum_to_mux;
  wire   [3:0] carry_sum_to_mux;

  RCA_N4_6 rca_nocarry ( .A(A), .B(B), .Ci(1'b0), .S(nocarry_sum_to_mux) );
  RCA_N4_5 rca_carry ( .A(A), .B(B), .Ci(1'b1), .S(carry_sum_to_mux) );
  mux21_SIZE4_3 outmux ( .IN0(nocarry_sum_to_mux), .IN1(carry_sum_to_mux), 
        .CTRL(Ci), .OUT1(S) );
endmodule


module carry_sel_gen_N4_2 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:0] nocarry_sum_to_mux;
  wire   [3:0] carry_sum_to_mux;

  RCA_N4_4 rca_nocarry ( .A(A), .B(B), .Ci(1'b0), .S(nocarry_sum_to_mux) );
  RCA_N4_3 rca_carry ( .A(A), .B(B), .Ci(1'b1), .S(carry_sum_to_mux) );
  mux21_SIZE4_2 outmux ( .IN0(nocarry_sum_to_mux), .IN1(carry_sum_to_mux), 
        .CTRL(Ci), .OUT1(S) );
endmodule


module carry_sel_gen_N4_1 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:0] nocarry_sum_to_mux;
  wire   [3:0] carry_sum_to_mux;

  RCA_N4_2 rca_nocarry ( .A(A), .B(B), .Ci(1'b0), .S(nocarry_sum_to_mux) );
  RCA_N4_1 rca_carry ( .A(A), .B(B), .Ci(1'b1), .S(carry_sum_to_mux) );
  mux21_SIZE4_1 outmux ( .IN0(nocarry_sum_to_mux), .IN1(carry_sum_to_mux), 
        .CTRL(Ci), .OUT1(S) );
endmodule


module pg_53 ( g, p, g_prec, p_prec, g_out, p_out );
  input g, p, g_prec, p_prec;
  output g_out, p_out;
  wire   n1;

  AOI21_X1 U3 ( .B1(g_prec), .B2(p), .A(g), .ZN(n1) );
  AND2_X1 U1 ( .A1(p), .A2(p_prec), .ZN(p_out) );
  INV_X1 U2 ( .A(n1), .ZN(g_out) );
endmodule


module pg_52 ( g, p, g_prec, p_prec, g_out, p_out );
  input g, p, g_prec, p_prec;
  output g_out, p_out;
  wire   n1;

  AOI21_X1 U3 ( .B1(g_prec), .B2(p), .A(g), .ZN(n1) );
  AND2_X1 U1 ( .A1(p), .A2(p_prec), .ZN(p_out) );
  INV_X1 U2 ( .A(n1), .ZN(g_out) );
endmodule


module pg_51 ( g, p, g_prec, p_prec, g_out, p_out );
  input g, p, g_prec, p_prec;
  output g_out, p_out;
  wire   n1;

  AOI21_X1 U3 ( .B1(g_prec), .B2(p), .A(g), .ZN(n1) );
  AND2_X1 U1 ( .A1(p), .A2(p_prec), .ZN(p_out) );
  INV_X1 U2 ( .A(n1), .ZN(g_out) );
endmodule


module pg_50 ( g, p, g_prec, p_prec, g_out, p_out );
  input g, p, g_prec, p_prec;
  output g_out, p_out;
  wire   n1;

  AOI21_X1 U3 ( .B1(g_prec), .B2(p), .A(g), .ZN(n1) );
  AND2_X1 U1 ( .A1(p), .A2(p_prec), .ZN(p_out) );
  INV_X1 U2 ( .A(n1), .ZN(g_out) );
endmodule


module pg_49 ( g, p, g_prec, p_prec, g_out, p_out );
  input g, p, g_prec, p_prec;
  output g_out, p_out;
  wire   n1;

  AOI21_X1 U3 ( .B1(g_prec), .B2(p), .A(g), .ZN(n1) );
  AND2_X1 U1 ( .A1(p), .A2(p_prec), .ZN(p_out) );
  INV_X1 U2 ( .A(n1), .ZN(g_out) );
endmodule


module pg_48 ( g, p, g_prec, p_prec, g_out, p_out );
  input g, p, g_prec, p_prec;
  output g_out, p_out;
  wire   n1;

  AOI21_X1 U3 ( .B1(g_prec), .B2(p), .A(g), .ZN(n1) );
  AND2_X1 U1 ( .A1(p), .A2(p_prec), .ZN(p_out) );
  INV_X1 U2 ( .A(n1), .ZN(g_out) );
endmodule


module pg_47 ( g, p, g_prec, p_prec, g_out, p_out );
  input g, p, g_prec, p_prec;
  output g_out, p_out;
  wire   n1;

  AOI21_X1 U3 ( .B1(g_prec), .B2(p), .A(g), .ZN(n1) );
  AND2_X1 U1 ( .A1(p), .A2(p_prec), .ZN(p_out) );
  INV_X1 U2 ( .A(n1), .ZN(g_out) );
endmodule


module pg_46 ( g, p, g_prec, p_prec, g_out, p_out );
  input g, p, g_prec, p_prec;
  output g_out, p_out;
  wire   n1;

  AOI21_X1 U3 ( .B1(g_prec), .B2(p), .A(g), .ZN(n1) );
  AND2_X1 U1 ( .A1(p), .A2(p_prec), .ZN(p_out) );
  INV_X1 U2 ( .A(n1), .ZN(g_out) );
endmodule


module pg_45 ( g, p, g_prec, p_prec, g_out, p_out );
  input g, p, g_prec, p_prec;
  output g_out, p_out;
  wire   n1;

  AOI21_X1 U3 ( .B1(g_prec), .B2(p), .A(g), .ZN(n1) );
  AND2_X1 U1 ( .A1(p), .A2(p_prec), .ZN(p_out) );
  INV_X1 U2 ( .A(n1), .ZN(g_out) );
endmodule


module pg_44 ( g, p, g_prec, p_prec, g_out, p_out );
  input g, p, g_prec, p_prec;
  output g_out, p_out;
  wire   n1;

  AOI21_X1 U3 ( .B1(g_prec), .B2(p), .A(g), .ZN(n1) );
  AND2_X1 U1 ( .A1(p), .A2(p_prec), .ZN(p_out) );
  INV_X1 U2 ( .A(n1), .ZN(g_out) );
endmodule


module pg_43 ( g, p, g_prec, p_prec, g_out, p_out );
  input g, p, g_prec, p_prec;
  output g_out, p_out;
  wire   n1;

  AOI21_X1 U3 ( .B1(g_prec), .B2(p), .A(g), .ZN(n1) );
  AND2_X1 U1 ( .A1(p), .A2(p_prec), .ZN(p_out) );
  INV_X1 U2 ( .A(n1), .ZN(g_out) );
endmodule


module pg_42 ( g, p, g_prec, p_prec, g_out, p_out );
  input g, p, g_prec, p_prec;
  output g_out, p_out;
  wire   n1;

  AOI21_X1 U3 ( .B1(g_prec), .B2(p), .A(g), .ZN(n1) );
  AND2_X1 U1 ( .A1(p), .A2(p_prec), .ZN(p_out) );
  INV_X1 U2 ( .A(n1), .ZN(g_out) );
endmodule


module pg_39 ( g, p, g_prec, p_prec, g_out, p_out );
  input g, p, g_prec, p_prec;
  output g_out, p_out;
  wire   n1;

  AOI21_X1 U3 ( .B1(g_prec), .B2(p), .A(g), .ZN(n1) );
  AND2_X1 U1 ( .A1(p), .A2(p_prec), .ZN(p_out) );
  INV_X1 U2 ( .A(n1), .ZN(g_out) );
endmodule


module pg_38 ( g, p, g_prec, p_prec, g_out, p_out );
  input g, p, g_prec, p_prec;
  output g_out, p_out;
  wire   n1;

  AOI21_X1 U3 ( .B1(g_prec), .B2(p), .A(g), .ZN(n1) );
  AND2_X1 U1 ( .A1(p), .A2(p_prec), .ZN(p_out) );
  INV_X1 U2 ( .A(n1), .ZN(g_out) );
endmodule


module pg_37 ( g, p, g_prec, p_prec, g_out, p_out );
  input g, p, g_prec, p_prec;
  output g_out, p_out;
  wire   n1;

  AOI21_X1 U3 ( .B1(g_prec), .B2(p), .A(g), .ZN(n1) );
  AND2_X1 U1 ( .A1(p), .A2(p_prec), .ZN(p_out) );
  INV_X1 U2 ( .A(n1), .ZN(g_out) );
endmodule


module pg_36 ( g, p, g_prec, p_prec, g_out, p_out );
  input g, p, g_prec, p_prec;
  output g_out, p_out;
  wire   n1;

  AOI21_X1 U3 ( .B1(g_prec), .B2(p), .A(g), .ZN(n1) );
  AND2_X1 U1 ( .A1(p), .A2(p_prec), .ZN(p_out) );
  INV_X1 U2 ( .A(n1), .ZN(g_out) );
endmodule


module pg_35 ( g, p, g_prec, p_prec, g_out, p_out );
  input g, p, g_prec, p_prec;
  output g_out, p_out;
  wire   n1;

  AOI21_X1 U3 ( .B1(g_prec), .B2(p), .A(g), .ZN(n1) );
  AND2_X1 U1 ( .A1(p), .A2(p_prec), .ZN(p_out) );
  INV_X1 U2 ( .A(n1), .ZN(g_out) );
endmodule


module pg_34 ( g, p, g_prec, p_prec, g_out, p_out );
  input g, p, g_prec, p_prec;
  output g_out, p_out;
  wire   n1;

  AOI21_X1 U3 ( .B1(g_prec), .B2(p), .A(g), .ZN(n1) );
  AND2_X1 U1 ( .A1(p), .A2(p_prec), .ZN(p_out) );
  INV_X1 U2 ( .A(n1), .ZN(g_out) );
endmodule


module pg_32 ( g, p, g_prec, p_prec, g_out, p_out );
  input g, p, g_prec, p_prec;
  output g_out, p_out;
  wire   n1;

  AOI21_X1 U3 ( .B1(g_prec), .B2(p), .A(g), .ZN(n1) );
  AND2_X1 U1 ( .A1(p), .A2(p_prec), .ZN(p_out) );
  INV_X1 U2 ( .A(n1), .ZN(g_out) );
endmodule


module pg_31 ( g, p, g_prec, p_prec, g_out, p_out );
  input g, p, g_prec, p_prec;
  output g_out, p_out;
  wire   n1;

  AOI21_X1 U3 ( .B1(g_prec), .B2(p), .A(g), .ZN(n1) );
  AND2_X1 U1 ( .A1(p), .A2(p_prec), .ZN(p_out) );
  INV_X1 U2 ( .A(n1), .ZN(g_out) );
endmodule


module pg_29 ( g, p, g_prec, p_prec, g_out, p_out );
  input g, p, g_prec, p_prec;
  output g_out, p_out;
  wire   n1;

  AOI21_X1 U3 ( .B1(g_prec), .B2(p), .A(g), .ZN(n1) );
  AND2_X1 U1 ( .A1(p), .A2(p_prec), .ZN(p_out) );
  INV_X1 U2 ( .A(n1), .ZN(g_out) );
endmodule


module pg_27 ( g, p, g_prec, p_prec, g_out, p_out );
  input g, p, g_prec, p_prec;
  output g_out, p_out;
  wire   n1;

  AOI21_X1 U3 ( .B1(g_prec), .B2(p), .A(g), .ZN(n1) );
  AND2_X1 U1 ( .A1(p), .A2(p_prec), .ZN(p_out) );
  INV_X1 U2 ( .A(n1), .ZN(g_out) );
endmodule


module pg_26 ( g, p, g_prec, p_prec, g_out, p_out );
  input g, p, g_prec, p_prec;
  output g_out, p_out;
  wire   n1;

  AOI21_X1 U3 ( .B1(g_prec), .B2(p), .A(g), .ZN(n1) );
  AND2_X1 U1 ( .A1(p), .A2(p_prec), .ZN(p_out) );
  INV_X1 U2 ( .A(n1), .ZN(g_out) );
endmodule


module pg_25 ( g, p, g_prec, p_prec, g_out, p_out );
  input g, p, g_prec, p_prec;
  output g_out, p_out;
  wire   n1;

  AOI21_X1 U3 ( .B1(g_prec), .B2(p), .A(g), .ZN(n1) );
  AND2_X1 U1 ( .A1(p), .A2(p_prec), .ZN(p_out) );
  INV_X1 U2 ( .A(n1), .ZN(g_out) );
endmodule


module pg_24 ( g, p, g_prec, p_prec, g_out, p_out );
  input g, p, g_prec, p_prec;
  output g_out, p_out;
  wire   n1;

  AOI21_X1 U3 ( .B1(g_prec), .B2(p), .A(g), .ZN(n1) );
  AND2_X1 U1 ( .A1(p), .A2(p_prec), .ZN(p_out) );
  INV_X1 U2 ( .A(n1), .ZN(g_out) );
endmodule


module pg_23 ( g, p, g_prec, p_prec, g_out, p_out );
  input g, p, g_prec, p_prec;
  output g_out, p_out;
  wire   n1;

  AOI21_X1 U3 ( .B1(g_prec), .B2(p), .A(g), .ZN(n1) );
  AND2_X1 U1 ( .A1(p), .A2(p_prec), .ZN(p_out) );
  INV_X1 U2 ( .A(n1), .ZN(g_out) );
endmodule


module pg_22 ( g, p, g_prec, p_prec, g_out, p_out );
  input g, p, g_prec, p_prec;
  output g_out, p_out;
  wire   n1;

  AOI21_X1 U3 ( .B1(g_prec), .B2(p), .A(g), .ZN(n1) );
  AND2_X1 U1 ( .A1(p), .A2(p_prec), .ZN(p_out) );
  INV_X1 U2 ( .A(n1), .ZN(g_out) );
endmodule


module pg_21 ( g, p, g_prec, p_prec, g_out, p_out );
  input g, p, g_prec, p_prec;
  output g_out, p_out;
  wire   n1;

  AOI21_X1 U3 ( .B1(g_prec), .B2(p), .A(g), .ZN(n1) );
  AND2_X1 U1 ( .A1(p), .A2(p_prec), .ZN(p_out) );
  INV_X1 U2 ( .A(n1), .ZN(g_out) );
endmodule


module pg_20 ( g, p, g_prec, p_prec, g_out, p_out );
  input g, p, g_prec, p_prec;
  output g_out, p_out;
  wire   n1;

  AOI21_X1 U3 ( .B1(g_prec), .B2(p), .A(g), .ZN(n1) );
  AND2_X1 U1 ( .A1(p), .A2(p_prec), .ZN(p_out) );
  INV_X1 U2 ( .A(n1), .ZN(g_out) );
endmodule


module pg_19 ( g, p, g_prec, p_prec, g_out, p_out );
  input g, p, g_prec, p_prec;
  output g_out, p_out;
  wire   n1;

  AOI21_X1 U3 ( .B1(g_prec), .B2(p), .A(g), .ZN(n1) );
  AND2_X1 U1 ( .A1(p), .A2(p_prec), .ZN(p_out) );
  INV_X1 U2 ( .A(n1), .ZN(g_out) );
endmodule


module pg_18 ( g, p, g_prec, p_prec, g_out, p_out );
  input g, p, g_prec, p_prec;
  output g_out, p_out;
  wire   n1;

  AOI21_X1 U3 ( .B1(g_prec), .B2(p), .A(g), .ZN(n1) );
  AND2_X1 U1 ( .A1(p), .A2(p_prec), .ZN(p_out) );
  INV_X1 U2 ( .A(n1), .ZN(g_out) );
endmodule


module pg_17 ( g, p, g_prec, p_prec, g_out, p_out );
  input g, p, g_prec, p_prec;
  output g_out, p_out;
  wire   n1;

  AOI21_X1 U3 ( .B1(g_prec), .B2(p), .A(g), .ZN(n1) );
  AND2_X1 U1 ( .A1(p), .A2(p_prec), .ZN(p_out) );
  INV_X1 U2 ( .A(n1), .ZN(g_out) );
endmodule


module pg_16 ( g, p, g_prec, p_prec, g_out, p_out );
  input g, p, g_prec, p_prec;
  output g_out, p_out;
  wire   n1;

  AOI21_X1 U3 ( .B1(g_prec), .B2(p), .A(g), .ZN(n1) );
  AND2_X1 U1 ( .A1(p), .A2(p_prec), .ZN(p_out) );
  INV_X1 U2 ( .A(n1), .ZN(g_out) );
endmodule


module pg_15 ( g, p, g_prec, p_prec, g_out, p_out );
  input g, p, g_prec, p_prec;
  output g_out, p_out;
  wire   n1;

  AOI21_X1 U3 ( .B1(g_prec), .B2(p), .A(g), .ZN(n1) );
  AND2_X1 U1 ( .A1(p), .A2(p_prec), .ZN(p_out) );
  INV_X1 U2 ( .A(n1), .ZN(g_out) );
endmodule


module pg_14 ( g, p, g_prec, p_prec, g_out, p_out );
  input g, p, g_prec, p_prec;
  output g_out, p_out;
  wire   n1;

  AOI21_X1 U3 ( .B1(g_prec), .B2(p), .A(g), .ZN(n1) );
  AND2_X1 U1 ( .A1(p), .A2(p_prec), .ZN(p_out) );
  INV_X1 U2 ( .A(n1), .ZN(g_out) );
endmodule


module pg_13 ( g, p, g_prec, p_prec, g_out, p_out );
  input g, p, g_prec, p_prec;
  output g_out, p_out;
  wire   n1;

  AOI21_X1 U3 ( .B1(g_prec), .B2(p), .A(g), .ZN(n1) );
  AND2_X1 U1 ( .A1(p), .A2(p_prec), .ZN(p_out) );
  INV_X1 U2 ( .A(n1), .ZN(g_out) );
endmodule


module pg_12 ( g, p, g_prec, p_prec, g_out, p_out );
  input g, p, g_prec, p_prec;
  output g_out, p_out;
  wire   n1;

  AOI21_X1 U3 ( .B1(g_prec), .B2(p), .A(g), .ZN(n1) );
  AND2_X1 U1 ( .A1(p), .A2(p_prec), .ZN(p_out) );
  INV_X1 U2 ( .A(n1), .ZN(g_out) );
endmodule


module pg_11 ( g, p, g_prec, p_prec, g_out, p_out );
  input g, p, g_prec, p_prec;
  output g_out, p_out;
  wire   n1;

  AOI21_X1 U3 ( .B1(g_prec), .B2(p), .A(g), .ZN(n1) );
  AND2_X1 U1 ( .A1(p), .A2(p_prec), .ZN(p_out) );
  INV_X1 U2 ( .A(n1), .ZN(g_out) );
endmodule


module pg_10 ( g, p, g_prec, p_prec, g_out, p_out );
  input g, p, g_prec, p_prec;
  output g_out, p_out;
  wire   n1;

  AOI21_X1 U3 ( .B1(g_prec), .B2(p), .A(g), .ZN(n1) );
  AND2_X1 U1 ( .A1(p), .A2(p_prec), .ZN(p_out) );
  INV_X1 U2 ( .A(n1), .ZN(g_out) );
endmodule


module pg_9 ( g, p, g_prec, p_prec, g_out, p_out );
  input g, p, g_prec, p_prec;
  output g_out, p_out;
  wire   n1;

  AOI21_X1 U3 ( .B1(g_prec), .B2(p), .A(g), .ZN(n1) );
  AND2_X1 U1 ( .A1(p), .A2(p_prec), .ZN(p_out) );
  INV_X1 U2 ( .A(n1), .ZN(g_out) );
endmodule


module pg_8 ( g, p, g_prec, p_prec, g_out, p_out );
  input g, p, g_prec, p_prec;
  output g_out, p_out;
  wire   n1;

  AOI21_X1 U3 ( .B1(g_prec), .B2(p), .A(g), .ZN(n1) );
  AND2_X1 U1 ( .A1(p), .A2(p_prec), .ZN(p_out) );
  INV_X1 U2 ( .A(n1), .ZN(g_out) );
endmodule


module pg_7 ( g, p, g_prec, p_prec, g_out, p_out );
  input g, p, g_prec, p_prec;
  output g_out, p_out;
  wire   n1;

  AOI21_X1 U3 ( .B1(g_prec), .B2(p), .A(g), .ZN(n1) );
  AND2_X1 U1 ( .A1(p), .A2(p_prec), .ZN(p_out) );
  INV_X1 U2 ( .A(n1), .ZN(g_out) );
endmodule


module pg_6 ( g, p, g_prec, p_prec, g_out, p_out );
  input g, p, g_prec, p_prec;
  output g_out, p_out;
  wire   n1;

  AOI21_X1 U3 ( .B1(g_prec), .B2(p), .A(g), .ZN(n1) );
  AND2_X1 U1 ( .A1(p), .A2(p_prec), .ZN(p_out) );
  INV_X1 U2 ( .A(n1), .ZN(g_out) );
endmodule


module pg_5 ( g, p, g_prec, p_prec, g_out, p_out );
  input g, p, g_prec, p_prec;
  output g_out, p_out;
  wire   n1;

  AOI21_X1 U3 ( .B1(g_prec), .B2(p), .A(g), .ZN(n1) );
  AND2_X1 U1 ( .A1(p), .A2(p_prec), .ZN(p_out) );
  INV_X1 U2 ( .A(n1), .ZN(g_out) );
endmodule


module pg_4 ( g, p, g_prec, p_prec, g_out, p_out );
  input g, p, g_prec, p_prec;
  output g_out, p_out;
  wire   n1;

  AOI21_X1 U3 ( .B1(g_prec), .B2(p), .A(g), .ZN(n1) );
  AND2_X1 U1 ( .A1(p), .A2(p_prec), .ZN(p_out) );
  INV_X1 U2 ( .A(n1), .ZN(g_out) );
endmodule


module pg_3 ( g, p, g_prec, p_prec, g_out, p_out );
  input g, p, g_prec, p_prec;
  output g_out, p_out;
  wire   n1;

  AOI21_X1 U3 ( .B1(g_prec), .B2(p), .A(g), .ZN(n1) );
  AND2_X1 U1 ( .A1(p), .A2(p_prec), .ZN(p_out) );
  INV_X1 U2 ( .A(n1), .ZN(g_out) );
endmodule


module pg_2 ( g, p, g_prec, p_prec, g_out, p_out );
  input g, p, g_prec, p_prec;
  output g_out, p_out;
  wire   n1;

  AOI21_X1 U3 ( .B1(g_prec), .B2(p), .A(g), .ZN(n1) );
  AND2_X1 U1 ( .A1(p), .A2(p_prec), .ZN(p_out) );
  INV_X1 U2 ( .A(n1), .ZN(g_out) );
endmodule


module pg_1 ( g, p, g_prec, p_prec, g_out, p_out );
  input g, p, g_prec, p_prec;
  output g_out, p_out;
  wire   n1;

  AOI21_X1 U3 ( .B1(g_prec), .B2(p), .A(g), .ZN(n1) );
  AND2_X1 U1 ( .A1(p), .A2(p_prec), .ZN(p_out) );
  INV_X1 U2 ( .A(n1), .ZN(g_out) );
endmodule


module g_19 ( g, p, g_prec, g_out );
  input g, p, g_prec;
  output g_out;
  wire   n1;

  AOI21_X1 U2 ( .B1(p), .B2(g_prec), .A(g), .ZN(n1) );
  INV_X1 U1 ( .A(n1), .ZN(g_out) );
endmodule


module g_18 ( g, p, g_prec, g_out );
  input g, p, g_prec;
  output g_out;
  wire   n1;

  AOI21_X1 U2 ( .B1(p), .B2(g_prec), .A(g), .ZN(n1) );
  INV_X1 U1 ( .A(n1), .ZN(g_out) );
endmodule


module g_17 ( g, p, g_prec, g_out );
  input g, p, g_prec;
  output g_out;
  wire   n1;

  AOI21_X1 U2 ( .B1(p), .B2(g_prec), .A(g), .ZN(n1) );
  INV_X1 U1 ( .A(n1), .ZN(g_out) );
endmodule


module g_16 ( g, p, g_prec, g_out );
  input g, p, g_prec;
  output g_out;
  wire   n1;

  AOI21_X1 U2 ( .B1(p), .B2(g_prec), .A(g), .ZN(n1) );
  INV_X1 U1 ( .A(n1), .ZN(g_out) );
endmodule


module g_15 ( g, p, g_prec, g_out );
  input g, p, g_prec;
  output g_out;
  wire   n1;

  AOI21_X1 U2 ( .B1(p), .B2(g_prec), .A(g), .ZN(n1) );
  INV_X1 U1 ( .A(n1), .ZN(g_out) );
endmodule


module g_14 ( g, p, g_prec, g_out );
  input g, p, g_prec;
  output g_out;
  wire   n1;

  AOI21_X1 U2 ( .B1(p), .B2(g_prec), .A(g), .ZN(n1) );
  INV_X1 U1 ( .A(n1), .ZN(g_out) );
endmodule


module g_13 ( g, p, g_prec, g_out );
  input g, p, g_prec;
  output g_out;
  wire   n1;

  AOI21_X1 U2 ( .B1(p), .B2(g_prec), .A(g), .ZN(n1) );
  INV_X1 U1 ( .A(n1), .ZN(g_out) );
endmodule


module g_12 ( g, p, g_prec, g_out );
  input g, p, g_prec;
  output g_out;
  wire   n1;

  AOI21_X1 U2 ( .B1(p), .B2(g_prec), .A(g), .ZN(n1) );
  INV_X1 U1 ( .A(n1), .ZN(g_out) );
endmodule


module g_10 ( g, p, g_prec, g_out );
  input g, p, g_prec;
  output g_out;
  wire   n1;

  AOI21_X1 U2 ( .B1(p), .B2(g_prec), .A(g), .ZN(n1) );
  INV_X1 U1 ( .A(n1), .ZN(g_out) );
endmodule


module g_9 ( g, p, g_prec, g_out );
  input g, p, g_prec;
  output g_out;
  wire   n1;

  AOI21_X1 U2 ( .B1(p), .B2(g_prec), .A(g), .ZN(n1) );
  INV_X1 U1 ( .A(n1), .ZN(g_out) );
endmodule


module g_8 ( g, p, g_prec, g_out );
  input g, p, g_prec;
  output g_out;
  wire   n1;

  AOI21_X1 U2 ( .B1(p), .B2(g_prec), .A(g), .ZN(n1) );
  INV_X1 U1 ( .A(n1), .ZN(g_out) );
endmodule


module g_7 ( g, p, g_prec, g_out );
  input g, p, g_prec;
  output g_out;
  wire   n1;

  AOI21_X1 U2 ( .B1(p), .B2(g_prec), .A(g), .ZN(n1) );
  INV_X1 U1 ( .A(n1), .ZN(g_out) );
endmodule


module g_6 ( g, p, g_prec, g_out );
  input g, p, g_prec;
  output g_out;
  wire   n1;

  AOI21_X1 U2 ( .B1(p), .B2(g_prec), .A(g), .ZN(n1) );
  INV_X1 U1 ( .A(n1), .ZN(g_out) );
endmodule


module g_5 ( g, p, g_prec, g_out );
  input g, p, g_prec;
  output g_out;
  wire   n1;

  AOI21_X1 U2 ( .B1(p), .B2(g_prec), .A(g), .ZN(n1) );
  INV_X1 U1 ( .A(n1), .ZN(g_out) );
endmodule


module g_4 ( g, p, g_prec, g_out );
  input g, p, g_prec;
  output g_out;
  wire   n1;

  AOI21_X1 U2 ( .B1(p), .B2(g_prec), .A(g), .ZN(n1) );
  INV_X1 U1 ( .A(n1), .ZN(g_out) );
endmodule


module g_3 ( g, p, g_prec, g_out );
  input g, p, g_prec;
  output g_out;
  wire   n1;

  AOI21_X1 U2 ( .B1(p), .B2(g_prec), .A(g), .ZN(n1) );
  INV_X1 U1 ( .A(n1), .ZN(g_out) );
endmodule


module g_2 ( g, p, g_prec, g_out );
  input g, p, g_prec;
  output g_out;
  wire   n1;

  AOI21_X1 U2 ( .B1(p), .B2(g_prec), .A(g), .ZN(n1) );
  INV_X1 U1 ( .A(n1), .ZN(g_out) );
endmodule


module g_1 ( g, p, g_prec, g_out );
  input g, p, g_prec;
  output g_out;
  wire   n1;

  AOI21_X1 U2 ( .B1(p), .B2(g_prec), .A(g), .ZN(n1) );
  INV_X1 U1 ( .A(n1), .ZN(g_out) );
endmodule


module pg_net_63 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p_out) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g_out) );
endmodule


module pg_net_62 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p_out) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g_out) );
endmodule


module pg_net_61 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p_out) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g_out) );
endmodule


module pg_net_60 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p_out) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g_out) );
endmodule


module pg_net_59 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p_out) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g_out) );
endmodule


module pg_net_58 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p_out) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g_out) );
endmodule


module pg_net_57 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p_out) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g_out) );
endmodule


module pg_net_56 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p_out) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g_out) );
endmodule


module pg_net_55 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p_out) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g_out) );
endmodule


module pg_net_54 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p_out) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g_out) );
endmodule


module pg_net_53 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p_out) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g_out) );
endmodule


module pg_net_52 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p_out) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g_out) );
endmodule


module pg_net_51 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p_out) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g_out) );
endmodule


module pg_net_50 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p_out) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g_out) );
endmodule


module pg_net_49 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p_out) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g_out) );
endmodule


module pg_net_48 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p_out) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g_out) );
endmodule


module pg_net_47 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p_out) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g_out) );
endmodule


module pg_net_46 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p_out) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g_out) );
endmodule


module pg_net_45 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p_out) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g_out) );
endmodule


module pg_net_44 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p_out) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g_out) );
endmodule


module pg_net_43 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p_out) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g_out) );
endmodule


module pg_net_42 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p_out) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g_out) );
endmodule


module pg_net_41 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p_out) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g_out) );
endmodule


module pg_net_40 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p_out) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g_out) );
endmodule


module pg_net_39 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p_out) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g_out) );
endmodule


module pg_net_38 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p_out) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g_out) );
endmodule


module pg_net_33 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g_out) );
endmodule


module pg_net_32 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p_out) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g_out) );
endmodule


module pg_net_31 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p_out) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g_out) );
endmodule


module pg_net_30 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p_out) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g_out) );
endmodule


module pg_net_29 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p_out) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g_out) );
endmodule


module pg_net_28 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p_out) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g_out) );
endmodule


module pg_net_27 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p_out) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g_out) );
endmodule


module pg_net_26 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p_out) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g_out) );
endmodule


module pg_net_25 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p_out) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g_out) );
endmodule


module pg_net_24 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p_out) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g_out) );
endmodule


module pg_net_23 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p_out) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g_out) );
endmodule


module pg_net_22 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p_out) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g_out) );
endmodule


module pg_net_21 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p_out) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g_out) );
endmodule


module pg_net_20 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p_out) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g_out) );
endmodule


module pg_net_19 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p_out) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g_out) );
endmodule


module pg_net_18 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p_out) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g_out) );
endmodule


module pg_net_17 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p_out) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g_out) );
endmodule


module pg_net_16 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p_out) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g_out) );
endmodule


module pg_net_15 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p_out) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g_out) );
endmodule


module pg_net_14 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p_out) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g_out) );
endmodule


module pg_net_13 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p_out) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g_out) );
endmodule


module pg_net_12 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p_out) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g_out) );
endmodule


module pg_net_11 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p_out) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g_out) );
endmodule


module pg_net_10 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p_out) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g_out) );
endmodule


module pg_net_9 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p_out) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g_out) );
endmodule


module pg_net_8 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p_out) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g_out) );
endmodule


module pg_net_7 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p_out) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g_out) );
endmodule


module pg_net_6 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p_out) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g_out) );
endmodule


module pg_net_5 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p_out) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g_out) );
endmodule


module pg_net_4 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p_out) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g_out) );
endmodule


module pg_net_3 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p_out) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g_out) );
endmodule


module pg_net_2 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p_out) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g_out) );
endmodule


module pg_net_1 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p_out) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g_out) );
endmodule


module sum_gen_N32_1 ( A, B, Cin, S );
  input [31:0] A;
  input [31:0] B;
  input [8:0] Cin;
  output [31:0] S;


  carry_sel_gen_N4_8 csel_N_0 ( .A(A[3:0]), .B(B[3:0]), .Ci(Cin[0]), .S(S[3:0]) );
  carry_sel_gen_N4_7 csel_N_1 ( .A(A[7:4]), .B(B[7:4]), .Ci(Cin[1]), .S(S[7:4]) );
  carry_sel_gen_N4_6 csel_N_2 ( .A(A[11:8]), .B(B[11:8]), .Ci(Cin[2]), .S(
        S[11:8]) );
  carry_sel_gen_N4_5 csel_N_3 ( .A(A[15:12]), .B(B[15:12]), .Ci(Cin[3]), .S(
        S[15:12]) );
  carry_sel_gen_N4_4 csel_N_4 ( .A(A[19:16]), .B(B[19:16]), .Ci(Cin[4]), .S(
        S[19:16]) );
  carry_sel_gen_N4_3 csel_N_5 ( .A(A[23:20]), .B(B[23:20]), .Ci(Cin[5]), .S(
        S[23:20]) );
  carry_sel_gen_N4_2 csel_N_6 ( .A(A[27:24]), .B(B[27:24]), .Ci(Cin[6]), .S(
        S[27:24]) );
  carry_sel_gen_N4_1 csel_N_7 ( .A(A[31:28]), .B(B[31:28]), .Ci(Cin[7]), .S(
        S[31:28]) );
endmodule


module carry_tree_N32_logN5_1 ( A, B, Cin, Cout );
  input [31:0] A;
  input [31:0] B;
  output [7:0] Cout;
  input Cin;
  wire   \pg_1[15][1] , \pg_1[15][0] , \pg_1[14][1] , \pg_1[14][0] ,
         \pg_1[13][1] , \pg_1[13][0] , \pg_1[12][1] , \pg_1[12][0] ,
         \pg_1[11][1] , \pg_1[11][0] , \pg_1[10][1] , \pg_1[10][0] ,
         \pg_1[9][1] , \pg_1[9][0] , \pg_1[8][1] , \pg_1[8][0] , \pg_1[7][1] ,
         \pg_1[7][0] , \pg_1[6][1] , \pg_1[6][0] , \pg_1[5][1] , \pg_1[5][0] ,
         \pg_1[4][1] , \pg_1[4][0] , \pg_1[3][1] , \pg_1[3][0] , \pg_1[2][1] ,
         \pg_1[2][0] , \pg_1[1][1] , \pg_1[1][0] , \pg_1[0][0] ,
         \pg_n[4][7][1] , \pg_n[4][7][0] , \pg_n[4][6][1] , \pg_n[4][6][0] ,
         \pg_n[3][7][1] , \pg_n[3][7][0] , \pg_n[3][5][1] , \pg_n[3][5][0] ,
         \pg_n[3][3][1] , \pg_n[3][3][0] , \pg_n[2][7][1] , \pg_n[2][7][0] ,
         \pg_n[2][6][1] , \pg_n[2][6][0] , \pg_n[2][5][1] , \pg_n[2][5][0] ,
         \pg_n[2][4][1] , \pg_n[2][4][0] , \pg_n[2][3][1] , \pg_n[2][3][0] ,
         \pg_n[2][2][1] , \pg_n[2][2][0] , \pg_n[2][1][1] , \pg_n[2][1][0] ;
  wire   [31:1] p_net;
  wire   [31:0] g_net;
  wire   [1:0] magic_pro;

  pg_net_32 pg_net_x_1 ( .a(A[1]), .b(B[1]), .g_out(g_net[1]), .p_out(p_net[1]) );
  pg_net_31 pg_net_x_2 ( .a(A[2]), .b(B[2]), .g_out(g_net[2]), .p_out(p_net[2]) );
  pg_net_30 pg_net_x_3 ( .a(A[3]), .b(B[3]), .g_out(g_net[3]), .p_out(p_net[3]) );
  pg_net_29 pg_net_x_4 ( .a(A[4]), .b(B[4]), .g_out(g_net[4]), .p_out(p_net[4]) );
  pg_net_28 pg_net_x_5 ( .a(A[5]), .b(B[5]), .g_out(g_net[5]), .p_out(p_net[5]) );
  pg_net_27 pg_net_x_6 ( .a(A[6]), .b(B[6]), .g_out(g_net[6]), .p_out(p_net[6]) );
  pg_net_26 pg_net_x_7 ( .a(A[7]), .b(B[7]), .g_out(g_net[7]), .p_out(p_net[7]) );
  pg_net_25 pg_net_x_8 ( .a(A[8]), .b(B[8]), .g_out(g_net[8]), .p_out(p_net[8]) );
  pg_net_24 pg_net_x_9 ( .a(A[9]), .b(B[9]), .g_out(g_net[9]), .p_out(p_net[9]) );
  pg_net_23 pg_net_x_10 ( .a(A[10]), .b(B[10]), .g_out(g_net[10]), .p_out(
        p_net[10]) );
  pg_net_22 pg_net_x_11 ( .a(A[11]), .b(B[11]), .g_out(g_net[11]), .p_out(
        p_net[11]) );
  pg_net_21 pg_net_x_12 ( .a(A[12]), .b(B[12]), .g_out(g_net[12]), .p_out(
        p_net[12]) );
  pg_net_20 pg_net_x_13 ( .a(A[13]), .b(B[13]), .g_out(g_net[13]), .p_out(
        p_net[13]) );
  pg_net_19 pg_net_x_14 ( .a(A[14]), .b(B[14]), .g_out(g_net[14]), .p_out(
        p_net[14]) );
  pg_net_18 pg_net_x_15 ( .a(A[15]), .b(B[15]), .g_out(g_net[15]), .p_out(
        p_net[15]) );
  pg_net_17 pg_net_x_16 ( .a(A[16]), .b(B[16]), .g_out(g_net[16]), .p_out(
        p_net[16]) );
  pg_net_16 pg_net_x_17 ( .a(A[17]), .b(B[17]), .g_out(g_net[17]), .p_out(
        p_net[17]) );
  pg_net_15 pg_net_x_18 ( .a(A[18]), .b(B[18]), .g_out(g_net[18]), .p_out(
        p_net[18]) );
  pg_net_14 pg_net_x_19 ( .a(A[19]), .b(B[19]), .g_out(g_net[19]), .p_out(
        p_net[19]) );
  pg_net_13 pg_net_x_20 ( .a(A[20]), .b(B[20]), .g_out(g_net[20]), .p_out(
        p_net[20]) );
  pg_net_12 pg_net_x_21 ( .a(A[21]), .b(B[21]), .g_out(g_net[21]), .p_out(
        p_net[21]) );
  pg_net_11 pg_net_x_22 ( .a(A[22]), .b(B[22]), .g_out(g_net[22]), .p_out(
        p_net[22]) );
  pg_net_10 pg_net_x_23 ( .a(A[23]), .b(B[23]), .g_out(g_net[23]), .p_out(
        p_net[23]) );
  pg_net_9 pg_net_x_24 ( .a(A[24]), .b(B[24]), .g_out(g_net[24]), .p_out(
        p_net[24]) );
  pg_net_8 pg_net_x_25 ( .a(A[25]), .b(B[25]), .g_out(g_net[25]), .p_out(
        p_net[25]) );
  pg_net_7 pg_net_x_26 ( .a(A[26]), .b(B[26]), .g_out(g_net[26]), .p_out(
        p_net[26]) );
  pg_net_6 pg_net_x_27 ( .a(A[27]), .b(B[27]), .g_out(g_net[27]), .p_out(
        p_net[27]) );
  pg_net_5 pg_net_x_28 ( .a(A[28]), .b(B[28]), .g_out(g_net[28]), .p_out(
        p_net[28]) );
  pg_net_4 pg_net_x_29 ( .a(A[29]), .b(B[29]), .g_out(g_net[29]), .p_out(
        p_net[29]) );
  pg_net_3 pg_net_x_30 ( .a(A[30]), .b(B[30]), .g_out(g_net[30]), .p_out(
        p_net[30]) );
  pg_net_2 pg_net_x_31 ( .a(A[31]), .b(B[31]), .g_out(g_net[31]), .p_out(
        p_net[31]) );
  pg_net_1 pg_net_0_MAGIC ( .a(A[0]), .b(B[0]), .g_out(magic_pro[0]), .p_out(
        magic_pro[1]) );
  g_10 xG_0_0_MAGIC ( .g(magic_pro[0]), .p(magic_pro[1]), .g_prec(Cin), 
        .g_out(g_net[0]) );
  g_9 xG_1_0 ( .g(g_net[1]), .p(p_net[1]), .g_prec(g_net[0]), .g_out(
        \pg_1[0][0] ) );
  pg_27 xPG_1_1 ( .g(g_net[3]), .p(p_net[3]), .g_prec(g_net[2]), .p_prec(
        p_net[2]), .g_out(\pg_1[1][0] ), .p_out(\pg_1[1][1] ) );
  pg_26 xPG_1_2 ( .g(g_net[5]), .p(p_net[5]), .g_prec(g_net[4]), .p_prec(
        p_net[4]), .g_out(\pg_1[2][0] ), .p_out(\pg_1[2][1] ) );
  pg_25 xPG_1_3 ( .g(g_net[7]), .p(p_net[7]), .g_prec(g_net[6]), .p_prec(
        p_net[6]), .g_out(\pg_1[3][0] ), .p_out(\pg_1[3][1] ) );
  pg_24 xPG_1_4 ( .g(g_net[9]), .p(p_net[9]), .g_prec(g_net[8]), .p_prec(
        p_net[8]), .g_out(\pg_1[4][0] ), .p_out(\pg_1[4][1] ) );
  pg_23 xPG_1_5 ( .g(g_net[11]), .p(p_net[11]), .g_prec(g_net[10]), .p_prec(
        p_net[10]), .g_out(\pg_1[5][0] ), .p_out(\pg_1[5][1] ) );
  pg_22 xPG_1_6 ( .g(g_net[13]), .p(p_net[13]), .g_prec(g_net[12]), .p_prec(
        p_net[12]), .g_out(\pg_1[6][0] ), .p_out(\pg_1[6][1] ) );
  pg_21 xPG_1_7 ( .g(g_net[15]), .p(p_net[15]), .g_prec(g_net[14]), .p_prec(
        p_net[14]), .g_out(\pg_1[7][0] ), .p_out(\pg_1[7][1] ) );
  pg_20 xPG_1_8 ( .g(g_net[17]), .p(p_net[17]), .g_prec(g_net[16]), .p_prec(
        p_net[16]), .g_out(\pg_1[8][0] ), .p_out(\pg_1[8][1] ) );
  pg_19 xPG_1_9 ( .g(g_net[19]), .p(p_net[19]), .g_prec(g_net[18]), .p_prec(
        p_net[18]), .g_out(\pg_1[9][0] ), .p_out(\pg_1[9][1] ) );
  pg_18 xPG_1_10 ( .g(g_net[21]), .p(p_net[21]), .g_prec(g_net[20]), .p_prec(
        p_net[20]), .g_out(\pg_1[10][0] ), .p_out(\pg_1[10][1] ) );
  pg_17 xPG_1_11 ( .g(g_net[23]), .p(p_net[23]), .g_prec(g_net[22]), .p_prec(
        p_net[22]), .g_out(\pg_1[11][0] ), .p_out(\pg_1[11][1] ) );
  pg_16 xPG_1_12 ( .g(g_net[25]), .p(p_net[25]), .g_prec(g_net[24]), .p_prec(
        p_net[24]), .g_out(\pg_1[12][0] ), .p_out(\pg_1[12][1] ) );
  pg_15 xPG_1_13 ( .g(g_net[27]), .p(p_net[27]), .g_prec(g_net[26]), .p_prec(
        p_net[26]), .g_out(\pg_1[13][0] ), .p_out(\pg_1[13][1] ) );
  pg_14 xPG_1_14 ( .g(g_net[29]), .p(p_net[29]), .g_prec(g_net[28]), .p_prec(
        p_net[28]), .g_out(\pg_1[14][0] ), .p_out(\pg_1[14][1] ) );
  pg_13 xPG_1_15 ( .g(g_net[31]), .p(p_net[31]), .g_prec(g_net[30]), .p_prec(
        p_net[30]), .g_out(\pg_1[15][0] ), .p_out(\pg_1[15][1] ) );
  g_8 xG_2_0 ( .g(\pg_1[1][0] ), .p(\pg_1[1][1] ), .g_prec(\pg_1[0][0] ), 
        .g_out(Cout[0]) );
  pg_12 xPG_2_1 ( .g(\pg_1[3][0] ), .p(\pg_1[3][1] ), .g_prec(\pg_1[2][0] ), 
        .p_prec(\pg_1[2][1] ), .g_out(\pg_n[2][1][0] ), .p_out(\pg_n[2][1][1] ) );
  pg_11 xPG_2_2 ( .g(\pg_1[5][0] ), .p(\pg_1[5][1] ), .g_prec(\pg_1[4][0] ), 
        .p_prec(\pg_1[4][1] ), .g_out(\pg_n[2][2][0] ), .p_out(\pg_n[2][2][1] ) );
  pg_10 xPG_2_3 ( .g(\pg_1[7][0] ), .p(\pg_1[7][1] ), .g_prec(\pg_1[6][0] ), 
        .p_prec(\pg_1[6][1] ), .g_out(\pg_n[2][3][0] ), .p_out(\pg_n[2][3][1] ) );
  pg_9 xPG_2_4 ( .g(\pg_1[9][0] ), .p(\pg_1[9][1] ), .g_prec(\pg_1[8][0] ), 
        .p_prec(\pg_1[8][1] ), .g_out(\pg_n[2][4][0] ), .p_out(\pg_n[2][4][1] ) );
  pg_8 xPG_2_5 ( .g(\pg_1[11][0] ), .p(\pg_1[11][1] ), .g_prec(\pg_1[10][0] ), 
        .p_prec(\pg_1[10][1] ), .g_out(\pg_n[2][5][0] ), .p_out(
        \pg_n[2][5][1] ) );
  pg_7 xPG_2_6 ( .g(\pg_1[13][0] ), .p(\pg_1[13][1] ), .g_prec(\pg_1[12][0] ), 
        .p_prec(\pg_1[12][1] ), .g_out(\pg_n[2][6][0] ), .p_out(
        \pg_n[2][6][1] ) );
  pg_6 xPG_2_7 ( .g(\pg_1[15][0] ), .p(\pg_1[15][1] ), .g_prec(\pg_1[14][0] ), 
        .p_prec(\pg_1[14][1] ), .g_out(\pg_n[2][7][0] ), .p_out(
        \pg_n[2][7][1] ) );
  g_7 xG_3_1 ( .g(\pg_n[2][1][0] ), .p(\pg_n[2][1][1] ), .g_prec(Cout[0]), 
        .g_out(Cout[1]) );
  g_6 xG_4_2 ( .g(\pg_n[2][2][0] ), .p(\pg_n[2][2][1] ), .g_prec(Cout[1]), 
        .g_out(Cout[2]) );
  g_5 xG_4_3 ( .g(\pg_n[3][3][0] ), .p(\pg_n[3][3][1] ), .g_prec(Cout[1]), 
        .g_out(Cout[3]) );
  g_4 xG_5_4 ( .g(\pg_n[2][4][0] ), .p(\pg_n[2][4][1] ), .g_prec(Cout[3]), 
        .g_out(Cout[4]) );
  g_3 xG_5_5 ( .g(\pg_n[3][5][0] ), .p(\pg_n[3][5][1] ), .g_prec(Cout[3]), 
        .g_out(Cout[5]) );
  g_2 xG_5_6 ( .g(\pg_n[4][6][0] ), .p(\pg_n[4][6][1] ), .g_prec(Cout[3]), 
        .g_out(Cout[6]) );
  g_1 xG_5_7 ( .g(\pg_n[4][7][0] ), .p(\pg_n[4][7][1] ), .g_prec(Cout[3]), 
        .g_out(Cout[7]) );
  pg_5 xPG_3_3 ( .g(\pg_n[2][3][0] ), .p(\pg_n[2][3][1] ), .g_prec(
        \pg_n[2][2][0] ), .p_prec(\pg_n[2][2][1] ), .g_out(\pg_n[3][3][0] ), 
        .p_out(\pg_n[3][3][1] ) );
  pg_4 xPG_3_5 ( .g(\pg_n[2][5][0] ), .p(\pg_n[2][5][1] ), .g_prec(
        \pg_n[2][4][0] ), .p_prec(\pg_n[2][4][1] ), .g_out(\pg_n[3][5][0] ), 
        .p_out(\pg_n[3][5][1] ) );
  pg_3 xPG_3_7 ( .g(\pg_n[2][7][0] ), .p(\pg_n[2][7][1] ), .g_prec(
        \pg_n[2][6][0] ), .p_prec(\pg_n[2][6][1] ), .g_out(\pg_n[3][7][0] ), 
        .p_out(\pg_n[3][7][1] ) );
  pg_2 xPG_4_6 ( .g(\pg_n[2][6][0] ), .p(\pg_n[2][6][1] ), .g_prec(
        \pg_n[3][5][0] ), .p_prec(\pg_n[3][5][1] ), .g_out(\pg_n[4][6][0] ), 
        .p_out(\pg_n[4][6][1] ) );
  pg_1 xPG_4_7 ( .g(\pg_n[3][7][0] ), .p(\pg_n[3][7][1] ), .g_prec(
        \pg_n[3][5][0] ), .p_prec(\pg_n[3][5][1] ), .g_out(\pg_n[4][7][0] ), 
        .p_out(\pg_n[4][7][1] ) );
endmodule


module xor_gen_N32_1 ( A, B, S );
  input [31:0] A;
  output [31:0] S;
  input B;


  XOR2_X1 U1 ( .A(B), .B(A[9]), .Z(S[9]) );
  XOR2_X1 U2 ( .A(B), .B(A[8]), .Z(S[8]) );
  XOR2_X1 U3 ( .A(B), .B(A[7]), .Z(S[7]) );
  XOR2_X1 U4 ( .A(B), .B(A[6]), .Z(S[6]) );
  XOR2_X1 U5 ( .A(B), .B(A[5]), .Z(S[5]) );
  XOR2_X1 U6 ( .A(B), .B(A[4]), .Z(S[4]) );
  XOR2_X1 U7 ( .A(B), .B(A[3]), .Z(S[3]) );
  XOR2_X1 U8 ( .A(B), .B(A[31]), .Z(S[31]) );
  XOR2_X1 U9 ( .A(B), .B(A[30]), .Z(S[30]) );
  XOR2_X1 U10 ( .A(B), .B(A[2]), .Z(S[2]) );
  XOR2_X1 U11 ( .A(B), .B(A[29]), .Z(S[29]) );
  XOR2_X1 U12 ( .A(B), .B(A[28]), .Z(S[28]) );
  XOR2_X1 U13 ( .A(B), .B(A[27]), .Z(S[27]) );
  XOR2_X1 U14 ( .A(B), .B(A[26]), .Z(S[26]) );
  XOR2_X1 U15 ( .A(B), .B(A[25]), .Z(S[25]) );
  XOR2_X1 U16 ( .A(B), .B(A[24]), .Z(S[24]) );
  XOR2_X1 U17 ( .A(B), .B(A[23]), .Z(S[23]) );
  XOR2_X1 U18 ( .A(B), .B(A[22]), .Z(S[22]) );
  XOR2_X1 U19 ( .A(B), .B(A[21]), .Z(S[21]) );
  XOR2_X1 U20 ( .A(B), .B(A[20]), .Z(S[20]) );
  XOR2_X1 U21 ( .A(B), .B(A[1]), .Z(S[1]) );
  XOR2_X1 U22 ( .A(B), .B(A[19]), .Z(S[19]) );
  XOR2_X1 U23 ( .A(B), .B(A[18]), .Z(S[18]) );
  XOR2_X1 U24 ( .A(B), .B(A[17]), .Z(S[17]) );
  XOR2_X1 U25 ( .A(B), .B(A[16]), .Z(S[16]) );
  XOR2_X1 U26 ( .A(B), .B(A[15]), .Z(S[15]) );
  XOR2_X1 U27 ( .A(B), .B(A[14]), .Z(S[14]) );
  XOR2_X1 U28 ( .A(B), .B(A[13]), .Z(S[13]) );
  XOR2_X1 U29 ( .A(B), .B(A[12]), .Z(S[12]) );
  XOR2_X1 U30 ( .A(B), .B(A[11]), .Z(S[11]) );
  XOR2_X1 U31 ( .A(B), .B(A[10]), .Z(S[10]) );
  XOR2_X1 U32 ( .A(B), .B(A[0]), .Z(S[0]) );
endmodule


module ff32_en_SIZE5_3 ( D, en, clk, rst, Q );
  input [4:0] D;
  output [4:0] Q;
  input en, clk, rst;
  wire   net338012, n5;

  DFFR_X1 \Q_reg[4]  ( .D(D[4]), .CK(net338012), .RN(n5), .Q(Q[4]) );
  DFFR_X1 \Q_reg[3]  ( .D(D[3]), .CK(net338012), .RN(n5), .Q(Q[3]) );
  DFFR_X1 \Q_reg[2]  ( .D(D[2]), .CK(net338012), .RN(n5), .Q(Q[2]) );
  DFFR_X1 \Q_reg[1]  ( .D(D[1]), .CK(net338012), .RN(n5), .Q(Q[1]) );
  DFFR_X1 \Q_reg[0]  ( .D(D[0]), .CK(net338012), .RN(n5), .Q(Q[0]) );
  SNPS_CLOCK_GATE_HIGH_ff32_en_SIZE5_3 clk_gate_Q_reg ( .CLK(clk), .EN(en), 
        .ENCLK(net338012) );
  INV_X1 U2 ( .A(rst), .ZN(n5) );
endmodule


module ff32_en_SIZE5_2 ( D, en, clk, rst, Q );
  input [4:0] D;
  output [4:0] Q;
  input en, clk, rst;
  wire   net338012, n5;

  DFFR_X1 \Q_reg[4]  ( .D(D[4]), .CK(net338012), .RN(n5), .Q(Q[4]) );
  DFFR_X1 \Q_reg[3]  ( .D(D[3]), .CK(net338012), .RN(n5), .Q(Q[3]) );
  DFFR_X1 \Q_reg[2]  ( .D(D[2]), .CK(net338012), .RN(n5), .Q(Q[2]) );
  DFFR_X1 \Q_reg[1]  ( .D(D[1]), .CK(net338012), .RN(n5), .Q(Q[1]) );
  DFFR_X1 \Q_reg[0]  ( .D(D[0]), .CK(net338012), .RN(n5), .Q(Q[0]) );
  SNPS_CLOCK_GATE_HIGH_ff32_en_SIZE5_2 clk_gate_Q_reg ( .CLK(clk), .EN(en), 
        .ENCLK(net338012) );
  INV_X1 U2 ( .A(rst), .ZN(n5) );
endmodule


module ff32_en_SIZE5_1 ( D, en, clk, rst, Q );
  input [4:0] D;
  output [4:0] Q;
  input en, clk, rst;
  wire   n5;

  DFFR_X1 \Q_reg[4]  ( .D(D[4]), .CK(clk), .RN(n5), .Q(Q[4]) );
  DFFR_X1 \Q_reg[3]  ( .D(D[3]), .CK(clk), .RN(n5), .Q(Q[3]) );
  DFFR_X1 \Q_reg[2]  ( .D(D[2]), .CK(clk), .RN(n5), .Q(Q[2]) );
  DFFR_X1 \Q_reg[1]  ( .D(D[1]), .CK(clk), .RN(n5), .Q(Q[1]) );
  DFFR_X1 \Q_reg[0]  ( .D(D[0]), .CK(clk), .RN(n5), .Q(Q[0]) );
  INV_X1 U2 ( .A(rst), .ZN(n5) );
endmodule


module ff32_en_SIZE32_5 ( D, en, clk, rst, Q );
  input [31:0] D;
  output [31:0] Q;
  input en, clk, rst;
  wire   net337997, n32, n34;

  DFFR_X1 \Q_reg[31]  ( .D(D[31]), .CK(net337997), .RN(n34), .Q(Q[31]) );
  DFFR_X1 \Q_reg[30]  ( .D(D[30]), .CK(net337997), .RN(n34), .Q(Q[30]) );
  DFFR_X1 \Q_reg[29]  ( .D(D[29]), .CK(net337997), .RN(n34), .Q(Q[29]) );
  DFFR_X1 \Q_reg[28]  ( .D(D[28]), .CK(net337997), .RN(n34), .Q(Q[28]) );
  DFFR_X1 \Q_reg[27]  ( .D(D[27]), .CK(net337997), .RN(n34), .Q(Q[27]) );
  DFFR_X1 \Q_reg[26]  ( .D(D[26]), .CK(net337997), .RN(n34), .Q(Q[26]) );
  DFFR_X1 \Q_reg[25]  ( .D(D[25]), .CK(net337997), .RN(n34), .Q(Q[25]) );
  DFFR_X1 \Q_reg[24]  ( .D(D[24]), .CK(net337997), .RN(n34), .Q(Q[24]) );
  DFFR_X1 \Q_reg[23]  ( .D(D[23]), .CK(net337997), .RN(n32), .Q(Q[23]) );
  DFFR_X1 \Q_reg[22]  ( .D(D[22]), .CK(net337997), .RN(n34), .Q(Q[22]) );
  DFFR_X1 \Q_reg[21]  ( .D(D[21]), .CK(net337997), .RN(n32), .Q(Q[21]) );
  DFFR_X1 \Q_reg[20]  ( .D(D[20]), .CK(net337997), .RN(n34), .Q(Q[20]) );
  DFFR_X1 \Q_reg[19]  ( .D(D[19]), .CK(net337997), .RN(n32), .Q(Q[19]) );
  DFFR_X1 \Q_reg[18]  ( .D(D[18]), .CK(net337997), .RN(n34), .Q(Q[18]) );
  DFFR_X1 \Q_reg[17]  ( .D(D[17]), .CK(net337997), .RN(n32), .Q(Q[17]) );
  DFFR_X1 \Q_reg[16]  ( .D(D[16]), .CK(net337997), .RN(n34), .Q(Q[16]) );
  DFFR_X1 \Q_reg[15]  ( .D(D[15]), .CK(net337997), .RN(n34), .Q(Q[15]) );
  DFFR_X1 \Q_reg[14]  ( .D(D[14]), .CK(net337997), .RN(n34), .Q(Q[14]) );
  DFFR_X1 \Q_reg[13]  ( .D(D[13]), .CK(net337997), .RN(n34), .Q(Q[13]) );
  DFFR_X1 \Q_reg[12]  ( .D(D[12]), .CK(net337997), .RN(n34), .Q(Q[12]) );
  DFFR_X1 \Q_reg[11]  ( .D(D[11]), .CK(net337997), .RN(n32), .Q(Q[11]) );
  DFFR_X1 \Q_reg[10]  ( .D(D[10]), .CK(net337997), .RN(n32), .Q(Q[10]) );
  DFFR_X1 \Q_reg[9]  ( .D(D[9]), .CK(net337997), .RN(n32), .Q(Q[9]) );
  DFFR_X1 \Q_reg[8]  ( .D(D[8]), .CK(net337997), .RN(n32), .Q(Q[8]) );
  DFFR_X1 \Q_reg[7]  ( .D(D[7]), .CK(net337997), .RN(n32), .Q(Q[7]) );
  DFFR_X1 \Q_reg[6]  ( .D(D[6]), .CK(net337997), .RN(n32), .Q(Q[6]) );
  DFFR_X1 \Q_reg[5]  ( .D(D[5]), .CK(net337997), .RN(n32), .Q(Q[5]) );
  DFFR_X1 \Q_reg[4]  ( .D(D[4]), .CK(net337997), .RN(n32), .Q(Q[4]) );
  DFFR_X1 \Q_reg[3]  ( .D(D[3]), .CK(net337997), .RN(n32), .Q(Q[3]) );
  DFFR_X1 \Q_reg[2]  ( .D(D[2]), .CK(net337997), .RN(n32), .Q(Q[2]) );
  DFFR_X1 \Q_reg[1]  ( .D(D[1]), .CK(net337997), .RN(n32), .Q(Q[1]) );
  DFFR_X1 \Q_reg[0]  ( .D(D[0]), .CK(net337997), .RN(n32), .Q(Q[0]) );
  SNPS_CLOCK_GATE_HIGH_ff32_en_SIZE32_5 clk_gate_Q_reg ( .CLK(clk), .EN(en), 
        .ENCLK(net337997) );
  CLKBUF_X1 U2 ( .A(n34), .Z(n32) );
  INV_X1 U3 ( .A(rst), .ZN(n34) );
endmodule


module ff32_en_SIZE32_4 ( D, en, clk, rst, Q );
  input [31:0] D;
  output [31:0] Q;
  input en, clk, rst;
  wire   net337997, n32, n34;

  DFFR_X1 \Q_reg[31]  ( .D(D[31]), .CK(net337997), .RN(n34), .Q(Q[31]) );
  DFFR_X1 \Q_reg[30]  ( .D(D[30]), .CK(net337997), .RN(n34), .Q(Q[30]) );
  DFFR_X1 \Q_reg[29]  ( .D(D[29]), .CK(net337997), .RN(n34), .Q(Q[29]) );
  DFFR_X1 \Q_reg[28]  ( .D(D[28]), .CK(net337997), .RN(n34), .Q(Q[28]) );
  DFFR_X1 \Q_reg[27]  ( .D(D[27]), .CK(net337997), .RN(n34), .Q(Q[27]) );
  DFFR_X1 \Q_reg[26]  ( .D(D[26]), .CK(net337997), .RN(n34), .Q(Q[26]) );
  DFFR_X1 \Q_reg[25]  ( .D(D[25]), .CK(net337997), .RN(n34), .Q(Q[25]) );
  DFFR_X1 \Q_reg[24]  ( .D(D[24]), .CK(net337997), .RN(n34), .Q(Q[24]) );
  DFFR_X1 \Q_reg[23]  ( .D(D[23]), .CK(net337997), .RN(n32), .Q(Q[23]) );
  DFFR_X1 \Q_reg[22]  ( .D(D[22]), .CK(net337997), .RN(n34), .Q(Q[22]) );
  DFFR_X1 \Q_reg[21]  ( .D(D[21]), .CK(net337997), .RN(n32), .Q(Q[21]) );
  DFFR_X1 \Q_reg[20]  ( .D(D[20]), .CK(net337997), .RN(n34), .Q(Q[20]) );
  DFFR_X1 \Q_reg[19]  ( .D(D[19]), .CK(net337997), .RN(n32), .Q(Q[19]) );
  DFFR_X1 \Q_reg[18]  ( .D(D[18]), .CK(net337997), .RN(n34), .Q(Q[18]) );
  DFFR_X1 \Q_reg[17]  ( .D(D[17]), .CK(net337997), .RN(n32), .Q(Q[17]) );
  DFFR_X1 \Q_reg[16]  ( .D(D[16]), .CK(net337997), .RN(n34), .Q(Q[16]) );
  DFFR_X1 \Q_reg[15]  ( .D(D[15]), .CK(net337997), .RN(n34), .Q(Q[15]) );
  DFFR_X1 \Q_reg[14]  ( .D(D[14]), .CK(net337997), .RN(n34), .Q(Q[14]) );
  DFFR_X1 \Q_reg[13]  ( .D(D[13]), .CK(net337997), .RN(n34), .Q(Q[13]) );
  DFFR_X1 \Q_reg[12]  ( .D(D[12]), .CK(net337997), .RN(n34), .Q(Q[12]) );
  DFFR_X1 \Q_reg[11]  ( .D(D[11]), .CK(net337997), .RN(n32), .Q(Q[11]) );
  DFFR_X1 \Q_reg[10]  ( .D(D[10]), .CK(net337997), .RN(n32), .Q(Q[10]) );
  DFFR_X1 \Q_reg[9]  ( .D(D[9]), .CK(net337997), .RN(n32), .Q(Q[9]) );
  DFFR_X1 \Q_reg[8]  ( .D(D[8]), .CK(net337997), .RN(n32), .Q(Q[8]) );
  DFFR_X1 \Q_reg[7]  ( .D(D[7]), .CK(net337997), .RN(n32), .Q(Q[7]) );
  DFFR_X1 \Q_reg[6]  ( .D(D[6]), .CK(net337997), .RN(n32), .Q(Q[6]) );
  DFFR_X1 \Q_reg[5]  ( .D(D[5]), .CK(net337997), .RN(n32), .Q(Q[5]) );
  DFFR_X1 \Q_reg[4]  ( .D(D[4]), .CK(net337997), .RN(n32), .Q(Q[4]) );
  DFFR_X1 \Q_reg[3]  ( .D(D[3]), .CK(net337997), .RN(n32), .Q(Q[3]) );
  DFFR_X1 \Q_reg[2]  ( .D(D[2]), .CK(net337997), .RN(n32), .Q(Q[2]) );
  DFFR_X1 \Q_reg[1]  ( .D(D[1]), .CK(net337997), .RN(n32), .Q(Q[1]) );
  DFFR_X1 \Q_reg[0]  ( .D(D[0]), .CK(net337997), .RN(n32), .Q(Q[0]) );
  SNPS_CLOCK_GATE_HIGH_ff32_en_SIZE32_4 clk_gate_Q_reg ( .CLK(clk), .EN(en), 
        .ENCLK(net337997) );
  CLKBUF_X1 U2 ( .A(n34), .Z(n32) );
  INV_X1 U3 ( .A(rst), .ZN(n34) );
endmodule


module ff32_en_SIZE32_3 ( D, en, clk, rst, Q );
  input [31:0] D;
  output [31:0] Q;
  input en, clk, rst;
  wire   n32, n34;

  DFFR_X1 \Q_reg[31]  ( .D(D[31]), .CK(clk), .RN(n34), .Q(Q[31]) );
  DFFR_X1 \Q_reg[30]  ( .D(D[30]), .CK(clk), .RN(n34), .Q(Q[30]) );
  DFFR_X1 \Q_reg[29]  ( .D(D[29]), .CK(clk), .RN(n34), .Q(Q[29]) );
  DFFR_X1 \Q_reg[28]  ( .D(D[28]), .CK(clk), .RN(n34), .Q(Q[28]) );
  DFFR_X1 \Q_reg[27]  ( .D(D[27]), .CK(clk), .RN(n34), .Q(Q[27]) );
  DFFR_X1 \Q_reg[26]  ( .D(D[26]), .CK(clk), .RN(n34), .Q(Q[26]) );
  DFFR_X1 \Q_reg[25]  ( .D(D[25]), .CK(clk), .RN(n34), .Q(Q[25]) );
  DFFR_X1 \Q_reg[24]  ( .D(D[24]), .CK(clk), .RN(n34), .Q(Q[24]) );
  DFFR_X1 \Q_reg[23]  ( .D(D[23]), .CK(clk), .RN(n32), .Q(Q[23]) );
  DFFR_X1 \Q_reg[22]  ( .D(D[22]), .CK(clk), .RN(n34), .Q(Q[22]) );
  DFFR_X1 \Q_reg[21]  ( .D(D[21]), .CK(clk), .RN(n32), .Q(Q[21]) );
  DFFR_X1 \Q_reg[20]  ( .D(D[20]), .CK(clk), .RN(n34), .Q(Q[20]) );
  DFFR_X1 \Q_reg[19]  ( .D(D[19]), .CK(clk), .RN(n32), .Q(Q[19]) );
  DFFR_X1 \Q_reg[18]  ( .D(D[18]), .CK(clk), .RN(n34), .Q(Q[18]) );
  DFFR_X1 \Q_reg[17]  ( .D(D[17]), .CK(clk), .RN(n32), .Q(Q[17]) );
  DFFR_X1 \Q_reg[16]  ( .D(D[16]), .CK(clk), .RN(n34), .Q(Q[16]) );
  DFFR_X1 \Q_reg[15]  ( .D(D[15]), .CK(clk), .RN(n34), .Q(Q[15]) );
  DFFR_X1 \Q_reg[14]  ( .D(D[14]), .CK(clk), .RN(n34), .Q(Q[14]) );
  DFFR_X1 \Q_reg[13]  ( .D(D[13]), .CK(clk), .RN(n34), .Q(Q[13]) );
  DFFR_X1 \Q_reg[12]  ( .D(D[12]), .CK(clk), .RN(n34), .Q(Q[12]) );
  DFFR_X1 \Q_reg[11]  ( .D(D[11]), .CK(clk), .RN(n32), .Q(Q[11]) );
  DFFR_X1 \Q_reg[10]  ( .D(D[10]), .CK(clk), .RN(n32), .Q(Q[10]) );
  DFFR_X1 \Q_reg[9]  ( .D(D[9]), .CK(clk), .RN(n32), .Q(Q[9]) );
  DFFR_X1 \Q_reg[8]  ( .D(D[8]), .CK(clk), .RN(n32), .Q(Q[8]) );
  DFFR_X1 \Q_reg[7]  ( .D(D[7]), .CK(clk), .RN(n32), .Q(Q[7]) );
  DFFR_X1 \Q_reg[6]  ( .D(D[6]), .CK(clk), .RN(n32), .Q(Q[6]) );
  DFFR_X1 \Q_reg[5]  ( .D(D[5]), .CK(clk), .RN(n32), .Q(Q[5]) );
  DFFR_X1 \Q_reg[4]  ( .D(D[4]), .CK(clk), .RN(n32), .Q(Q[4]) );
  DFFR_X1 \Q_reg[3]  ( .D(D[3]), .CK(clk), .RN(n32), .Q(Q[3]) );
  DFFR_X1 \Q_reg[2]  ( .D(D[2]), .CK(clk), .RN(n32), .Q(Q[2]) );
  DFFR_X1 \Q_reg[1]  ( .D(D[1]), .CK(clk), .RN(n32), .Q(Q[1]) );
  DFFR_X1 \Q_reg[0]  ( .D(D[0]), .CK(clk), .RN(n32), .Q(Q[0]) );
  CLKBUF_X1 U2 ( .A(n34), .Z(n32) );
  INV_X1 U3 ( .A(rst), .ZN(n34) );
endmodule


module ff32_en_SIZE32_2 ( D, en, clk, rst, Q );
  input [31:0] D;
  output [31:0] Q;
  input en, clk, rst;
  wire   n32, n34;

  DFFR_X1 \Q_reg[31]  ( .D(D[31]), .CK(clk), .RN(n34), .Q(Q[31]) );
  DFFR_X1 \Q_reg[30]  ( .D(D[30]), .CK(clk), .RN(n34), .Q(Q[30]) );
  DFFR_X1 \Q_reg[29]  ( .D(D[29]), .CK(clk), .RN(n34), .Q(Q[29]) );
  DFFR_X1 \Q_reg[28]  ( .D(D[28]), .CK(clk), .RN(n34), .Q(Q[28]) );
  DFFR_X1 \Q_reg[27]  ( .D(D[27]), .CK(clk), .RN(n34), .Q(Q[27]) );
  DFFR_X1 \Q_reg[26]  ( .D(D[26]), .CK(clk), .RN(n34), .Q(Q[26]) );
  DFFR_X1 \Q_reg[25]  ( .D(D[25]), .CK(clk), .RN(n34), .Q(Q[25]) );
  DFFR_X1 \Q_reg[24]  ( .D(D[24]), .CK(clk), .RN(n34), .Q(Q[24]) );
  DFFR_X1 \Q_reg[23]  ( .D(D[23]), .CK(clk), .RN(n32), .Q(Q[23]) );
  DFFR_X1 \Q_reg[22]  ( .D(D[22]), .CK(clk), .RN(n34), .Q(Q[22]) );
  DFFR_X1 \Q_reg[21]  ( .D(D[21]), .CK(clk), .RN(n32), .Q(Q[21]) );
  DFFR_X1 \Q_reg[20]  ( .D(D[20]), .CK(clk), .RN(n34), .Q(Q[20]) );
  DFFR_X1 \Q_reg[19]  ( .D(D[19]), .CK(clk), .RN(n32), .Q(Q[19]) );
  DFFR_X1 \Q_reg[18]  ( .D(D[18]), .CK(clk), .RN(n34), .Q(Q[18]) );
  DFFR_X1 \Q_reg[17]  ( .D(D[17]), .CK(clk), .RN(n32), .Q(Q[17]) );
  DFFR_X1 \Q_reg[16]  ( .D(D[16]), .CK(clk), .RN(n34), .Q(Q[16]) );
  DFFR_X1 \Q_reg[15]  ( .D(D[15]), .CK(clk), .RN(n34), .Q(Q[15]) );
  DFFR_X1 \Q_reg[14]  ( .D(D[14]), .CK(clk), .RN(n34), .Q(Q[14]) );
  DFFR_X1 \Q_reg[13]  ( .D(D[13]), .CK(clk), .RN(n34), .Q(Q[13]) );
  DFFR_X1 \Q_reg[12]  ( .D(D[12]), .CK(clk), .RN(n34), .Q(Q[12]) );
  DFFR_X1 \Q_reg[11]  ( .D(D[11]), .CK(clk), .RN(n32), .Q(Q[11]) );
  DFFR_X1 \Q_reg[10]  ( .D(D[10]), .CK(clk), .RN(n32), .Q(Q[10]) );
  DFFR_X1 \Q_reg[9]  ( .D(D[9]), .CK(clk), .RN(n32), .Q(Q[9]) );
  DFFR_X1 \Q_reg[8]  ( .D(D[8]), .CK(clk), .RN(n32), .Q(Q[8]) );
  DFFR_X1 \Q_reg[7]  ( .D(D[7]), .CK(clk), .RN(n32), .Q(Q[7]) );
  DFFR_X1 \Q_reg[6]  ( .D(D[6]), .CK(clk), .RN(n32), .Q(Q[6]) );
  DFFR_X1 \Q_reg[5]  ( .D(D[5]), .CK(clk), .RN(n32), .Q(Q[5]) );
  DFFR_X1 \Q_reg[4]  ( .D(D[4]), .CK(clk), .RN(n32), .Q(Q[4]) );
  DFFR_X1 \Q_reg[3]  ( .D(D[3]), .CK(clk), .RN(n32), .Q(Q[3]) );
  DFFR_X1 \Q_reg[2]  ( .D(D[2]), .CK(clk), .RN(n32), .Q(Q[2]) );
  DFFR_X1 \Q_reg[1]  ( .D(D[1]), .CK(clk), .RN(n32), .Q(Q[1]) );
  DFFR_X1 \Q_reg[0]  ( .D(D[0]), .CK(clk), .RN(n32), .Q(Q[0]) );
  CLKBUF_X1 U2 ( .A(n34), .Z(n32) );
  INV_X1 U3 ( .A(rst), .ZN(n34) );
endmodule


module ff32_en_SIZE32_1 ( D, en, clk, rst, Q );
  input [31:0] D;
  output [31:0] Q;
  input en, clk, rst;
  wire   net337997, n32, n34;

  DFFR_X1 \Q_reg[31]  ( .D(D[31]), .CK(net337997), .RN(n34), .Q(Q[31]) );
  DFFR_X1 \Q_reg[30]  ( .D(D[30]), .CK(net337997), .RN(n34), .Q(Q[30]) );
  DFFR_X1 \Q_reg[29]  ( .D(D[29]), .CK(net337997), .RN(n34), .Q(Q[29]) );
  DFFR_X1 \Q_reg[28]  ( .D(D[28]), .CK(net337997), .RN(n34), .Q(Q[28]) );
  DFFR_X1 \Q_reg[27]  ( .D(D[27]), .CK(net337997), .RN(n34), .Q(Q[27]) );
  DFFR_X1 \Q_reg[26]  ( .D(D[26]), .CK(net337997), .RN(n34), .Q(Q[26]) );
  DFFR_X1 \Q_reg[25]  ( .D(D[25]), .CK(net337997), .RN(n34), .Q(Q[25]) );
  DFFR_X1 \Q_reg[24]  ( .D(D[24]), .CK(net337997), .RN(n34), .Q(Q[24]) );
  DFFR_X1 \Q_reg[23]  ( .D(D[23]), .CK(net337997), .RN(n32), .Q(Q[23]) );
  DFFR_X1 \Q_reg[22]  ( .D(D[22]), .CK(net337997), .RN(n34), .Q(Q[22]) );
  DFFR_X1 \Q_reg[21]  ( .D(D[21]), .CK(net337997), .RN(n32), .Q(Q[21]) );
  DFFR_X1 \Q_reg[20]  ( .D(D[20]), .CK(net337997), .RN(n34), .Q(Q[20]) );
  DFFR_X1 \Q_reg[19]  ( .D(D[19]), .CK(net337997), .RN(n32), .Q(Q[19]) );
  DFFR_X1 \Q_reg[18]  ( .D(D[18]), .CK(net337997), .RN(n34), .Q(Q[18]) );
  DFFR_X1 \Q_reg[17]  ( .D(D[17]), .CK(net337997), .RN(n32), .Q(Q[17]) );
  DFFR_X1 \Q_reg[16]  ( .D(D[16]), .CK(net337997), .RN(n34), .Q(Q[16]) );
  DFFR_X1 \Q_reg[15]  ( .D(D[15]), .CK(net337997), .RN(n34), .Q(Q[15]) );
  DFFR_X1 \Q_reg[14]  ( .D(D[14]), .CK(net337997), .RN(n34), .Q(Q[14]) );
  DFFR_X1 \Q_reg[13]  ( .D(D[13]), .CK(net337997), .RN(n34), .Q(Q[13]) );
  DFFR_X1 \Q_reg[12]  ( .D(D[12]), .CK(net337997), .RN(n34), .Q(Q[12]) );
  DFFR_X1 \Q_reg[11]  ( .D(D[11]), .CK(net337997), .RN(n32), .Q(Q[11]) );
  DFFR_X1 \Q_reg[10]  ( .D(D[10]), .CK(net337997), .RN(n32), .Q(Q[10]) );
  DFFR_X1 \Q_reg[9]  ( .D(D[9]), .CK(net337997), .RN(n32), .Q(Q[9]) );
  DFFR_X1 \Q_reg[8]  ( .D(D[8]), .CK(net337997), .RN(n32), .Q(Q[8]) );
  DFFR_X1 \Q_reg[7]  ( .D(D[7]), .CK(net337997), .RN(n32), .Q(Q[7]) );
  DFFR_X1 \Q_reg[6]  ( .D(D[6]), .CK(net337997), .RN(n32), .Q(Q[6]) );
  DFFR_X1 \Q_reg[5]  ( .D(D[5]), .CK(net337997), .RN(n32), .Q(Q[5]) );
  DFFR_X1 \Q_reg[4]  ( .D(D[4]), .CK(net337997), .RN(n32), .Q(Q[4]) );
  DFFR_X1 \Q_reg[3]  ( .D(D[3]), .CK(net337997), .RN(n32), .Q(Q[3]) );
  DFFR_X1 \Q_reg[2]  ( .D(D[2]), .CK(net337997), .RN(n32), .Q(Q[2]) );
  DFFR_X1 \Q_reg[1]  ( .D(D[1]), .CK(net337997), .RN(n32), .Q(Q[1]) );
  DFFR_X1 \Q_reg[0]  ( .D(D[0]), .CK(net337997), .RN(n32), .Q(Q[0]) );
  SNPS_CLOCK_GATE_HIGH_ff32_en_SIZE32_1 clk_gate_Q_reg ( .CLK(clk), .EN(en), 
        .ENCLK(net337997) );
  CLKBUF_X1 U2 ( .A(n34), .Z(n32) );
  INV_X1 U3 ( .A(rst), .ZN(n34) );
endmodule


module mux41_MUX_SIZE32_2 ( IN0, IN1, IN2, IN3, CTRL, OUT1 );
  input [31:0] IN0;
  input [31:0] IN1;
  input [31:0] IN2;
  input [31:0] IN3;
  input [1:0] CTRL;
  output [31:0] OUT1;
  wire   n1, n2, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141;

  NOR2_X1 U99 ( .A1(CTRL[0]), .A2(CTRL[1]), .ZN(n136) );
  AOI22_X1 U98 ( .A1(n137), .A2(IN1[0]), .B1(n1), .B2(IN0[0]), .ZN(n75) );
  AOI22_X1 U95 ( .A1(n72), .A2(IN3[0]), .B1(n2), .B2(IN2[0]), .ZN(n74) );
  NAND2_X1 U94 ( .A1(n75), .A2(n74), .ZN(OUT1[0]) );
  AOI22_X1 U63 ( .A1(n137), .A2(IN1[1]), .B1(n1), .B2(IN0[1]), .ZN(n97) );
  AOI22_X1 U62 ( .A1(n72), .A2(IN3[1]), .B1(n2), .B2(IN2[1]), .ZN(n96) );
  NAND2_X1 U61 ( .A1(n97), .A2(n96), .ZN(OUT1[1]) );
  AOI22_X1 U66 ( .A1(n137), .A2(IN1[19]), .B1(n1), .B2(IN0[19]), .ZN(n95) );
  AOI22_X1 U65 ( .A1(n72), .A2(IN3[19]), .B1(n2), .B2(IN2[19]), .ZN(n94) );
  NAND2_X1 U64 ( .A1(n95), .A2(n94), .ZN(OUT1[19]) );
  AOI22_X1 U75 ( .A1(n137), .A2(IN1[16]), .B1(n1), .B2(IN0[16]), .ZN(n89) );
  AOI22_X1 U74 ( .A1(n72), .A2(IN3[16]), .B1(n2), .B2(IN2[16]), .ZN(n88) );
  NAND2_X1 U73 ( .A1(n89), .A2(n88), .ZN(OUT1[16]) );
  AOI22_X1 U72 ( .A1(n137), .A2(IN1[17]), .B1(n1), .B2(IN0[17]), .ZN(n91) );
  AOI22_X1 U71 ( .A1(n72), .A2(IN3[17]), .B1(n2), .B2(IN2[17]), .ZN(n90) );
  NAND2_X1 U70 ( .A1(n91), .A2(n90), .ZN(OUT1[17]) );
  AOI22_X1 U69 ( .A1(n137), .A2(IN1[18]), .B1(n1), .B2(IN0[18]), .ZN(n93) );
  AOI22_X1 U68 ( .A1(n72), .A2(IN3[18]), .B1(n2), .B2(IN2[18]), .ZN(n92) );
  NAND2_X1 U67 ( .A1(n93), .A2(n92), .ZN(OUT1[18]) );
  AOI22_X1 U78 ( .A1(n137), .A2(IN1[15]), .B1(n1), .B2(IN0[15]), .ZN(n87) );
  AOI22_X1 U77 ( .A1(n72), .A2(IN3[15]), .B1(n2), .B2(IN2[15]), .ZN(n86) );
  AOI22_X1 U81 ( .A1(n137), .A2(IN1[14]), .B1(n1), .B2(IN0[14]), .ZN(n85) );
  AOI22_X1 U80 ( .A1(n72), .A2(IN3[14]), .B1(n2), .B2(IN2[14]), .ZN(n84) );
  AOI22_X1 U84 ( .A1(n137), .A2(IN1[13]), .B1(n1), .B2(IN0[13]), .ZN(n83) );
  AOI22_X1 U83 ( .A1(n72), .A2(IN3[13]), .B1(n2), .B2(IN2[13]), .ZN(n82) );
  AOI22_X1 U87 ( .A1(n137), .A2(IN1[12]), .B1(n1), .B2(IN0[12]), .ZN(n81) );
  AOI22_X1 U86 ( .A1(n72), .A2(IN3[12]), .B1(n2), .B2(IN2[12]), .ZN(n80) );
  AOI22_X1 U90 ( .A1(n137), .A2(IN1[11]), .B1(n1), .B2(IN0[11]), .ZN(n79) );
  AOI22_X1 U89 ( .A1(n72), .A2(IN3[11]), .B1(n2), .B2(IN2[11]), .ZN(n78) );
  AOI22_X1 U93 ( .A1(n137), .A2(IN1[10]), .B1(n1), .B2(IN0[10]), .ZN(n77) );
  AOI22_X1 U92 ( .A1(n72), .A2(IN3[10]), .B1(n2), .B2(IN2[10]), .ZN(n76) );
  AOI22_X1 U3 ( .A1(n137), .A2(IN1[9]), .B1(n136), .B2(IN0[9]), .ZN(n141) );
  AOI22_X1 U2 ( .A1(n139), .A2(IN3[9]), .B1(n138), .B2(IN2[9]), .ZN(n140) );
  AOI22_X1 U6 ( .A1(n137), .A2(IN1[8]), .B1(n136), .B2(IN0[8]), .ZN(n135) );
  AOI22_X1 U5 ( .A1(n139), .A2(IN3[8]), .B1(n2), .B2(IN2[8]), .ZN(n134) );
  AOI22_X1 U9 ( .A1(n137), .A2(IN1[7]), .B1(n1), .B2(IN0[7]), .ZN(n133) );
  AOI22_X1 U8 ( .A1(n139), .A2(IN3[7]), .B1(n138), .B2(IN2[7]), .ZN(n132) );
  AOI22_X1 U12 ( .A1(n137), .A2(IN1[6]), .B1(n136), .B2(IN0[6]), .ZN(n131) );
  AOI22_X1 U11 ( .A1(n139), .A2(IN3[6]), .B1(n138), .B2(IN2[6]), .ZN(n130) );
  AOI22_X1 U15 ( .A1(n137), .A2(IN1[5]), .B1(n1), .B2(IN0[5]), .ZN(n129) );
  AOI22_X1 U14 ( .A1(n72), .A2(IN3[5]), .B1(n138), .B2(IN2[5]), .ZN(n128) );
  NAND2_X1 U13 ( .A1(n129), .A2(n128), .ZN(OUT1[5]) );
  AOI22_X1 U18 ( .A1(n137), .A2(IN1[4]), .B1(n136), .B2(IN0[4]), .ZN(n127) );
  AOI22_X1 U17 ( .A1(n139), .A2(IN3[4]), .B1(n2), .B2(IN2[4]), .ZN(n126) );
  AOI22_X1 U21 ( .A1(n137), .A2(IN1[3]), .B1(n1), .B2(IN0[3]), .ZN(n125) );
  AOI22_X1 U20 ( .A1(n72), .A2(IN3[3]), .B1(n2), .B2(IN2[3]), .ZN(n124) );
  NAND2_X1 U19 ( .A1(n125), .A2(n124), .ZN(OUT1[3]) );
  AOI22_X1 U30 ( .A1(n137), .A2(IN1[2]), .B1(n136), .B2(IN0[2]), .ZN(n119) );
  AOI22_X1 U29 ( .A1(n139), .A2(IN3[2]), .B1(n138), .B2(IN2[2]), .ZN(n118) );
  AOI22_X1 U51 ( .A1(n137), .A2(IN1[23]), .B1(n136), .B2(IN0[23]), .ZN(n105)
         );
  AOI22_X1 U50 ( .A1(n139), .A2(IN3[23]), .B1(n138), .B2(IN2[23]), .ZN(n104)
         );
  NAND2_X1 U49 ( .A1(n105), .A2(n104), .ZN(OUT1[23]) );
  AOI22_X1 U60 ( .A1(n137), .A2(IN1[20]), .B1(n1), .B2(IN0[20]), .ZN(n99) );
  AOI22_X1 U59 ( .A1(n139), .A2(IN3[20]), .B1(n2), .B2(IN2[20]), .ZN(n98) );
  NAND2_X1 U58 ( .A1(n99), .A2(n98), .ZN(OUT1[20]) );
  AOI22_X1 U57 ( .A1(n137), .A2(IN1[21]), .B1(n136), .B2(IN0[21]), .ZN(n101)
         );
  AOI22_X1 U56 ( .A1(n139), .A2(IN3[21]), .B1(n138), .B2(IN2[21]), .ZN(n100)
         );
  NAND2_X1 U55 ( .A1(n101), .A2(n100), .ZN(OUT1[21]) );
  AOI22_X1 U54 ( .A1(n137), .A2(IN1[22]), .B1(n1), .B2(IN0[22]), .ZN(n103) );
  AOI22_X1 U53 ( .A1(n139), .A2(IN3[22]), .B1(n2), .B2(IN2[22]), .ZN(n102) );
  NAND2_X1 U52 ( .A1(n103), .A2(n102), .ZN(OUT1[22]) );
  AOI22_X1 U24 ( .A1(n137), .A2(IN1[31]), .B1(n1), .B2(IN0[31]), .ZN(n123) );
  AOI22_X1 U23 ( .A1(n72), .A2(IN3[31]), .B1(n2), .B2(IN2[31]), .ZN(n122) );
  NAND2_X1 U22 ( .A1(n123), .A2(n122), .ZN(OUT1[31]) );
  AOI22_X1 U36 ( .A1(n137), .A2(IN1[28]), .B1(n1), .B2(IN0[28]), .ZN(n115) );
  AOI22_X1 U35 ( .A1(n139), .A2(IN3[28]), .B1(n2), .B2(IN2[28]), .ZN(n114) );
  NAND2_X1 U34 ( .A1(n115), .A2(n114), .ZN(OUT1[28]) );
  AOI22_X1 U33 ( .A1(n137), .A2(IN1[29]), .B1(n1), .B2(IN0[29]), .ZN(n117) );
  AOI22_X1 U32 ( .A1(n72), .A2(IN3[29]), .B1(n2), .B2(IN2[29]), .ZN(n116) );
  NAND2_X1 U31 ( .A1(n117), .A2(n116), .ZN(OUT1[29]) );
  AOI22_X1 U27 ( .A1(n137), .A2(IN1[30]), .B1(n1), .B2(IN0[30]), .ZN(n121) );
  AOI22_X1 U26 ( .A1(n72), .A2(IN3[30]), .B1(n2), .B2(IN2[30]), .ZN(n120) );
  NAND2_X1 U25 ( .A1(n121), .A2(n120), .ZN(OUT1[30]) );
  AOI22_X1 U39 ( .A1(n137), .A2(IN1[27]), .B1(n1), .B2(IN0[27]), .ZN(n113) );
  AOI22_X1 U38 ( .A1(n139), .A2(IN3[27]), .B1(n2), .B2(IN2[27]), .ZN(n112) );
  NAND2_X1 U37 ( .A1(n113), .A2(n112), .ZN(OUT1[27]) );
  AOI22_X1 U42 ( .A1(n137), .A2(IN1[26]), .B1(n1), .B2(IN0[26]), .ZN(n111) );
  AOI22_X1 U41 ( .A1(n139), .A2(IN3[26]), .B1(n2), .B2(IN2[26]), .ZN(n110) );
  NAND2_X1 U40 ( .A1(n111), .A2(n110), .ZN(OUT1[26]) );
  AOI22_X1 U45 ( .A1(n137), .A2(IN1[25]), .B1(n1), .B2(IN0[25]), .ZN(n109) );
  AOI22_X1 U44 ( .A1(n139), .A2(IN3[25]), .B1(n2), .B2(IN2[25]), .ZN(n108) );
  NAND2_X1 U43 ( .A1(n109), .A2(n108), .ZN(OUT1[25]) );
  AOI22_X1 U48 ( .A1(n137), .A2(IN1[24]), .B1(n1), .B2(IN0[24]), .ZN(n107) );
  AOI22_X1 U47 ( .A1(n139), .A2(IN3[24]), .B1(n2), .B2(IN2[24]), .ZN(n106) );
  NAND2_X1 U46 ( .A1(n107), .A2(n106), .ZN(OUT1[24]) );
  NAND2_X1 U79 ( .A1(n85), .A2(n84), .ZN(OUT1[14]) );
  NAND2_X1 U82 ( .A1(n83), .A2(n82), .ZN(OUT1[13]) );
  NAND2_X1 U85 ( .A1(n81), .A2(n80), .ZN(OUT1[12]) );
  NAND2_X1 U88 ( .A1(n79), .A2(n78), .ZN(OUT1[11]) );
  NAND2_X1 U91 ( .A1(n77), .A2(n76), .ZN(OUT1[10]) );
  NAND2_X1 U1 ( .A1(n141), .A2(n140), .ZN(OUT1[9]) );
  NAND2_X1 U4 ( .A1(n135), .A2(n134), .ZN(OUT1[8]) );
  NAND2_X1 U7 ( .A1(n133), .A2(n132), .ZN(OUT1[7]) );
  NAND2_X1 U10 ( .A1(n131), .A2(n130), .ZN(OUT1[6]) );
  NAND2_X1 U16 ( .A1(n127), .A2(n126), .ZN(OUT1[4]) );
  NAND2_X1 U28 ( .A1(n119), .A2(n118), .ZN(OUT1[2]) );
  NAND2_X1 U76 ( .A1(n87), .A2(n86), .ZN(OUT1[15]) );
  NOR2_X1 U96 ( .A1(CTRL[0]), .A2(n73), .ZN(n138) );
  INV_X1 U101 ( .A(CTRL[1]), .ZN(n73) );
  BUF_X1 U97 ( .A(n138), .Z(n2) );
  BUF_X1 U100 ( .A(n136), .Z(n1) );
  BUF_X1 U102 ( .A(n139), .Z(n72) );
  AND2_X2 U103 ( .A1(n73), .A2(CTRL[0]), .ZN(n137) );
  AND2_X1 U104 ( .A1(CTRL[0]), .A2(CTRL[1]), .ZN(n139) );
endmodule


module mux41_MUX_SIZE32_1 ( IN0, IN1, IN2, IN3, CTRL, OUT1 );
  input [31:0] IN0;
  input [31:0] IN1;
  input [31:0] IN2;
  input [31:0] IN3;
  input [1:0] CTRL;
  output [31:0] OUT1;
  wire   n1, n2, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141;

  AOI22_X1 U98 ( .A1(n137), .A2(IN1[0]), .B1(n136), .B2(IN0[0]), .ZN(n75) );
  AOI22_X1 U95 ( .A1(n1), .A2(IN3[0]), .B1(n72), .B2(IN2[0]), .ZN(n74) );
  NAND2_X1 U94 ( .A1(n75), .A2(n74), .ZN(OUT1[0]) );
  AOI22_X1 U63 ( .A1(n137), .A2(IN1[1]), .B1(n2), .B2(IN0[1]), .ZN(n97) );
  AOI22_X1 U62 ( .A1(n1), .A2(IN3[1]), .B1(n72), .B2(IN2[1]), .ZN(n96) );
  NAND2_X1 U61 ( .A1(n97), .A2(n96), .ZN(OUT1[1]) );
  AOI22_X1 U75 ( .A1(n137), .A2(IN1[16]), .B1(n2), .B2(IN0[16]), .ZN(n89) );
  AOI22_X1 U74 ( .A1(n1), .A2(IN3[16]), .B1(n72), .B2(IN2[16]), .ZN(n88) );
  NAND2_X1 U73 ( .A1(n89), .A2(n88), .ZN(OUT1[16]) );
  AOI22_X1 U72 ( .A1(n137), .A2(IN1[17]), .B1(n136), .B2(IN0[17]), .ZN(n91) );
  AOI22_X1 U71 ( .A1(n1), .A2(IN3[17]), .B1(n72), .B2(IN2[17]), .ZN(n90) );
  NAND2_X1 U70 ( .A1(n91), .A2(n90), .ZN(OUT1[17]) );
  AOI22_X1 U69 ( .A1(n137), .A2(IN1[18]), .B1(n136), .B2(IN0[18]), .ZN(n93) );
  AOI22_X1 U68 ( .A1(n1), .A2(IN3[18]), .B1(n72), .B2(IN2[18]), .ZN(n92) );
  NAND2_X1 U67 ( .A1(n93), .A2(n92), .ZN(OUT1[18]) );
  AOI22_X1 U66 ( .A1(n137), .A2(IN1[19]), .B1(n136), .B2(IN0[19]), .ZN(n95) );
  AOI22_X1 U65 ( .A1(n1), .A2(IN3[19]), .B1(n72), .B2(IN2[19]), .ZN(n94) );
  NAND2_X1 U64 ( .A1(n95), .A2(n94), .ZN(OUT1[19]) );
  AOI22_X1 U78 ( .A1(n137), .A2(IN1[15]), .B1(n2), .B2(IN0[15]), .ZN(n87) );
  AOI22_X1 U77 ( .A1(n1), .A2(IN3[15]), .B1(n72), .B2(IN2[15]), .ZN(n86) );
  NAND2_X1 U76 ( .A1(n87), .A2(n86), .ZN(OUT1[15]) );
  AOI22_X1 U81 ( .A1(n137), .A2(IN1[14]), .B1(n2), .B2(IN0[14]), .ZN(n85) );
  AOI22_X1 U80 ( .A1(n1), .A2(IN3[14]), .B1(n72), .B2(IN2[14]), .ZN(n84) );
  NAND2_X1 U79 ( .A1(n85), .A2(n84), .ZN(OUT1[14]) );
  AOI22_X1 U84 ( .A1(n137), .A2(IN1[13]), .B1(n2), .B2(IN0[13]), .ZN(n83) );
  AOI22_X1 U83 ( .A1(n1), .A2(IN3[13]), .B1(n72), .B2(IN2[13]), .ZN(n82) );
  NAND2_X1 U82 ( .A1(n83), .A2(n82), .ZN(OUT1[13]) );
  AOI22_X1 U87 ( .A1(n137), .A2(IN1[12]), .B1(n136), .B2(IN0[12]), .ZN(n81) );
  AOI22_X1 U86 ( .A1(n1), .A2(IN3[12]), .B1(n72), .B2(IN2[12]), .ZN(n80) );
  NAND2_X1 U85 ( .A1(n81), .A2(n80), .ZN(OUT1[12]) );
  AOI22_X1 U90 ( .A1(n137), .A2(IN1[11]), .B1(n136), .B2(IN0[11]), .ZN(n79) );
  AOI22_X1 U89 ( .A1(n1), .A2(IN3[11]), .B1(n72), .B2(IN2[11]), .ZN(n78) );
  NAND2_X1 U88 ( .A1(n79), .A2(n78), .ZN(OUT1[11]) );
  AOI22_X1 U93 ( .A1(n137), .A2(IN1[10]), .B1(n2), .B2(IN0[10]), .ZN(n77) );
  AOI22_X1 U92 ( .A1(n1), .A2(IN3[10]), .B1(n72), .B2(IN2[10]), .ZN(n76) );
  NAND2_X1 U91 ( .A1(n77), .A2(n76), .ZN(OUT1[10]) );
  AOI22_X1 U3 ( .A1(n137), .A2(IN1[9]), .B1(n2), .B2(IN0[9]), .ZN(n141) );
  AOI22_X1 U2 ( .A1(n1), .A2(IN3[9]), .B1(n138), .B2(IN2[9]), .ZN(n140) );
  NAND2_X1 U1 ( .A1(n141), .A2(n140), .ZN(OUT1[9]) );
  AOI22_X1 U6 ( .A1(n137), .A2(IN1[8]), .B1(n2), .B2(IN0[8]), .ZN(n135) );
  AOI22_X1 U5 ( .A1(n1), .A2(IN3[8]), .B1(n72), .B2(IN2[8]), .ZN(n134) );
  NAND2_X1 U4 ( .A1(n135), .A2(n134), .ZN(OUT1[8]) );
  AOI22_X1 U9 ( .A1(n137), .A2(IN1[7]), .B1(n2), .B2(IN0[7]), .ZN(n133) );
  AOI22_X1 U8 ( .A1(n1), .A2(IN3[7]), .B1(n138), .B2(IN2[7]), .ZN(n132) );
  NAND2_X1 U7 ( .A1(n133), .A2(n132), .ZN(OUT1[7]) );
  AOI22_X1 U12 ( .A1(n137), .A2(IN1[6]), .B1(n2), .B2(IN0[6]), .ZN(n131) );
  AOI22_X1 U11 ( .A1(n1), .A2(IN3[6]), .B1(n138), .B2(IN2[6]), .ZN(n130) );
  NAND2_X1 U10 ( .A1(n131), .A2(n130), .ZN(OUT1[6]) );
  AOI22_X1 U15 ( .A1(n137), .A2(IN1[5]), .B1(n2), .B2(IN0[5]), .ZN(n129) );
  AOI22_X1 U14 ( .A1(n1), .A2(IN3[5]), .B1(n138), .B2(IN2[5]), .ZN(n128) );
  NAND2_X1 U13 ( .A1(n129), .A2(n128), .ZN(OUT1[5]) );
  AOI22_X1 U18 ( .A1(n137), .A2(IN1[4]), .B1(n2), .B2(IN0[4]), .ZN(n127) );
  AOI22_X1 U17 ( .A1(n1), .A2(IN3[4]), .B1(n72), .B2(IN2[4]), .ZN(n126) );
  NAND2_X1 U16 ( .A1(n127), .A2(n126), .ZN(OUT1[4]) );
  AOI22_X1 U21 ( .A1(n137), .A2(IN1[3]), .B1(n2), .B2(IN0[3]), .ZN(n125) );
  AOI22_X1 U20 ( .A1(n1), .A2(IN3[3]), .B1(n138), .B2(IN2[3]), .ZN(n124) );
  NAND2_X1 U19 ( .A1(n125), .A2(n124), .ZN(OUT1[3]) );
  AOI22_X1 U30 ( .A1(n137), .A2(IN1[2]), .B1(n2), .B2(IN0[2]), .ZN(n119) );
  AOI22_X1 U29 ( .A1(n1), .A2(IN3[2]), .B1(n138), .B2(IN2[2]), .ZN(n118) );
  NAND2_X1 U28 ( .A1(n119), .A2(n118), .ZN(OUT1[2]) );
  AOI22_X1 U60 ( .A1(n137), .A2(IN1[20]), .B1(n2), .B2(IN0[20]), .ZN(n99) );
  AOI22_X1 U59 ( .A1(n1), .A2(IN3[20]), .B1(n72), .B2(IN2[20]), .ZN(n98) );
  NAND2_X1 U58 ( .A1(n99), .A2(n98), .ZN(OUT1[20]) );
  AOI22_X1 U57 ( .A1(n137), .A2(IN1[21]), .B1(n2), .B2(IN0[21]), .ZN(n101) );
  AOI22_X1 U56 ( .A1(n1), .A2(IN3[21]), .B1(n72), .B2(IN2[21]), .ZN(n100) );
  NAND2_X1 U55 ( .A1(n101), .A2(n100), .ZN(OUT1[21]) );
  AOI22_X1 U54 ( .A1(n137), .A2(IN1[22]), .B1(n2), .B2(IN0[22]), .ZN(n103) );
  AOI22_X1 U53 ( .A1(n1), .A2(IN3[22]), .B1(n72), .B2(IN2[22]), .ZN(n102) );
  NAND2_X1 U52 ( .A1(n103), .A2(n102), .ZN(OUT1[22]) );
  AOI22_X1 U51 ( .A1(n137), .A2(IN1[23]), .B1(n2), .B2(IN0[23]), .ZN(n105) );
  AOI22_X1 U50 ( .A1(n1), .A2(IN3[23]), .B1(n72), .B2(IN2[23]), .ZN(n104) );
  NAND2_X1 U49 ( .A1(n105), .A2(n104), .ZN(OUT1[23]) );
  AOI22_X1 U36 ( .A1(n137), .A2(IN1[28]), .B1(n2), .B2(IN0[28]), .ZN(n115) );
  AOI22_X1 U35 ( .A1(n139), .A2(IN3[28]), .B1(n72), .B2(IN2[28]), .ZN(n114) );
  NAND2_X1 U34 ( .A1(n115), .A2(n114), .ZN(OUT1[28]) );
  AOI22_X1 U33 ( .A1(n137), .A2(IN1[29]), .B1(n2), .B2(IN0[29]), .ZN(n117) );
  AOI22_X1 U32 ( .A1(n139), .A2(IN3[29]), .B1(n72), .B2(IN2[29]), .ZN(n116) );
  NAND2_X1 U31 ( .A1(n117), .A2(n116), .ZN(OUT1[29]) );
  AOI22_X1 U27 ( .A1(n137), .A2(IN1[30]), .B1(n2), .B2(IN0[30]), .ZN(n121) );
  AOI22_X1 U26 ( .A1(n139), .A2(IN3[30]), .B1(n138), .B2(IN2[30]), .ZN(n120)
         );
  NAND2_X1 U25 ( .A1(n121), .A2(n120), .ZN(OUT1[30]) );
  AOI22_X1 U24 ( .A1(n137), .A2(IN1[31]), .B1(n2), .B2(IN0[31]), .ZN(n123) );
  AOI22_X1 U23 ( .A1(n1), .A2(IN3[31]), .B1(n72), .B2(IN2[31]), .ZN(n122) );
  NAND2_X1 U22 ( .A1(n123), .A2(n122), .ZN(OUT1[31]) );
  AOI22_X1 U39 ( .A1(n137), .A2(IN1[27]), .B1(n2), .B2(IN0[27]), .ZN(n113) );
  AOI22_X1 U38 ( .A1(n139), .A2(IN3[27]), .B1(n72), .B2(IN2[27]), .ZN(n112) );
  NAND2_X1 U37 ( .A1(n113), .A2(n112), .ZN(OUT1[27]) );
  AOI22_X1 U42 ( .A1(n137), .A2(IN1[26]), .B1(n2), .B2(IN0[26]), .ZN(n111) );
  AOI22_X1 U41 ( .A1(n1), .A2(IN3[26]), .B1(n72), .B2(IN2[26]), .ZN(n110) );
  NAND2_X1 U40 ( .A1(n111), .A2(n110), .ZN(OUT1[26]) );
  AOI22_X1 U45 ( .A1(n137), .A2(IN1[25]), .B1(n2), .B2(IN0[25]), .ZN(n109) );
  AOI22_X1 U44 ( .A1(n1), .A2(IN3[25]), .B1(n72), .B2(IN2[25]), .ZN(n108) );
  NAND2_X1 U43 ( .A1(n109), .A2(n108), .ZN(OUT1[25]) );
  AOI22_X1 U48 ( .A1(n137), .A2(IN1[24]), .B1(n2), .B2(IN0[24]), .ZN(n107) );
  AOI22_X1 U47 ( .A1(n139), .A2(IN3[24]), .B1(n72), .B2(IN2[24]), .ZN(n106) );
  NAND2_X1 U46 ( .A1(n107), .A2(n106), .ZN(OUT1[24]) );
  NOR2_X1 U99 ( .A1(CTRL[0]), .A2(CTRL[1]), .ZN(n136) );
  NOR2_X1 U96 ( .A1(CTRL[0]), .A2(n73), .ZN(n138) );
  INV_X1 U101 ( .A(CTRL[1]), .ZN(n73) );
  BUF_X1 U97 ( .A(n138), .Z(n72) );
  BUF_X1 U100 ( .A(n136), .Z(n2) );
  BUF_X2 U102 ( .A(n139), .Z(n1) );
  AND2_X2 U103 ( .A1(n73), .A2(CTRL[0]), .ZN(n137) );
  AND2_X1 U104 ( .A1(CTRL[0]), .A2(CTRL[1]), .ZN(n139) );
endmodule


module mux21_4 ( IN0, IN1, CTRL, OUT1 );
  input [31:0] IN0;
  input [31:0] IN1;
  output [31:0] OUT1;
  input CTRL;


  MUX2_X1 U1 ( .A(IN0[9]), .B(IN1[9]), .S(CTRL), .Z(OUT1[9]) );
  MUX2_X1 U2 ( .A(IN0[8]), .B(IN1[8]), .S(CTRL), .Z(OUT1[8]) );
  MUX2_X1 U3 ( .A(IN0[7]), .B(IN1[7]), .S(CTRL), .Z(OUT1[7]) );
  MUX2_X1 U4 ( .A(IN0[6]), .B(IN1[6]), .S(CTRL), .Z(OUT1[6]) );
  MUX2_X1 U5 ( .A(IN0[5]), .B(IN1[5]), .S(CTRL), .Z(OUT1[5]) );
  MUX2_X1 U6 ( .A(IN0[4]), .B(IN1[4]), .S(CTRL), .Z(OUT1[4]) );
  MUX2_X1 U7 ( .A(IN0[3]), .B(IN1[3]), .S(CTRL), .Z(OUT1[3]) );
  MUX2_X1 U8 ( .A(IN0[31]), .B(IN1[31]), .S(CTRL), .Z(OUT1[31]) );
  MUX2_X1 U9 ( .A(IN0[30]), .B(IN1[30]), .S(CTRL), .Z(OUT1[30]) );
  MUX2_X1 U10 ( .A(IN0[2]), .B(IN1[2]), .S(CTRL), .Z(OUT1[2]) );
  MUX2_X1 U11 ( .A(IN0[29]), .B(IN1[29]), .S(CTRL), .Z(OUT1[29]) );
  MUX2_X1 U12 ( .A(IN0[28]), .B(IN1[28]), .S(CTRL), .Z(OUT1[28]) );
  MUX2_X1 U13 ( .A(IN0[27]), .B(IN1[27]), .S(CTRL), .Z(OUT1[27]) );
  MUX2_X1 U14 ( .A(IN0[26]), .B(IN1[26]), .S(CTRL), .Z(OUT1[26]) );
  MUX2_X1 U15 ( .A(IN0[25]), .B(IN1[25]), .S(CTRL), .Z(OUT1[25]) );
  MUX2_X1 U16 ( .A(IN0[24]), .B(IN1[24]), .S(CTRL), .Z(OUT1[24]) );
  MUX2_X1 U17 ( .A(IN0[23]), .B(IN1[23]), .S(CTRL), .Z(OUT1[23]) );
  MUX2_X1 U18 ( .A(IN0[22]), .B(IN1[22]), .S(CTRL), .Z(OUT1[22]) );
  MUX2_X1 U19 ( .A(IN0[21]), .B(IN1[21]), .S(CTRL), .Z(OUT1[21]) );
  MUX2_X1 U20 ( .A(IN0[20]), .B(IN1[20]), .S(CTRL), .Z(OUT1[20]) );
  MUX2_X1 U21 ( .A(IN0[1]), .B(IN1[1]), .S(CTRL), .Z(OUT1[1]) );
  MUX2_X1 U22 ( .A(IN0[19]), .B(IN1[19]), .S(CTRL), .Z(OUT1[19]) );
  MUX2_X1 U23 ( .A(IN0[18]), .B(IN1[18]), .S(CTRL), .Z(OUT1[18]) );
  MUX2_X1 U24 ( .A(IN0[17]), .B(IN1[17]), .S(CTRL), .Z(OUT1[17]) );
  MUX2_X1 U25 ( .A(IN0[16]), .B(IN1[16]), .S(CTRL), .Z(OUT1[16]) );
  MUX2_X1 U26 ( .A(IN0[15]), .B(IN1[15]), .S(CTRL), .Z(OUT1[15]) );
  MUX2_X1 U27 ( .A(IN0[14]), .B(IN1[14]), .S(CTRL), .Z(OUT1[14]) );
  MUX2_X1 U28 ( .A(IN0[13]), .B(IN1[13]), .S(CTRL), .Z(OUT1[13]) );
  MUX2_X1 U29 ( .A(IN0[12]), .B(IN1[12]), .S(CTRL), .Z(OUT1[12]) );
  MUX2_X1 U30 ( .A(IN0[11]), .B(IN1[11]), .S(CTRL), .Z(OUT1[11]) );
  MUX2_X1 U31 ( .A(IN0[10]), .B(IN1[10]), .S(CTRL), .Z(OUT1[10]) );
  MUX2_X1 U32 ( .A(IN0[0]), .B(IN1[0]), .S(CTRL), .Z(OUT1[0]) );
endmodule


module mux21_3 ( IN0, IN1, CTRL, OUT1 );
  input [31:0] IN0;
  input [31:0] IN1;
  output [31:0] OUT1;
  input CTRL;
  wire   n1;

  MUX2_X1 U2 ( .A(IN0[8]), .B(IN1[8]), .S(n1), .Z(OUT1[8]) );
  MUX2_X1 U4 ( .A(IN0[6]), .B(IN1[6]), .S(n1), .Z(OUT1[6]) );
  MUX2_X1 U8 ( .A(IN0[31]), .B(IN1[31]), .S(CTRL), .Z(OUT1[31]) );
  MUX2_X1 U9 ( .A(IN0[30]), .B(IN1[30]), .S(CTRL), .Z(OUT1[30]) );
  MUX2_X1 U10 ( .A(IN0[2]), .B(IN1[2]), .S(CTRL), .Z(OUT1[2]) );
  MUX2_X1 U11 ( .A(IN0[29]), .B(IN1[29]), .S(n1), .Z(OUT1[29]) );
  MUX2_X1 U12 ( .A(IN0[28]), .B(IN1[28]), .S(CTRL), .Z(OUT1[28]) );
  MUX2_X1 U13 ( .A(IN0[27]), .B(IN1[27]), .S(CTRL), .Z(OUT1[27]) );
  MUX2_X1 U14 ( .A(IN0[26]), .B(IN1[26]), .S(CTRL), .Z(OUT1[26]) );
  MUX2_X1 U15 ( .A(IN0[25]), .B(IN1[25]), .S(CTRL), .Z(OUT1[25]) );
  MUX2_X1 U16 ( .A(IN0[24]), .B(IN1[24]), .S(CTRL), .Z(OUT1[24]) );
  MUX2_X1 U17 ( .A(IN0[23]), .B(IN1[23]), .S(CTRL), .Z(OUT1[23]) );
  MUX2_X1 U18 ( .A(IN0[22]), .B(IN1[22]), .S(CTRL), .Z(OUT1[22]) );
  MUX2_X1 U19 ( .A(IN0[21]), .B(IN1[21]), .S(CTRL), .Z(OUT1[21]) );
  MUX2_X1 U20 ( .A(IN0[20]), .B(IN1[20]), .S(CTRL), .Z(OUT1[20]) );
  MUX2_X1 U22 ( .A(IN0[19]), .B(IN1[19]), .S(CTRL), .Z(OUT1[19]) );
  MUX2_X1 U23 ( .A(IN0[18]), .B(IN1[18]), .S(CTRL), .Z(OUT1[18]) );
  MUX2_X1 U24 ( .A(IN0[17]), .B(IN1[17]), .S(CTRL), .Z(OUT1[17]) );
  MUX2_X1 U25 ( .A(IN0[16]), .B(IN1[16]), .S(n1), .Z(OUT1[16]) );
  MUX2_X1 U27 ( .A(IN0[14]), .B(IN1[14]), .S(n1), .Z(OUT1[14]) );
  MUX2_X1 U29 ( .A(IN0[12]), .B(IN1[12]), .S(n1), .Z(OUT1[12]) );
  MUX2_X1 U31 ( .A(IN0[10]), .B(IN1[10]), .S(n1), .Z(OUT1[10]) );
  MUX2_X1 U32 ( .A(IN0[0]), .B(IN1[0]), .S(n1), .Z(OUT1[0]) );
  MUX2_X1 U1 ( .A(IN0[9]), .B(IN1[9]), .S(CTRL), .Z(OUT1[9]) );
  MUX2_X1 U3 ( .A(IN0[7]), .B(IN1[7]), .S(CTRL), .Z(OUT1[7]) );
  MUX2_X1 U5 ( .A(IN0[5]), .B(IN1[5]), .S(CTRL), .Z(OUT1[5]) );
  MUX2_X1 U21 ( .A(IN0[1]), .B(IN1[1]), .S(CTRL), .Z(OUT1[1]) );
  MUX2_X1 U28 ( .A(IN0[13]), .B(IN1[13]), .S(n1), .Z(OUT1[13]) );
  MUX2_X1 U30 ( .A(IN0[11]), .B(IN1[11]), .S(n1), .Z(OUT1[11]) );
  MUX2_X1 U6 ( .A(IN0[4]), .B(IN1[4]), .S(n1), .Z(OUT1[4]) );
  MUX2_X1 U7 ( .A(IN0[3]), .B(IN1[3]), .S(CTRL), .Z(OUT1[3]) );
  MUX2_X1 U26 ( .A(IN0[15]), .B(IN1[15]), .S(n1), .Z(OUT1[15]) );
  BUF_X1 U33 ( .A(CTRL), .Z(n1) );
endmodule


module mux21_2 ( IN0, IN1, CTRL, OUT1 );
  input [31:0] IN0;
  input [31:0] IN1;
  output [31:0] OUT1;
  input CTRL;


  MUX2_X1 U1 ( .A(IN0[9]), .B(IN1[9]), .S(CTRL), .Z(OUT1[9]) );
  MUX2_X1 U2 ( .A(IN0[8]), .B(IN1[8]), .S(CTRL), .Z(OUT1[8]) );
  MUX2_X1 U3 ( .A(IN0[7]), .B(IN1[7]), .S(CTRL), .Z(OUT1[7]) );
  MUX2_X1 U4 ( .A(IN0[6]), .B(IN1[6]), .S(CTRL), .Z(OUT1[6]) );
  MUX2_X1 U5 ( .A(IN0[5]), .B(IN1[5]), .S(CTRL), .Z(OUT1[5]) );
  MUX2_X1 U6 ( .A(IN0[4]), .B(IN1[4]), .S(CTRL), .Z(OUT1[4]) );
  MUX2_X1 U7 ( .A(IN0[3]), .B(IN1[3]), .S(CTRL), .Z(OUT1[3]) );
  MUX2_X1 U8 ( .A(IN0[31]), .B(IN1[31]), .S(CTRL), .Z(OUT1[31]) );
  MUX2_X1 U9 ( .A(IN0[30]), .B(IN1[30]), .S(CTRL), .Z(OUT1[30]) );
  MUX2_X1 U10 ( .A(IN0[2]), .B(IN1[2]), .S(CTRL), .Z(OUT1[2]) );
  MUX2_X1 U11 ( .A(IN0[29]), .B(IN1[29]), .S(CTRL), .Z(OUT1[29]) );
  MUX2_X1 U12 ( .A(IN0[28]), .B(IN1[28]), .S(CTRL), .Z(OUT1[28]) );
  MUX2_X1 U13 ( .A(IN0[27]), .B(IN1[27]), .S(CTRL), .Z(OUT1[27]) );
  MUX2_X1 U14 ( .A(IN0[26]), .B(IN1[26]), .S(CTRL), .Z(OUT1[26]) );
  MUX2_X1 U15 ( .A(IN0[25]), .B(IN1[25]), .S(CTRL), .Z(OUT1[25]) );
  MUX2_X1 U16 ( .A(IN0[24]), .B(IN1[24]), .S(CTRL), .Z(OUT1[24]) );
  MUX2_X1 U17 ( .A(IN0[23]), .B(IN1[23]), .S(CTRL), .Z(OUT1[23]) );
  MUX2_X1 U18 ( .A(IN0[22]), .B(IN1[22]), .S(CTRL), .Z(OUT1[22]) );
  MUX2_X1 U19 ( .A(IN0[21]), .B(IN1[21]), .S(CTRL), .Z(OUT1[21]) );
  MUX2_X1 U20 ( .A(IN0[20]), .B(IN1[20]), .S(CTRL), .Z(OUT1[20]) );
  MUX2_X1 U21 ( .A(IN0[1]), .B(IN1[1]), .S(CTRL), .Z(OUT1[1]) );
  MUX2_X1 U22 ( .A(IN0[19]), .B(IN1[19]), .S(CTRL), .Z(OUT1[19]) );
  MUX2_X1 U23 ( .A(IN0[18]), .B(IN1[18]), .S(CTRL), .Z(OUT1[18]) );
  MUX2_X1 U24 ( .A(IN0[17]), .B(IN1[17]), .S(CTRL), .Z(OUT1[17]) );
  MUX2_X1 U25 ( .A(IN0[16]), .B(IN1[16]), .S(CTRL), .Z(OUT1[16]) );
  MUX2_X1 U26 ( .A(IN0[15]), .B(IN1[15]), .S(CTRL), .Z(OUT1[15]) );
  MUX2_X1 U27 ( .A(IN0[14]), .B(IN1[14]), .S(CTRL), .Z(OUT1[14]) );
  MUX2_X1 U28 ( .A(IN0[13]), .B(IN1[13]), .S(CTRL), .Z(OUT1[13]) );
  MUX2_X1 U29 ( .A(IN0[12]), .B(IN1[12]), .S(CTRL), .Z(OUT1[12]) );
  MUX2_X1 U30 ( .A(IN0[11]), .B(IN1[11]), .S(CTRL), .Z(OUT1[11]) );
  MUX2_X1 U31 ( .A(IN0[10]), .B(IN1[10]), .S(CTRL), .Z(OUT1[10]) );
  MUX2_X1 U32 ( .A(IN0[0]), .B(IN1[0]), .S(CTRL), .Z(OUT1[0]) );
endmodule


module mux21_1 ( IN0, IN1, CTRL, OUT1 );
  input [31:0] IN0;
  input [31:0] IN1;
  output [31:0] OUT1;
  input CTRL;
  wire   n1, n2;

  MUX2_X1 U1 ( .A(IN0[9]), .B(IN1[9]), .S(n1), .Z(OUT1[9]) );
  MUX2_X1 U2 ( .A(IN0[8]), .B(IN1[8]), .S(n1), .Z(OUT1[8]) );
  MUX2_X1 U3 ( .A(IN0[7]), .B(IN1[7]), .S(n1), .Z(OUT1[7]) );
  MUX2_X1 U4 ( .A(IN0[6]), .B(IN1[6]), .S(n1), .Z(OUT1[6]) );
  MUX2_X1 U5 ( .A(IN0[5]), .B(IN1[5]), .S(n1), .Z(OUT1[5]) );
  MUX2_X1 U6 ( .A(IN0[4]), .B(IN1[4]), .S(n1), .Z(OUT1[4]) );
  MUX2_X1 U7 ( .A(IN0[3]), .B(IN1[3]), .S(n1), .Z(OUT1[3]) );
  MUX2_X1 U8 ( .A(IN0[31]), .B(IN1[31]), .S(n1), .Z(OUT1[31]) );
  MUX2_X1 U9 ( .A(IN0[30]), .B(IN1[30]), .S(n1), .Z(OUT1[30]) );
  MUX2_X1 U10 ( .A(IN0[2]), .B(IN1[2]), .S(n1), .Z(OUT1[2]) );
  MUX2_X1 U11 ( .A(IN0[29]), .B(IN1[29]), .S(n1), .Z(OUT1[29]) );
  MUX2_X1 U12 ( .A(IN0[28]), .B(IN1[28]), .S(n1), .Z(OUT1[28]) );
  MUX2_X1 U13 ( .A(IN0[27]), .B(IN1[27]), .S(n1), .Z(OUT1[27]) );
  MUX2_X1 U14 ( .A(IN0[26]), .B(IN1[26]), .S(n1), .Z(OUT1[26]) );
  MUX2_X1 U15 ( .A(IN0[25]), .B(IN1[25]), .S(n1), .Z(OUT1[25]) );
  MUX2_X1 U16 ( .A(IN0[24]), .B(IN1[24]), .S(n1), .Z(OUT1[24]) );
  MUX2_X1 U17 ( .A(IN0[23]), .B(IN1[23]), .S(CTRL), .Z(OUT1[23]) );
  MUX2_X1 U18 ( .A(IN0[22]), .B(IN1[22]), .S(CTRL), .Z(OUT1[22]) );
  MUX2_X1 U19 ( .A(IN0[21]), .B(IN1[21]), .S(n1), .Z(OUT1[21]) );
  MUX2_X1 U20 ( .A(IN0[20]), .B(IN1[20]), .S(CTRL), .Z(OUT1[20]) );
  MUX2_X1 U21 ( .A(IN0[1]), .B(IN1[1]), .S(n1), .Z(OUT1[1]) );
  MUX2_X1 U22 ( .A(IN0[19]), .B(IN1[19]), .S(CTRL), .Z(OUT1[19]) );
  MUX2_X1 U23 ( .A(IN0[18]), .B(IN1[18]), .S(CTRL), .Z(OUT1[18]) );
  MUX2_X1 U24 ( .A(IN0[17]), .B(IN1[17]), .S(CTRL), .Z(OUT1[17]) );
  MUX2_X1 U25 ( .A(IN0[16]), .B(IN1[16]), .S(CTRL), .Z(OUT1[16]) );
  MUX2_X1 U26 ( .A(IN0[15]), .B(IN1[15]), .S(CTRL), .Z(OUT1[15]) );
  MUX2_X1 U27 ( .A(IN0[14]), .B(IN1[14]), .S(CTRL), .Z(OUT1[14]) );
  MUX2_X1 U28 ( .A(IN0[13]), .B(IN1[13]), .S(n1), .Z(OUT1[13]) );
  MUX2_X1 U29 ( .A(IN0[12]), .B(IN1[12]), .S(CTRL), .Z(OUT1[12]) );
  MUX2_X1 U30 ( .A(IN0[11]), .B(IN1[11]), .S(CTRL), .Z(OUT1[11]) );
  MUX2_X1 U31 ( .A(IN0[10]), .B(IN1[10]), .S(CTRL), .Z(OUT1[10]) );
  BUF_X1 U32 ( .A(CTRL), .Z(n1) );
  INV_X1 U33 ( .A(IN0[0]), .ZN(n2) );
  NOR2_X1 U34 ( .A1(n1), .A2(n2), .ZN(OUT1[0]) );
endmodule


module p4add_N32_logN5_1 ( A, B, Cin, sign, S, Cout );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input Cin, sign;
  output Cout;

  wire   [31:0] new_B;
  wire   [7:0] carry_pro;
  assign carry_pro[0] = sign;

  xor_gen_N32_1 xor32 ( .A(B), .B(carry_pro[0]), .S(new_B) );
  carry_tree_N32_logN5_1 ct ( .A(A), .B(new_B), .Cin(carry_pro[0]), .Cout({
        Cout, carry_pro[7:1]}) );
  sum_gen_N32_1 add ( .A(A), .B(new_B), .Cin({1'b0, carry_pro}), .S(S) );
endmodule


module predictor_2_15 ( clock, reset, enable, taken_i, prediction_o );
  input clock, reset, enable, taken_i;
  output prediction_o;
  wire   N11, N12, n1, n2, n5, n7, n8, n9, n10;
  wire   [1:0] next_STATE;

  DLH_X1 \next_STATE_reg[0]  ( .G(enable), .D(N11), .Q(next_STATE[0]) );
  DFFR_X1 \STATE_reg[0]  ( .D(n7), .CK(clock), .RN(n2), .Q(n1), .QN(n5) );
  DLH_X1 \next_STATE_reg[1]  ( .G(enable), .D(N12), .Q(next_STATE[1]) );
  DFFR_X1 \STATE_reg[1]  ( .D(n8), .CK(clock), .RN(n2), .Q(prediction_o) );
  MUX2_X1 U2 ( .A(prediction_o), .B(next_STATE[1]), .S(enable), .Z(n8) );
  MUX2_X1 U4 ( .A(n1), .B(next_STATE[0]), .S(enable), .Z(n7) );
  NOR2_X1 U9 ( .A1(prediction_o), .A2(taken_i), .ZN(n10) );
  NAND2_X1 U7 ( .A1(prediction_o), .A2(taken_i), .ZN(n9) );
  OAI21_X1 U6 ( .B1(n10), .B2(n1), .A(n9), .ZN(N11) );
  OAI21_X1 U5 ( .B1(n5), .B2(n10), .A(n9), .ZN(N12) );
  INV_X1 U3 ( .A(reset), .ZN(n2) );
endmodule


module predictor_2_14 ( clock, reset, enable, taken_i, prediction_o );
  input clock, reset, enable, taken_i;
  output prediction_o;
  wire   N11, N12, n1, n2, n5, n7, n8, n9, n10;
  wire   [1:0] next_STATE;

  DLH_X1 \next_STATE_reg[0]  ( .G(enable), .D(N11), .Q(next_STATE[0]) );
  DFFR_X1 \STATE_reg[0]  ( .D(n7), .CK(clock), .RN(n2), .Q(n1), .QN(n5) );
  DLH_X1 \next_STATE_reg[1]  ( .G(enable), .D(N12), .Q(next_STATE[1]) );
  DFFR_X1 \STATE_reg[1]  ( .D(n8), .CK(clock), .RN(n2), .Q(prediction_o) );
  MUX2_X1 U2 ( .A(prediction_o), .B(next_STATE[1]), .S(enable), .Z(n8) );
  MUX2_X1 U4 ( .A(n1), .B(next_STATE[0]), .S(enable), .Z(n7) );
  NOR2_X1 U9 ( .A1(prediction_o), .A2(taken_i), .ZN(n10) );
  NAND2_X1 U7 ( .A1(prediction_o), .A2(taken_i), .ZN(n9) );
  OAI21_X1 U6 ( .B1(n10), .B2(n1), .A(n9), .ZN(N11) );
  OAI21_X1 U5 ( .B1(n5), .B2(n10), .A(n9), .ZN(N12) );
  INV_X1 U3 ( .A(reset), .ZN(n2) );
endmodule


module predictor_2_13 ( clock, reset, enable, taken_i, prediction_o );
  input clock, reset, enable, taken_i;
  output prediction_o;
  wire   N11, N12, n1, n2, n5, n7, n8, n9, n10;
  wire   [1:0] next_STATE;

  DLH_X1 \next_STATE_reg[0]  ( .G(enable), .D(N11), .Q(next_STATE[0]) );
  DFFR_X1 \STATE_reg[0]  ( .D(n7), .CK(clock), .RN(n2), .Q(n1), .QN(n5) );
  DLH_X1 \next_STATE_reg[1]  ( .G(enable), .D(N12), .Q(next_STATE[1]) );
  DFFR_X1 \STATE_reg[1]  ( .D(n8), .CK(clock), .RN(n2), .Q(prediction_o) );
  MUX2_X1 U2 ( .A(prediction_o), .B(next_STATE[1]), .S(enable), .Z(n8) );
  MUX2_X1 U4 ( .A(n1), .B(next_STATE[0]), .S(enable), .Z(n7) );
  NOR2_X1 U9 ( .A1(prediction_o), .A2(taken_i), .ZN(n10) );
  NAND2_X1 U7 ( .A1(prediction_o), .A2(taken_i), .ZN(n9) );
  OAI21_X1 U6 ( .B1(n10), .B2(n1), .A(n9), .ZN(N11) );
  OAI21_X1 U5 ( .B1(n5), .B2(n10), .A(n9), .ZN(N12) );
  INV_X1 U3 ( .A(reset), .ZN(n2) );
endmodule


module predictor_2_12 ( clock, reset, enable, taken_i, prediction_o );
  input clock, reset, enable, taken_i;
  output prediction_o;
  wire   N11, N12, n1, n2, n5, n7, n8, n9, n10;
  wire   [1:0] next_STATE;

  DLH_X1 \next_STATE_reg[0]  ( .G(enable), .D(N11), .Q(next_STATE[0]) );
  DFFR_X1 \STATE_reg[0]  ( .D(n7), .CK(clock), .RN(n2), .Q(n1), .QN(n5) );
  DLH_X1 \next_STATE_reg[1]  ( .G(enable), .D(N12), .Q(next_STATE[1]) );
  DFFR_X1 \STATE_reg[1]  ( .D(n8), .CK(clock), .RN(n2), .Q(prediction_o) );
  MUX2_X1 U2 ( .A(prediction_o), .B(next_STATE[1]), .S(enable), .Z(n8) );
  MUX2_X1 U4 ( .A(n1), .B(next_STATE[0]), .S(enable), .Z(n7) );
  NOR2_X1 U9 ( .A1(prediction_o), .A2(taken_i), .ZN(n10) );
  NAND2_X1 U7 ( .A1(prediction_o), .A2(taken_i), .ZN(n9) );
  OAI21_X1 U6 ( .B1(n10), .B2(n1), .A(n9), .ZN(N11) );
  OAI21_X1 U5 ( .B1(n5), .B2(n10), .A(n9), .ZN(N12) );
  INV_X1 U3 ( .A(reset), .ZN(n2) );
endmodule


module predictor_2_11 ( clock, reset, enable, taken_i, prediction_o );
  input clock, reset, enable, taken_i;
  output prediction_o;
  wire   N11, N12, n1, n2, n5, n7, n8, n9, n10;
  wire   [1:0] next_STATE;

  DLH_X1 \next_STATE_reg[0]  ( .G(enable), .D(N11), .Q(next_STATE[0]) );
  DFFR_X1 \STATE_reg[0]  ( .D(n7), .CK(clock), .RN(n2), .Q(n1), .QN(n5) );
  DLH_X1 \next_STATE_reg[1]  ( .G(enable), .D(N12), .Q(next_STATE[1]) );
  DFFR_X1 \STATE_reg[1]  ( .D(n8), .CK(clock), .RN(n2), .Q(prediction_o) );
  MUX2_X1 U2 ( .A(prediction_o), .B(next_STATE[1]), .S(enable), .Z(n8) );
  MUX2_X1 U4 ( .A(n1), .B(next_STATE[0]), .S(enable), .Z(n7) );
  NOR2_X1 U9 ( .A1(prediction_o), .A2(taken_i), .ZN(n10) );
  NAND2_X1 U7 ( .A1(prediction_o), .A2(taken_i), .ZN(n9) );
  OAI21_X1 U6 ( .B1(n10), .B2(n1), .A(n9), .ZN(N11) );
  OAI21_X1 U5 ( .B1(n5), .B2(n10), .A(n9), .ZN(N12) );
  INV_X1 U3 ( .A(reset), .ZN(n2) );
endmodule


module predictor_2_10 ( clock, reset, enable, taken_i, prediction_o );
  input clock, reset, enable, taken_i;
  output prediction_o;
  wire   N11, N12, n1, n2, n5, n7, n8, n9, n10;
  wire   [1:0] next_STATE;

  DLH_X1 \next_STATE_reg[0]  ( .G(enable), .D(N11), .Q(next_STATE[0]) );
  DFFR_X1 \STATE_reg[0]  ( .D(n7), .CK(clock), .RN(n2), .Q(n1), .QN(n5) );
  DLH_X1 \next_STATE_reg[1]  ( .G(enable), .D(N12), .Q(next_STATE[1]) );
  DFFR_X1 \STATE_reg[1]  ( .D(n8), .CK(clock), .RN(n2), .Q(prediction_o) );
  MUX2_X1 U2 ( .A(prediction_o), .B(next_STATE[1]), .S(enable), .Z(n8) );
  MUX2_X1 U4 ( .A(n1), .B(next_STATE[0]), .S(enable), .Z(n7) );
  NOR2_X1 U9 ( .A1(prediction_o), .A2(taken_i), .ZN(n10) );
  NAND2_X1 U7 ( .A1(prediction_o), .A2(taken_i), .ZN(n9) );
  OAI21_X1 U6 ( .B1(n10), .B2(n1), .A(n9), .ZN(N11) );
  OAI21_X1 U5 ( .B1(n5), .B2(n10), .A(n9), .ZN(N12) );
  INV_X1 U3 ( .A(reset), .ZN(n2) );
endmodule


module predictor_2_9 ( clock, reset, enable, taken_i, prediction_o );
  input clock, reset, enable, taken_i;
  output prediction_o;
  wire   N11, N12, n1, n2, n5, n7, n8, n9, n10;
  wire   [1:0] next_STATE;

  DLH_X1 \next_STATE_reg[0]  ( .G(enable), .D(N11), .Q(next_STATE[0]) );
  DFFR_X1 \STATE_reg[0]  ( .D(n7), .CK(clock), .RN(n2), .Q(n1), .QN(n5) );
  DLH_X1 \next_STATE_reg[1]  ( .G(enable), .D(N12), .Q(next_STATE[1]) );
  DFFR_X1 \STATE_reg[1]  ( .D(n8), .CK(clock), .RN(n2), .Q(prediction_o) );
  MUX2_X1 U2 ( .A(prediction_o), .B(next_STATE[1]), .S(enable), .Z(n8) );
  MUX2_X1 U4 ( .A(n1), .B(next_STATE[0]), .S(enable), .Z(n7) );
  NOR2_X1 U9 ( .A1(prediction_o), .A2(taken_i), .ZN(n10) );
  NAND2_X1 U7 ( .A1(prediction_o), .A2(taken_i), .ZN(n9) );
  OAI21_X1 U6 ( .B1(n10), .B2(n1), .A(n9), .ZN(N11) );
  OAI21_X1 U5 ( .B1(n5), .B2(n10), .A(n9), .ZN(N12) );
  INV_X1 U3 ( .A(reset), .ZN(n2) );
endmodule


module predictor_2_8 ( clock, reset, enable, taken_i, prediction_o );
  input clock, reset, enable, taken_i;
  output prediction_o;
  wire   N11, N12, n1, n2, n5, n7, n8, n9, n10;
  wire   [1:0] next_STATE;

  DLH_X1 \next_STATE_reg[0]  ( .G(enable), .D(N11), .Q(next_STATE[0]) );
  DFFR_X1 \STATE_reg[0]  ( .D(n7), .CK(clock), .RN(n2), .Q(n1), .QN(n5) );
  DLH_X1 \next_STATE_reg[1]  ( .G(enable), .D(N12), .Q(next_STATE[1]) );
  DFFR_X1 \STATE_reg[1]  ( .D(n8), .CK(clock), .RN(n2), .Q(prediction_o) );
  MUX2_X1 U2 ( .A(prediction_o), .B(next_STATE[1]), .S(enable), .Z(n8) );
  MUX2_X1 U4 ( .A(n1), .B(next_STATE[0]), .S(enable), .Z(n7) );
  NOR2_X1 U9 ( .A1(prediction_o), .A2(taken_i), .ZN(n10) );
  NAND2_X1 U7 ( .A1(prediction_o), .A2(taken_i), .ZN(n9) );
  OAI21_X1 U6 ( .B1(n10), .B2(n1), .A(n9), .ZN(N11) );
  OAI21_X1 U5 ( .B1(n5), .B2(n10), .A(n9), .ZN(N12) );
  INV_X1 U3 ( .A(reset), .ZN(n2) );
endmodule


module predictor_2_7 ( clock, reset, enable, taken_i, prediction_o );
  input clock, reset, enable, taken_i;
  output prediction_o;
  wire   N11, N12, n1, n2, n5, n7, n8, n9, n10;
  wire   [1:0] next_STATE;

  DLH_X1 \next_STATE_reg[0]  ( .G(enable), .D(N11), .Q(next_STATE[0]) );
  DFFR_X1 \STATE_reg[0]  ( .D(n7), .CK(clock), .RN(n2), .Q(n1), .QN(n5) );
  DLH_X1 \next_STATE_reg[1]  ( .G(enable), .D(N12), .Q(next_STATE[1]) );
  DFFR_X1 \STATE_reg[1]  ( .D(n8), .CK(clock), .RN(n2), .Q(prediction_o) );
  MUX2_X1 U2 ( .A(prediction_o), .B(next_STATE[1]), .S(enable), .Z(n8) );
  MUX2_X1 U4 ( .A(n1), .B(next_STATE[0]), .S(enable), .Z(n7) );
  NOR2_X1 U9 ( .A1(prediction_o), .A2(taken_i), .ZN(n10) );
  NAND2_X1 U7 ( .A1(prediction_o), .A2(taken_i), .ZN(n9) );
  OAI21_X1 U6 ( .B1(n10), .B2(n1), .A(n9), .ZN(N11) );
  OAI21_X1 U5 ( .B1(n5), .B2(n10), .A(n9), .ZN(N12) );
  INV_X1 U3 ( .A(reset), .ZN(n2) );
endmodule


module predictor_2_6 ( clock, reset, enable, taken_i, prediction_o );
  input clock, reset, enable, taken_i;
  output prediction_o;
  wire   N11, N12, n1, n2, n5, n7, n8, n9, n10;
  wire   [1:0] next_STATE;

  DLH_X1 \next_STATE_reg[0]  ( .G(enable), .D(N11), .Q(next_STATE[0]) );
  DFFR_X1 \STATE_reg[0]  ( .D(n7), .CK(clock), .RN(n2), .Q(n1), .QN(n5) );
  DLH_X1 \next_STATE_reg[1]  ( .G(enable), .D(N12), .Q(next_STATE[1]) );
  DFFR_X1 \STATE_reg[1]  ( .D(n8), .CK(clock), .RN(n2), .Q(prediction_o) );
  MUX2_X1 U2 ( .A(prediction_o), .B(next_STATE[1]), .S(enable), .Z(n8) );
  MUX2_X1 U4 ( .A(n1), .B(next_STATE[0]), .S(enable), .Z(n7) );
  NOR2_X1 U9 ( .A1(prediction_o), .A2(taken_i), .ZN(n10) );
  NAND2_X1 U7 ( .A1(prediction_o), .A2(taken_i), .ZN(n9) );
  OAI21_X1 U5 ( .B1(n5), .B2(n10), .A(n9), .ZN(N12) );
  OAI21_X1 U6 ( .B1(n10), .B2(n1), .A(n9), .ZN(N11) );
  INV_X1 U3 ( .A(reset), .ZN(n2) );
endmodule


module predictor_2_5 ( clock, reset, enable, taken_i, prediction_o );
  input clock, reset, enable, taken_i;
  output prediction_o;
  wire   N11, N12, n1, n2, n5, n7, n8, n9, n10;
  wire   [1:0] next_STATE;

  DLH_X1 \next_STATE_reg[0]  ( .G(enable), .D(N11), .Q(next_STATE[0]) );
  DFFR_X1 \STATE_reg[0]  ( .D(n7), .CK(clock), .RN(n2), .Q(n1), .QN(n5) );
  DLH_X1 \next_STATE_reg[1]  ( .G(enable), .D(N12), .Q(next_STATE[1]) );
  DFFR_X1 \STATE_reg[1]  ( .D(n8), .CK(clock), .RN(n2), .Q(prediction_o) );
  MUX2_X1 U2 ( .A(prediction_o), .B(next_STATE[1]), .S(enable), .Z(n8) );
  MUX2_X1 U4 ( .A(n1), .B(next_STATE[0]), .S(enable), .Z(n7) );
  NOR2_X1 U9 ( .A1(prediction_o), .A2(taken_i), .ZN(n10) );
  NAND2_X1 U7 ( .A1(prediction_o), .A2(taken_i), .ZN(n9) );
  OAI21_X1 U5 ( .B1(n5), .B2(n10), .A(n9), .ZN(N12) );
  OAI21_X1 U6 ( .B1(n10), .B2(n1), .A(n9), .ZN(N11) );
  INV_X1 U3 ( .A(reset), .ZN(n2) );
endmodule


module predictor_2_4 ( clock, reset, enable, taken_i, prediction_o );
  input clock, reset, enable, taken_i;
  output prediction_o;
  wire   N11, N12, n1, n2, n5, n7, n8, n9, n10;
  wire   [1:0] next_STATE;

  DLH_X1 \next_STATE_reg[0]  ( .G(enable), .D(N11), .Q(next_STATE[0]) );
  DFFR_X1 \STATE_reg[0]  ( .D(n7), .CK(clock), .RN(n2), .Q(n1), .QN(n5) );
  DLH_X1 \next_STATE_reg[1]  ( .G(enable), .D(N12), .Q(next_STATE[1]) );
  DFFR_X1 \STATE_reg[1]  ( .D(n8), .CK(clock), .RN(n2), .Q(prediction_o) );
  MUX2_X1 U2 ( .A(prediction_o), .B(next_STATE[1]), .S(enable), .Z(n8) );
  MUX2_X1 U4 ( .A(n1), .B(next_STATE[0]), .S(enable), .Z(n7) );
  NOR2_X1 U9 ( .A1(prediction_o), .A2(taken_i), .ZN(n10) );
  NAND2_X1 U7 ( .A1(prediction_o), .A2(taken_i), .ZN(n9) );
  OAI21_X1 U6 ( .B1(n10), .B2(n1), .A(n9), .ZN(N11) );
  OAI21_X1 U5 ( .B1(n5), .B2(n10), .A(n9), .ZN(N12) );
  INV_X1 U3 ( .A(reset), .ZN(n2) );
endmodule


module predictor_2_3 ( clock, reset, enable, taken_i, prediction_o );
  input clock, reset, enable, taken_i;
  output prediction_o;
  wire   N11, N12, n1, n2, n5, n7, n8, n9, n10;
  wire   [1:0] next_STATE;

  DLH_X1 \next_STATE_reg[0]  ( .G(enable), .D(N11), .Q(next_STATE[0]) );
  DFFR_X1 \STATE_reg[0]  ( .D(n7), .CK(clock), .RN(n2), .Q(n1), .QN(n5) );
  DLH_X1 \next_STATE_reg[1]  ( .G(enable), .D(N12), .Q(next_STATE[1]) );
  DFFR_X1 \STATE_reg[1]  ( .D(n8), .CK(clock), .RN(n2), .Q(prediction_o) );
  MUX2_X1 U2 ( .A(prediction_o), .B(next_STATE[1]), .S(enable), .Z(n8) );
  MUX2_X1 U4 ( .A(n1), .B(next_STATE[0]), .S(enable), .Z(n7) );
  NOR2_X1 U9 ( .A1(prediction_o), .A2(taken_i), .ZN(n10) );
  NAND2_X1 U7 ( .A1(prediction_o), .A2(taken_i), .ZN(n9) );
  OAI21_X1 U5 ( .B1(n5), .B2(n10), .A(n9), .ZN(N12) );
  OAI21_X1 U6 ( .B1(n10), .B2(n1), .A(n9), .ZN(N11) );
  INV_X1 U3 ( .A(reset), .ZN(n2) );
endmodule


module predictor_2_2 ( clock, reset, enable, taken_i, prediction_o );
  input clock, reset, enable, taken_i;
  output prediction_o;
  wire   N11, N12, n1, n2, n5, n7, n8, n9, n10;
  wire   [1:0] next_STATE;

  DLH_X1 \next_STATE_reg[0]  ( .G(enable), .D(N11), .Q(next_STATE[0]) );
  DFFR_X1 \STATE_reg[0]  ( .D(n7), .CK(clock), .RN(n2), .Q(n1), .QN(n5) );
  DLH_X1 \next_STATE_reg[1]  ( .G(enable), .D(N12), .Q(next_STATE[1]) );
  DFFR_X1 \STATE_reg[1]  ( .D(n8), .CK(clock), .RN(n2), .Q(prediction_o) );
  MUX2_X1 U2 ( .A(prediction_o), .B(next_STATE[1]), .S(enable), .Z(n8) );
  MUX2_X1 U4 ( .A(n1), .B(next_STATE[0]), .S(enable), .Z(n7) );
  NOR2_X1 U9 ( .A1(prediction_o), .A2(taken_i), .ZN(n10) );
  NAND2_X1 U7 ( .A1(prediction_o), .A2(taken_i), .ZN(n9) );
  OAI21_X1 U6 ( .B1(n10), .B2(n1), .A(n9), .ZN(N11) );
  OAI21_X1 U5 ( .B1(n5), .B2(n10), .A(n9), .ZN(N12) );
  INV_X1 U3 ( .A(reset), .ZN(n2) );
endmodule


module predictor_2_1 ( clock, reset, enable, taken_i, prediction_o );
  input clock, reset, enable, taken_i;
  output prediction_o;
  wire   N11, N12, n1, n2, n5, n7, n8, n9, n10;
  wire   [1:0] next_STATE;

  DLH_X1 \next_STATE_reg[0]  ( .G(enable), .D(N11), .Q(next_STATE[0]) );
  DFFR_X1 \STATE_reg[0]  ( .D(n7), .CK(clock), .RN(n2), .Q(n1), .QN(n5) );
  DLH_X1 \next_STATE_reg[1]  ( .G(enable), .D(N12), .Q(next_STATE[1]) );
  DFFR_X1 \STATE_reg[1]  ( .D(n8), .CK(clock), .RN(n2), .Q(prediction_o) );
  MUX2_X1 U2 ( .A(prediction_o), .B(next_STATE[1]), .S(enable), .Z(n8) );
  MUX2_X1 U4 ( .A(n1), .B(next_STATE[0]), .S(enable), .Z(n7) );
  NOR2_X1 U9 ( .A1(prediction_o), .A2(taken_i), .ZN(n10) );
  NAND2_X1 U7 ( .A1(prediction_o), .A2(taken_i), .ZN(n9) );
  OAI21_X1 U5 ( .B1(n5), .B2(n10), .A(n9), .ZN(N12) );
  OAI21_X1 U6 ( .B1(n10), .B2(n1), .A(n9), .ZN(N11) );
  INV_X1 U3 ( .A(reset), .ZN(n2) );
endmodule


module mux41_1 ( IN0, IN1, IN2, IN3, CTRL, OUT1 );
  input [31:0] IN0;
  input [31:0] IN1;
  input [31:0] IN2;
  input [31:0] IN3;
  input [1:0] CTRL;
  output [31:0] OUT1;
  wire   n1, n2, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141;

  AOI22_X1 U45 ( .A1(n2), .A2(IN1[25]), .B1(n72), .B2(IN0[25]), .ZN(n109) );
  AOI22_X1 U44 ( .A1(n139), .A2(IN3[25]), .B1(n1), .B2(IN2[25]), .ZN(n108) );
  NAND2_X1 U43 ( .A1(n109), .A2(n108), .ZN(OUT1[25]) );
  AOI22_X1 U87 ( .A1(n2), .A2(IN1[12]), .B1(n72), .B2(IN0[12]), .ZN(n81) );
  AOI22_X1 U86 ( .A1(n139), .A2(IN3[12]), .B1(n1), .B2(IN2[12]), .ZN(n80) );
  NAND2_X1 U85 ( .A1(n81), .A2(n80), .ZN(OUT1[12]) );
  AOI22_X1 U39 ( .A1(n2), .A2(IN1[27]), .B1(n72), .B2(IN0[27]), .ZN(n113) );
  AOI22_X1 U38 ( .A1(n139), .A2(IN3[27]), .B1(n1), .B2(IN2[27]), .ZN(n112) );
  NAND2_X1 U37 ( .A1(n113), .A2(n112), .ZN(OUT1[27]) );
  AOI22_X1 U93 ( .A1(n2), .A2(IN1[10]), .B1(n72), .B2(IN0[10]), .ZN(n77) );
  AOI22_X1 U92 ( .A1(n139), .A2(IN3[10]), .B1(n1), .B2(IN2[10]), .ZN(n76) );
  NAND2_X1 U91 ( .A1(n77), .A2(n76), .ZN(OUT1[10]) );
  AOI22_X1 U30 ( .A1(n2), .A2(IN1[2]), .B1(n72), .B2(IN0[2]), .ZN(n119) );
  AOI22_X1 U29 ( .A1(n139), .A2(IN3[2]), .B1(n1), .B2(IN2[2]), .ZN(n118) );
  NAND2_X1 U28 ( .A1(n119), .A2(n118), .ZN(OUT1[2]) );
  AOI22_X1 U78 ( .A1(n2), .A2(IN1[15]), .B1(n72), .B2(IN0[15]), .ZN(n87) );
  AOI22_X1 U77 ( .A1(n139), .A2(IN3[15]), .B1(n1), .B2(IN2[15]), .ZN(n86) );
  NAND2_X1 U76 ( .A1(n87), .A2(n86), .ZN(OUT1[15]) );
  AOI22_X1 U21 ( .A1(n2), .A2(IN1[3]), .B1(n72), .B2(IN0[3]), .ZN(n125) );
  AOI22_X1 U20 ( .A1(n139), .A2(IN3[3]), .B1(n138), .B2(IN2[3]), .ZN(n124) );
  NAND2_X1 U19 ( .A1(n125), .A2(n124), .ZN(OUT1[3]) );
  AOI22_X1 U51 ( .A1(n2), .A2(IN1[23]), .B1(n72), .B2(IN0[23]), .ZN(n105) );
  AOI22_X1 U50 ( .A1(n139), .A2(IN3[23]), .B1(n1), .B2(IN2[23]), .ZN(n104) );
  NAND2_X1 U49 ( .A1(n105), .A2(n104), .ZN(OUT1[23]) );
  AOI22_X1 U15 ( .A1(n2), .A2(IN1[5]), .B1(n72), .B2(IN0[5]), .ZN(n129) );
  AOI22_X1 U14 ( .A1(n139), .A2(IN3[5]), .B1(n138), .B2(IN2[5]), .ZN(n128) );
  NAND2_X1 U13 ( .A1(n129), .A2(n128), .ZN(OUT1[5]) );
  AOI22_X1 U57 ( .A1(n2), .A2(IN1[21]), .B1(n72), .B2(IN0[21]), .ZN(n101) );
  AOI22_X1 U56 ( .A1(n139), .A2(IN3[21]), .B1(n1), .B2(IN2[21]), .ZN(n100) );
  NAND2_X1 U55 ( .A1(n101), .A2(n100), .ZN(OUT1[21]) );
  AOI22_X1 U75 ( .A1(n2), .A2(IN1[16]), .B1(n72), .B2(IN0[16]), .ZN(n89) );
  AOI22_X1 U74 ( .A1(n139), .A2(IN3[16]), .B1(n1), .B2(IN2[16]), .ZN(n88) );
  NAND2_X1 U73 ( .A1(n89), .A2(n88), .ZN(OUT1[16]) );
  AOI22_X1 U66 ( .A1(n2), .A2(IN1[19]), .B1(n72), .B2(IN0[19]), .ZN(n95) );
  AOI22_X1 U65 ( .A1(n139), .A2(IN3[19]), .B1(n1), .B2(IN2[19]), .ZN(n94) );
  NAND2_X1 U64 ( .A1(n95), .A2(n94), .ZN(OUT1[19]) );
  AOI22_X1 U54 ( .A1(n2), .A2(IN1[22]), .B1(n72), .B2(IN0[22]), .ZN(n103) );
  AOI22_X1 U53 ( .A1(n139), .A2(IN3[22]), .B1(n1), .B2(IN2[22]), .ZN(n102) );
  NAND2_X1 U52 ( .A1(n103), .A2(n102), .ZN(OUT1[22]) );
  AOI22_X1 U72 ( .A1(n2), .A2(IN1[17]), .B1(n72), .B2(IN0[17]), .ZN(n91) );
  AOI22_X1 U71 ( .A1(n139), .A2(IN3[17]), .B1(n1), .B2(IN2[17]), .ZN(n90) );
  NAND2_X1 U70 ( .A1(n91), .A2(n90), .ZN(OUT1[17]) );
  AOI22_X1 U69 ( .A1(n2), .A2(IN1[18]), .B1(n72), .B2(IN0[18]), .ZN(n93) );
  AOI22_X1 U68 ( .A1(n139), .A2(IN3[18]), .B1(n1), .B2(IN2[18]), .ZN(n92) );
  NAND2_X1 U67 ( .A1(n93), .A2(n92), .ZN(OUT1[18]) );
  AOI22_X1 U90 ( .A1(n2), .A2(IN1[11]), .B1(n72), .B2(IN0[11]), .ZN(n79) );
  AOI22_X1 U89 ( .A1(n139), .A2(IN3[11]), .B1(n1), .B2(IN2[11]), .ZN(n78) );
  NAND2_X1 U88 ( .A1(n79), .A2(n78), .ZN(OUT1[11]) );
  AOI22_X1 U33 ( .A1(n2), .A2(IN1[29]), .B1(n72), .B2(IN0[29]), .ZN(n117) );
  AOI22_X1 U32 ( .A1(n139), .A2(IN3[29]), .B1(n1), .B2(IN2[29]), .ZN(n116) );
  NAND2_X1 U31 ( .A1(n117), .A2(n116), .ZN(OUT1[29]) );
  AOI22_X1 U84 ( .A1(n2), .A2(IN1[13]), .B1(n72), .B2(IN0[13]), .ZN(n83) );
  AOI22_X1 U83 ( .A1(n139), .A2(IN3[13]), .B1(n1), .B2(IN2[13]), .ZN(n82) );
  NAND2_X1 U82 ( .A1(n83), .A2(n82), .ZN(OUT1[13]) );
  AOI22_X1 U81 ( .A1(n2), .A2(IN1[14]), .B1(n72), .B2(IN0[14]), .ZN(n85) );
  AOI22_X1 U80 ( .A1(n139), .A2(IN3[14]), .B1(n1), .B2(IN2[14]), .ZN(n84) );
  NAND2_X1 U79 ( .A1(n85), .A2(n84), .ZN(OUT1[14]) );
  AOI22_X1 U60 ( .A1(n2), .A2(IN1[20]), .B1(n72), .B2(IN0[20]), .ZN(n99) );
  AOI22_X1 U59 ( .A1(n139), .A2(IN3[20]), .B1(n1), .B2(IN2[20]), .ZN(n98) );
  NAND2_X1 U58 ( .A1(n99), .A2(n98), .ZN(OUT1[20]) );
  AOI22_X1 U48 ( .A1(n2), .A2(IN1[24]), .B1(n72), .B2(IN0[24]), .ZN(n107) );
  AOI22_X1 U47 ( .A1(n139), .A2(IN3[24]), .B1(n1), .B2(IN2[24]), .ZN(n106) );
  NAND2_X1 U46 ( .A1(n107), .A2(n106), .ZN(OUT1[24]) );
  AOI22_X1 U36 ( .A1(n2), .A2(IN1[28]), .B1(n72), .B2(IN0[28]), .ZN(n115) );
  AOI22_X1 U35 ( .A1(n139), .A2(IN3[28]), .B1(n1), .B2(IN2[28]), .ZN(n114) );
  NAND2_X1 U34 ( .A1(n115), .A2(n114), .ZN(OUT1[28]) );
  AOI22_X1 U42 ( .A1(n2), .A2(IN1[26]), .B1(n72), .B2(IN0[26]), .ZN(n111) );
  AOI22_X1 U41 ( .A1(n139), .A2(IN3[26]), .B1(n1), .B2(IN2[26]), .ZN(n110) );
  NAND2_X1 U40 ( .A1(n111), .A2(n110), .ZN(OUT1[26]) );
  AOI22_X1 U98 ( .A1(n2), .A2(IN1[0]), .B1(n72), .B2(IN0[0]), .ZN(n75) );
  AOI22_X1 U95 ( .A1(n139), .A2(IN3[0]), .B1(n1), .B2(IN2[0]), .ZN(n74) );
  NAND2_X1 U94 ( .A1(n75), .A2(n74), .ZN(OUT1[0]) );
  AOI22_X1 U63 ( .A1(n2), .A2(IN1[1]), .B1(n72), .B2(IN0[1]), .ZN(n97) );
  AOI22_X1 U62 ( .A1(n139), .A2(IN3[1]), .B1(n1), .B2(IN2[1]), .ZN(n96) );
  NAND2_X1 U61 ( .A1(n97), .A2(n96), .ZN(OUT1[1]) );
  AOI22_X1 U27 ( .A1(n2), .A2(IN1[30]), .B1(n72), .B2(IN0[30]), .ZN(n121) );
  AOI22_X1 U26 ( .A1(n139), .A2(IN3[30]), .B1(n1), .B2(IN2[30]), .ZN(n120) );
  NAND2_X1 U25 ( .A1(n121), .A2(n120), .ZN(OUT1[30]) );
  AOI22_X1 U6 ( .A1(n137), .A2(IN1[8]), .B1(n136), .B2(IN0[8]), .ZN(n135) );
  AOI22_X1 U5 ( .A1(n139), .A2(IN3[8]), .B1(n138), .B2(IN2[8]), .ZN(n134) );
  NAND2_X1 U4 ( .A1(n135), .A2(n134), .ZN(OUT1[8]) );
  AOI22_X1 U24 ( .A1(n137), .A2(IN1[31]), .B1(n136), .B2(IN0[31]), .ZN(n123)
         );
  AOI22_X1 U23 ( .A1(n139), .A2(IN3[31]), .B1(n138), .B2(IN2[31]), .ZN(n122)
         );
  NAND2_X1 U22 ( .A1(n123), .A2(n122), .ZN(OUT1[31]) );
  AOI22_X1 U9 ( .A1(n137), .A2(IN1[7]), .B1(n136), .B2(IN0[7]), .ZN(n133) );
  AOI22_X1 U8 ( .A1(n139), .A2(IN3[7]), .B1(n138), .B2(IN2[7]), .ZN(n132) );
  NAND2_X1 U7 ( .A1(n133), .A2(n132), .ZN(OUT1[7]) );
  AOI22_X1 U12 ( .A1(n137), .A2(IN1[6]), .B1(n136), .B2(IN0[6]), .ZN(n131) );
  AOI22_X1 U11 ( .A1(n139), .A2(IN3[6]), .B1(n138), .B2(IN2[6]), .ZN(n130) );
  NAND2_X1 U10 ( .A1(n131), .A2(n130), .ZN(OUT1[6]) );
  AOI22_X1 U3 ( .A1(n137), .A2(IN1[9]), .B1(n136), .B2(IN0[9]), .ZN(n141) );
  AOI22_X1 U2 ( .A1(n139), .A2(IN3[9]), .B1(n138), .B2(IN2[9]), .ZN(n140) );
  NAND2_X1 U1 ( .A1(n141), .A2(n140), .ZN(OUT1[9]) );
  AOI22_X1 U18 ( .A1(n137), .A2(IN1[4]), .B1(n136), .B2(IN0[4]), .ZN(n127) );
  AOI22_X1 U17 ( .A1(n139), .A2(IN3[4]), .B1(n138), .B2(IN2[4]), .ZN(n126) );
  NAND2_X1 U16 ( .A1(n127), .A2(n126), .ZN(OUT1[4]) );
  INV_X1 U101 ( .A(CTRL[1]), .ZN(n73) );
  NOR2_X1 U96 ( .A1(CTRL[0]), .A2(n73), .ZN(n138) );
  AND2_X2 U97 ( .A1(CTRL[0]), .A2(CTRL[1]), .ZN(n139) );
  BUF_X1 U99 ( .A(n138), .Z(n1) );
  BUF_X1 U100 ( .A(n136), .Z(n72) );
  BUF_X2 U102 ( .A(n137), .Z(n2) );
  AND2_X1 U103 ( .A1(n73), .A2(CTRL[0]), .ZN(n137) );
  NOR2_X1 U104 ( .A1(CTRL[0]), .A2(CTRL[1]), .ZN(n136) );
endmodule


module ff32_en_1 ( D, en, clk, rst, Q );
  input [31:0] D;
  output [31:0] Q;
  input en, clk, rst;
  wire   net338257, n32, n34;

  DFFR_X1 \Q_reg[31]  ( .D(D[31]), .CK(net338257), .RN(n34), .Q(Q[31]) );
  DFFR_X1 \Q_reg[30]  ( .D(D[30]), .CK(net338257), .RN(n34), .Q(Q[30]) );
  DFFR_X1 \Q_reg[29]  ( .D(D[29]), .CK(net338257), .RN(n34), .Q(Q[29]) );
  DFFR_X1 \Q_reg[28]  ( .D(D[28]), .CK(net338257), .RN(n34), .Q(Q[28]) );
  DFFR_X1 \Q_reg[27]  ( .D(D[27]), .CK(net338257), .RN(n34), .Q(Q[27]) );
  DFFR_X1 \Q_reg[26]  ( .D(D[26]), .CK(net338257), .RN(n34), .Q(Q[26]) );
  DFFR_X1 \Q_reg[25]  ( .D(D[25]), .CK(net338257), .RN(n34), .Q(Q[25]) );
  DFFR_X1 \Q_reg[24]  ( .D(D[24]), .CK(net338257), .RN(n34), .Q(Q[24]) );
  DFFR_X1 \Q_reg[23]  ( .D(D[23]), .CK(net338257), .RN(n32), .Q(Q[23]) );
  DFFR_X1 \Q_reg[22]  ( .D(D[22]), .CK(net338257), .RN(n34), .Q(Q[22]) );
  DFFR_X1 \Q_reg[21]  ( .D(D[21]), .CK(net338257), .RN(n32), .Q(Q[21]) );
  DFFR_X1 \Q_reg[20]  ( .D(D[20]), .CK(net338257), .RN(n34), .Q(Q[20]) );
  DFFR_X1 \Q_reg[19]  ( .D(D[19]), .CK(net338257), .RN(n32), .Q(Q[19]) );
  DFFR_X1 \Q_reg[18]  ( .D(D[18]), .CK(net338257), .RN(n34), .Q(Q[18]) );
  DFFR_X1 \Q_reg[17]  ( .D(D[17]), .CK(net338257), .RN(n32), .Q(Q[17]) );
  DFFR_X1 \Q_reg[16]  ( .D(D[16]), .CK(net338257), .RN(n34), .Q(Q[16]) );
  DFFR_X1 \Q_reg[15]  ( .D(D[15]), .CK(net338257), .RN(n34), .Q(Q[15]) );
  DFFR_X1 \Q_reg[14]  ( .D(D[14]), .CK(net338257), .RN(n34), .Q(Q[14]) );
  DFFR_X1 \Q_reg[13]  ( .D(D[13]), .CK(net338257), .RN(n34), .Q(Q[13]) );
  DFFR_X1 \Q_reg[12]  ( .D(D[12]), .CK(net338257), .RN(n34), .Q(Q[12]) );
  DFFR_X1 \Q_reg[11]  ( .D(D[11]), .CK(net338257), .RN(n32), .Q(Q[11]) );
  DFFR_X1 \Q_reg[10]  ( .D(D[10]), .CK(net338257), .RN(n32), .Q(Q[10]) );
  DFFR_X1 \Q_reg[9]  ( .D(D[9]), .CK(net338257), .RN(n32), .Q(Q[9]) );
  DFFR_X1 \Q_reg[8]  ( .D(D[8]), .CK(net338257), .RN(n32), .Q(Q[8]) );
  DFFR_X1 \Q_reg[7]  ( .D(D[7]), .CK(net338257), .RN(n32), .Q(Q[7]) );
  DFFR_X1 \Q_reg[6]  ( .D(D[6]), .CK(net338257), .RN(n32), .Q(Q[6]) );
  DFFR_X1 \Q_reg[5]  ( .D(D[5]), .CK(net338257), .RN(n32), .Q(Q[5]) );
  DFFR_X1 \Q_reg[4]  ( .D(D[4]), .CK(net338257), .RN(n32), .Q(Q[4]) );
  DFFR_X1 \Q_reg[3]  ( .D(D[3]), .CK(net338257), .RN(n32), .Q(Q[3]) );
  DFFR_X1 \Q_reg[2]  ( .D(D[2]), .CK(net338257), .RN(n32), .Q(Q[2]) );
  DFFR_X1 \Q_reg[1]  ( .D(D[1]), .CK(net338257), .RN(n32), .Q(Q[1]) );
  DFFR_X1 \Q_reg[0]  ( .D(D[0]), .CK(net338257), .RN(n32), .Q(Q[0]) );
  SNPS_CLOCK_GATE_HIGH_ff32_en_1 clk_gate_Q_reg ( .CLK(clk), .EN(en), .ENCLK(
        net338257) );
  CLKBUF_X1 U2 ( .A(n34), .Z(n32) );
  INV_X1 U3 ( .A(rst), .ZN(n34) );
endmodule


module FA_0 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(S) );
  AND2_X1 U2 ( .A1(B), .A2(A), .ZN(Co) );
endmodule


module mux21_SIZE4_0 ( IN0, IN1, CTRL, OUT1 );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] OUT1;
  input CTRL;

  assign OUT1[3] = IN0[3];
  assign OUT1[2] = IN0[2];
  assign OUT1[1] = IN0[1];
  assign OUT1[0] = IN0[0];

endmodule


module RCA_N4_0 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_0 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(1'b0), .S(S[0]), .Co(CTMP[1]) );
  FA_127 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_126 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_125 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module shift_thirdLevel ( sel, A, Y );
  input [2:0] sel;
  input [38:0] A;
  output [31:0] Y;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n1, n3, n71,
         n72, n73, n74, n75;

  MUX2_X1 U7 ( .A(n7), .B(n6), .S(n3), .Z(Y[30]) );
  MUX2_X1 U10 ( .A(n6), .B(n9), .S(n3), .Z(Y[29]) );
  MUX2_X1 U13 ( .A(n9), .B(n11), .S(sel[0]), .Z(Y[28]) );
  MUX2_X1 U16 ( .A(n11), .B(n13), .S(n3), .Z(Y[27]) );
  MUX2_X1 U19 ( .A(n13), .B(n15), .S(n3), .Z(Y[26]) );
  MUX2_X1 U22 ( .A(n15), .B(n17), .S(n3), .Z(Y[25]) );
  MUX2_X1 U25 ( .A(n17), .B(n19), .S(n3), .Z(Y[24]) );
  MUX2_X1 U28 ( .A(n19), .B(n21), .S(n3), .Z(Y[23]) );
  MUX2_X1 U31 ( .A(n21), .B(n23), .S(n3), .Z(Y[22]) );
  MUX2_X1 U34 ( .A(n23), .B(n25), .S(n3), .Z(Y[21]) );
  MUX2_X1 U37 ( .A(n25), .B(n27), .S(n3), .Z(Y[20]) );
  MUX2_X1 U40 ( .A(n27), .B(n29), .S(n3), .Z(Y[19]) );
  MUX2_X1 U43 ( .A(n29), .B(n31), .S(n3), .Z(Y[18]) );
  MUX2_X1 U46 ( .A(n31), .B(n33), .S(n3), .Z(Y[17]) );
  MUX2_X1 U49 ( .A(n33), .B(n35), .S(sel[0]), .Z(Y[16]) );
  MUX2_X1 U52 ( .A(n35), .B(n37), .S(sel[0]), .Z(Y[15]) );
  MUX2_X1 U55 ( .A(n37), .B(n39), .S(n3), .Z(Y[14]) );
  MUX2_X1 U58 ( .A(n39), .B(n41), .S(sel[0]), .Z(Y[13]) );
  MUX2_X1 U61 ( .A(n41), .B(n43), .S(sel[0]), .Z(Y[12]) );
  MUX2_X1 U64 ( .A(n43), .B(n45), .S(sel[0]), .Z(Y[11]) );
  MUX2_X1 U67 ( .A(n45), .B(n47), .S(sel[0]), .Z(Y[10]) );
  MUX2_X1 U70 ( .A(n47), .B(n49), .S(sel[0]), .Z(Y[9]) );
  MUX2_X1 U73 ( .A(n49), .B(n51), .S(sel[0]), .Z(Y[8]) );
  MUX2_X1 U76 ( .A(n51), .B(n53), .S(n3), .Z(Y[7]) );
  MUX2_X1 U79 ( .A(n53), .B(n55), .S(n3), .Z(Y[6]) );
  MUX2_X1 U82 ( .A(n55), .B(n57), .S(n3), .Z(Y[5]) );
  MUX2_X1 U85 ( .A(n57), .B(n59), .S(n3), .Z(Y[4]) );
  MUX2_X1 U88 ( .A(n59), .B(n61), .S(n3), .Z(Y[3]) );
  MUX2_X1 U91 ( .A(n61), .B(n63), .S(n3), .Z(Y[2]) );
  MUX2_X1 U92 ( .A(n63), .B(n64), .S(n3), .Z(Y[1]) );
  MUX2_X1 U97 ( .A(n64), .B(n67), .S(n3), .Z(Y[0]) );
  MUX2_X1 U102 ( .A(n70), .B(n7), .S(n3), .Z(Y[31]) );
  AOI22_X1 U93 ( .A1(n74), .A2(A[1]), .B1(A[5]), .B2(n72), .ZN(n65) );
  AOI22_X1 U86 ( .A1(n75), .A2(A[3]), .B1(A[7]), .B2(n73), .ZN(n60) );
  AOI22_X1 U94 ( .A1(sel[1]), .A2(n65), .B1(n60), .B2(n1), .ZN(n64) );
  AOI22_X1 U95 ( .A1(n74), .A2(A[0]), .B1(A[4]), .B2(n73), .ZN(n66) );
  AOI22_X1 U89 ( .A1(n75), .A2(A[2]), .B1(A[6]), .B2(n72), .ZN(n62) );
  AOI22_X1 U96 ( .A1(n71), .A2(n66), .B1(n62), .B2(n1), .ZN(n67) );
  AOI22_X1 U20 ( .A1(sel[2]), .A2(A[25]), .B1(A[29]), .B2(n72), .ZN(n16) );
  AOI22_X1 U14 ( .A1(sel[2]), .A2(A[27]), .B1(A[31]), .B2(n72), .ZN(n12) );
  AOI22_X1 U21 ( .A1(n71), .A2(n16), .B1(n12), .B2(n1), .ZN(n17) );
  AOI22_X1 U23 ( .A1(sel[2]), .A2(A[24]), .B1(A[28]), .B2(n72), .ZN(n18) );
  AOI22_X1 U17 ( .A1(n75), .A2(A[26]), .B1(A[30]), .B2(n72), .ZN(n14) );
  AOI22_X1 U24 ( .A1(sel[1]), .A2(n18), .B1(n14), .B2(n1), .ZN(n19) );
  AOI22_X1 U8 ( .A1(sel[2]), .A2(A[29]), .B1(A[33]), .B2(n72), .ZN(n8) );
  AOI22_X1 U4 ( .A1(sel[2]), .A2(A[31]), .B1(A[35]), .B2(n72), .ZN(n4) );
  AOI22_X1 U9 ( .A1(n71), .A2(n8), .B1(n4), .B2(n1), .ZN(n9) );
  AOI22_X1 U11 ( .A1(sel[2]), .A2(A[28]), .B1(A[32]), .B2(n72), .ZN(n10) );
  AOI22_X1 U5 ( .A1(n74), .A2(A[30]), .B1(A[34]), .B2(n72), .ZN(n5) );
  AOI22_X1 U12 ( .A1(n71), .A2(n10), .B1(n5), .B2(n1), .ZN(n11) );
  AOI22_X1 U32 ( .A1(n74), .A2(A[21]), .B1(A[25]), .B2(n72), .ZN(n24) );
  AOI22_X1 U26 ( .A1(n74), .A2(A[23]), .B1(A[27]), .B2(n72), .ZN(n20) );
  AOI22_X1 U33 ( .A1(n71), .A2(n24), .B1(n20), .B2(n1), .ZN(n25) );
  AOI22_X1 U35 ( .A1(n74), .A2(A[20]), .B1(A[24]), .B2(n73), .ZN(n26) );
  AOI22_X1 U29 ( .A1(n74), .A2(A[22]), .B1(A[26]), .B2(n72), .ZN(n22) );
  AOI22_X1 U36 ( .A1(sel[1]), .A2(n26), .B1(n22), .B2(n1), .ZN(n27) );
  AOI22_X1 U2 ( .A1(sel[2]), .A2(A[32]), .B1(A[36]), .B2(n72), .ZN(n2) );
  AOI22_X1 U6 ( .A1(n71), .A2(n5), .B1(n2), .B2(n1), .ZN(n6) );
  AOI22_X1 U30 ( .A1(n71), .A2(n22), .B1(n18), .B2(n1), .ZN(n23) );
  AOI22_X1 U18 ( .A1(n71), .A2(n14), .B1(n10), .B2(n1), .ZN(n15) );
  AOI22_X1 U15 ( .A1(n71), .A2(n12), .B1(n8), .B2(n1), .ZN(n13) );
  AOI22_X1 U27 ( .A1(n71), .A2(n20), .B1(n16), .B2(n1), .ZN(n21) );
  AOI22_X1 U98 ( .A1(sel[2]), .A2(A[33]), .B1(A[37]), .B2(n72), .ZN(n68) );
  AOI22_X1 U99 ( .A1(n71), .A2(n4), .B1(n68), .B2(n1), .ZN(n7) );
  AOI22_X1 U100 ( .A1(sel[2]), .A2(A[34]), .B1(A[38]), .B2(n73), .ZN(n69) );
  AOI22_X1 U101 ( .A1(sel[1]), .A2(n2), .B1(n69), .B2(n1), .ZN(n70) );
  AOI22_X1 U41 ( .A1(n74), .A2(A[18]), .B1(A[22]), .B2(n73), .ZN(n30) );
  AOI22_X1 U42 ( .A1(n71), .A2(n30), .B1(n26), .B2(n1), .ZN(n31) );
  AOI22_X1 U44 ( .A1(n75), .A2(A[17]), .B1(A[21]), .B2(n73), .ZN(n32) );
  AOI22_X1 U38 ( .A1(n75), .A2(A[19]), .B1(A[23]), .B2(n73), .ZN(n28) );
  AOI22_X1 U45 ( .A1(n71), .A2(n32), .B1(n28), .B2(n1), .ZN(n33) );
  AOI22_X1 U39 ( .A1(n71), .A2(n28), .B1(n24), .B2(n1), .ZN(n29) );
  AOI22_X1 U47 ( .A1(n75), .A2(A[16]), .B1(A[20]), .B2(n73), .ZN(n34) );
  AOI22_X1 U48 ( .A1(sel[1]), .A2(n34), .B1(n30), .B2(n1), .ZN(n35) );
  AOI22_X1 U53 ( .A1(n75), .A2(A[14]), .B1(A[18]), .B2(n73), .ZN(n38) );
  AOI22_X1 U54 ( .A1(n71), .A2(n38), .B1(n34), .B2(n1), .ZN(n39) );
  AOI22_X1 U56 ( .A1(n75), .A2(A[13]), .B1(A[17]), .B2(n73), .ZN(n40) );
  AOI22_X1 U50 ( .A1(n75), .A2(A[15]), .B1(A[19]), .B2(n73), .ZN(n36) );
  AOI22_X1 U57 ( .A1(n71), .A2(n40), .B1(n36), .B2(n1), .ZN(n41) );
  AOI22_X1 U59 ( .A1(n74), .A2(A[12]), .B1(A[16]), .B2(n73), .ZN(n42) );
  AOI22_X1 U60 ( .A1(sel[1]), .A2(n42), .B1(n38), .B2(n1), .ZN(n43) );
  AOI22_X1 U51 ( .A1(n71), .A2(n36), .B1(n32), .B2(n1), .ZN(n37) );
  AOI22_X1 U62 ( .A1(n74), .A2(A[11]), .B1(A[15]), .B2(n73), .ZN(n44) );
  AOI22_X1 U63 ( .A1(n71), .A2(n44), .B1(n40), .B2(n1), .ZN(n45) );
  AOI22_X1 U65 ( .A1(n74), .A2(A[10]), .B1(A[14]), .B2(n73), .ZN(n46) );
  AOI22_X1 U66 ( .A1(sel[1]), .A2(n46), .B1(n42), .B2(n1), .ZN(n47) );
  AOI22_X1 U68 ( .A1(n74), .A2(A[9]), .B1(A[13]), .B2(n73), .ZN(n48) );
  AOI22_X1 U69 ( .A1(sel[1]), .A2(n48), .B1(n44), .B2(n1), .ZN(n49) );
  AOI22_X1 U71 ( .A1(n74), .A2(A[8]), .B1(A[12]), .B2(n73), .ZN(n50) );
  AOI22_X1 U72 ( .A1(n71), .A2(n50), .B1(n46), .B2(n1), .ZN(n51) );
  AOI22_X1 U74 ( .A1(n75), .A2(A[7]), .B1(A[11]), .B2(n72), .ZN(n52) );
  AOI22_X1 U75 ( .A1(sel[1]), .A2(n52), .B1(n48), .B2(n1), .ZN(n53) );
  AOI22_X1 U83 ( .A1(n75), .A2(A[4]), .B1(A[8]), .B2(n72), .ZN(n58) );
  AOI22_X1 U77 ( .A1(n75), .A2(A[6]), .B1(A[10]), .B2(n73), .ZN(n54) );
  AOI22_X1 U84 ( .A1(n71), .A2(n58), .B1(n54), .B2(n1), .ZN(n59) );
  AOI22_X1 U80 ( .A1(sel[2]), .A2(A[5]), .B1(A[9]), .B2(n73), .ZN(n56) );
  AOI22_X1 U87 ( .A1(sel[1]), .A2(n60), .B1(n56), .B2(n1), .ZN(n61) );
  AOI22_X1 U78 ( .A1(n71), .A2(n54), .B1(n50), .B2(n1), .ZN(n55) );
  AOI22_X1 U81 ( .A1(n71), .A2(n56), .B1(n52), .B2(n1), .ZN(n57) );
  AOI22_X1 U90 ( .A1(n71), .A2(n62), .B1(n58), .B2(n1), .ZN(n63) );
  INV_X2 U1 ( .A(n71), .ZN(n1) );
  BUF_X1 U3 ( .A(sel[1]), .Z(n71) );
  BUF_X1 U103 ( .A(sel[0]), .Z(n3) );
  BUF_X1 U104 ( .A(sel[2]), .Z(n74) );
  BUF_X1 U105 ( .A(sel[2]), .Z(n75) );
  INV_X1 U106 ( .A(n75), .ZN(n73) );
  INV_X1 U107 ( .A(n75), .ZN(n72) );
endmodule


module shift_secondLevel ( sel, mask00, mask08, mask16, Y );
  input [1:0] sel;
  input [38:0] mask00;
  input [38:0] mask08;
  input [38:0] mask16;
  output [38:0] Y;
  wire   n42, n43, n44, n45, n46, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n1, n2, n3, n4, n5;

  AOI222_X1 U57 ( .A1(n2), .A2(mask00[1]), .B1(n5), .B2(mask16[1]), .C1(n4), 
        .C2(mask08[1]), .ZN(n72) );
  AOI222_X1 U11 ( .A1(n2), .A2(mask00[5]), .B1(n5), .B2(mask16[5]), .C1(n4), 
        .C2(mask08[5]), .ZN(n49) );
  AOI222_X1 U15 ( .A1(n2), .A2(mask00[3]), .B1(n5), .B2(mask16[3]), .C1(n4), 
        .C2(mask08[3]), .ZN(n51) );
  AOI222_X1 U79 ( .A1(n2), .A2(mask00[0]), .B1(n5), .B2(mask16[0]), .C1(n4), 
        .C2(mask08[0]), .ZN(n83) );
  AOI222_X1 U13 ( .A1(n2), .A2(mask00[4]), .B1(n5), .B2(mask16[4]), .C1(n4), 
        .C2(mask08[4]), .ZN(n50) );
  AOI222_X1 U35 ( .A1(n2), .A2(mask00[2]), .B1(n44), .B2(mask16[2]), .C1(n3), 
        .C2(mask08[2]), .ZN(n61) );
  AOI222_X1 U9 ( .A1(n2), .A2(mask00[6]), .B1(n5), .B2(mask16[6]), .C1(n4), 
        .C2(mask08[6]), .ZN(n48) );
  AOI222_X1 U45 ( .A1(n2), .A2(mask00[25]), .B1(n44), .B2(mask16[25]), .C1(n3), 
        .C2(mask08[25]), .ZN(n66) );
  AOI222_X1 U37 ( .A1(n2), .A2(mask00[29]), .B1(n44), .B2(mask16[29]), .C1(n3), 
        .C2(mask08[29]), .ZN(n62) );
  AOI222_X1 U41 ( .A1(n2), .A2(mask00[27]), .B1(n44), .B2(mask16[27]), .C1(n3), 
        .C2(mask08[27]), .ZN(n64) );
  AOI222_X1 U31 ( .A1(n2), .A2(mask00[31]), .B1(n5), .B2(mask16[31]), .C1(n4), 
        .C2(mask08[31]), .ZN(n59) );
  AOI222_X1 U47 ( .A1(n2), .A2(mask00[24]), .B1(n44), .B2(mask16[24]), .C1(n3), 
        .C2(mask08[24]), .ZN(n67) );
  AOI222_X1 U39 ( .A1(n2), .A2(mask00[28]), .B1(n44), .B2(mask16[28]), .C1(n3), 
        .C2(mask08[28]), .ZN(n63) );
  AOI222_X1 U43 ( .A1(n2), .A2(mask00[26]), .B1(n5), .B2(mask16[26]), .C1(n3), 
        .C2(mask08[26]), .ZN(n65) );
  AOI222_X1 U33 ( .A1(n2), .A2(mask00[30]), .B1(n44), .B2(mask16[30]), .C1(n3), 
        .C2(mask08[30]), .ZN(n60) );
  AOI222_X1 U27 ( .A1(n2), .A2(mask00[33]), .B1(n5), .B2(mask16[33]), .C1(n4), 
        .C2(mask08[33]), .ZN(n57) );
  AOI222_X1 U23 ( .A1(n2), .A2(mask00[35]), .B1(n5), .B2(mask16[35]), .C1(n4), 
        .C2(mask08[35]), .ZN(n55) );
  AOI222_X1 U29 ( .A1(n2), .A2(mask00[32]), .B1(n5), .B2(mask16[32]), .C1(n4), 
        .C2(mask08[32]), .ZN(n58) );
  AOI222_X1 U25 ( .A1(n2), .A2(mask00[34]), .B1(n5), .B2(mask16[34]), .C1(n4), 
        .C2(mask08[34]), .ZN(n56) );
  AOI222_X1 U53 ( .A1(n2), .A2(mask00[21]), .B1(n44), .B2(mask16[21]), .C1(n3), 
        .C2(mask08[21]), .ZN(n70) );
  AOI222_X1 U49 ( .A1(n2), .A2(mask00[23]), .B1(n44), .B2(mask16[23]), .C1(n3), 
        .C2(mask08[23]), .ZN(n68) );
  AOI222_X1 U55 ( .A1(n2), .A2(mask00[20]), .B1(n5), .B2(mask16[20]), .C1(n3), 
        .C2(mask08[20]), .ZN(n71) );
  AOI222_X1 U51 ( .A1(n2), .A2(mask00[22]), .B1(n44), .B2(mask16[22]), .C1(n3), 
        .C2(mask08[22]), .ZN(n69) );
  AOI222_X1 U21 ( .A1(n2), .A2(mask00[36]), .B1(n5), .B2(mask16[36]), .C1(n4), 
        .C2(mask08[36]), .ZN(n54) );
  AOI222_X1 U19 ( .A1(n2), .A2(mask00[37]), .B1(n5), .B2(mask16[37]), .C1(n4), 
        .C2(mask08[37]), .ZN(n53) );
  AOI222_X1 U17 ( .A1(n2), .A2(mask00[38]), .B1(n5), .B2(mask16[38]), .C1(n4), 
        .C2(mask08[38]), .ZN(n52) );
  AOI222_X1 U61 ( .A1(n2), .A2(mask00[18]), .B1(n5), .B2(mask16[18]), .C1(n4), 
        .C2(mask08[18]), .ZN(n74) );
  AOI222_X1 U63 ( .A1(n2), .A2(mask00[17]), .B1(n5), .B2(mask16[17]), .C1(n4), 
        .C2(mask08[17]), .ZN(n75) );
  AOI222_X1 U59 ( .A1(n2), .A2(mask00[19]), .B1(n5), .B2(mask16[19]), .C1(n4), 
        .C2(mask08[19]), .ZN(n73) );
  AOI222_X1 U65 ( .A1(n2), .A2(mask00[16]), .B1(n5), .B2(mask16[16]), .C1(n4), 
        .C2(mask08[16]), .ZN(n76) );
  AOI222_X1 U69 ( .A1(n2), .A2(mask00[14]), .B1(n5), .B2(mask16[14]), .C1(n4), 
        .C2(mask08[14]), .ZN(n78) );
  AOI222_X1 U71 ( .A1(n2), .A2(mask00[13]), .B1(n5), .B2(mask16[13]), .C1(n4), 
        .C2(mask08[13]), .ZN(n79) );
  AOI222_X1 U67 ( .A1(n2), .A2(mask00[15]), .B1(n5), .B2(mask16[15]), .C1(n4), 
        .C2(mask08[15]), .ZN(n77) );
  AOI222_X1 U73 ( .A1(n2), .A2(mask00[12]), .B1(n5), .B2(mask16[12]), .C1(n4), 
        .C2(mask08[12]), .ZN(n80) );
  AOI222_X1 U75 ( .A1(n2), .A2(mask00[11]), .B1(n5), .B2(mask16[11]), .C1(n4), 
        .C2(mask08[11]), .ZN(n81) );
  AOI222_X1 U77 ( .A1(n2), .A2(mask00[10]), .B1(n5), .B2(mask16[10]), .C1(n4), 
        .C2(mask08[10]), .ZN(n82) );
  AOI222_X1 U3 ( .A1(n2), .A2(mask00[9]), .B1(n44), .B2(mask16[9]), .C1(n4), 
        .C2(mask08[9]), .ZN(n42) );
  AOI222_X1 U5 ( .A1(n2), .A2(mask00[8]), .B1(n5), .B2(mask16[8]), .C1(n3), 
        .C2(mask08[8]), .ZN(n46) );
  INV_X1 U82 ( .A(sel[0]), .ZN(n84) );
  INV_X1 U56 ( .A(n72), .ZN(Y[1]) );
  INV_X1 U10 ( .A(n49), .ZN(Y[5]) );
  INV_X1 U14 ( .A(n51), .ZN(Y[3]) );
  INV_X1 U78 ( .A(n83), .ZN(Y[0]) );
  INV_X1 U12 ( .A(n50), .ZN(Y[4]) );
  INV_X1 U34 ( .A(n61), .ZN(Y[2]) );
  INV_X1 U8 ( .A(n48), .ZN(Y[6]) );
  INV_X1 U44 ( .A(n66), .ZN(Y[25]) );
  INV_X1 U36 ( .A(n62), .ZN(Y[29]) );
  INV_X1 U40 ( .A(n64), .ZN(Y[27]) );
  INV_X1 U30 ( .A(n59), .ZN(Y[31]) );
  INV_X1 U46 ( .A(n67), .ZN(Y[24]) );
  INV_X1 U38 ( .A(n63), .ZN(Y[28]) );
  INV_X1 U42 ( .A(n65), .ZN(Y[26]) );
  INV_X1 U32 ( .A(n60), .ZN(Y[30]) );
  INV_X1 U26 ( .A(n57), .ZN(Y[33]) );
  INV_X1 U22 ( .A(n55), .ZN(Y[35]) );
  INV_X1 U28 ( .A(n58), .ZN(Y[32]) );
  INV_X1 U24 ( .A(n56), .ZN(Y[34]) );
  INV_X1 U52 ( .A(n70), .ZN(Y[21]) );
  INV_X1 U48 ( .A(n68), .ZN(Y[23]) );
  INV_X1 U54 ( .A(n71), .ZN(Y[20]) );
  INV_X1 U50 ( .A(n69), .ZN(Y[22]) );
  INV_X1 U20 ( .A(n54), .ZN(Y[36]) );
  INV_X1 U18 ( .A(n53), .ZN(Y[37]) );
  INV_X1 U16 ( .A(n52), .ZN(Y[38]) );
  INV_X1 U60 ( .A(n74), .ZN(Y[18]) );
  INV_X1 U62 ( .A(n75), .ZN(Y[17]) );
  INV_X1 U58 ( .A(n73), .ZN(Y[19]) );
  INV_X1 U64 ( .A(n76), .ZN(Y[16]) );
  INV_X1 U68 ( .A(n78), .ZN(Y[14]) );
  INV_X1 U70 ( .A(n79), .ZN(Y[13]) );
  INV_X1 U66 ( .A(n77), .ZN(Y[15]) );
  INV_X1 U72 ( .A(n80), .ZN(Y[12]) );
  INV_X1 U74 ( .A(n81), .ZN(Y[11]) );
  INV_X1 U76 ( .A(n82), .ZN(Y[10]) );
  INV_X1 U2 ( .A(n42), .ZN(Y[9]) );
  INV_X1 U4 ( .A(n46), .ZN(Y[8]) );
  AOI222_X1 U6 ( .A1(n44), .A2(mask16[7]), .B1(n4), .B2(mask08[7]), .C1(
        mask00[7]), .C2(n2), .ZN(n1) );
  INV_X1 U7 ( .A(n1), .ZN(Y[7]) );
  BUF_X2 U80 ( .A(n43), .Z(n2) );
  BUF_X1 U81 ( .A(n45), .Z(n3) );
  BUF_X2 U83 ( .A(n44), .Z(n5) );
  BUF_X1 U84 ( .A(n45), .Z(n4) );
  AND2_X1 U85 ( .A1(n84), .A2(sel[1]), .ZN(n44) );
  NOR2_X1 U86 ( .A1(sel[1]), .A2(n84), .ZN(n45) );
  NOR2_X1 U87 ( .A1(sel[1]), .A2(sel[0]), .ZN(n43) );
endmodule


module shift_firstLevel ( A, sel, mask00, mask08, mask16 );
  input [31:0] A;
  input [1:0] sel;
  output [38:0] mask00;
  output [38:0] mask08;
  output [38:0] mask16;
  wire   n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n89, n90, n91, n92, n93, n94,
         n95, n96, n1, n2, \mask16[17] , n4;
  assign mask08[30] = mask16[38];
  assign mask08[29] = mask16[37];
  assign mask08[28] = mask16[36];
  assign mask08[27] = mask16[35];
  assign mask08[26] = mask16[34];
  assign mask08[25] = mask16[33];
  assign mask08[24] = mask16[32];
  assign mask08[14] = mask16[6];
  assign mask08[13] = mask16[5];
  assign mask08[12] = mask16[4];
  assign mask08[11] = mask16[3];
  assign mask08[10] = mask16[2];
  assign mask08[9] = mask16[1];
  assign mask08[8] = mask16[0];
  assign mask16[18] = \mask16[17] ;
  assign mask16[19] = \mask16[17] ;
  assign mask16[20] = \mask16[17] ;
  assign mask16[22] = \mask16[17] ;
  assign mask16[21] = \mask16[17] ;
  assign mask16[16] = \mask16[17] ;
  assign mask16[17] = \mask16[17] ;

  NAND2_X1 U134 ( .A1(n4), .A2(A[17]), .ZN(n55) );
  NAND2_X1 U59 ( .A1(sel[0]), .A2(A[9]), .ZN(n79) );
  NAND2_X1 U122 ( .A1(sel[0]), .A2(A[21]), .ZN(n81) );
  NAND2_X1 U146 ( .A1(sel[0]), .A2(A[13]), .ZN(n59) );
  NAND2_X1 U129 ( .A1(sel[0]), .A2(A[19]), .ZN(n83) );
  NAND2_X1 U152 ( .A1(sel[0]), .A2(A[11]), .ZN(n61) );
  NAND2_X1 U67 ( .A1(n2), .A2(A[0]), .ZN(n49) );
  NAND2_X1 U116 ( .A1(n4), .A2(A[23]), .ZN(n39) );
  NAND2_X1 U140 ( .A1(sel[0]), .A2(A[15]), .ZN(n57) );
  NAND2_X1 U137 ( .A1(sel[0]), .A2(A[16]), .ZN(n56) );
  NAND2_X1 U62 ( .A1(n4), .A2(A[8]), .ZN(n85) );
  NAND2_X1 U125 ( .A1(sel[0]), .A2(A[20]), .ZN(n82) );
  NAND2_X1 U149 ( .A1(sel[0]), .A2(A[12]), .ZN(n60) );
  NAND2_X1 U131 ( .A1(n4), .A2(A[18]), .ZN(n84) );
  NAND2_X1 U155 ( .A1(sel[0]), .A2(A[10]), .ZN(n71) );
  NAND2_X1 U119 ( .A1(n4), .A2(A[22]), .ZN(n80) );
  NAND2_X1 U143 ( .A1(sel[0]), .A2(A[14]), .ZN(n58) );
  NAND2_X1 U110 ( .A1(n4), .A2(A[25]), .ZN(n37) );
  NAND2_X1 U109 ( .A1(n2), .A2(A[18]), .ZN(n67) );
  NAND2_X1 U108 ( .A1(n37), .A2(n67), .ZN(mask00[25]) );
  NAND2_X1 U91 ( .A1(n4), .A2(A[31]), .ZN(n78) );
  NAND2_X1 U60 ( .A1(n2), .A2(A[2]), .ZN(n47) );
  NAND2_X1 U11 ( .A1(n41), .A2(n47), .ZN(mask16[25]) );
  NAND2_X1 U135 ( .A1(n2), .A2(A[10]), .ZN(n76) );
  NAND2_X1 U40 ( .A1(n76), .A2(n41), .ZN(mask16[33]) );
  NAND2_X1 U98 ( .A1(n4), .A2(A[29]), .ZN(n51) );
  NAND2_X1 U97 ( .A1(n2), .A2(A[22]), .ZN(n63) );
  NAND2_X1 U96 ( .A1(n51), .A2(n63), .ZN(mask00[29]) );
  NAND2_X1 U147 ( .A1(n86), .A2(A[6]), .ZN(n43) );
  NAND2_X1 U7 ( .A1(n43), .A2(n41), .ZN(mask16[29]) );
  NAND2_X1 U121 ( .A1(n86), .A2(A[14]), .ZN(n72) );
  NAND2_X1 U36 ( .A1(n72), .A2(n41), .ZN(mask16[37]) );
  NAND2_X1 U104 ( .A1(n4), .A2(A[27]), .ZN(n53) );
  NAND2_X1 U103 ( .A1(n2), .A2(A[20]), .ZN(n65) );
  NAND2_X1 U102 ( .A1(n53), .A2(n65), .ZN(mask00[27]) );
  NAND2_X1 U153 ( .A1(n2), .A2(A[4]), .ZN(n45) );
  NAND2_X1 U9 ( .A1(n45), .A2(n41), .ZN(mask16[27]) );
  NAND2_X1 U128 ( .A1(n86), .A2(A[12]), .ZN(n74) );
  NAND2_X1 U38 ( .A1(n74), .A2(n41), .ZN(mask16[35]) );
  AOI21_X1 U89 ( .B1(A[24]), .B2(n2), .A(mask16[15]), .ZN(n96) );
  NAND2_X1 U141 ( .A1(n2), .A2(A[8]), .ZN(n40) );
  NAND2_X1 U5 ( .A1(n40), .A2(n41), .ZN(mask16[31]) );
  NAND2_X1 U115 ( .A1(n2), .A2(A[16]), .ZN(n69) );
  NAND2_X1 U33 ( .A1(n69), .A2(n41), .ZN(mask08[31]) );
  NAND2_X1 U113 ( .A1(n4), .A2(A[24]), .ZN(n38) );
  NAND2_X1 U112 ( .A1(n2), .A2(A[17]), .ZN(n68) );
  NAND2_X1 U111 ( .A1(n38), .A2(n68), .ZN(mask00[24]) );
  NAND2_X1 U63 ( .A1(n2), .A2(A[1]), .ZN(n48) );
  NAND2_X1 U12 ( .A1(n41), .A2(n48), .ZN(mask16[24]) );
  NAND2_X1 U138 ( .A1(n2), .A2(A[9]), .ZN(n77) );
  NAND2_X1 U41 ( .A1(n77), .A2(n41), .ZN(mask16[32]) );
  NAND2_X1 U101 ( .A1(n4), .A2(A[28]), .ZN(n52) );
  NAND2_X1 U100 ( .A1(n2), .A2(A[21]), .ZN(n64) );
  NAND2_X1 U99 ( .A1(n52), .A2(n64), .ZN(mask00[28]) );
  NAND2_X1 U150 ( .A1(n2), .A2(A[5]), .ZN(n44) );
  NAND2_X1 U8 ( .A1(n44), .A2(n41), .ZN(mask16[28]) );
  NAND2_X1 U124 ( .A1(n86), .A2(A[13]), .ZN(n73) );
  NAND2_X1 U37 ( .A1(n73), .A2(n41), .ZN(mask16[36]) );
  NAND2_X1 U107 ( .A1(n4), .A2(A[26]), .ZN(n54) );
  NAND2_X1 U106 ( .A1(n2), .A2(A[19]), .ZN(n66) );
  NAND2_X1 U105 ( .A1(n54), .A2(n66), .ZN(mask00[26]) );
  NAND2_X1 U156 ( .A1(n2), .A2(A[3]), .ZN(n46) );
  NAND2_X1 U10 ( .A1(n46), .A2(n41), .ZN(mask16[26]) );
  NAND2_X1 U132 ( .A1(n86), .A2(A[11]), .ZN(n75) );
  NAND2_X1 U39 ( .A1(n75), .A2(n41), .ZN(mask16[34]) );
  NAND2_X1 U94 ( .A1(n4), .A2(A[30]), .ZN(n50) );
  NAND2_X1 U93 ( .A1(n2), .A2(A[23]), .ZN(n62) );
  NAND2_X1 U92 ( .A1(n50), .A2(n62), .ZN(mask00[30]) );
  NAND2_X1 U144 ( .A1(n2), .A2(A[7]), .ZN(n42) );
  NAND2_X1 U6 ( .A1(n42), .A2(n41), .ZN(mask16[30]) );
  NAND2_X1 U118 ( .A1(n86), .A2(A[15]), .ZN(n70) );
  NAND2_X1 U34 ( .A1(n70), .A2(n41), .ZN(mask16[38]) );
  AOI21_X1 U83 ( .B1(A[26]), .B2(n2), .A(\mask16[17] ), .ZN(n94) );
  NAND2_X1 U31 ( .A1(n67), .A2(n41), .ZN(mask08[33]) );
  AOI21_X1 U79 ( .B1(A[28]), .B2(n2), .A(\mask16[17] ), .ZN(n92) );
  NAND2_X1 U29 ( .A1(n65), .A2(n41), .ZN(mask08[35]) );
  AOI21_X1 U85 ( .B1(A[25]), .B2(n2), .A(\mask16[17] ), .ZN(n95) );
  NAND2_X1 U32 ( .A1(n68), .A2(n41), .ZN(mask08[32]) );
  AOI21_X1 U81 ( .B1(A[27]), .B2(n2), .A(\mask16[17] ), .ZN(n93) );
  NAND2_X1 U30 ( .A1(n66), .A2(n41), .ZN(mask08[34]) );
  NAND2_X1 U120 ( .A1(n81), .A2(n72), .ZN(mask00[21]) );
  NAND2_X1 U44 ( .A1(n43), .A2(n51), .ZN(mask08[21]) );
  NAND2_X1 U114 ( .A1(n39), .A2(n69), .ZN(mask00[23]) );
  NAND2_X1 U13 ( .A1(n41), .A2(n49), .ZN(mask16[23]) );
  NAND2_X1 U42 ( .A1(n40), .A2(n78), .ZN(mask08[23]) );
  NAND2_X1 U123 ( .A1(n82), .A2(n73), .ZN(mask00[20]) );
  NAND2_X1 U45 ( .A1(n44), .A2(n52), .ZN(mask08[20]) );
  NAND2_X1 U117 ( .A1(n80), .A2(n70), .ZN(mask00[22]) );
  NAND2_X1 U43 ( .A1(n42), .A2(n50), .ZN(mask08[22]) );
  AOI21_X1 U77 ( .B1(A[29]), .B2(n2), .A(\mask16[17] ), .ZN(n91) );
  NAND2_X1 U28 ( .A1(n64), .A2(n41), .ZN(mask08[36]) );
  AOI21_X1 U75 ( .B1(A[30]), .B2(n2), .A(\mask16[17] ), .ZN(n90) );
  NAND2_X1 U27 ( .A1(n63), .A2(n41), .ZN(mask08[37]) );
  AOI21_X1 U73 ( .B1(A[31]), .B2(n2), .A(\mask16[17] ), .ZN(n89) );
  NAND2_X1 U26 ( .A1(n62), .A2(n41), .ZN(mask08[38]) );
  NAND2_X1 U130 ( .A1(n75), .A2(n84), .ZN(mask00[18]) );
  NAND2_X1 U48 ( .A1(n46), .A2(n54), .ZN(mask08[18]) );
  NAND2_X1 U133 ( .A1(n76), .A2(n55), .ZN(mask00[17]) );
  NAND2_X1 U49 ( .A1(n37), .A2(n47), .ZN(mask08[17]) );
  NAND2_X1 U127 ( .A1(n83), .A2(n74), .ZN(mask00[19]) );
  NAND2_X1 U47 ( .A1(n45), .A2(n53), .ZN(mask08[19]) );
  NAND2_X1 U136 ( .A1(n77), .A2(n56), .ZN(mask00[16]) );
  NAND2_X1 U50 ( .A1(n38), .A2(n48), .ZN(mask08[16]) );
  NAND2_X1 U142 ( .A1(n42), .A2(n58), .ZN(mask00[14]) );
  NAND2_X1 U145 ( .A1(n43), .A2(n59), .ZN(mask00[13]) );
  NAND2_X1 U139 ( .A1(n40), .A2(n57), .ZN(mask00[15]) );
  NAND2_X1 U51 ( .A1(n39), .A2(n49), .ZN(mask08[15]) );
  NAND2_X1 U148 ( .A1(n44), .A2(n60), .ZN(mask00[12]) );
  NAND2_X1 U151 ( .A1(n45), .A2(n61), .ZN(mask00[11]) );
  NAND2_X1 U154 ( .A1(n46), .A2(n71), .ZN(mask00[10]) );
  NAND2_X1 U58 ( .A1(n47), .A2(n79), .ZN(mask00[9]) );
  NAND2_X1 U61 ( .A1(n48), .A2(n85), .ZN(mask00[8]) );
  AND2_X1 U126 ( .A1(n4), .A2(A[1]), .ZN(mask00[1]) );
  INV_X1 U19 ( .A(n55), .ZN(mask16[1]) );
  INV_X1 U46 ( .A(n79), .ZN(mask08[1]) );
  AND2_X1 U69 ( .A1(sel[0]), .A2(A[5]), .ZN(mask00[5]) );
  INV_X1 U53 ( .A(n81), .ZN(mask16[5]) );
  INV_X1 U23 ( .A(n59), .ZN(mask08[5]) );
  AND2_X1 U71 ( .A1(sel[0]), .A2(A[3]), .ZN(mask00[3]) );
  INV_X1 U55 ( .A(n83), .ZN(mask16[3]) );
  INV_X1 U25 ( .A(n61), .ZN(mask08[3]) );
  AND2_X1 U158 ( .A1(n4), .A2(A[0]), .ZN(mask00[0]) );
  INV_X1 U20 ( .A(n56), .ZN(mask16[0]) );
  INV_X1 U57 ( .A(n85), .ZN(mask08[0]) );
  AND2_X1 U70 ( .A1(sel[0]), .A2(A[4]), .ZN(mask00[4]) );
  INV_X1 U54 ( .A(n82), .ZN(mask16[4]) );
  INV_X1 U24 ( .A(n60), .ZN(mask08[4]) );
  AND2_X1 U95 ( .A1(sel[0]), .A2(A[2]), .ZN(mask00[2]) );
  INV_X1 U56 ( .A(n84), .ZN(mask16[2]) );
  INV_X1 U35 ( .A(n71), .ZN(mask08[2]) );
  AND2_X1 U68 ( .A1(sel[0]), .A2(A[6]), .ZN(mask00[6]) );
  INV_X1 U52 ( .A(n80), .ZN(mask16[6]) );
  INV_X1 U22 ( .A(n58), .ZN(mask08[6]) );
  INV_X1 U90 ( .A(n78), .ZN(mask16[15]) );
  INV_X1 U88 ( .A(n96), .ZN(mask00[31]) );
  INV_X1 U82 ( .A(n94), .ZN(mask00[33]) );
  INV_X1 U78 ( .A(n92), .ZN(mask00[35]) );
  INV_X1 U84 ( .A(n95), .ZN(mask00[32]) );
  INV_X1 U80 ( .A(n93), .ZN(mask00[34]) );
  INV_X1 U76 ( .A(n91), .ZN(mask00[36]) );
  INV_X1 U74 ( .A(n90), .ZN(mask00[37]) );
  INV_X1 U72 ( .A(n89), .ZN(mask00[38]) );
  INV_X1 U14 ( .A(n50), .ZN(mask16[14]) );
  INV_X1 U15 ( .A(n51), .ZN(mask16[13]) );
  INV_X1 U16 ( .A(n52), .ZN(mask16[12]) );
  INV_X1 U17 ( .A(n53), .ZN(mask16[11]) );
  INV_X1 U18 ( .A(n54), .ZN(mask16[10]) );
  INV_X1 U2 ( .A(n37), .ZN(mask16[9]) );
  INV_X1 U3 ( .A(n38), .ZN(mask16[8]) );
  INV_X1 U4 ( .A(n57), .ZN(mask08[7]) );
  INV_X1 U21 ( .A(n39), .ZN(mask16[7]) );
  NAND2_X1 U64 ( .A1(n4), .A2(A[7]), .ZN(n1) );
  NAND2_X1 U65 ( .A1(n49), .A2(n1), .ZN(mask00[7]) );
  BUF_X1 U66 ( .A(n86), .Z(n2) );
  BUF_X1 U86 ( .A(sel[0]), .Z(n4) );
  INV_X1 U87 ( .A(n41), .ZN(\mask16[17] ) );
  NOR2_X1 U157 ( .A1(n4), .A2(sel[1]), .ZN(n86) );
  NAND2_X1 U159 ( .A1(sel[1]), .A2(mask16[15]), .ZN(n41) );
endmodule


module SNPS_CLOCK_GATE_HIGH_simple_booth_add_ext_N16 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net337970, net337972, net337973, net337976;
  assign net337970 = CLK;
  assign ENCLK = net337972;
  assign net337973 = EN;

  DLL_X1 latch ( .D(net337973), .GN(net337970), .Q(net337976) );
  AND2_X1 main_gate ( .A1(net337976), .A2(net337970), .ZN(net337972) );
endmodule


module piso_r_2_N32 ( Clock, ALOAD, D, SO );
  input [31:0] D;
  output [31:0] SO;
  input Clock, ALOAD;
  wire   N3, N4;

  DFF_X1 \tmp_reg[1]  ( .D(N4), .CK(Clock), .Q(SO[1]) );
  SDFF_X1 \tmp_reg[3]  ( .D(SO[1]), .SI(D[3]), .SE(ALOAD), .CK(Clock), .Q(
        SO[3]) );
  SDFF_X1 \tmp_reg[5]  ( .D(SO[3]), .SI(D[5]), .SE(ALOAD), .CK(Clock), .Q(
        SO[5]) );
  SDFF_X1 \tmp_reg[7]  ( .D(SO[5]), .SI(D[7]), .SE(ALOAD), .CK(Clock), .Q(
        SO[7]) );
  SDFF_X1 \tmp_reg[9]  ( .D(SO[7]), .SI(D[9]), .SE(ALOAD), .CK(Clock), .Q(
        SO[9]) );
  SDFF_X1 \tmp_reg[11]  ( .D(SO[9]), .SI(D[11]), .SE(ALOAD), .CK(Clock), .Q(
        SO[11]) );
  SDFF_X1 \tmp_reg[13]  ( .D(SO[11]), .SI(D[13]), .SE(ALOAD), .CK(Clock), .Q(
        SO[13]) );
  SDFF_X1 \tmp_reg[15]  ( .D(SO[13]), .SI(D[15]), .SE(ALOAD), .CK(Clock), .Q(
        SO[15]) );
  SDFF_X1 \tmp_reg[17]  ( .D(SO[15]), .SI(D[17]), .SE(ALOAD), .CK(Clock), .Q(
        SO[17]) );
  SDFF_X1 \tmp_reg[19]  ( .D(SO[17]), .SI(D[19]), .SE(ALOAD), .CK(Clock), .Q(
        SO[19]) );
  SDFF_X1 \tmp_reg[21]  ( .D(SO[19]), .SI(D[21]), .SE(ALOAD), .CK(Clock), .Q(
        SO[21]) );
  SDFF_X1 \tmp_reg[23]  ( .D(SO[21]), .SI(D[23]), .SE(ALOAD), .CK(Clock), .Q(
        SO[23]) );
  SDFF_X1 \tmp_reg[25]  ( .D(SO[23]), .SI(D[25]), .SE(ALOAD), .CK(Clock), .Q(
        SO[25]) );
  SDFF_X1 \tmp_reg[27]  ( .D(SO[25]), .SI(D[27]), .SE(ALOAD), .CK(Clock), .Q(
        SO[27]) );
  SDFF_X1 \tmp_reg[29]  ( .D(SO[27]), .SI(D[29]), .SE(ALOAD), .CK(Clock), .Q(
        SO[29]) );
  SDFF_X1 \tmp_reg[31]  ( .D(SO[29]), .SI(D[31]), .SE(ALOAD), .CK(Clock), .Q(
        SO[31]) );
  DFF_X1 \tmp_reg[0]  ( .D(N3), .CK(Clock), .Q(SO[0]) );
  SDFF_X1 \tmp_reg[2]  ( .D(SO[0]), .SI(D[2]), .SE(ALOAD), .CK(Clock), .Q(
        SO[2]) );
  SDFF_X1 \tmp_reg[4]  ( .D(SO[2]), .SI(D[4]), .SE(ALOAD), .CK(Clock), .Q(
        SO[4]) );
  SDFF_X1 \tmp_reg[6]  ( .D(SO[4]), .SI(D[6]), .SE(ALOAD), .CK(Clock), .Q(
        SO[6]) );
  SDFF_X1 \tmp_reg[8]  ( .D(SO[6]), .SI(D[8]), .SE(ALOAD), .CK(Clock), .Q(
        SO[8]) );
  SDFF_X1 \tmp_reg[10]  ( .D(SO[8]), .SI(D[10]), .SE(ALOAD), .CK(Clock), .Q(
        SO[10]) );
  SDFF_X1 \tmp_reg[12]  ( .D(SO[10]), .SI(D[12]), .SE(ALOAD), .CK(Clock), .Q(
        SO[12]) );
  SDFF_X1 \tmp_reg[14]  ( .D(SO[12]), .SI(D[14]), .SE(ALOAD), .CK(Clock), .Q(
        SO[14]) );
  SDFF_X1 \tmp_reg[16]  ( .D(SO[14]), .SI(D[16]), .SE(ALOAD), .CK(Clock), .Q(
        SO[16]) );
  SDFF_X1 \tmp_reg[18]  ( .D(SO[16]), .SI(D[18]), .SE(ALOAD), .CK(Clock), .Q(
        SO[18]) );
  SDFF_X1 \tmp_reg[20]  ( .D(SO[18]), .SI(D[20]), .SE(ALOAD), .CK(Clock), .Q(
        SO[20]) );
  SDFF_X1 \tmp_reg[22]  ( .D(SO[20]), .SI(D[22]), .SE(ALOAD), .CK(Clock), .Q(
        SO[22]) );
  SDFF_X1 \tmp_reg[24]  ( .D(SO[22]), .SI(D[24]), .SE(ALOAD), .CK(Clock), .Q(
        SO[24]) );
  SDFF_X1 \tmp_reg[26]  ( .D(SO[24]), .SI(D[26]), .SE(ALOAD), .CK(Clock), .Q(
        SO[26]) );
  SDFF_X1 \tmp_reg[28]  ( .D(SO[26]), .SI(D[28]), .SE(ALOAD), .CK(Clock), .Q(
        SO[28]) );
  SDFF_X1 \tmp_reg[30]  ( .D(SO[28]), .SI(D[30]), .SE(ALOAD), .CK(Clock), .Q(
        SO[30]) );
  AND2_X1 U4 ( .A1(ALOAD), .A2(D[0]), .ZN(N3) );
  AND2_X1 U3 ( .A1(ALOAD), .A2(D[1]), .ZN(N4) );
endmodule


module shift_N9_0 ( Clock, ALOAD, D, SO );
  input [8:0] D;
  input Clock, ALOAD;
  output SO;
  wire   N11;
  wire   [8:1] tmp;

  DFF_X1 \tmp_reg[8]  ( .D(N11), .CK(Clock), .Q(tmp[8]) );
  SDFF_X1 \tmp_reg[7]  ( .D(tmp[8]), .SI(D[7]), .SE(ALOAD), .CK(Clock), .Q(
        tmp[7]) );
  SDFF_X1 \tmp_reg[6]  ( .D(tmp[7]), .SI(D[6]), .SE(ALOAD), .CK(Clock), .Q(
        tmp[6]) );
  SDFF_X1 \tmp_reg[5]  ( .D(tmp[6]), .SI(D[5]), .SE(ALOAD), .CK(Clock), .Q(
        tmp[5]) );
  SDFF_X1 \tmp_reg[4]  ( .D(tmp[5]), .SI(D[4]), .SE(ALOAD), .CK(Clock), .Q(
        tmp[4]) );
  SDFF_X1 \tmp_reg[3]  ( .D(tmp[4]), .SI(D[3]), .SE(ALOAD), .CK(Clock), .Q(
        tmp[3]) );
  SDFF_X1 \tmp_reg[2]  ( .D(tmp[3]), .SI(D[2]), .SE(ALOAD), .CK(Clock), .Q(
        tmp[2]) );
  SDFF_X1 \tmp_reg[1]  ( .D(tmp[2]), .SI(D[1]), .SE(ALOAD), .CK(Clock), .Q(
        tmp[1]) );
  SDFF_X1 \tmp_reg[0]  ( .D(tmp[1]), .SI(D[0]), .SE(ALOAD), .CK(Clock), .Q(SO)
         );
  AND2_X1 U3 ( .A1(ALOAD), .A2(D[8]), .ZN(N11) );
endmodule


module booth_encoder_0 ( B_in, A_out );
  input [2:0] B_in;
  output [2:0] A_out;
  wire   N53, N57, n3, n4;
  assign A_out[1] = B_in[2];
  assign A_out[0] = N53;
  assign A_out[2] = N57;

  INV_X1 U7 ( .A(B_in[1]), .ZN(n3) );
  INV_X1 U3 ( .A(B_in[2]), .ZN(n4) );
  NAND2_X1 U4 ( .A1(n4), .A2(n3), .ZN(N57) );
  NOR2_X1 U5 ( .A1(B_in[1]), .A2(n4), .ZN(N53) );
endmodule


module carry_sel_gen_N4_0 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:0] nocarry_sum_to_mux;

  RCA_N4_0 rca_nocarry ( .A(A), .B(B), .Ci(1'b0), .S(nocarry_sum_to_mux) );
  mux21_SIZE4_0 outmux ( .IN0(nocarry_sum_to_mux), .IN1({1'b0, 1'b0, 1'b0, 
        1'b0}), .CTRL(1'b0), .OUT1(S) );
endmodule


module pg_0 ( g, p, g_prec, p_prec, g_out, p_out );
  input g, p, g_prec, p_prec;
  output g_out, p_out;
  wire   n2;

  AOI21_X1 U3 ( .B1(g_prec), .B2(p), .A(g), .ZN(n2) );
  AND2_X1 U1 ( .A1(p), .A2(p_prec), .ZN(p_out) );
  INV_X1 U2 ( .A(n2), .ZN(g_out) );
endmodule


module g_0 ( g, p, g_prec, g_out );
  input g, p, g_prec;
  output g_out;
  wire   g;
  assign g_out = g;

endmodule


module pg_net_0 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p_out) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g_out) );
endmodule


module logic_unit_SIZE32 ( IN1, IN2, CTRL, OUT1 );
  input [31:0] IN1;
  input [31:0] IN2;
  input [1:0] CTRL;
  output [31:0] OUT1;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n1, n2;

  AOI21_X1 U97 ( .B1(IN2[0]), .B2(IN1[0]), .A(CTRL[0]), .ZN(n66) );
  OAI22_X1 U96 ( .A1(IN1[0]), .A2(IN2[0]), .B1(n1), .B2(n66), .ZN(n67) );
  AOI21_X1 U95 ( .B1(n1), .B2(n66), .A(n67), .ZN(OUT1[0]) );
  AOI21_X1 U49 ( .B1(IN2[24]), .B2(IN1[24]), .A(n2), .ZN(n34) );
  OAI22_X1 U48 ( .A1(IN1[24]), .A2(IN2[24]), .B1(n3), .B2(n34), .ZN(n35) );
  AOI21_X1 U47 ( .B1(n1), .B2(n34), .A(n35), .ZN(OUT1[24]) );
  AOI21_X1 U37 ( .B1(IN2[28]), .B2(IN1[28]), .A(n2), .ZN(n26) );
  OAI22_X1 U36 ( .A1(IN1[28]), .A2(IN2[28]), .B1(n3), .B2(n26), .ZN(n27) );
  AOI21_X1 U35 ( .B1(n3), .B2(n26), .A(n27), .ZN(OUT1[28]) );
  AOI21_X1 U61 ( .B1(IN2[20]), .B2(IN1[20]), .A(n2), .ZN(n42) );
  OAI22_X1 U60 ( .A1(IN1[20]), .A2(IN2[20]), .B1(n1), .B2(n42), .ZN(n43) );
  AOI21_X1 U59 ( .B1(n3), .B2(n42), .A(n43), .ZN(OUT1[20]) );
  AOI21_X1 U34 ( .B1(IN2[29]), .B2(IN1[29]), .A(n2), .ZN(n24) );
  OAI22_X1 U33 ( .A1(IN1[29]), .A2(IN2[29]), .B1(n3), .B2(n24), .ZN(n25) );
  AOI21_X1 U32 ( .B1(n1), .B2(n24), .A(n25), .ZN(OUT1[29]) );
  AOI21_X1 U58 ( .B1(IN2[21]), .B2(IN1[21]), .A(n2), .ZN(n40) );
  OAI22_X1 U57 ( .A1(IN1[21]), .A2(IN2[21]), .B1(n1), .B2(n40), .ZN(n41) );
  AOI21_X1 U56 ( .B1(n3), .B2(n40), .A(n41), .ZN(OUT1[21]) );
  AOI21_X1 U46 ( .B1(IN2[25]), .B2(IN1[25]), .A(n2), .ZN(n32) );
  OAI22_X1 U45 ( .A1(IN1[25]), .A2(IN2[25]), .B1(n1), .B2(n32), .ZN(n33) );
  AOI21_X1 U44 ( .B1(n1), .B2(n32), .A(n33), .ZN(OUT1[25]) );
  AOI21_X1 U43 ( .B1(IN2[26]), .B2(IN1[26]), .A(n2), .ZN(n30) );
  OAI22_X1 U42 ( .A1(IN1[26]), .A2(IN2[26]), .B1(n1), .B2(n30), .ZN(n31) );
  AOI21_X1 U41 ( .B1(n1), .B2(n30), .A(n31), .ZN(OUT1[26]) );
  AOI21_X1 U55 ( .B1(IN2[22]), .B2(IN1[22]), .A(n2), .ZN(n38) );
  OAI22_X1 U54 ( .A1(IN1[22]), .A2(IN2[22]), .B1(n1), .B2(n38), .ZN(n39) );
  AOI21_X1 U53 ( .B1(n3), .B2(n38), .A(n39), .ZN(OUT1[22]) );
  AOI21_X1 U40 ( .B1(IN2[27]), .B2(IN1[27]), .A(n2), .ZN(n28) );
  OAI22_X1 U39 ( .A1(IN1[27]), .A2(IN2[27]), .B1(n3), .B2(n28), .ZN(n29) );
  AOI21_X1 U38 ( .B1(n3), .B2(n28), .A(n29), .ZN(OUT1[27]) );
  AOI21_X1 U52 ( .B1(IN2[23]), .B2(IN1[23]), .A(n2), .ZN(n36) );
  OAI22_X1 U51 ( .A1(IN1[23]), .A2(IN2[23]), .B1(n1), .B2(n36), .ZN(n37) );
  AOI21_X1 U50 ( .B1(n3), .B2(n36), .A(n37), .ZN(OUT1[23]) );
  AOI21_X1 U28 ( .B1(IN2[30]), .B2(IN1[30]), .A(n2), .ZN(n20) );
  OAI22_X1 U27 ( .A1(IN1[30]), .A2(IN2[30]), .B1(n1), .B2(n20), .ZN(n21) );
  AOI21_X1 U26 ( .B1(n1), .B2(n20), .A(n21), .ZN(OUT1[30]) );
  AOI21_X1 U25 ( .B1(IN2[31]), .B2(IN1[31]), .A(CTRL[0]), .ZN(n18) );
  OAI22_X1 U24 ( .A1(IN1[31]), .A2(IN2[31]), .B1(n3), .B2(n18), .ZN(n19) );
  AOI21_X1 U23 ( .B1(n3), .B2(n18), .A(n19), .ZN(OUT1[31]) );
  AOI21_X1 U73 ( .B1(IN2[17]), .B2(IN1[17]), .A(CTRL[0]), .ZN(n50) );
  OAI22_X1 U72 ( .A1(IN1[17]), .A2(IN2[17]), .B1(n1), .B2(n50), .ZN(n51) );
  AOI21_X1 U71 ( .B1(n3), .B2(n50), .A(n51), .ZN(OUT1[17]) );
  AOI21_X1 U70 ( .B1(IN2[18]), .B2(IN1[18]), .A(CTRL[0]), .ZN(n48) );
  OAI22_X1 U69 ( .A1(IN1[18]), .A2(IN2[18]), .B1(n1), .B2(n48), .ZN(n49) );
  AOI21_X1 U68 ( .B1(n1), .B2(n48), .A(n49), .ZN(OUT1[18]) );
  AOI21_X1 U67 ( .B1(IN2[19]), .B2(IN1[19]), .A(CTRL[0]), .ZN(n46) );
  OAI22_X1 U66 ( .A1(IN1[19]), .A2(IN2[19]), .B1(n1), .B2(n46), .ZN(n47) );
  AOI21_X1 U65 ( .B1(n3), .B2(n46), .A(n47), .ZN(OUT1[19]) );
  AOI21_X1 U76 ( .B1(IN2[16]), .B2(IN1[16]), .A(CTRL[0]), .ZN(n52) );
  OAI22_X1 U75 ( .A1(IN1[16]), .A2(IN2[16]), .B1(n1), .B2(n52), .ZN(n53) );
  AOI21_X1 U74 ( .B1(n3), .B2(n52), .A(n53), .ZN(OUT1[16]) );
  AOI21_X1 U85 ( .B1(IN2[13]), .B2(IN1[13]), .A(CTRL[0]), .ZN(n58) );
  OAI22_X1 U84 ( .A1(IN1[13]), .A2(IN2[13]), .B1(n1), .B2(n58), .ZN(n59) );
  AOI21_X1 U83 ( .B1(n3), .B2(n58), .A(n59), .ZN(OUT1[13]) );
  AOI21_X1 U88 ( .B1(IN2[12]), .B2(IN1[12]), .A(CTRL[0]), .ZN(n60) );
  OAI22_X1 U87 ( .A1(IN1[12]), .A2(IN2[12]), .B1(n1), .B2(n60), .ZN(n61) );
  AOI21_X1 U86 ( .B1(n3), .B2(n60), .A(n61), .ZN(OUT1[12]) );
  AOI21_X1 U82 ( .B1(IN2[14]), .B2(IN1[14]), .A(CTRL[0]), .ZN(n56) );
  OAI22_X1 U81 ( .A1(IN1[14]), .A2(IN2[14]), .B1(n1), .B2(n56), .ZN(n57) );
  AOI21_X1 U80 ( .B1(n1), .B2(n56), .A(n57), .ZN(OUT1[14]) );
  AOI21_X1 U79 ( .B1(IN2[15]), .B2(IN1[15]), .A(CTRL[0]), .ZN(n54) );
  OAI22_X1 U78 ( .A1(IN1[15]), .A2(IN2[15]), .B1(n1), .B2(n54), .ZN(n55) );
  AOI21_X1 U77 ( .B1(n3), .B2(n54), .A(n55), .ZN(OUT1[15]) );
  AOI21_X1 U94 ( .B1(IN2[10]), .B2(IN1[10]), .A(CTRL[0]), .ZN(n64) );
  OAI22_X1 U93 ( .A1(IN1[10]), .A2(IN2[10]), .B1(n1), .B2(n64), .ZN(n65) );
  AOI21_X1 U92 ( .B1(n1), .B2(n64), .A(n65), .ZN(OUT1[10]) );
  AOI21_X1 U91 ( .B1(IN2[11]), .B2(IN1[11]), .A(CTRL[0]), .ZN(n62) );
  OAI22_X1 U90 ( .A1(IN1[11]), .A2(IN2[11]), .B1(n1), .B2(n62), .ZN(n63) );
  AOI21_X1 U89 ( .B1(n1), .B2(n62), .A(n63), .ZN(OUT1[11]) );
  AOI21_X1 U7 ( .B1(IN2[8]), .B2(IN1[8]), .A(CTRL[0]), .ZN(n6) );
  OAI22_X1 U6 ( .A1(IN1[8]), .A2(IN2[8]), .B1(n1), .B2(n6), .ZN(n7) );
  AOI21_X1 U5 ( .B1(n3), .B2(n6), .A(n7), .ZN(OUT1[8]) );
  AOI21_X1 U4 ( .B1(IN2[9]), .B2(IN1[9]), .A(CTRL[0]), .ZN(n4) );
  OAI22_X1 U3 ( .A1(IN1[9]), .A2(IN2[9]), .B1(n1), .B2(n4), .ZN(n5) );
  AOI21_X1 U2 ( .B1(n1), .B2(n4), .A(n5), .ZN(OUT1[9]) );
  AOI21_X1 U10 ( .B1(IN2[7]), .B2(IN1[7]), .A(CTRL[0]), .ZN(n8) );
  OAI22_X1 U9 ( .A1(IN1[7]), .A2(IN2[7]), .B1(n1), .B2(n8), .ZN(n9) );
  AOI21_X1 U8 ( .B1(n1), .B2(n8), .A(n9), .ZN(OUT1[7]) );
  AOI21_X1 U22 ( .B1(IN2[3]), .B2(IN1[3]), .A(CTRL[0]), .ZN(n16) );
  OAI22_X1 U21 ( .A1(IN1[3]), .A2(IN2[3]), .B1(n1), .B2(n16), .ZN(n17) );
  AOI21_X1 U20 ( .B1(n3), .B2(n16), .A(n17), .ZN(OUT1[3]) );
  AOI21_X1 U13 ( .B1(IN2[6]), .B2(IN1[6]), .A(CTRL[0]), .ZN(n10) );
  OAI22_X1 U12 ( .A1(IN1[6]), .A2(IN2[6]), .B1(n1), .B2(n10), .ZN(n11) );
  AOI21_X1 U11 ( .B1(n3), .B2(n10), .A(n11), .ZN(OUT1[6]) );
  AOI21_X1 U19 ( .B1(IN2[4]), .B2(IN1[4]), .A(n2), .ZN(n14) );
  OAI22_X1 U18 ( .A1(IN1[4]), .A2(IN2[4]), .B1(n1), .B2(n14), .ZN(n15) );
  AOI21_X1 U17 ( .B1(n1), .B2(n14), .A(n15), .ZN(OUT1[4]) );
  AOI21_X1 U16 ( .B1(IN2[5]), .B2(IN1[5]), .A(n2), .ZN(n12) );
  OAI22_X1 U15 ( .A1(IN1[5]), .A2(IN2[5]), .B1(n1), .B2(n12), .ZN(n13) );
  AOI21_X1 U14 ( .B1(n1), .B2(n12), .A(n13), .ZN(OUT1[5]) );
  AOI21_X1 U31 ( .B1(IN2[2]), .B2(IN1[2]), .A(n2), .ZN(n22) );
  OAI22_X1 U30 ( .A1(IN1[2]), .A2(IN2[2]), .B1(n3), .B2(n22), .ZN(n23) );
  AOI21_X1 U29 ( .B1(n3), .B2(n22), .A(n23), .ZN(OUT1[2]) );
  AOI21_X1 U64 ( .B1(IN2[1]), .B2(IN1[1]), .A(CTRL[0]), .ZN(n44) );
  OAI22_X1 U63 ( .A1(IN1[1]), .A2(IN2[1]), .B1(n1), .B2(n44), .ZN(n45) );
  AOI21_X1 U62 ( .B1(n3), .B2(n44), .A(n45), .ZN(OUT1[1]) );
  BUF_X2 U98 ( .A(n3), .Z(n1) );
  BUF_X1 U99 ( .A(CTRL[0]), .Z(n2) );
  INV_X1 U100 ( .A(CTRL[1]), .ZN(n3) );
endmodule


module shifter ( A, B, LOGIC_ARITH, LEFT_RIGHT, OUTPUT );
  input [31:0] A;
  input [4:0] B;
  output [31:0] OUTPUT;
  input LOGIC_ARITH, LEFT_RIGHT;
  wire   n6, n8, n9, n10, n1;
  wire   [2:0] s3;
  wire   [38:0] m0;
  wire   [38:0] m8;
  wire   [38:0] m16;
  wire   [38:0] y;

  shift_firstLevel IL ( .A(A), .sel({LOGIC_ARITH, LEFT_RIGHT}), .mask00(m0), 
        .mask08(m8), .mask16(m16) );
  shift_secondLevel IIL ( .sel(B[4:3]), .mask00(m0), .mask08(m8), .mask16(m16), 
        .Y(y) );
  shift_thirdLevel IIIL ( .sel(s3), .A(y), .Y(OUTPUT) );
  OR2_X1 U8 ( .A1(LOGIC_ARITH), .A2(LEFT_RIGHT), .ZN(n6) );
  INV_X1 U4 ( .A(B[1]), .ZN(n9) );
  INV_X1 U2 ( .A(B[2]), .ZN(n8) );
  INV_X1 U6 ( .A(B[0]), .ZN(n10) );
  INV_X1 U1 ( .A(LEFT_RIGHT), .ZN(n1) );
  AOI22_X1 U3 ( .A1(B[0]), .A2(n6), .B1(n1), .B2(n10), .ZN(s3[0]) );
  AOI22_X1 U5 ( .A1(B[1]), .A2(n6), .B1(n1), .B2(n9), .ZN(s3[1]) );
  AOI22_X1 U7 ( .A1(B[2]), .A2(n6), .B1(n1), .B2(n8), .ZN(s3[2]) );
endmodule


module comparator_M32 ( C, V, SUM, sel, sign, S );
  input [31:0] SUM;
  input [2:0] sel;
  input C, V, sign;
  output S;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24;

  XOR2_X1 U23 ( .A(n6), .B(n14), .Z(n10) );
  NOR2_X1 U22 ( .A1(sel[2]), .A2(sel[1]), .ZN(n3) );
  NOR4_X1 U20 ( .A1(SUM[1]), .A2(SUM[19]), .A3(SUM[18]), .A4(SUM[17]), .ZN(n21) );
  NOR4_X1 U19 ( .A1(SUM[23]), .A2(SUM[22]), .A3(SUM[21]), .A4(SUM[20]), .ZN(
        n22) );
  NOR4_X1 U18 ( .A1(SUM[12]), .A2(SUM[11]), .A3(SUM[10]), .A4(SUM[0]), .ZN(n23) );
  NOR4_X1 U17 ( .A1(SUM[16]), .A2(SUM[15]), .A3(SUM[14]), .A4(SUM[13]), .ZN(
        n24) );
  NAND4_X1 U16 ( .A1(n21), .A2(n22), .A3(n23), .A4(n24), .ZN(n15) );
  NOR4_X1 U15 ( .A1(SUM[6]), .A2(SUM[5]), .A3(SUM[4]), .A4(SUM[3]), .ZN(n17)
         );
  NOR4_X1 U14 ( .A1(SUM[31]), .A2(SUM[9]), .A3(SUM[8]), .A4(SUM[7]), .ZN(n18)
         );
  NOR4_X1 U13 ( .A1(SUM[27]), .A2(SUM[26]), .A3(SUM[25]), .A4(SUM[24]), .ZN(
        n19) );
  NOR4_X1 U12 ( .A1(SUM[30]), .A2(SUM[2]), .A3(SUM[29]), .A4(SUM[28]), .ZN(n20) );
  NAND4_X1 U11 ( .A1(n17), .A2(n18), .A3(n19), .A4(n20), .ZN(n16) );
  OAI21_X1 U9 ( .B1(sel[1]), .B2(sel[0]), .A(sel[2]), .ZN(n14) );
  NAND2_X1 U7 ( .A1(SUM[31]), .A2(V), .ZN(n13) );
  OAI211_X1 U6 ( .C1(V), .C2(SUM[31]), .A(n13), .B(sign), .ZN(n12) );
  OAI21_X1 U5 ( .B1(sign), .B2(C), .A(n12), .ZN(n8) );
  AOI22_X1 U4 ( .A1(n9), .A2(n10), .B1(n11), .B2(n8), .ZN(n4) );
  NOR3_X1 U3 ( .A1(n8), .A2(sel[2]), .A3(sel[1]), .ZN(n7) );
  OAI21_X1 U2 ( .B1(sel[0]), .B2(n6), .A(n7), .ZN(n5) );
  OAI21_X1 U1 ( .B1(n3), .B2(n4), .A(n5), .ZN(S) );
  OR2_X1 U21 ( .A1(sel[2]), .A2(sel[0]), .ZN(n9) );
  OR2_X1 U10 ( .A1(n15), .A2(n16), .ZN(n6) );
  INV_X1 U8 ( .A(sel[2]), .ZN(n11) );
endmodule


module simple_booth_add_ext_N16 ( Clock, Reset, sign, enable, valid, A, B, 
        A_to_add, B_to_add, sign_to_add, final_out, ACC_from_add );
  input [15:0] A;
  input [15:0] B;
  output [31:0] A_to_add;
  output [31:0] B_to_add;
  output [31:0] final_out;
  input [31:0] ACC_from_add;
  input Clock, Reset, sign, enable;
  output valid, sign_to_add;
  wire   \enc_N2_in[2] , \extend_vector[15] , \input_mux_sel[2] ,
         input_mux_sel_0, reg_enable, N23, N37, N39, N41, N43, N44, N45,
         net337982, n8, n9, n10, n11, n1, n4, n6, n7, n12, n13, n14, n15, n16,
         n17, n18, n19;
  wire   [8:0] piso_0_in;
  wire   [8:0] piso_1_in;
  wire   [8:0] piso_2_in;
  wire   [31:0] A_to_mux;
  wire   [31:0] next_accumulate;
  wire   [4:0] count;

  DFFS_X1 \count_reg[0]  ( .D(N37), .CK(net337982), .SN(n19), .Q(count[0]), 
        .QN(n13) );
  DFFR_X1 \count_reg[1]  ( .D(N39), .CK(net337982), .RN(n19), .Q(count[1]) );
  DFFR_X1 \count_reg[2]  ( .D(N41), .CK(net337982), .RN(n19), .Q(count[2]), 
        .QN(n14) );
  DFFS_X1 \count_reg[3]  ( .D(N43), .CK(net337982), .SN(n19), .Q(count[3]) );
  DFFR_X1 \count_reg[4]  ( .D(N45), .CK(net337982), .RN(n19), .Q(count[4]) );
  MUX2_X1 U51 ( .A(A_to_add[9]), .B(ACC_from_add[9]), .S(n18), .Z(final_out[9]) );
  MUX2_X1 U52 ( .A(A_to_add[8]), .B(ACC_from_add[8]), .S(n18), .Z(final_out[8]) );
  MUX2_X1 U53 ( .A(A_to_add[7]), .B(ACC_from_add[7]), .S(n18), .Z(final_out[7]) );
  MUX2_X1 U54 ( .A(A_to_add[6]), .B(ACC_from_add[6]), .S(n18), .Z(final_out[6]) );
  MUX2_X1 U55 ( .A(A_to_add[5]), .B(ACC_from_add[5]), .S(n18), .Z(final_out[5]) );
  MUX2_X1 U56 ( .A(A_to_add[4]), .B(ACC_from_add[4]), .S(n18), .Z(final_out[4]) );
  MUX2_X1 U57 ( .A(A_to_add[3]), .B(ACC_from_add[3]), .S(n18), .Z(final_out[3]) );
  MUX2_X1 U58 ( .A(A_to_add[31]), .B(ACC_from_add[31]), .S(n18), .Z(
        final_out[31]) );
  MUX2_X1 U59 ( .A(A_to_add[30]), .B(ACC_from_add[30]), .S(\input_mux_sel[2] ), 
        .Z(final_out[30]) );
  MUX2_X1 U60 ( .A(A_to_add[2]), .B(ACC_from_add[2]), .S(\input_mux_sel[2] ), 
        .Z(final_out[2]) );
  MUX2_X1 U61 ( .A(A_to_add[29]), .B(ACC_from_add[29]), .S(\input_mux_sel[2] ), 
        .Z(final_out[29]) );
  MUX2_X1 U62 ( .A(A_to_add[28]), .B(ACC_from_add[28]), .S(\input_mux_sel[2] ), 
        .Z(final_out[28]) );
  MUX2_X1 U63 ( .A(A_to_add[27]), .B(ACC_from_add[27]), .S(\input_mux_sel[2] ), 
        .Z(final_out[27]) );
  MUX2_X1 U64 ( .A(A_to_add[26]), .B(ACC_from_add[26]), .S(\input_mux_sel[2] ), 
        .Z(final_out[26]) );
  MUX2_X1 U65 ( .A(A_to_add[25]), .B(ACC_from_add[25]), .S(\input_mux_sel[2] ), 
        .Z(final_out[25]) );
  MUX2_X1 U66 ( .A(A_to_add[24]), .B(ACC_from_add[24]), .S(\input_mux_sel[2] ), 
        .Z(final_out[24]) );
  MUX2_X1 U67 ( .A(A_to_add[23]), .B(ACC_from_add[23]), .S(\input_mux_sel[2] ), 
        .Z(final_out[23]) );
  MUX2_X1 U68 ( .A(A_to_add[22]), .B(ACC_from_add[22]), .S(\input_mux_sel[2] ), 
        .Z(final_out[22]) );
  MUX2_X1 U69 ( .A(A_to_add[21]), .B(ACC_from_add[21]), .S(\input_mux_sel[2] ), 
        .Z(final_out[21]) );
  MUX2_X1 U70 ( .A(A_to_add[20]), .B(ACC_from_add[20]), .S(\input_mux_sel[2] ), 
        .Z(final_out[20]) );
  MUX2_X1 U71 ( .A(A_to_add[1]), .B(ACC_from_add[1]), .S(n18), .Z(final_out[1]) );
  MUX2_X1 U72 ( .A(A_to_add[19]), .B(ACC_from_add[19]), .S(\input_mux_sel[2] ), 
        .Z(final_out[19]) );
  MUX2_X1 U73 ( .A(A_to_add[18]), .B(ACC_from_add[18]), .S(\input_mux_sel[2] ), 
        .Z(final_out[18]) );
  MUX2_X1 U74 ( .A(A_to_add[17]), .B(ACC_from_add[17]), .S(\input_mux_sel[2] ), 
        .Z(final_out[17]) );
  MUX2_X1 U75 ( .A(A_to_add[16]), .B(ACC_from_add[16]), .S(\input_mux_sel[2] ), 
        .Z(final_out[16]) );
  MUX2_X1 U76 ( .A(A_to_add[15]), .B(ACC_from_add[15]), .S(n18), .Z(
        final_out[15]) );
  MUX2_X1 U77 ( .A(A_to_add[14]), .B(ACC_from_add[14]), .S(n18), .Z(
        final_out[14]) );
  MUX2_X1 U78 ( .A(A_to_add[13]), .B(ACC_from_add[13]), .S(\input_mux_sel[2] ), 
        .Z(final_out[13]) );
  MUX2_X1 U79 ( .A(A_to_add[12]), .B(ACC_from_add[12]), .S(\input_mux_sel[2] ), 
        .Z(final_out[12]) );
  MUX2_X1 U80 ( .A(A_to_add[11]), .B(ACC_from_add[11]), .S(\input_mux_sel[2] ), 
        .Z(final_out[11]) );
  MUX2_X1 U81 ( .A(A_to_add[10]), .B(ACC_from_add[10]), .S(\input_mux_sel[2] ), 
        .Z(final_out[10]) );
  MUX2_X1 U82 ( .A(A_to_add[0]), .B(ACC_from_add[0]), .S(\input_mux_sel[2] ), 
        .Z(final_out[0]) );
  booth_encoder_0 encod_0_0 ( .B_in({B[1:0], 1'b0}), .A_out({piso_2_in[0], 
        piso_1_in[0], piso_0_in[0]}) );
  booth_encoder_8 encod_i_1 ( .B_in(B[3:1]), .A_out({piso_2_in[1], 
        piso_1_in[1], piso_0_in[1]}) );
  booth_encoder_7 encod_i_2 ( .B_in(B[5:3]), .A_out({piso_2_in[2], 
        piso_1_in[2], piso_0_in[2]}) );
  booth_encoder_6 encod_i_3 ( .B_in(B[7:5]), .A_out({piso_2_in[3], 
        piso_1_in[3], piso_0_in[3]}) );
  booth_encoder_5 encod_i_4 ( .B_in(B[9:7]), .A_out({piso_2_in[4], 
        piso_1_in[4], piso_0_in[4]}) );
  booth_encoder_4 encod_i_5 ( .B_in(B[11:9]), .A_out({piso_2_in[5], 
        piso_1_in[5], piso_0_in[5]}) );
  booth_encoder_3 encod_i_6 ( .B_in(B[13:11]), .A_out({piso_2_in[6], 
        piso_1_in[6], piso_0_in[6]}) );
  booth_encoder_2 encod_i_7 ( .B_in(B[15:13]), .A_out({piso_2_in[7], 
        piso_1_in[7], piso_0_in[7]}) );
  booth_encoder_1 encod_i_8 ( .B_in({\enc_N2_in[2] , \enc_N2_in[2] , B[15]}), 
        .A_out({piso_2_in[8], piso_1_in[8], piso_0_in[8]}) );
  shift_N9_0 piso_0 ( .Clock(Clock), .ALOAD(n17), .D(piso_0_in), .SO(
        input_mux_sel_0) );
  shift_N9_2 piso_1 ( .Clock(Clock), .ALOAD(n17), .D(piso_1_in), .SO(
        sign_to_add) );
  shift_N9_1 piso_2 ( .Clock(Clock), .ALOAD(n17), .D(piso_2_in), .SO(
        \input_mux_sel[2] ) );
  piso_r_2_N32 A_reg ( .Clock(Clock), .ALOAD(n17), .D({\extend_vector[15] , 
        \extend_vector[15] , \extend_vector[15] , \extend_vector[15] , 
        \extend_vector[15] , \extend_vector[15] , \extend_vector[15] , 
        \extend_vector[15] , \extend_vector[15] , \extend_vector[15] , 
        \extend_vector[15] , \extend_vector[15] , \extend_vector[15] , 
        \extend_vector[15] , \extend_vector[15] , \extend_vector[15] , A}), 
        .SO(A_to_mux) );
  mux21_1 INPUTMUX ( .IN0(A_to_mux), .IN1({A_to_mux[30:0], 1'b0}), .CTRL(
        input_mux_sel_0), .OUT1(B_to_add) );
  ff32_en_SIZE32_1 ACCUMULATOR ( .D(next_accumulate), .en(reg_enable), .clk(
        Clock), .rst(Reset), .Q(A_to_add) );
  SNPS_CLOCK_GATE_HIGH_simple_booth_add_ext_N16 clk_gate_count_reg ( .CLK(
        Clock), .EN(N44), .ENCLK(net337982) );
  OR2_X1 U41 ( .A1(valid), .A2(enable), .ZN(N44) );
  INV_X1 U48 ( .A(n9), .ZN(n11) );
  OR2_X1 U4 ( .A1(n17), .A2(n18), .ZN(reg_enable) );
  AND2_X1 U12 ( .A1(n8), .A2(ACC_from_add[31]), .ZN(next_accumulate[31]) );
  AND2_X1 U24 ( .A1(n8), .A2(ACC_from_add[20]), .ZN(next_accumulate[20]) );
  AND2_X1 U20 ( .A1(n8), .A2(ACC_from_add[24]), .ZN(next_accumulate[24]) );
  AND2_X1 U16 ( .A1(n8), .A2(ACC_from_add[28]), .ZN(next_accumulate[28]) );
  AND2_X1 U19 ( .A1(n8), .A2(ACC_from_add[25]), .ZN(next_accumulate[25]) );
  AND2_X1 U23 ( .A1(n8), .A2(ACC_from_add[21]), .ZN(next_accumulate[21]) );
  AND2_X1 U15 ( .A1(n8), .A2(ACC_from_add[29]), .ZN(next_accumulate[29]) );
  AND2_X1 U22 ( .A1(n8), .A2(ACC_from_add[22]), .ZN(next_accumulate[22]) );
  AND2_X1 U18 ( .A1(n8), .A2(ACC_from_add[26]), .ZN(next_accumulate[26]) );
  AND2_X1 U17 ( .A1(n8), .A2(ACC_from_add[27]), .ZN(next_accumulate[27]) );
  AND2_X1 U21 ( .A1(n8), .A2(ACC_from_add[23]), .ZN(next_accumulate[23]) );
  AND2_X1 U13 ( .A1(n8), .A2(ACC_from_add[30]), .ZN(next_accumulate[30]) );
  AND2_X1 U28 ( .A1(n8), .A2(ACC_from_add[17]), .ZN(next_accumulate[17]) );
  AND2_X1 U27 ( .A1(n8), .A2(ACC_from_add[18]), .ZN(next_accumulate[18]) );
  AND2_X1 U26 ( .A1(n8), .A2(ACC_from_add[19]), .ZN(next_accumulate[19]) );
  AND2_X1 U29 ( .A1(n8), .A2(ACC_from_add[16]), .ZN(next_accumulate[16]) );
  AND2_X1 U32 ( .A1(n8), .A2(ACC_from_add[13]), .ZN(next_accumulate[13]) );
  AND2_X1 U31 ( .A1(n8), .A2(ACC_from_add[14]), .ZN(next_accumulate[14]) );
  AND2_X1 U30 ( .A1(n8), .A2(ACC_from_add[15]), .ZN(next_accumulate[15]) );
  AND2_X1 U33 ( .A1(n8), .A2(ACC_from_add[12]), .ZN(next_accumulate[12]) );
  AND2_X1 U6 ( .A1(n8), .A2(ACC_from_add[8]), .ZN(next_accumulate[8]) );
  AND2_X1 U35 ( .A1(n8), .A2(ACC_from_add[10]), .ZN(next_accumulate[10]) );
  AND2_X1 U5 ( .A1(n8), .A2(ACC_from_add[9]), .ZN(next_accumulate[9]) );
  AND2_X1 U34 ( .A1(n8), .A2(ACC_from_add[11]), .ZN(next_accumulate[11]) );
  AND2_X1 U7 ( .A1(n8), .A2(ACC_from_add[7]), .ZN(next_accumulate[7]) );
  AND2_X1 U11 ( .A1(n8), .A2(ACC_from_add[3]), .ZN(next_accumulate[3]) );
  AND2_X1 U8 ( .A1(n8), .A2(ACC_from_add[6]), .ZN(next_accumulate[6]) );
  AND2_X1 U10 ( .A1(n8), .A2(ACC_from_add[4]), .ZN(next_accumulate[4]) );
  AND2_X1 U9 ( .A1(n8), .A2(ACC_from_add[5]), .ZN(next_accumulate[5]) );
  AND2_X1 U14 ( .A1(n8), .A2(ACC_from_add[2]), .ZN(next_accumulate[2]) );
  AND2_X1 U25 ( .A1(n8), .A2(ACC_from_add[1]), .ZN(next_accumulate[1]) );
  AND2_X1 U36 ( .A1(n8), .A2(ACC_from_add[0]), .ZN(next_accumulate[0]) );
  AND2_X1 U38 ( .A1(sign), .A2(A[15]), .ZN(\extend_vector[15] ) );
  INV_X1 U45 ( .A(valid), .ZN(n10) );
  AND2_X1 U43 ( .A1(N23), .A2(n10), .ZN(N41) );
  OR2_X1 U46 ( .A1(valid), .A2(n13), .ZN(N37) );
  NOR3_X1 U49 ( .A1(count[1]), .A2(count[4]), .A3(count[2]), .ZN(n9) );
  NOR3_X1 U47 ( .A1(count[3]), .A2(count[0]), .A3(n11), .ZN(valid) );
  NOR2_X1 U3 ( .A1(count[3]), .A2(n16), .ZN(n1) );
  OAI21_X1 U37 ( .B1(count[4]), .B2(n1), .A(n10), .ZN(n4) );
  AOI21_X1 U39 ( .B1(count[4]), .B2(n1), .A(n4), .ZN(N45) );
  AOI21_X1 U40 ( .B1(n16), .B2(count[3]), .A(valid), .ZN(n6) );
  OAI21_X1 U42 ( .B1(n16), .B2(count[3]), .A(n6), .ZN(N43) );
  INV_X1 U44 ( .A(n10), .ZN(n7) );
  AOI21_X1 U50 ( .B1(count[1]), .B2(count[0]), .A(n15), .ZN(n12) );
  NOR2_X1 U83 ( .A1(n12), .A2(n7), .ZN(N39) );
  BUF_X1 U84 ( .A(\input_mux_sel[2] ), .Z(n18) );
  NOR2_X1 U85 ( .A1(count[0]), .A2(count[1]), .ZN(n15) );
  OR3_X1 U86 ( .A1(count[2]), .A2(count[0]), .A3(count[1]), .ZN(n16) );
  OAI21_X1 U87 ( .B1(n15), .B2(n14), .A(n16), .ZN(N23) );
  INV_X1 U88 ( .A(Reset), .ZN(n19) );
  AND2_X1 U89 ( .A1(sign), .A2(B[15]), .ZN(\enc_N2_in[2] ) );
  INV_X4 U90 ( .A(n8), .ZN(n17) );
  NAND3_X2 U91 ( .A1(n9), .A2(count[3]), .A3(count[0]), .ZN(n8) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ff32_en_SIZE13 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net338015, net338017, net338018, net338021;
  assign net338015 = CLK;
  assign ENCLK = net338017;
  assign net338018 = EN;

  DLL_X1 latch ( .D(net338018), .GN(net338015), .Q(net338021) );
  AND2_X1 main_gate ( .A1(net338021), .A2(net338015), .ZN(net338017) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ff32_en_SIZE5_0 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net338000, net338002, net338003, net338006;
  assign net338000 = CLK;
  assign ENCLK = net338002;
  assign net338003 = EN;

  DLL_X1 latch ( .D(net338003), .GN(net338000), .Q(net338006) );
  AND2_X1 main_gate ( .A1(net338006), .A2(net338000), .ZN(net338002) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ff32_en_SIZE32_0 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net337985, net337987, net337988, net337991;
  assign net337985 = CLK;
  assign ENCLK = net337987;
  assign net337988 = EN;

  DLL_X1 latch ( .D(net337988), .GN(net337985), .Q(net337991) );
  AND2_X1 main_gate ( .A1(net337991), .A2(net337985), .ZN(net337987) );
endmodule


module sum_gen_N32_0 ( A, B, Cin, S );
  input [31:0] A;
  input [31:0] B;
  input [8:0] Cin;
  output [31:0] S;


  carry_sel_gen_N4_0 csel_N_0 ( .A(A[3:0]), .B(B[3:0]), .Ci(1'b0), .S(S[3:0])
         );
  carry_sel_gen_N4_15 csel_N_1 ( .A(A[7:4]), .B(B[7:4]), .Ci(Cin[1]), .S(
        S[7:4]) );
  carry_sel_gen_N4_14 csel_N_2 ( .A(A[11:8]), .B(B[11:8]), .Ci(Cin[2]), .S(
        S[11:8]) );
  carry_sel_gen_N4_13 csel_N_3 ( .A(A[15:12]), .B(B[15:12]), .Ci(Cin[3]), .S(
        S[15:12]) );
  carry_sel_gen_N4_12 csel_N_4 ( .A(A[19:16]), .B(B[19:16]), .Ci(Cin[4]), .S(
        S[19:16]) );
  carry_sel_gen_N4_11 csel_N_5 ( .A(A[23:20]), .B(B[23:20]), .Ci(Cin[5]), .S(
        S[23:20]) );
  carry_sel_gen_N4_10 csel_N_6 ( .A(A[27:24]), .B(B[27:24]), .Ci(Cin[6]), .S(
        S[27:24]) );
  carry_sel_gen_N4_9 csel_N_7 ( .A(A[31:28]), .B(B[31:28]), .Ci(Cin[7]), .S(
        S[31:28]) );
endmodule


module carry_tree_N32_logN5_0 ( A, B, Cin, Cout );
  input [31:0] A;
  input [31:0] B;
  output [7:0] Cout;
  input Cin;
  wire   \magic_pro[0] , \pg_1[13][1] , \pg_1[13][0] , \pg_1[12][1] ,
         \pg_1[12][0] , \pg_1[11][1] , \pg_1[11][0] , \pg_1[10][1] ,
         \pg_1[10][0] , \pg_1[9][1] , \pg_1[9][0] , \pg_1[8][1] , \pg_1[8][0] ,
         \pg_1[7][1] , \pg_1[7][0] , \pg_1[6][1] , \pg_1[6][0] , \pg_1[5][1] ,
         \pg_1[5][0] , \pg_1[4][1] , \pg_1[4][0] , \pg_1[3][1] , \pg_1[3][0] ,
         \pg_1[2][1] , \pg_1[2][0] , \pg_1[1][1] , \pg_1[1][0] , \pg_1[0][0] ,
         \pg_n[4][6][1] , \pg_n[4][6][0] , \pg_n[3][5][1] , \pg_n[3][5][0] ,
         \pg_n[3][3][1] , \pg_n[3][3][0] , \pg_n[2][6][1] , \pg_n[2][6][0] ,
         \pg_n[2][5][1] , \pg_n[2][5][0] , \pg_n[2][4][1] , \pg_n[2][4][0] ,
         \pg_n[2][3][1] , \pg_n[2][3][0] , \pg_n[2][2][1] , \pg_n[2][2][0] ,
         \pg_n[2][1][1] , \pg_n[2][1][0] ;
  wire   [31:1] p_net;
  wire   [31:0] g_net;

  pg_net_0 pg_net_x_1 ( .a(A[1]), .b(B[1]), .g_out(g_net[1]), .p_out(p_net[1])
         );
  pg_net_63 pg_net_x_2 ( .a(A[2]), .b(B[2]), .g_out(g_net[2]), .p_out(p_net[2]) );
  pg_net_62 pg_net_x_3 ( .a(A[3]), .b(B[3]), .g_out(g_net[3]), .p_out(p_net[3]) );
  pg_net_61 pg_net_x_4 ( .a(A[4]), .b(B[4]), .g_out(g_net[4]), .p_out(p_net[4]) );
  pg_net_60 pg_net_x_5 ( .a(A[5]), .b(B[5]), .g_out(g_net[5]), .p_out(p_net[5]) );
  pg_net_59 pg_net_x_6 ( .a(A[6]), .b(B[6]), .g_out(g_net[6]), .p_out(p_net[6]) );
  pg_net_58 pg_net_x_7 ( .a(A[7]), .b(B[7]), .g_out(g_net[7]), .p_out(p_net[7]) );
  pg_net_57 pg_net_x_8 ( .a(A[8]), .b(B[8]), .g_out(g_net[8]), .p_out(p_net[8]) );
  pg_net_56 pg_net_x_9 ( .a(A[9]), .b(B[9]), .g_out(g_net[9]), .p_out(p_net[9]) );
  pg_net_55 pg_net_x_10 ( .a(A[10]), .b(B[10]), .g_out(g_net[10]), .p_out(
        p_net[10]) );
  pg_net_54 pg_net_x_11 ( .a(A[11]), .b(B[11]), .g_out(g_net[11]), .p_out(
        p_net[11]) );
  pg_net_53 pg_net_x_12 ( .a(A[12]), .b(B[12]), .g_out(g_net[12]), .p_out(
        p_net[12]) );
  pg_net_52 pg_net_x_13 ( .a(A[13]), .b(B[13]), .g_out(g_net[13]), .p_out(
        p_net[13]) );
  pg_net_51 pg_net_x_14 ( .a(A[14]), .b(B[14]), .g_out(g_net[14]), .p_out(
        p_net[14]) );
  pg_net_50 pg_net_x_15 ( .a(A[15]), .b(B[15]), .g_out(g_net[15]), .p_out(
        p_net[15]) );
  pg_net_49 pg_net_x_16 ( .a(A[16]), .b(B[16]), .g_out(g_net[16]), .p_out(
        p_net[16]) );
  pg_net_48 pg_net_x_17 ( .a(A[17]), .b(B[17]), .g_out(g_net[17]), .p_out(
        p_net[17]) );
  pg_net_47 pg_net_x_18 ( .a(A[18]), .b(B[18]), .g_out(g_net[18]), .p_out(
        p_net[18]) );
  pg_net_46 pg_net_x_19 ( .a(A[19]), .b(B[19]), .g_out(g_net[19]), .p_out(
        p_net[19]) );
  pg_net_45 pg_net_x_20 ( .a(A[20]), .b(B[20]), .g_out(g_net[20]), .p_out(
        p_net[20]) );
  pg_net_44 pg_net_x_21 ( .a(A[21]), .b(B[21]), .g_out(g_net[21]), .p_out(
        p_net[21]) );
  pg_net_43 pg_net_x_22 ( .a(A[22]), .b(B[22]), .g_out(g_net[22]), .p_out(
        p_net[22]) );
  pg_net_42 pg_net_x_23 ( .a(A[23]), .b(B[23]), .g_out(g_net[23]), .p_out(
        p_net[23]) );
  pg_net_41 pg_net_x_24 ( .a(A[24]), .b(B[24]), .g_out(g_net[24]), .p_out(
        p_net[24]) );
  pg_net_40 pg_net_x_25 ( .a(A[25]), .b(B[25]), .g_out(g_net[25]), .p_out(
        p_net[25]) );
  pg_net_39 pg_net_x_26 ( .a(A[26]), .b(B[26]), .g_out(g_net[26]), .p_out(
        p_net[26]) );
  pg_net_38 pg_net_x_27 ( .a(A[27]), .b(B[27]), .g_out(g_net[27]), .p_out(
        p_net[27]) );
  pg_net_33 pg_net_0_MAGIC ( .a(A[0]), .b(B[0]), .g_out(\magic_pro[0] ) );
  g_0 xG_0_0_MAGIC ( .g(\magic_pro[0] ), .p(1'b0), .g_prec(1'b0), .g_out(
        g_net[0]) );
  g_19 xG_1_0 ( .g(g_net[1]), .p(p_net[1]), .g_prec(g_net[0]), .g_out(
        \pg_1[0][0] ) );
  pg_0 xPG_1_1 ( .g(g_net[3]), .p(p_net[3]), .g_prec(g_net[2]), .p_prec(
        p_net[2]), .g_out(\pg_1[1][0] ), .p_out(\pg_1[1][1] ) );
  pg_53 xPG_1_2 ( .g(g_net[5]), .p(p_net[5]), .g_prec(g_net[4]), .p_prec(
        p_net[4]), .g_out(\pg_1[2][0] ), .p_out(\pg_1[2][1] ) );
  pg_52 xPG_1_3 ( .g(g_net[7]), .p(p_net[7]), .g_prec(g_net[6]), .p_prec(
        p_net[6]), .g_out(\pg_1[3][0] ), .p_out(\pg_1[3][1] ) );
  pg_51 xPG_1_4 ( .g(g_net[9]), .p(p_net[9]), .g_prec(g_net[8]), .p_prec(
        p_net[8]), .g_out(\pg_1[4][0] ), .p_out(\pg_1[4][1] ) );
  pg_50 xPG_1_5 ( .g(g_net[11]), .p(p_net[11]), .g_prec(g_net[10]), .p_prec(
        p_net[10]), .g_out(\pg_1[5][0] ), .p_out(\pg_1[5][1] ) );
  pg_49 xPG_1_6 ( .g(g_net[13]), .p(p_net[13]), .g_prec(g_net[12]), .p_prec(
        p_net[12]), .g_out(\pg_1[6][0] ), .p_out(\pg_1[6][1] ) );
  pg_48 xPG_1_7 ( .g(g_net[15]), .p(p_net[15]), .g_prec(g_net[14]), .p_prec(
        p_net[14]), .g_out(\pg_1[7][0] ), .p_out(\pg_1[7][1] ) );
  pg_47 xPG_1_8 ( .g(g_net[17]), .p(p_net[17]), .g_prec(g_net[16]), .p_prec(
        p_net[16]), .g_out(\pg_1[8][0] ), .p_out(\pg_1[8][1] ) );
  pg_46 xPG_1_9 ( .g(g_net[19]), .p(p_net[19]), .g_prec(g_net[18]), .p_prec(
        p_net[18]), .g_out(\pg_1[9][0] ), .p_out(\pg_1[9][1] ) );
  pg_45 xPG_1_10 ( .g(g_net[21]), .p(p_net[21]), .g_prec(g_net[20]), .p_prec(
        p_net[20]), .g_out(\pg_1[10][0] ), .p_out(\pg_1[10][1] ) );
  pg_44 xPG_1_11 ( .g(g_net[23]), .p(p_net[23]), .g_prec(g_net[22]), .p_prec(
        p_net[22]), .g_out(\pg_1[11][0] ), .p_out(\pg_1[11][1] ) );
  pg_43 xPG_1_12 ( .g(g_net[25]), .p(p_net[25]), .g_prec(g_net[24]), .p_prec(
        p_net[24]), .g_out(\pg_1[12][0] ), .p_out(\pg_1[12][1] ) );
  pg_42 xPG_1_13 ( .g(g_net[27]), .p(p_net[27]), .g_prec(g_net[26]), .p_prec(
        p_net[26]), .g_out(\pg_1[13][0] ), .p_out(\pg_1[13][1] ) );
  g_18 xG_2_0 ( .g(\pg_1[1][0] ), .p(\pg_1[1][1] ), .g_prec(\pg_1[0][0] ), 
        .g_out(Cout[0]) );
  pg_39 xPG_2_1 ( .g(\pg_1[3][0] ), .p(\pg_1[3][1] ), .g_prec(\pg_1[2][0] ), 
        .p_prec(\pg_1[2][1] ), .g_out(\pg_n[2][1][0] ), .p_out(\pg_n[2][1][1] ) );
  pg_38 xPG_2_2 ( .g(\pg_1[5][0] ), .p(\pg_1[5][1] ), .g_prec(\pg_1[4][0] ), 
        .p_prec(\pg_1[4][1] ), .g_out(\pg_n[2][2][0] ), .p_out(\pg_n[2][2][1] ) );
  pg_37 xPG_2_3 ( .g(\pg_1[7][0] ), .p(\pg_1[7][1] ), .g_prec(\pg_1[6][0] ), 
        .p_prec(\pg_1[6][1] ), .g_out(\pg_n[2][3][0] ), .p_out(\pg_n[2][3][1] ) );
  pg_36 xPG_2_4 ( .g(\pg_1[9][0] ), .p(\pg_1[9][1] ), .g_prec(\pg_1[8][0] ), 
        .p_prec(\pg_1[8][1] ), .g_out(\pg_n[2][4][0] ), .p_out(\pg_n[2][4][1] ) );
  pg_35 xPG_2_5 ( .g(\pg_1[11][0] ), .p(\pg_1[11][1] ), .g_prec(\pg_1[10][0] ), 
        .p_prec(\pg_1[10][1] ), .g_out(\pg_n[2][5][0] ), .p_out(
        \pg_n[2][5][1] ) );
  pg_34 xPG_2_6 ( .g(\pg_1[13][0] ), .p(\pg_1[13][1] ), .g_prec(\pg_1[12][0] ), 
        .p_prec(\pg_1[12][1] ), .g_out(\pg_n[2][6][0] ), .p_out(
        \pg_n[2][6][1] ) );
  g_17 xG_3_1 ( .g(\pg_n[2][1][0] ), .p(\pg_n[2][1][1] ), .g_prec(Cout[0]), 
        .g_out(Cout[1]) );
  g_16 xG_4_2 ( .g(\pg_n[2][2][0] ), .p(\pg_n[2][2][1] ), .g_prec(Cout[1]), 
        .g_out(Cout[2]) );
  g_15 xG_4_3 ( .g(\pg_n[3][3][0] ), .p(\pg_n[3][3][1] ), .g_prec(Cout[1]), 
        .g_out(Cout[3]) );
  g_14 xG_5_4 ( .g(\pg_n[2][4][0] ), .p(\pg_n[2][4][1] ), .g_prec(Cout[3]), 
        .g_out(Cout[4]) );
  g_13 xG_5_5 ( .g(\pg_n[3][5][0] ), .p(\pg_n[3][5][1] ), .g_prec(Cout[3]), 
        .g_out(Cout[5]) );
  g_12 xG_5_6 ( .g(\pg_n[4][6][0] ), .p(\pg_n[4][6][1] ), .g_prec(Cout[3]), 
        .g_out(Cout[6]) );
  pg_32 xPG_3_3 ( .g(\pg_n[2][3][0] ), .p(\pg_n[2][3][1] ), .g_prec(
        \pg_n[2][2][0] ), .p_prec(\pg_n[2][2][1] ), .g_out(\pg_n[3][3][0] ), 
        .p_out(\pg_n[3][3][1] ) );
  pg_31 xPG_3_5 ( .g(\pg_n[2][5][0] ), .p(\pg_n[2][5][1] ), .g_prec(
        \pg_n[2][4][0] ), .p_prec(\pg_n[2][4][1] ), .g_out(\pg_n[3][5][0] ), 
        .p_out(\pg_n[3][5][1] ) );
  pg_29 xPG_4_6 ( .g(\pg_n[2][6][0] ), .p(\pg_n[2][6][1] ), .g_prec(
        \pg_n[3][5][0] ), .p_prec(\pg_n[3][5][1] ), .g_out(\pg_n[4][6][0] ), 
        .p_out(\pg_n[4][6][1] ) );
endmodule


module xor_gen_N32_0 ( A, B, S );
  input [31:0] A;
  output [31:0] S;
  input B;

  assign S[31] = A[31];
  assign S[30] = A[30];
  assign S[29] = A[29];
  assign S[28] = A[28];
  assign S[27] = A[27];
  assign S[26] = A[26];
  assign S[25] = A[25];
  assign S[24] = A[24];
  assign S[23] = A[23];
  assign S[22] = A[22];
  assign S[21] = A[21];
  assign S[20] = A[20];
  assign S[19] = A[19];
  assign S[18] = A[18];
  assign S[17] = A[17];
  assign S[16] = A[16];
  assign S[15] = A[15];
  assign S[14] = A[14];
  assign S[13] = A[13];
  assign S[12] = A[12];
  assign S[11] = A[11];
  assign S[10] = A[10];
  assign S[9] = A[9];
  assign S[8] = A[8];
  assign S[7] = A[7];
  assign S[6] = A[6];
  assign S[5] = A[5];
  assign S[4] = A[4];
  assign S[3] = A[3];
  assign S[2] = A[2];
  assign S[1] = A[1];
  assign S[0] = A[0];

endmodule


module SNPS_CLOCK_GATE_HIGH_ff32_en_IR ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net338230, net338232, net338233, net338236;
  assign net338230 = CLK;
  assign ENCLK = net338232;
  assign net338233 = EN;

  DLL_X1 latch ( .D(net338233), .GN(net338230), .Q(net338236) );
  AND2_X1 main_gate ( .A1(net338236), .A2(net338230), .ZN(net338232) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ff32_en_0 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net338245, net338247, net338248, net338251;
  assign net338245 = CLK;
  assign ENCLK = net338247;
  assign net338248 = EN;

  DLL_X1 latch ( .D(net338248), .GN(net338245), .Q(net338251) );
  AND2_X1 main_gate ( .A1(net338251), .A2(net338245), .ZN(net338247) );
endmodule


module ff32_SIZE5 ( D, clk, rst, Q );
  input [4:0] D;
  output [4:0] Q;
  input clk, rst;
  wire   n5;

  DFFR_X1 \Q_reg[4]  ( .D(D[4]), .CK(clk), .RN(n5), .Q(Q[4]) );
  DFFR_X1 \Q_reg[3]  ( .D(D[3]), .CK(clk), .RN(n5), .Q(Q[3]) );
  DFFR_X1 \Q_reg[2]  ( .D(D[2]), .CK(clk), .RN(n5), .Q(Q[2]) );
  DFFR_X1 \Q_reg[1]  ( .D(D[1]), .CK(clk), .RN(n5), .Q(Q[1]) );
  DFFR_X1 \Q_reg[0]  ( .D(D[0]), .CK(clk), .RN(n5), .Q(Q[0]) );
  INV_X1 U3 ( .A(rst), .ZN(n5) );
endmodule


module ff32_SIZE32 ( D, clk, rst, Q );
  input [31:0] D;
  output [31:0] Q;
  input clk, rst;
  wire   n32;

  DFFR_X1 \Q_reg[31]  ( .D(D[31]), .CK(clk), .RN(n32), .Q(Q[31]) );
  DFFR_X1 \Q_reg[30]  ( .D(D[30]), .CK(clk), .RN(n32), .Q(Q[30]) );
  DFFR_X1 \Q_reg[29]  ( .D(D[29]), .CK(clk), .RN(n32), .Q(Q[29]) );
  DFFR_X1 \Q_reg[28]  ( .D(D[28]), .CK(clk), .RN(n32), .Q(Q[28]) );
  DFFR_X1 \Q_reg[27]  ( .D(D[27]), .CK(clk), .RN(n32), .Q(Q[27]) );
  DFFR_X1 \Q_reg[26]  ( .D(D[26]), .CK(clk), .RN(n32), .Q(Q[26]) );
  DFFR_X1 \Q_reg[25]  ( .D(D[25]), .CK(clk), .RN(n32), .Q(Q[25]) );
  DFFR_X1 \Q_reg[24]  ( .D(D[24]), .CK(clk), .RN(n32), .Q(Q[24]) );
  DFFR_X1 \Q_reg[23]  ( .D(D[23]), .CK(clk), .RN(n32), .Q(Q[23]) );
  DFFR_X1 \Q_reg[22]  ( .D(D[22]), .CK(clk), .RN(n32), .Q(Q[22]) );
  DFFR_X1 \Q_reg[21]  ( .D(D[21]), .CK(clk), .RN(n32), .Q(Q[21]) );
  DFFR_X1 \Q_reg[20]  ( .D(D[20]), .CK(clk), .RN(n32), .Q(Q[20]) );
  DFFR_X1 \Q_reg[19]  ( .D(D[19]), .CK(clk), .RN(n32), .Q(Q[19]) );
  DFFR_X1 \Q_reg[18]  ( .D(D[18]), .CK(clk), .RN(n32), .Q(Q[18]) );
  DFFR_X1 \Q_reg[17]  ( .D(D[17]), .CK(clk), .RN(n32), .Q(Q[17]) );
  DFFR_X1 \Q_reg[16]  ( .D(D[16]), .CK(clk), .RN(n32), .Q(Q[16]) );
  DFFR_X1 \Q_reg[15]  ( .D(D[15]), .CK(clk), .RN(n32), .Q(Q[15]) );
  DFFR_X1 \Q_reg[14]  ( .D(D[14]), .CK(clk), .RN(n32), .Q(Q[14]) );
  DFFR_X1 \Q_reg[13]  ( .D(D[13]), .CK(clk), .RN(n32), .Q(Q[13]) );
  DFFR_X1 \Q_reg[12]  ( .D(D[12]), .CK(clk), .RN(n32), .Q(Q[12]) );
  DFFR_X1 \Q_reg[11]  ( .D(D[11]), .CK(clk), .RN(n32), .Q(Q[11]) );
  DFFR_X1 \Q_reg[10]  ( .D(D[10]), .CK(clk), .RN(n32), .Q(Q[10]) );
  DFFR_X1 \Q_reg[9]  ( .D(D[9]), .CK(clk), .RN(n32), .Q(Q[9]) );
  DFFR_X1 \Q_reg[8]  ( .D(D[8]), .CK(clk), .RN(n32), .Q(Q[8]) );
  DFFR_X1 \Q_reg[7]  ( .D(D[7]), .CK(clk), .RN(n32), .Q(Q[7]) );
  DFFR_X1 \Q_reg[6]  ( .D(D[6]), .CK(clk), .RN(n32), .Q(Q[6]) );
  DFFR_X1 \Q_reg[5]  ( .D(D[5]), .CK(clk), .RN(n32), .Q(Q[5]) );
  DFFR_X1 \Q_reg[4]  ( .D(D[4]), .CK(clk), .RN(n32), .Q(Q[4]) );
  DFFR_X1 \Q_reg[3]  ( .D(D[3]), .CK(clk), .RN(n32), .Q(Q[3]) );
  DFFR_X1 \Q_reg[2]  ( .D(D[2]), .CK(clk), .RN(n32), .Q(Q[2]) );
  DFFR_X1 \Q_reg[1]  ( .D(D[1]), .CK(clk), .RN(n32), .Q(Q[1]) );
  DFFR_X1 \Q_reg[0]  ( .D(D[0]), .CK(clk), .RN(n32), .Q(Q[0]) );
  INV_X2 U3 ( .A(rst), .ZN(n32) );
endmodule


module mux41_MUX_SIZE5 ( IN0, IN1, IN2, IN3, CTRL, OUT1 );
  input [4:0] IN0;
  input [4:0] IN1;
  input [4:0] IN2;
  input [4:0] IN3;
  input [1:0] CTRL;
  output [4:0] OUT1;
  wire   n3, n4, n5, n6, n7, n9, n10, n11, n12, n13, n14, n15, n16, n17;

  NAND2_X1 U1 ( .A1(n3), .A2(n4), .ZN(OUT1[4]) );
  NAND2_X1 U4 ( .A1(n9), .A2(n10), .ZN(OUT1[3]) );
  NAND2_X1 U7 ( .A1(n11), .A2(n12), .ZN(OUT1[2]) );
  AOI22_X1 U17 ( .A1(n6), .A2(IN2[0]), .B1(n7), .B2(IN1[0]), .ZN(n15) );
  NOR2_X1 U19 ( .A1(CTRL[0]), .A2(n17), .ZN(n6) );
  NAND2_X1 U10 ( .A1(n13), .A2(n14), .ZN(OUT1[1]) );
  NAND2_X1 U13 ( .A1(n15), .A2(n16), .ZN(OUT1[0]) );
  INV_X1 U20 ( .A(CTRL[1]), .ZN(n17) );
  AND2_X1 U18 ( .A1(n17), .A2(CTRL[0]), .ZN(n7) );
  AND2_X1 U16 ( .A1(CTRL[0]), .A2(CTRL[1]), .ZN(n5) );
  INV_X1 U2 ( .A(n5), .ZN(n16) );
  AOI21_X1 U3 ( .B1(n6), .B2(IN2[1]), .A(n5), .ZN(n14) );
  NAND2_X1 U5 ( .A1(n7), .A2(IN1[1]), .ZN(n13) );
  AOI21_X1 U6 ( .B1(n6), .B2(IN2[2]), .A(n5), .ZN(n12) );
  NAND2_X1 U8 ( .A1(n7), .A2(IN1[2]), .ZN(n11) );
  AOI21_X1 U9 ( .B1(n6), .B2(IN2[3]), .A(n5), .ZN(n10) );
  NAND2_X1 U11 ( .A1(n7), .A2(IN1[3]), .ZN(n9) );
  AOI21_X1 U12 ( .B1(n6), .B2(IN2[4]), .A(n5), .ZN(n4) );
  NAND2_X1 U14 ( .A1(n7), .A2(IN1[4]), .ZN(n3) );
endmodule


module real_alu_DATA_SIZE32 ( IN1, IN2, ALUW_i, DOUT, stall_o, Clock, Reset );
  input [31:0] IN1;
  input [31:0] IN2;
  input [12:0] ALUW_i;
  output [31:0] DOUT;
  input Clock, Reset;
  output stall_o;
  wire   mux_sign, sign_booth_to_add, valid_from_booth, carry_from_adder,
         overflow, comp_out, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n1, n2,
         n3, n4, n5;
  wire   [31:0] mux_A;
  wire   [31:0] A_booth_to_add;
  wire   [31:0] mux_B;
  wire   [31:0] B_booth_to_add;
  wire   [31:0] mult_out;
  wire   [31:0] sum_out;
  wire   [31:0] shift_out;
  wire   [31:0] lu_out;

  OAI33_X1 U111 ( .A1(IN2[31]), .A2(sum_out[31]), .A3(n10), .B1(n11), .B2(n12), 
        .B3(IN1[31]), .ZN(overflow) );
  MUX2_X1 U113 ( .A(B_booth_to_add[9]), .B(IN2[9]), .S(n5), .Z(mux_B[9]) );
  MUX2_X1 U114 ( .A(B_booth_to_add[8]), .B(IN2[8]), .S(n5), .Z(mux_B[8]) );
  MUX2_X1 U115 ( .A(B_booth_to_add[7]), .B(IN2[7]), .S(n5), .Z(mux_B[7]) );
  MUX2_X1 U116 ( .A(B_booth_to_add[6]), .B(IN2[6]), .S(n5), .Z(mux_B[6]) );
  MUX2_X1 U117 ( .A(B_booth_to_add[5]), .B(IN2[5]), .S(n5), .Z(mux_B[5]) );
  MUX2_X1 U118 ( .A(B_booth_to_add[4]), .B(IN2[4]), .S(n5), .Z(mux_B[4]) );
  MUX2_X1 U119 ( .A(B_booth_to_add[3]), .B(IN2[3]), .S(n5), .Z(mux_B[3]) );
  MUX2_X1 U120 ( .A(B_booth_to_add[31]), .B(IN2[31]), .S(n5), .Z(mux_B[31]) );
  MUX2_X1 U121 ( .A(B_booth_to_add[30]), .B(IN2[30]), .S(n5), .Z(mux_B[30]) );
  MUX2_X1 U122 ( .A(B_booth_to_add[2]), .B(IN2[2]), .S(n5), .Z(mux_B[2]) );
  MUX2_X1 U123 ( .A(B_booth_to_add[29]), .B(IN2[29]), .S(n5), .Z(mux_B[29]) );
  MUX2_X1 U124 ( .A(B_booth_to_add[28]), .B(IN2[28]), .S(n5), .Z(mux_B[28]) );
  MUX2_X1 U125 ( .A(B_booth_to_add[27]), .B(IN2[27]), .S(n4), .Z(mux_B[27]) );
  MUX2_X1 U126 ( .A(B_booth_to_add[26]), .B(IN2[26]), .S(n4), .Z(mux_B[26]) );
  MUX2_X1 U127 ( .A(B_booth_to_add[25]), .B(IN2[25]), .S(n4), .Z(mux_B[25]) );
  MUX2_X1 U128 ( .A(B_booth_to_add[24]), .B(IN2[24]), .S(n4), .Z(mux_B[24]) );
  MUX2_X1 U129 ( .A(B_booth_to_add[23]), .B(IN2[23]), .S(n4), .Z(mux_B[23]) );
  MUX2_X1 U130 ( .A(B_booth_to_add[22]), .B(IN2[22]), .S(n4), .Z(mux_B[22]) );
  MUX2_X1 U131 ( .A(B_booth_to_add[21]), .B(IN2[21]), .S(n4), .Z(mux_B[21]) );
  MUX2_X1 U132 ( .A(B_booth_to_add[20]), .B(IN2[20]), .S(n4), .Z(mux_B[20]) );
  MUX2_X1 U133 ( .A(B_booth_to_add[1]), .B(IN2[1]), .S(n4), .Z(mux_B[1]) );
  MUX2_X1 U134 ( .A(B_booth_to_add[19]), .B(IN2[19]), .S(n4), .Z(mux_B[19]) );
  MUX2_X1 U135 ( .A(B_booth_to_add[18]), .B(IN2[18]), .S(n4), .Z(mux_B[18]) );
  MUX2_X1 U136 ( .A(B_booth_to_add[17]), .B(IN2[17]), .S(n4), .Z(mux_B[17]) );
  MUX2_X1 U137 ( .A(B_booth_to_add[16]), .B(IN2[16]), .S(n4), .Z(mux_B[16]) );
  MUX2_X1 U138 ( .A(B_booth_to_add[15]), .B(IN2[15]), .S(n4), .Z(mux_B[15]) );
  MUX2_X1 U139 ( .A(B_booth_to_add[14]), .B(IN2[14]), .S(n4), .Z(mux_B[14]) );
  MUX2_X1 U140 ( .A(B_booth_to_add[13]), .B(IN2[13]), .S(n4), .Z(mux_B[13]) );
  MUX2_X1 U141 ( .A(B_booth_to_add[12]), .B(IN2[12]), .S(n4), .Z(mux_B[12]) );
  MUX2_X1 U142 ( .A(B_booth_to_add[11]), .B(IN2[11]), .S(n4), .Z(mux_B[11]) );
  MUX2_X1 U143 ( .A(B_booth_to_add[10]), .B(IN2[10]), .S(n4), .Z(mux_B[10]) );
  MUX2_X1 U144 ( .A(B_booth_to_add[0]), .B(IN2[0]), .S(n4), .Z(mux_B[0]) );
  MUX2_X1 U145 ( .A(A_booth_to_add[9]), .B(IN1[9]), .S(n4), .Z(mux_A[9]) );
  MUX2_X1 U146 ( .A(A_booth_to_add[8]), .B(IN1[8]), .S(n4), .Z(mux_A[8]) );
  MUX2_X1 U147 ( .A(A_booth_to_add[7]), .B(IN1[7]), .S(n4), .Z(mux_A[7]) );
  MUX2_X1 U148 ( .A(A_booth_to_add[6]), .B(IN1[6]), .S(n4), .Z(mux_A[6]) );
  MUX2_X1 U149 ( .A(A_booth_to_add[5]), .B(IN1[5]), .S(n4), .Z(mux_A[5]) );
  MUX2_X1 U150 ( .A(A_booth_to_add[4]), .B(IN1[4]), .S(n4), .Z(mux_A[4]) );
  MUX2_X1 U151 ( .A(A_booth_to_add[3]), .B(IN1[3]), .S(n4), .Z(mux_A[3]) );
  MUX2_X1 U152 ( .A(A_booth_to_add[31]), .B(IN1[31]), .S(n4), .Z(mux_A[31]) );
  MUX2_X1 U153 ( .A(A_booth_to_add[30]), .B(IN1[30]), .S(n4), .Z(mux_A[30]) );
  MUX2_X1 U154 ( .A(A_booth_to_add[2]), .B(IN1[2]), .S(n4), .Z(mux_A[2]) );
  MUX2_X1 U155 ( .A(A_booth_to_add[29]), .B(IN1[29]), .S(n4), .Z(mux_A[29]) );
  MUX2_X1 U156 ( .A(A_booth_to_add[28]), .B(IN1[28]), .S(n4), .Z(mux_A[28]) );
  MUX2_X1 U157 ( .A(A_booth_to_add[27]), .B(IN1[27]), .S(n4), .Z(mux_A[27]) );
  MUX2_X1 U158 ( .A(A_booth_to_add[26]), .B(IN1[26]), .S(n4), .Z(mux_A[26]) );
  MUX2_X1 U159 ( .A(A_booth_to_add[25]), .B(IN1[25]), .S(n4), .Z(mux_A[25]) );
  MUX2_X1 U160 ( .A(A_booth_to_add[24]), .B(IN1[24]), .S(n4), .Z(mux_A[24]) );
  MUX2_X1 U161 ( .A(A_booth_to_add[23]), .B(IN1[23]), .S(n9), .Z(mux_A[23]) );
  MUX2_X1 U162 ( .A(A_booth_to_add[22]), .B(IN1[22]), .S(n9), .Z(mux_A[22]) );
  MUX2_X1 U163 ( .A(A_booth_to_add[21]), .B(IN1[21]), .S(n9), .Z(mux_A[21]) );
  MUX2_X1 U164 ( .A(A_booth_to_add[20]), .B(IN1[20]), .S(n9), .Z(mux_A[20]) );
  MUX2_X1 U165 ( .A(A_booth_to_add[1]), .B(IN1[1]), .S(n9), .Z(mux_A[1]) );
  MUX2_X1 U166 ( .A(A_booth_to_add[19]), .B(IN1[19]), .S(n9), .Z(mux_A[19]) );
  MUX2_X1 U167 ( .A(A_booth_to_add[18]), .B(IN1[18]), .S(n9), .Z(mux_A[18]) );
  MUX2_X1 U168 ( .A(A_booth_to_add[17]), .B(IN1[17]), .S(n9), .Z(mux_A[17]) );
  MUX2_X1 U169 ( .A(A_booth_to_add[16]), .B(IN1[16]), .S(n9), .Z(mux_A[16]) );
  MUX2_X1 U170 ( .A(A_booth_to_add[15]), .B(IN1[15]), .S(n9), .Z(mux_A[15]) );
  MUX2_X1 U171 ( .A(A_booth_to_add[14]), .B(IN1[14]), .S(n9), .Z(mux_A[14]) );
  MUX2_X1 U172 ( .A(A_booth_to_add[13]), .B(IN1[13]), .S(n9), .Z(mux_A[13]) );
  MUX2_X1 U173 ( .A(A_booth_to_add[12]), .B(IN1[12]), .S(n9), .Z(mux_A[12]) );
  MUX2_X1 U174 ( .A(A_booth_to_add[11]), .B(IN1[11]), .S(n9), .Z(mux_A[11]) );
  MUX2_X1 U175 ( .A(A_booth_to_add[10]), .B(IN1[10]), .S(n9), .Z(mux_A[10]) );
  MUX2_X1 U176 ( .A(A_booth_to_add[0]), .B(IN1[0]), .S(n4), .Z(mux_A[0]) );
  NAND3_X1 U177 ( .A1(n81), .A2(n82), .A3(n83), .ZN(DOUT[0]) );
  NAND3_X1 U178 ( .A1(n84), .A2(n85), .A3(ALUW_i[12]), .ZN(n32) );
  simple_booth_add_ext_N16 MULT ( .Clock(Clock), .Reset(Reset), .sign(
        ALUW_i[0]), .enable(ALUW_i[1]), .valid(valid_from_booth), .A(IN1[15:0]), .B(IN2[15:0]), .A_to_add(A_booth_to_add), .B_to_add(B_booth_to_add), 
        .sign_to_add(sign_booth_to_add), .final_out(mult_out), .ACC_from_add(
        sum_out) );
  p4add_N32_logN5_1 ADDER ( .A(mux_A), .B(mux_B), .Cin(1'b0), .sign(mux_sign), 
        .S(sum_out), .Cout(carry_from_adder) );
  comparator_M32 COMP ( .C(carry_from_adder), .V(overflow), .SUM(sum_out), 
        .sel(ALUW_i[4:2]), .sign(ALUW_i[0]), .S(comp_out) );
  shifter SHIFT ( .A(IN1), .B(IN2[4:0]), .LOGIC_ARITH(ALUW_i[8]), .LEFT_RIGHT(
        ALUW_i[9]), .OUTPUT(shift_out) );
  logic_unit_SIZE32 LU ( .IN1(IN1), .IN2(IN2), .CTRL(ALUW_i[6:5]), .OUT1(
        lu_out) );
  NOR3_X1 U107 ( .A1(ALUW_i[12]), .A2(n84), .A3(n85), .ZN(n86) );
  AOI22_X1 U106 ( .A1(n1), .A2(lu_out[0]), .B1(n86), .B2(comp_out), .ZN(n81)
         );
  AOI22_X1 U103 ( .A1(n17), .A2(IN2[0]), .B1(n3), .B2(sum_out[0]), .ZN(n82) );
  AOI22_X1 U100 ( .A1(n2), .A2(shift_out[0]), .B1(n19), .B2(mult_out[0]), .ZN(
        n83) );
  AOI222_X1 U54 ( .A1(IN2[24]), .A2(n17), .B1(n1), .B2(lu_out[24]), .C1(n19), 
        .C2(mult_out[24]), .ZN(n49) );
  AOI22_X1 U53 ( .A1(n2), .A2(shift_out[24]), .B1(n3), .B2(sum_out[24]), .ZN(
        n50) );
  NAND2_X1 U52 ( .A1(n49), .A2(n50), .ZN(DOUT[24]) );
  AOI222_X1 U42 ( .A1(IN2[28]), .A2(n17), .B1(n1), .B2(lu_out[28]), .C1(n19), 
        .C2(mult_out[28]), .ZN(n41) );
  AOI22_X1 U41 ( .A1(n2), .A2(shift_out[28]), .B1(n3), .B2(sum_out[28]), .ZN(
        n42) );
  NAND2_X1 U40 ( .A1(n41), .A2(n42), .ZN(DOUT[28]) );
  AOI222_X1 U66 ( .A1(IN2[20]), .A2(n17), .B1(n1), .B2(lu_out[20]), .C1(n19), 
        .C2(mult_out[20]), .ZN(n57) );
  AOI22_X1 U65 ( .A1(n2), .A2(shift_out[20]), .B1(n3), .B2(sum_out[20]), .ZN(
        n58) );
  NAND2_X1 U64 ( .A1(n57), .A2(n58), .ZN(DOUT[20]) );
  AOI222_X1 U39 ( .A1(IN2[29]), .A2(n17), .B1(n1), .B2(lu_out[29]), .C1(n19), 
        .C2(mult_out[29]), .ZN(n39) );
  AOI22_X1 U38 ( .A1(n2), .A2(shift_out[29]), .B1(n3), .B2(sum_out[29]), .ZN(
        n40) );
  NAND2_X1 U37 ( .A1(n39), .A2(n40), .ZN(DOUT[29]) );
  AOI222_X1 U63 ( .A1(IN2[21]), .A2(n17), .B1(n1), .B2(lu_out[21]), .C1(n19), 
        .C2(mult_out[21]), .ZN(n55) );
  AOI22_X1 U62 ( .A1(n2), .A2(shift_out[21]), .B1(n3), .B2(sum_out[21]), .ZN(
        n56) );
  NAND2_X1 U61 ( .A1(n55), .A2(n56), .ZN(DOUT[21]) );
  AOI222_X1 U51 ( .A1(IN2[25]), .A2(n17), .B1(n1), .B2(lu_out[25]), .C1(n19), 
        .C2(mult_out[25]), .ZN(n47) );
  AOI22_X1 U50 ( .A1(n2), .A2(shift_out[25]), .B1(n3), .B2(sum_out[25]), .ZN(
        n48) );
  NAND2_X1 U49 ( .A1(n47), .A2(n48), .ZN(DOUT[25]) );
  AOI222_X1 U48 ( .A1(IN2[26]), .A2(n17), .B1(n1), .B2(lu_out[26]), .C1(n19), 
        .C2(mult_out[26]), .ZN(n45) );
  AOI22_X1 U47 ( .A1(n2), .A2(shift_out[26]), .B1(n3), .B2(sum_out[26]), .ZN(
        n46) );
  NAND2_X1 U46 ( .A1(n45), .A2(n46), .ZN(DOUT[26]) );
  AOI222_X1 U60 ( .A1(IN2[22]), .A2(n17), .B1(n1), .B2(lu_out[22]), .C1(n19), 
        .C2(mult_out[22]), .ZN(n53) );
  AOI22_X1 U59 ( .A1(n2), .A2(shift_out[22]), .B1(n3), .B2(sum_out[22]), .ZN(
        n54) );
  NAND2_X1 U58 ( .A1(n53), .A2(n54), .ZN(DOUT[22]) );
  AOI222_X1 U45 ( .A1(IN2[27]), .A2(n17), .B1(n1), .B2(lu_out[27]), .C1(n19), 
        .C2(mult_out[27]), .ZN(n43) );
  AOI22_X1 U44 ( .A1(n2), .A2(shift_out[27]), .B1(n3), .B2(sum_out[27]), .ZN(
        n44) );
  NAND2_X1 U43 ( .A1(n43), .A2(n44), .ZN(DOUT[27]) );
  AOI222_X1 U57 ( .A1(IN2[23]), .A2(n17), .B1(n1), .B2(lu_out[23]), .C1(n19), 
        .C2(mult_out[23]), .ZN(n51) );
  AOI22_X1 U56 ( .A1(n2), .A2(shift_out[23]), .B1(n3), .B2(sum_out[23]), .ZN(
        n52) );
  NAND2_X1 U55 ( .A1(n51), .A2(n52), .ZN(DOUT[23]) );
  AOI222_X1 U33 ( .A1(IN2[30]), .A2(n17), .B1(n1), .B2(lu_out[30]), .C1(n19), 
        .C2(mult_out[30]), .ZN(n35) );
  AOI22_X1 U32 ( .A1(n2), .A2(shift_out[30]), .B1(n3), .B2(sum_out[30]), .ZN(
        n36) );
  NAND2_X1 U31 ( .A1(n35), .A2(n36), .ZN(DOUT[30]) );
  AOI22_X1 U29 ( .A1(n2), .A2(shift_out[31]), .B1(n16), .B2(sum_out[31]), .ZN(
        n33) );
  AOI22_X1 U28 ( .A1(n1), .A2(lu_out[31]), .B1(n19), .B2(mult_out[31]), .ZN(
        n34) );
  OAI211_X1 U27 ( .C1(n32), .C2(n11), .A(n33), .B(n34), .ZN(DOUT[31]) );
  AOI222_X1 U78 ( .A1(IN2[17]), .A2(n17), .B1(n18), .B2(lu_out[17]), .C1(n19), 
        .C2(mult_out[17]), .ZN(n65) );
  AOI22_X1 U77 ( .A1(n2), .A2(shift_out[17]), .B1(n3), .B2(sum_out[17]), .ZN(
        n66) );
  NAND2_X1 U76 ( .A1(n65), .A2(n66), .ZN(DOUT[17]) );
  AOI222_X1 U75 ( .A1(IN2[18]), .A2(n17), .B1(n18), .B2(lu_out[18]), .C1(n19), 
        .C2(mult_out[18]), .ZN(n63) );
  AOI22_X1 U74 ( .A1(n2), .A2(shift_out[18]), .B1(n3), .B2(sum_out[18]), .ZN(
        n64) );
  NAND2_X1 U73 ( .A1(n63), .A2(n64), .ZN(DOUT[18]) );
  AOI222_X1 U72 ( .A1(IN2[19]), .A2(n17), .B1(n1), .B2(lu_out[19]), .C1(n19), 
        .C2(mult_out[19]), .ZN(n61) );
  AOI22_X1 U71 ( .A1(n2), .A2(shift_out[19]), .B1(n3), .B2(sum_out[19]), .ZN(
        n62) );
  NAND2_X1 U70 ( .A1(n61), .A2(n62), .ZN(DOUT[19]) );
  AOI222_X1 U81 ( .A1(IN2[16]), .A2(n17), .B1(n18), .B2(lu_out[16]), .C1(n19), 
        .C2(mult_out[16]), .ZN(n67) );
  AOI22_X1 U80 ( .A1(n2), .A2(shift_out[16]), .B1(n3), .B2(sum_out[16]), .ZN(
        n68) );
  NAND2_X1 U79 ( .A1(n67), .A2(n68), .ZN(DOUT[16]) );
  AOI222_X1 U90 ( .A1(IN2[13]), .A2(n17), .B1(n18), .B2(lu_out[13]), .C1(n19), 
        .C2(mult_out[13]), .ZN(n73) );
  AOI22_X1 U89 ( .A1(n2), .A2(shift_out[13]), .B1(n3), .B2(sum_out[13]), .ZN(
        n74) );
  NAND2_X1 U88 ( .A1(n73), .A2(n74), .ZN(DOUT[13]) );
  AOI222_X1 U93 ( .A1(IN2[12]), .A2(n17), .B1(n18), .B2(lu_out[12]), .C1(n19), 
        .C2(mult_out[12]), .ZN(n75) );
  AOI22_X1 U92 ( .A1(n2), .A2(shift_out[12]), .B1(n3), .B2(sum_out[12]), .ZN(
        n76) );
  NAND2_X1 U91 ( .A1(n75), .A2(n76), .ZN(DOUT[12]) );
  AOI222_X1 U87 ( .A1(IN2[14]), .A2(n17), .B1(n1), .B2(lu_out[14]), .C1(n19), 
        .C2(mult_out[14]), .ZN(n71) );
  AOI22_X1 U86 ( .A1(n2), .A2(shift_out[14]), .B1(n3), .B2(sum_out[14]), .ZN(
        n72) );
  NAND2_X1 U85 ( .A1(n71), .A2(n72), .ZN(DOUT[14]) );
  AOI222_X1 U84 ( .A1(IN2[15]), .A2(n17), .B1(n1), .B2(lu_out[15]), .C1(n19), 
        .C2(mult_out[15]), .ZN(n69) );
  AOI22_X1 U83 ( .A1(n2), .A2(shift_out[15]), .B1(n3), .B2(sum_out[15]), .ZN(
        n70) );
  NAND2_X1 U82 ( .A1(n69), .A2(n70), .ZN(DOUT[15]) );
  AOI222_X1 U99 ( .A1(IN2[10]), .A2(n17), .B1(n1), .B2(lu_out[10]), .C1(n19), 
        .C2(mult_out[10]), .ZN(n79) );
  AOI22_X1 U98 ( .A1(n2), .A2(shift_out[10]), .B1(n3), .B2(sum_out[10]), .ZN(
        n80) );
  NAND2_X1 U97 ( .A1(n79), .A2(n80), .ZN(DOUT[10]) );
  AOI222_X1 U96 ( .A1(IN2[11]), .A2(n17), .B1(n1), .B2(lu_out[11]), .C1(n19), 
        .C2(mult_out[11]), .ZN(n77) );
  AOI22_X1 U95 ( .A1(n2), .A2(shift_out[11]), .B1(n3), .B2(sum_out[11]), .ZN(
        n78) );
  NAND2_X1 U94 ( .A1(n77), .A2(n78), .ZN(DOUT[11]) );
  AOI222_X1 U11 ( .A1(IN2[8]), .A2(n17), .B1(n1), .B2(lu_out[8]), .C1(n19), 
        .C2(mult_out[8]), .ZN(n20) );
  AOI22_X1 U10 ( .A1(n15), .A2(shift_out[8]), .B1(n3), .B2(sum_out[8]), .ZN(
        n21) );
  NAND2_X1 U9 ( .A1(n20), .A2(n21), .ZN(DOUT[8]) );
  AOI222_X1 U8 ( .A1(IN2[9]), .A2(n17), .B1(n1), .B2(lu_out[9]), .C1(n19), 
        .C2(mult_out[9]), .ZN(n13) );
  AOI22_X1 U7 ( .A1(n15), .A2(shift_out[9]), .B1(n16), .B2(sum_out[9]), .ZN(
        n14) );
  NAND2_X1 U6 ( .A1(n13), .A2(n14), .ZN(DOUT[9]) );
  AOI222_X1 U14 ( .A1(IN2[7]), .A2(n17), .B1(n1), .B2(lu_out[7]), .C1(n19), 
        .C2(mult_out[7]), .ZN(n22) );
  AOI22_X1 U13 ( .A1(n2), .A2(shift_out[7]), .B1(n3), .B2(sum_out[7]), .ZN(n23) );
  NAND2_X1 U12 ( .A1(n22), .A2(n23), .ZN(DOUT[7]) );
  AOI222_X1 U26 ( .A1(IN2[3]), .A2(n17), .B1(n1), .B2(lu_out[3]), .C1(n19), 
        .C2(mult_out[3]), .ZN(n30) );
  AOI22_X1 U25 ( .A1(n2), .A2(shift_out[3]), .B1(n16), .B2(sum_out[3]), .ZN(
        n31) );
  NAND2_X1 U24 ( .A1(n30), .A2(n31), .ZN(DOUT[3]) );
  AOI222_X1 U17 ( .A1(IN2[6]), .A2(n17), .B1(n1), .B2(lu_out[6]), .C1(n19), 
        .C2(mult_out[6]), .ZN(n24) );
  AOI22_X1 U16 ( .A1(n15), .A2(shift_out[6]), .B1(n16), .B2(sum_out[6]), .ZN(
        n25) );
  NAND2_X1 U15 ( .A1(n24), .A2(n25), .ZN(DOUT[6]) );
  AOI222_X1 U23 ( .A1(IN2[4]), .A2(n17), .B1(n1), .B2(lu_out[4]), .C1(n19), 
        .C2(mult_out[4]), .ZN(n28) );
  AOI22_X1 U22 ( .A1(n15), .A2(shift_out[4]), .B1(n16), .B2(sum_out[4]), .ZN(
        n29) );
  NAND2_X1 U21 ( .A1(n28), .A2(n29), .ZN(DOUT[4]) );
  AOI222_X1 U20 ( .A1(IN2[5]), .A2(n17), .B1(n1), .B2(lu_out[5]), .C1(n19), 
        .C2(mult_out[5]), .ZN(n26) );
  AOI22_X1 U19 ( .A1(n15), .A2(shift_out[5]), .B1(n16), .B2(sum_out[5]), .ZN(
        n27) );
  NAND2_X1 U18 ( .A1(n26), .A2(n27), .ZN(DOUT[5]) );
  AOI222_X1 U36 ( .A1(IN2[2]), .A2(n17), .B1(n1), .B2(lu_out[2]), .C1(n19), 
        .C2(mult_out[2]), .ZN(n37) );
  AOI22_X1 U35 ( .A1(n2), .A2(shift_out[2]), .B1(n3), .B2(sum_out[2]), .ZN(n38) );
  NAND2_X1 U34 ( .A1(n37), .A2(n38), .ZN(DOUT[2]) );
  AOI222_X1 U69 ( .A1(IN2[1]), .A2(n17), .B1(n1), .B2(lu_out[1]), .C1(n19), 
        .C2(mult_out[1]), .ZN(n59) );
  AOI22_X1 U68 ( .A1(n2), .A2(shift_out[1]), .B1(n3), .B2(sum_out[1]), .ZN(n60) );
  NAND2_X1 U67 ( .A1(n59), .A2(n60), .ZN(DOUT[1]) );
  NOR3_X1 U109 ( .A1(ALUW_i[11]), .A2(ALUW_i[12]), .A3(n85), .ZN(n18) );
  NOR3_X1 U104 ( .A1(ALUW_i[11]), .A2(ALUW_i[12]), .A3(ALUW_i[10]), .ZN(n16)
         );
  NOR3_X1 U102 ( .A1(ALUW_i[12]), .A2(ALUW_i[10]), .A3(n84), .ZN(n15) );
  INV_X1 U110 ( .A(ALUW_i[10]), .ZN(n85) );
  INV_X1 U108 ( .A(ALUW_i[11]), .ZN(n84) );
  INV_X1 U4 ( .A(IN1[31]), .ZN(n10) );
  INV_X1 U30 ( .A(IN2[31]), .ZN(n11) );
  INV_X1 U3 ( .A(sum_out[31]), .ZN(n12) );
  NOR2_X1 U2 ( .A1(valid_from_booth), .A2(n9), .ZN(stall_o) );
  INV_X2 U5 ( .A(n32), .ZN(n17) );
  BUF_X1 U101 ( .A(n16), .Z(n3) );
  INV_X1 U105 ( .A(ALUW_i[1]), .ZN(n9) );
  BUF_X2 U112 ( .A(n5), .Z(n4) );
  AND2_X2 U179 ( .A1(n32), .A2(ALUW_i[12]), .ZN(n19) );
  BUF_X2 U180 ( .A(n18), .Z(n1) );
  BUF_X2 U181 ( .A(n15), .Z(n2) );
  BUF_X1 U182 ( .A(n9), .Z(n5) );
  MUX2_X2 U183 ( .A(sign_booth_to_add), .B(ALUW_i[7]), .S(n5), .Z(mux_sign) );
endmodule


module ff32_en_SIZE13 ( D, en, clk, rst, Q );
  input [12:0] D;
  output [12:0] Q;
  input en, clk, rst;
  wire   net338027, n13;

  DFFR_X1 \Q_reg[12]  ( .D(D[12]), .CK(net338027), .RN(n13), .Q(Q[12]) );
  DFFR_X1 \Q_reg[11]  ( .D(D[11]), .CK(net338027), .RN(n13), .Q(Q[11]) );
  DFFR_X1 \Q_reg[10]  ( .D(D[10]), .CK(net338027), .RN(n13), .Q(Q[10]) );
  DFFR_X1 \Q_reg[9]  ( .D(D[9]), .CK(net338027), .RN(n13), .Q(Q[9]) );
  DFFR_X1 \Q_reg[8]  ( .D(D[8]), .CK(net338027), .RN(n13), .Q(Q[8]) );
  DFFR_X1 \Q_reg[7]  ( .D(D[7]), .CK(net338027), .RN(n13), .Q(Q[7]) );
  DFFR_X1 \Q_reg[6]  ( .D(D[6]), .CK(net338027), .RN(n13), .Q(Q[6]) );
  DFFR_X1 \Q_reg[5]  ( .D(D[5]), .CK(net338027), .RN(n13), .Q(Q[5]) );
  DFFR_X1 \Q_reg[4]  ( .D(D[4]), .CK(net338027), .RN(n13), .Q(Q[4]) );
  DFFR_X1 \Q_reg[3]  ( .D(D[3]), .CK(net338027), .RN(n13), .Q(Q[3]) );
  DFFR_X1 \Q_reg[2]  ( .D(D[2]), .CK(net338027), .RN(n13), .Q(Q[2]) );
  DFFR_X1 \Q_reg[1]  ( .D(D[1]), .CK(net338027), .RN(n13), .Q(Q[1]) );
  DFFR_X1 \Q_reg[0]  ( .D(D[0]), .CK(net338027), .RN(n13), .Q(Q[0]) );
  SNPS_CLOCK_GATE_HIGH_ff32_en_SIZE13 clk_gate_Q_reg ( .CLK(clk), .EN(en), 
        .ENCLK(net338027) );
  INV_X1 U2 ( .A(rst), .ZN(n13) );
endmodule


module ff32_en_SIZE5_0 ( D, en, clk, rst, Q );
  input [4:0] D;
  output [4:0] Q;
  input en, clk, rst;
  wire   net338012, n5;

  DFFR_X1 \Q_reg[4]  ( .D(D[4]), .CK(net338012), .RN(n5), .Q(Q[4]) );
  DFFR_X1 \Q_reg[3]  ( .D(D[3]), .CK(net338012), .RN(n5), .Q(Q[3]) );
  DFFR_X1 \Q_reg[2]  ( .D(D[2]), .CK(net338012), .RN(n5), .Q(Q[2]) );
  DFFR_X1 \Q_reg[1]  ( .D(D[1]), .CK(net338012), .RN(n5), .Q(Q[1]) );
  DFFR_X1 \Q_reg[0]  ( .D(D[0]), .CK(net338012), .RN(n5), .Q(Q[0]) );
  SNPS_CLOCK_GATE_HIGH_ff32_en_SIZE5_0 clk_gate_Q_reg ( .CLK(clk), .EN(en), 
        .ENCLK(net338012) );
  INV_X1 U2 ( .A(rst), .ZN(n5) );
endmodule


module ff32_en_SIZE32_0 ( D, en, clk, rst, Q );
  input [31:0] D;
  output [31:0] Q;
  input en, clk, rst;
  wire   net337997, n32, n34;

  DFFR_X1 \Q_reg[31]  ( .D(D[31]), .CK(net337997), .RN(n34), .Q(Q[31]) );
  DFFR_X1 \Q_reg[30]  ( .D(D[30]), .CK(net337997), .RN(n34), .Q(Q[30]) );
  DFFR_X1 \Q_reg[29]  ( .D(D[29]), .CK(net337997), .RN(n34), .Q(Q[29]) );
  DFFR_X1 \Q_reg[28]  ( .D(D[28]), .CK(net337997), .RN(n34), .Q(Q[28]) );
  DFFR_X1 \Q_reg[27]  ( .D(D[27]), .CK(net337997), .RN(n34), .Q(Q[27]) );
  DFFR_X1 \Q_reg[26]  ( .D(D[26]), .CK(net337997), .RN(n34), .Q(Q[26]) );
  DFFR_X1 \Q_reg[25]  ( .D(D[25]), .CK(net337997), .RN(n34), .Q(Q[25]) );
  DFFR_X1 \Q_reg[24]  ( .D(D[24]), .CK(net337997), .RN(n34), .Q(Q[24]) );
  DFFR_X1 \Q_reg[23]  ( .D(D[23]), .CK(net337997), .RN(n32), .Q(Q[23]) );
  DFFR_X1 \Q_reg[22]  ( .D(D[22]), .CK(net337997), .RN(n34), .Q(Q[22]) );
  DFFR_X1 \Q_reg[21]  ( .D(D[21]), .CK(net337997), .RN(n32), .Q(Q[21]) );
  DFFR_X1 \Q_reg[20]  ( .D(D[20]), .CK(net337997), .RN(n34), .Q(Q[20]) );
  DFFR_X1 \Q_reg[19]  ( .D(D[19]), .CK(net337997), .RN(n32), .Q(Q[19]) );
  DFFR_X1 \Q_reg[18]  ( .D(D[18]), .CK(net337997), .RN(n34), .Q(Q[18]) );
  DFFR_X1 \Q_reg[17]  ( .D(D[17]), .CK(net337997), .RN(n32), .Q(Q[17]) );
  DFFR_X1 \Q_reg[16]  ( .D(D[16]), .CK(net337997), .RN(n34), .Q(Q[16]) );
  DFFR_X1 \Q_reg[15]  ( .D(D[15]), .CK(net337997), .RN(n34), .Q(Q[15]) );
  DFFR_X1 \Q_reg[14]  ( .D(D[14]), .CK(net337997), .RN(n34), .Q(Q[14]) );
  DFFR_X1 \Q_reg[13]  ( .D(D[13]), .CK(net337997), .RN(n34), .Q(Q[13]) );
  DFFR_X1 \Q_reg[12]  ( .D(D[12]), .CK(net337997), .RN(n34), .Q(Q[12]) );
  DFFR_X1 \Q_reg[11]  ( .D(D[11]), .CK(net337997), .RN(n32), .Q(Q[11]) );
  DFFR_X1 \Q_reg[10]  ( .D(D[10]), .CK(net337997), .RN(n32), .Q(Q[10]) );
  DFFR_X1 \Q_reg[9]  ( .D(D[9]), .CK(net337997), .RN(n32), .Q(Q[9]) );
  DFFR_X1 \Q_reg[8]  ( .D(D[8]), .CK(net337997), .RN(n32), .Q(Q[8]) );
  DFFR_X1 \Q_reg[7]  ( .D(D[7]), .CK(net337997), .RN(n32), .Q(Q[7]) );
  DFFR_X1 \Q_reg[6]  ( .D(D[6]), .CK(net337997), .RN(n32), .Q(Q[6]) );
  DFFR_X1 \Q_reg[5]  ( .D(D[5]), .CK(net337997), .RN(n32), .Q(Q[5]) );
  DFFR_X1 \Q_reg[4]  ( .D(D[4]), .CK(net337997), .RN(n32), .Q(Q[4]) );
  DFFR_X1 \Q_reg[3]  ( .D(D[3]), .CK(net337997), .RN(n32), .Q(Q[3]) );
  DFFR_X1 \Q_reg[2]  ( .D(D[2]), .CK(net337997), .RN(n32), .Q(Q[2]) );
  DFFR_X1 \Q_reg[1]  ( .D(D[1]), .CK(net337997), .RN(n32), .Q(Q[1]) );
  DFFR_X1 \Q_reg[0]  ( .D(D[0]), .CK(net337997), .RN(n32), .Q(Q[0]) );
  SNPS_CLOCK_GATE_HIGH_ff32_en_SIZE32_0 clk_gate_Q_reg ( .CLK(clk), .EN(en), 
        .ENCLK(net337997) );
  CLKBUF_X1 U2 ( .A(n34), .Z(n32) );
  INV_X1 U3 ( .A(rst), .ZN(n34) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dlx_regfile_0 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net338030, net338032, net338033, net338036;
  assign net338030 = CLK;
  assign ENCLK = net338032;
  assign net338033 = EN;

  DLL_X1 latch ( .D(net338033), .GN(net338030), .Q(net338036) );
  AND2_X1 main_gate ( .A1(net338036), .A2(net338030), .ZN(net338032) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_dlx_cu_MICROCODE_MEM_SIZE64_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE13_0 ( 
        CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net338210, net338212, net338213, net338216;
  assign net338210 = CLK;
  assign ENCLK = net338212;
  assign net338213 = EN;

  DLL_X1 latch ( .D(net338213), .GN(net338210), .Q(net338216) );
  AND2_X1 main_gate ( .A1(net338216), .A2(net338210), .ZN(net338212) );
endmodule


module alu_ctrl ( .OP({\OP[4] , \OP[3] , \OP[2] , \OP[1] , \OP[0] }), ALU_WORD
 );
  output [12:0] ALU_WORD;
  input \OP[4] , \OP[3] , \OP[2] , \OP[1] , \OP[0] ;
  wire   N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32, N33,
         n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35;

  DLH_X1 \comp_sel_reg[2]  ( .G(N32), .D(N33), .Q(ALU_WORD[4]) );
  DLH_X1 \comp_sel_reg[1]  ( .G(N32), .D(N31), .Q(ALU_WORD[3]) );
  DLH_X1 \comp_sel_reg[0]  ( .G(N32), .D(N30), .Q(ALU_WORD[2]) );
  DLH_X1 sign_to_booth_reg ( .G(N20), .D(N21), .Q(ALU_WORD[0]) );
  DLH_X1 left_right_reg ( .G(N23), .D(N22), .Q(ALU_WORD[9]) );
  DLH_X1 logic_arith_reg ( .G(N23), .D(N24), .Q(ALU_WORD[8]) );
  DLH_X1 sign_to_adder_reg ( .G(N25), .D(N26), .Q(ALU_WORD[7]) );
  DLH_X1 \lu_ctrl_reg[1]  ( .G(N28), .D(N29), .Q(ALU_WORD[6]) );
  DLH_X1 \lu_ctrl_reg[0]  ( .G(N28), .D(N27), .Q(ALU_WORD[5]) );
  NAND3_X1 U53 ( .A1(n9), .A2(OP[1]), .A3(n28), .ZN(n30) );
  NAND3_X1 U54 ( .A1(n15), .A2(n35), .A3(n22), .ZN(n19) );
  NOR3_X1 U48 ( .A1(OP[2]), .A2(OP[0]), .A3(n22), .ZN(n10) );
  NOR3_X1 U45 ( .A1(OP[2]), .A2(n35), .A3(n22), .ZN(n33) );
  NOR2_X1 U43 ( .A1(n3), .A2(n2), .ZN(n32) );
  NOR2_X1 U41 ( .A1(OP[0]), .A2(n15), .ZN(n28) );
  NAND2_X1 U40 ( .A1(n28), .A2(n22), .ZN(n1) );
  NOR2_X1 U39 ( .A1(n19), .A2(OP[3]), .ZN(n34) );
  NOR4_X1 U38 ( .A1(n15), .A2(n3), .A3(n35), .A4(n22), .ZN(n8) );
  AOI21_X1 U37 ( .B1(n34), .B2(OP[4]), .A(n8), .ZN(n18) );
  NAND2_X1 U36 ( .A1(n33), .A2(n26), .ZN(n6) );
  OAI211_X1 U35 ( .C1(n1), .C2(n16), .A(n18), .B(n6), .ZN(N30) );
  AOI211_X1 U34 ( .C1(n26), .C2(n10), .A(n32), .B(N30), .ZN(n29) );
  NAND2_X1 U33 ( .A1(OP[0]), .A2(n22), .ZN(n27) );
  NOR2_X1 U32 ( .A1(n3), .A2(n27), .ZN(n31) );
  NAND2_X1 U31 ( .A1(OP[2]), .A2(n31), .ZN(n4) );
  NOR2_X1 U29 ( .A1(OP[2]), .A2(n27), .ZN(n24) );
  NAND2_X1 U28 ( .A1(n26), .A2(n24), .ZN(n7) );
  NAND4_X1 U27 ( .A1(n29), .A2(n4), .A3(n30), .A4(n7), .ZN(N32) );
  AOI211_X1 U26 ( .C1(OP[0]), .C2(OP[1]), .A(OP[2]), .B(n3), .ZN(N28) );
  NAND2_X1 U25 ( .A1(OP[1]), .A2(n28), .ZN(n17) );
  OAI21_X1 U24 ( .B1(n27), .B2(n15), .A(n17), .ZN(n25) );
  NAND2_X1 U23 ( .A1(n25), .A2(n26), .ZN(n20) );
  NOR3_X1 U18 ( .A1(OP[2]), .A2(n22), .A3(n13), .ZN(N22) );
  OAI21_X1 U16 ( .B1(n11), .B2(n13), .A(n21), .ZN(N23) );
  OAI21_X1 U14 ( .B1(n19), .B2(n13), .A(n20), .ZN(ALU_WORD[12]) );
  NOR2_X1 U6 ( .A1(n3), .A2(n11), .ZN(N27) );
  NAND2_X1 U8 ( .A1(OP[2]), .A2(OP[1]), .ZN(n12) );
  OAI21_X1 U7 ( .B1(n12), .B2(n13), .A(n14), .ZN(N26) );
  NOR2_X1 U11 ( .A1(n2), .A2(n13), .ZN(N24) );
  OAI211_X1 U12 ( .C1(n16), .C2(n17), .A(n18), .B(n4), .ZN(N21) );
  NAND4_X1 U3 ( .A1(n4), .A2(n5), .A3(n6), .A4(n7), .ZN(N31) );
  AOI21_X1 U2 ( .B1(n1), .B2(n2), .A(n3), .ZN(N33) );
  OAI21_X1 U9 ( .B1(n15), .B2(n13), .A(n14), .ZN(N25) );
  NAND2_X1 U47 ( .A1(OP[3]), .A2(n23), .ZN(n3) );
  NAND2_X1 U19 ( .A1(n23), .A2(n16), .ZN(n13) );
  NOR2_X1 U50 ( .A1(n23), .A2(n16), .ZN(n26) );
  INV_X1 U52 ( .A(OP[4]), .ZN(n23) );
  INV_X1 U51 ( .A(OP[3]), .ZN(n16) );
  INV_X1 U49 ( .A(OP[1]), .ZN(n22) );
  INV_X1 U46 ( .A(OP[0]), .ZN(n35) );
  INV_X1 U44 ( .A(n33), .ZN(n2) );
  INV_X1 U42 ( .A(OP[2]), .ZN(n15) );
  INV_X1 U30 ( .A(n3), .ZN(n9) );
  INV_X1 U22 ( .A(n20), .ZN(ALU_WORD[1]) );
  OR3_X1 U21 ( .A1(N32), .A2(N28), .A3(ALU_WORD[1]), .ZN(ALU_WORD[10]) );
  INV_X1 U20 ( .A(n24), .ZN(n11) );
  INV_X1 U17 ( .A(N22), .ZN(n21) );
  OR2_X1 U15 ( .A1(N32), .A2(N23), .ZN(ALU_WORD[11]) );
  AND2_X1 U5 ( .A1(n9), .A2(n10), .ZN(N29) );
  INV_X1 U10 ( .A(N32), .ZN(n14) );
  INV_X1 U4 ( .A(n8), .ZN(n5) );
  OR2_X1 U13 ( .A1(N32), .A2(ALU_WORD[12]), .ZN(N20) );
endmodule


module cw_mem_MICROCODE_MEM_SIZE64_OP_CODE_SIZE6_CW_SIZE13 ( OPCODE_IN, CW_OUT
 );
  input [5:0] OPCODE_IN;
  output [12:0] CW_OUT;
  wire   \CW_OUT[5] , CW_OUT_4, CW_OUT_3, CW_OUT_2, CW_OUT_1, CW_OUT_0, n6, n7,
         n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29;
  assign CW_OUT[6] = \CW_OUT[5] ;
  assign CW_OUT[5] = \CW_OUT[5] ;
  assign CW_OUT[4] = CW_OUT_4;
  assign CW_OUT[3] = CW_OUT_3;
  assign CW_OUT[2] = CW_OUT_2;
  assign CW_OUT[1] = CW_OUT_1;
  assign CW_OUT[0] = CW_OUT_0;

  NAND3_X1 U34 ( .A1(OPCODE_IN[3]), .A2(n13), .A3(n14), .ZN(n15) );
  NAND3_X1 U35 ( .A1(OPCODE_IN[3]), .A2(n23), .A3(n24), .ZN(n22) );
  NAND3_X1 U36 ( .A1(OPCODE_IN[4]), .A2(n14), .A3(n25), .ZN(n29) );
  NAND2_X1 U26 ( .A1(OPCODE_IN[2]), .A2(n13), .ZN(n17) );
  OAI21_X1 U23 ( .B1(OPCODE_IN[3]), .B2(n17), .A(n29), .ZN(CW_OUT[11]) );
  OAI221_X1 U6 ( .B1(OPCODE_IN[0]), .B2(n12), .C1(OPCODE_IN[0]), .C2(n15), .A(
        n16), .ZN(CW_OUT[9]) );
  NOR2_X1 U28 ( .A1(OPCODE_IN[3]), .A2(n12), .ZN(CW_OUT[10]) );
  NOR2_X1 U8 ( .A1(n10), .A2(n17), .ZN(CW_OUT[8]) );
  NAND2_X1 U5 ( .A1(n13), .A2(n14), .ZN(n11) );
  OAI22_X1 U4 ( .A1(OPCODE_IN[3]), .A2(n11), .B1(n12), .B2(n10), .ZN(CW_OUT_4)
         );
  NAND2_X1 U20 ( .A1(OPCODE_IN[5]), .A2(n28), .ZN(n8) );
  NOR2_X1 U3 ( .A1(n8), .A2(n10), .ZN(CW_OUT_1) );
  NOR2_X1 U19 ( .A1(n7), .A2(n8), .ZN(CW_OUT_3) );
  NAND2_X1 U16 ( .A1(OPCODE_IN[3]), .A2(OPCODE_IN[4]), .ZN(n20) );
  NAND2_X1 U15 ( .A1(n23), .A2(n7), .ZN(n27) );
  AOI21_X1 U14 ( .B1(n6), .B2(n27), .A(OPCODE_IN[1]), .ZN(n26) );
  OAI211_X1 U13 ( .C1(n25), .C2(n26), .A(OPCODE_IN[2]), .B(OPCODE_IN[4]), .ZN(
        n21) );
  OAI211_X1 U12 ( .C1(OPCODE_IN[4]), .C2(OPCODE_IN[0]), .A(OPCODE_IN[1]), .B(
        OPCODE_IN[2]), .ZN(n24) );
  OAI211_X1 U11 ( .C1(n19), .C2(n20), .A(n21), .B(n22), .ZN(n18) );
  NOR3_X1 U1 ( .A1(n6), .A2(n7), .A3(n8), .ZN(CW_OUT_2) );
  NOR3_X1 U27 ( .A1(OPCODE_IN[5]), .A2(OPCODE_IN[1]), .A3(OPCODE_IN[4]), .ZN(
        n13) );
  AOI21_X1 U22 ( .B1(n12), .B2(n17), .A(OPCODE_IN[3]), .ZN(CW_OUT[12]) );
  INV_X1 U21 ( .A(OPCODE_IN[0]), .ZN(n7) );
  NAND2_X1 U18 ( .A1(OPCODE_IN[0]), .A2(n6), .ZN(n10) );
  NOR3_X1 U17 ( .A1(OPCODE_IN[5]), .A2(n19), .A3(n10), .ZN(CW_OUT[7]) );
  NAND2_X1 U32 ( .A1(OPCODE_IN[1]), .A2(n14), .ZN(n19) );
  INV_X1 U30 ( .A(OPCODE_IN[5]), .ZN(n23) );
  NOR2_X1 U31 ( .A1(OPCODE_IN[4]), .A2(n19), .ZN(n28) );
  NAND2_X1 U29 ( .A1(n28), .A2(n23), .ZN(n12) );
  AND3_X1 U24 ( .A1(n23), .A2(n6), .A3(OPCODE_IN[1]), .ZN(n25) );
  INV_X1 U7 ( .A(CW_OUT[12]), .ZN(n16) );
  OR2_X1 U10 ( .A1(CW_OUT[7]), .A2(n18), .ZN(n9) );
  OR2_X1 U9 ( .A1(CW_OUT_3), .A2(n9), .ZN(\CW_OUT[5] ) );
  OR3_X1 U2 ( .A1(n9), .A2(CW_OUT_4), .A3(CW_OUT_1), .ZN(CW_OUT_0) );
  INV_X1 U33 ( .A(OPCODE_IN[2]), .ZN(n14) );
  INV_X1 U25 ( .A(OPCODE_IN[3]), .ZN(n6) );
endmodule


module stall_logic_FUNC_SIZE11_OP_CODE_SIZE6 ( OPCODE_i, FUNC_i, rA_i, rB_i, 
        D1_i, D2_i, S_mem_LOAD_i, S_exe_LOAD_i, S_exe_WRITE_i, S_MUX_PC_BUS_i, 
        mispredict_i, bubble_dec_o, bubble_exe_o, stall_exe_o, stall_dec_o, 
        stall_btb_o, stall_fetch_o );
  input [5:0] OPCODE_i;
  input [10:0] FUNC_i;
  input [4:0] rA_i;
  input [4:0] rB_i;
  input [4:0] D1_i;
  input [4:0] D2_i;
  input [1:0] S_MUX_PC_BUS_i;
  input S_mem_LOAD_i, S_exe_LOAD_i, S_exe_WRITE_i, mispredict_i;
  output bubble_dec_o, bubble_exe_o, stall_exe_o, stall_dec_o, stall_btb_o,
         stall_fetch_o;
  wire   stall_fetch_o, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58;
  assign stall_dec_o = stall_fetch_o;
  assign stall_btb_o = stall_fetch_o;

  OAI33_X1 U46 ( .A1(OPCODE_i[2]), .A2(n52), .A3(n53), .B1(n50), .B2(
        OPCODE_i[4]), .B3(OPCODE_i[1]), .ZN(n51) );
  OAI22_X1 U43 ( .A1(n43), .A2(D2_i[3]), .B1(n40), .B2(D2_i[1]), .ZN(n58) );
  AOI221_X1 U42 ( .B1(n43), .B2(D2_i[3]), .C1(D2_i[1]), .C2(n40), .A(n58), 
        .ZN(n54) );
  OAI22_X1 U39 ( .A1(n41), .A2(D2_i[0]), .B1(n44), .B2(D2_i[2]), .ZN(n57) );
  AOI221_X1 U38 ( .B1(n41), .B2(D2_i[0]), .C1(D2_i[2]), .C2(n44), .A(n57), 
        .ZN(n55) );
  XNOR2_X1 U37 ( .A(rA_i[4]), .B(D2_i[4]), .ZN(n56) );
  NAND4_X1 U36 ( .A1(S_mem_LOAD_i), .A2(n54), .A3(n55), .A4(n56), .ZN(n17) );
  NOR2_X1 U35 ( .A1(OPCODE_i[5]), .A2(OPCODE_i[3]), .ZN(n27) );
  INV_X1 U32 ( .A(OPCODE_i[2]), .ZN(n50) );
  NAND2_X1 U31 ( .A1(n27), .A2(n51), .ZN(n18) );
  OAI21_X1 U30 ( .B1(OPCODE_i[0]), .B2(n50), .A(OPCODE_i[4]), .ZN(n48) );
  NAND2_X1 U29 ( .A1(OPCODE_i[1]), .A2(n50), .ZN(n49) );
  OAI22_X1 U28 ( .A1(OPCODE_i[1]), .A2(n48), .B1(OPCODE_i[4]), .B2(n49), .ZN(
        n46) );
  AOI21_X1 U26 ( .B1(n27), .B2(n46), .A(n47), .ZN(n34) );
  XNOR2_X1 U23 ( .A(n31), .B(rA_i[4]), .ZN(n37) );
  AOI22_X1 U22 ( .A1(n43), .A2(D1_i[3]), .B1(D1_i[2]), .B2(n44), .ZN(n45) );
  OAI221_X1 U21 ( .B1(n43), .B2(D1_i[3]), .C1(n44), .C2(D1_i[2]), .A(n45), 
        .ZN(n38) );
  AOI22_X1 U20 ( .A1(n40), .A2(D1_i[1]), .B1(D1_i[0]), .B2(n41), .ZN(n42) );
  OAI221_X1 U19 ( .B1(n40), .B2(D1_i[1]), .C1(n41), .C2(D1_i[0]), .A(n42), 
        .ZN(n39) );
  NOR3_X1 U18 ( .A1(n37), .A2(n38), .A3(n39), .ZN(n36) );
  OAI221_X1 U17 ( .B1(n34), .B2(n35), .C1(n34), .C2(S_exe_WRITE_i), .A(n36), 
        .ZN(n19) );
  OAI22_X1 U15 ( .A1(n31), .A2(rB_i[4]), .B1(n32), .B2(rB_i[2]), .ZN(n33) );
  AOI221_X1 U14 ( .B1(n31), .B2(rB_i[4]), .C1(rB_i[2]), .C2(n32), .A(n33), 
        .ZN(n21) );
  OAI22_X1 U11 ( .A1(n28), .A2(rB_i[0]), .B1(n29), .B2(rB_i[3]), .ZN(n30) );
  AOI221_X1 U10 ( .B1(n28), .B2(rB_i[0]), .C1(rB_i[3]), .C2(n29), .A(n30), 
        .ZN(n22) );
  NOR4_X1 U9 ( .A1(OPCODE_i[2]), .A2(OPCODE_i[4]), .A3(OPCODE_i[1]), .A4(
        OPCODE_i[0]), .ZN(n23) );
  OAI211_X1 U7 ( .C1(n25), .C2(rB_i[1]), .A(S_exe_LOAD_i), .B(n27), .ZN(n26)
         );
  AOI21_X1 U6 ( .B1(n25), .B2(rB_i[1]), .A(n26), .ZN(n24) );
  NAND4_X1 U5 ( .A1(n21), .A2(n22), .A3(n23), .A4(n24), .ZN(n20) );
  NOR2_X1 U2 ( .A1(stall_fetch_o), .A2(n16), .ZN(bubble_dec_o) );
  OAI211_X1 U4 ( .C1(n17), .C2(n18), .A(n19), .B(n20), .ZN(stall_fetch_o) );
  INV_X1 U33 ( .A(OPCODE_i[1]), .ZN(n53) );
  INV_X1 U45 ( .A(rA_i[3]), .ZN(n43) );
  INV_X1 U44 ( .A(rA_i[1]), .ZN(n40) );
  INV_X1 U41 ( .A(rA_i[0]), .ZN(n41) );
  INV_X1 U40 ( .A(rA_i[2]), .ZN(n44) );
  INV_X1 U34 ( .A(OPCODE_i[4]), .ZN(n52) );
  INV_X1 U27 ( .A(S_exe_LOAD_i), .ZN(n47) );
  INV_X1 U25 ( .A(n18), .ZN(n35) );
  INV_X1 U24 ( .A(D1_i[4]), .ZN(n31) );
  INV_X1 U16 ( .A(D1_i[2]), .ZN(n32) );
  INV_X1 U13 ( .A(D1_i[0]), .ZN(n28) );
  INV_X1 U12 ( .A(D1_i[3]), .ZN(n29) );
  INV_X1 U8 ( .A(D1_i[1]), .ZN(n25) );
  INV_X1 U3 ( .A(mispredict_i), .ZN(n16) );
endmodule


module mux41_MUX_SIZE32_0 ( IN0, IN1, IN2, IN3, CTRL, OUT1 );
  input [31:0] IN0;
  input [31:0] IN1;
  input [31:0] IN2;
  input [31:0] IN3;
  input [1:0] CTRL;
  output [31:0] OUT1;
  wire   n3, n4, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n25, n26, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n1, n2, n5, n21, n22, n23, n24;

  AOI22_X1 U63 ( .A1(n7), .A2(IN1[1]), .B1(n23), .B2(IN0[1]), .ZN(n47) );
  NAND2_X1 U61 ( .A1(n47), .A2(n48), .ZN(OUT1[1]) );
  AOI22_X1 U66 ( .A1(n7), .A2(IN1[19]), .B1(n23), .B2(IN0[19]), .ZN(n49) );
  NAND2_X1 U64 ( .A1(n49), .A2(n50), .ZN(OUT1[19]) );
  AOI22_X1 U69 ( .A1(n7), .A2(IN1[18]), .B1(n23), .B2(IN0[18]), .ZN(n51) );
  NAND2_X1 U67 ( .A1(n51), .A2(n52), .ZN(OUT1[18]) );
  AOI22_X1 U72 ( .A1(n7), .A2(IN1[17]), .B1(n23), .B2(IN0[17]), .ZN(n53) );
  NAND2_X1 U70 ( .A1(n53), .A2(n54), .ZN(OUT1[17]) );
  AOI22_X1 U51 ( .A1(n7), .A2(IN1[23]), .B1(n23), .B2(IN0[23]), .ZN(n39) );
  NAND2_X1 U49 ( .A1(n39), .A2(n40), .ZN(OUT1[23]) );
  AOI22_X1 U54 ( .A1(n7), .A2(IN1[22]), .B1(n23), .B2(IN0[22]), .ZN(n41) );
  NAND2_X1 U52 ( .A1(n41), .A2(n42), .ZN(OUT1[22]) );
  AOI22_X1 U57 ( .A1(n7), .A2(IN1[21]), .B1(n23), .B2(IN0[21]), .ZN(n43) );
  NAND2_X1 U55 ( .A1(n43), .A2(n44), .ZN(OUT1[21]) );
  AOI22_X1 U60 ( .A1(n7), .A2(IN1[20]), .B1(n23), .B2(IN0[20]), .ZN(n45) );
  NAND2_X1 U58 ( .A1(n45), .A2(n46), .ZN(OUT1[20]) );
  AOI22_X1 U87 ( .A1(n7), .A2(IN1[12]), .B1(n23), .B2(IN0[12]), .ZN(n63) );
  NAND2_X1 U85 ( .A1(n63), .A2(n64), .ZN(OUT1[12]) );
  AOI22_X1 U90 ( .A1(n7), .A2(IN1[11]), .B1(n23), .B2(IN0[11]), .ZN(n65) );
  NAND2_X1 U88 ( .A1(n65), .A2(n66), .ZN(OUT1[11]) );
  AOI22_X1 U93 ( .A1(n7), .A2(IN1[10]), .B1(n23), .B2(IN0[10]), .ZN(n67) );
  NAND2_X1 U91 ( .A1(n67), .A2(n68), .ZN(OUT1[10]) );
  AOI22_X1 U98 ( .A1(n7), .A2(IN1[0]), .B1(n23), .B2(IN0[0]), .ZN(n69) );
  NAND2_X1 U94 ( .A1(n69), .A2(n70), .ZN(OUT1[0]) );
  AOI22_X1 U75 ( .A1(n7), .A2(IN1[16]), .B1(n23), .B2(IN0[16]), .ZN(n55) );
  NAND2_X1 U73 ( .A1(n55), .A2(n56), .ZN(OUT1[16]) );
  AOI22_X1 U78 ( .A1(n7), .A2(IN1[15]), .B1(n23), .B2(IN0[15]), .ZN(n57) );
  NAND2_X1 U76 ( .A1(n57), .A2(n58), .ZN(OUT1[15]) );
  AOI22_X1 U81 ( .A1(n7), .A2(IN1[14]), .B1(n23), .B2(IN0[14]), .ZN(n59) );
  NAND2_X1 U79 ( .A1(n59), .A2(n60), .ZN(OUT1[14]) );
  AOI22_X1 U84 ( .A1(n7), .A2(IN1[13]), .B1(n23), .B2(IN0[13]), .ZN(n61) );
  NAND2_X1 U82 ( .A1(n61), .A2(n62), .ZN(OUT1[13]) );
  AOI22_X1 U15 ( .A1(n7), .A2(IN1[5]), .B1(n8), .B2(IN0[5]), .ZN(n15) );
  NAND2_X1 U13 ( .A1(n15), .A2(n16), .ZN(OUT1[5]) );
  AOI22_X1 U18 ( .A1(n7), .A2(IN1[4]), .B1(n8), .B2(IN0[4]), .ZN(n17) );
  NAND2_X1 U16 ( .A1(n17), .A2(n18), .ZN(OUT1[4]) );
  AOI22_X1 U21 ( .A1(n7), .A2(IN1[3]), .B1(n8), .B2(IN0[3]), .ZN(n19) );
  NAND2_X1 U19 ( .A1(n19), .A2(n20), .ZN(OUT1[3]) );
  AOI22_X1 U3 ( .A1(n7), .A2(IN1[9]), .B1(n8), .B2(IN0[9]), .ZN(n3) );
  NAND2_X1 U1 ( .A1(n3), .A2(n4), .ZN(OUT1[9]) );
  AOI22_X1 U6 ( .A1(n7), .A2(IN1[8]), .B1(n8), .B2(IN0[8]), .ZN(n9) );
  NAND2_X1 U4 ( .A1(n9), .A2(n10), .ZN(OUT1[8]) );
  AOI22_X1 U9 ( .A1(n7), .A2(IN1[7]), .B1(n23), .B2(IN0[7]), .ZN(n11) );
  NAND2_X1 U7 ( .A1(n11), .A2(n12), .ZN(OUT1[7]) );
  AOI22_X1 U12 ( .A1(n7), .A2(IN1[6]), .B1(n23), .B2(IN0[6]), .ZN(n13) );
  NAND2_X1 U10 ( .A1(n13), .A2(n14), .ZN(OUT1[6]) );
  AOI22_X1 U42 ( .A1(n7), .A2(IN1[26]), .B1(n23), .B2(IN0[26]), .ZN(n33) );
  NAND2_X1 U40 ( .A1(n33), .A2(n34), .ZN(OUT1[26]) );
  AOI22_X1 U45 ( .A1(n7), .A2(IN1[25]), .B1(n23), .B2(IN0[25]), .ZN(n35) );
  NAND2_X1 U43 ( .A1(n35), .A2(n36), .ZN(OUT1[25]) );
  AOI22_X1 U48 ( .A1(n7), .A2(IN1[24]), .B1(n23), .B2(IN0[24]), .ZN(n37) );
  NAND2_X1 U46 ( .A1(n37), .A2(n38), .ZN(OUT1[24]) );
  AOI22_X1 U30 ( .A1(n7), .A2(IN1[2]), .B1(n23), .B2(IN0[2]), .ZN(n25) );
  NAND2_X1 U28 ( .A1(n25), .A2(n26), .ZN(OUT1[2]) );
  INV_X1 U101 ( .A(CTRL[1]), .ZN(n71) );
  AOI222_X1 U2 ( .A1(n6), .A2(IN2[27]), .B1(n23), .B2(IN0[27]), .C1(IN1[27]), 
        .C2(n7), .ZN(n1) );
  INV_X1 U5 ( .A(n1), .ZN(OUT1[27]) );
  AOI222_X1 U8 ( .A1(n6), .A2(IN2[28]), .B1(n23), .B2(IN0[28]), .C1(IN1[28]), 
        .C2(n7), .ZN(n2) );
  INV_X1 U11 ( .A(n2), .ZN(OUT1[28]) );
  AOI222_X1 U14 ( .A1(n6), .A2(IN2[29]), .B1(n23), .B2(IN0[29]), .C1(IN1[29]), 
        .C2(n7), .ZN(n5) );
  INV_X1 U17 ( .A(n5), .ZN(OUT1[29]) );
  AOI222_X1 U20 ( .A1(n6), .A2(IN2[30]), .B1(n23), .B2(IN0[30]), .C1(IN1[30]), 
        .C2(n7), .ZN(n21) );
  INV_X1 U22 ( .A(n21), .ZN(OUT1[30]) );
  AOI222_X1 U23 ( .A1(n6), .A2(IN2[31]), .B1(n23), .B2(IN0[31]), .C1(IN1[31]), 
        .C2(n7), .ZN(n22) );
  INV_X1 U24 ( .A(n22), .ZN(OUT1[31]) );
  AND2_X2 U25 ( .A1(n71), .A2(CTRL[0]), .ZN(n7) );
  BUF_X1 U26 ( .A(n6), .Z(n24) );
  BUF_X2 U27 ( .A(n8), .Z(n23) );
  NOR2_X2 U29 ( .A1(CTRL[0]), .A2(n71), .ZN(n6) );
  NAND2_X1 U31 ( .A1(n6), .A2(IN2[2]), .ZN(n26) );
  NAND2_X1 U32 ( .A1(n6), .A2(IN2[24]), .ZN(n38) );
  NAND2_X1 U33 ( .A1(n6), .A2(IN2[25]), .ZN(n36) );
  NAND2_X1 U34 ( .A1(n6), .A2(IN2[26]), .ZN(n34) );
  NAND2_X1 U35 ( .A1(n24), .A2(IN2[6]), .ZN(n14) );
  NAND2_X1 U36 ( .A1(n24), .A2(IN2[7]), .ZN(n12) );
  NAND2_X1 U37 ( .A1(n24), .A2(IN2[8]), .ZN(n10) );
  NAND2_X1 U38 ( .A1(n24), .A2(IN2[9]), .ZN(n4) );
  NAND2_X1 U39 ( .A1(n24), .A2(IN2[3]), .ZN(n20) );
  NAND2_X1 U41 ( .A1(n24), .A2(IN2[4]), .ZN(n18) );
  NAND2_X1 U44 ( .A1(n24), .A2(IN2[5]), .ZN(n16) );
  NAND2_X1 U47 ( .A1(n24), .A2(IN2[13]), .ZN(n62) );
  NAND2_X1 U50 ( .A1(n24), .A2(IN2[14]), .ZN(n60) );
  NAND2_X1 U53 ( .A1(n24), .A2(IN2[15]), .ZN(n58) );
  NAND2_X1 U56 ( .A1(n24), .A2(IN2[16]), .ZN(n56) );
  NAND2_X1 U59 ( .A1(n24), .A2(IN2[0]), .ZN(n70) );
  NAND2_X1 U62 ( .A1(n6), .A2(IN2[10]), .ZN(n68) );
  NAND2_X1 U65 ( .A1(n24), .A2(IN2[11]), .ZN(n66) );
  NAND2_X1 U68 ( .A1(n24), .A2(IN2[12]), .ZN(n64) );
  NAND2_X1 U71 ( .A1(n6), .A2(IN2[20]), .ZN(n46) );
  NAND2_X1 U74 ( .A1(n6), .A2(IN2[21]), .ZN(n44) );
  NAND2_X1 U77 ( .A1(n24), .A2(IN2[22]), .ZN(n42) );
  NAND2_X1 U80 ( .A1(n24), .A2(IN2[23]), .ZN(n40) );
  NAND2_X1 U83 ( .A1(n6), .A2(IN2[17]), .ZN(n54) );
  NAND2_X1 U86 ( .A1(n6), .A2(IN2[18]), .ZN(n52) );
  NAND2_X1 U89 ( .A1(n24), .A2(IN2[19]), .ZN(n50) );
  NAND2_X1 U92 ( .A1(n24), .A2(IN2[1]), .ZN(n48) );
  NOR2_X1 U95 ( .A1(CTRL[0]), .A2(CTRL[1]), .ZN(n8) );
endmodule


module zerocheck ( IN0, CTRL, OUT1 );
  input [31:0] IN0;
  input CTRL;
  output OUT1;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12;

  NOR4_X1 U12 ( .A1(IN0[1]), .A2(IN0[19]), .A3(IN0[18]), .A4(IN0[17]), .ZN(n9)
         );
  NOR4_X1 U11 ( .A1(IN0[23]), .A2(IN0[22]), .A3(IN0[21]), .A4(IN0[20]), .ZN(
        n10) );
  NOR4_X1 U10 ( .A1(IN0[12]), .A2(IN0[11]), .A3(IN0[10]), .A4(IN0[0]), .ZN(n11) );
  NOR4_X1 U9 ( .A1(IN0[16]), .A2(IN0[15]), .A3(IN0[14]), .A4(IN0[13]), .ZN(n12) );
  NAND4_X1 U8 ( .A1(n9), .A2(n10), .A3(n11), .A4(n12), .ZN(n3) );
  NOR4_X1 U7 ( .A1(IN0[5]), .A2(IN0[4]), .A3(IN0[3]), .A4(IN0[31]), .ZN(n5) );
  NOR4_X1 U6 ( .A1(IN0[9]), .A2(IN0[8]), .A3(IN0[7]), .A4(IN0[6]), .ZN(n6) );
  NOR4_X1 U5 ( .A1(IN0[27]), .A2(IN0[26]), .A3(IN0[25]), .A4(IN0[24]), .ZN(n7)
         );
  NOR4_X1 U4 ( .A1(IN0[30]), .A2(IN0[2]), .A3(IN0[29]), .A4(IN0[28]), .ZN(n8)
         );
  NAND4_X1 U3 ( .A1(n5), .A2(n6), .A3(n7), .A4(n8), .ZN(n4) );
  NOR2_X1 U2 ( .A1(n3), .A2(n4), .ZN(n2) );
  XNOR2_X1 U1 ( .A(CTRL), .B(n2), .ZN(OUT1) );
endmodule


module mux21_0 ( IN0, IN1, CTRL, OUT1 );
  input [31:0] IN0;
  input [31:0] IN1;
  output [31:0] OUT1;
  input CTRL;
  wire   n1;

  MUX2_X1 U1 ( .A(IN0[9]), .B(IN1[9]), .S(n1), .Z(OUT1[9]) );
  MUX2_X1 U2 ( .A(IN0[8]), .B(IN1[8]), .S(n1), .Z(OUT1[8]) );
  MUX2_X1 U3 ( .A(IN0[7]), .B(IN1[7]), .S(n1), .Z(OUT1[7]) );
  MUX2_X1 U4 ( .A(IN0[6]), .B(IN1[6]), .S(n1), .Z(OUT1[6]) );
  MUX2_X1 U5 ( .A(IN0[5]), .B(IN1[5]), .S(CTRL), .Z(OUT1[5]) );
  MUX2_X1 U6 ( .A(IN0[4]), .B(IN1[4]), .S(n1), .Z(OUT1[4]) );
  MUX2_X1 U7 ( .A(IN0[3]), .B(IN1[3]), .S(n1), .Z(OUT1[3]) );
  MUX2_X1 U8 ( .A(IN0[31]), .B(IN1[31]), .S(n1), .Z(OUT1[31]) );
  MUX2_X1 U9 ( .A(IN0[30]), .B(IN1[30]), .S(n1), .Z(OUT1[30]) );
  MUX2_X1 U10 ( .A(IN0[2]), .B(IN1[2]), .S(n1), .Z(OUT1[2]) );
  MUX2_X1 U11 ( .A(IN0[29]), .B(IN1[29]), .S(n1), .Z(OUT1[29]) );
  MUX2_X1 U12 ( .A(IN0[28]), .B(IN1[28]), .S(n1), .Z(OUT1[28]) );
  MUX2_X1 U13 ( .A(IN0[27]), .B(IN1[27]), .S(n1), .Z(OUT1[27]) );
  MUX2_X1 U14 ( .A(IN0[26]), .B(IN1[26]), .S(n1), .Z(OUT1[26]) );
  MUX2_X1 U15 ( .A(IN0[25]), .B(IN1[25]), .S(n1), .Z(OUT1[25]) );
  MUX2_X1 U16 ( .A(IN0[24]), .B(IN1[24]), .S(n1), .Z(OUT1[24]) );
  MUX2_X1 U17 ( .A(IN0[23]), .B(IN1[23]), .S(n1), .Z(OUT1[23]) );
  MUX2_X1 U18 ( .A(IN0[22]), .B(IN1[22]), .S(n1), .Z(OUT1[22]) );
  MUX2_X1 U19 ( .A(IN0[21]), .B(IN1[21]), .S(n1), .Z(OUT1[21]) );
  MUX2_X1 U20 ( .A(IN0[20]), .B(IN1[20]), .S(n1), .Z(OUT1[20]) );
  MUX2_X1 U21 ( .A(IN0[1]), .B(IN1[1]), .S(n1), .Z(OUT1[1]) );
  MUX2_X1 U22 ( .A(IN0[19]), .B(IN1[19]), .S(n1), .Z(OUT1[19]) );
  MUX2_X1 U23 ( .A(IN0[18]), .B(IN1[18]), .S(n1), .Z(OUT1[18]) );
  MUX2_X1 U24 ( .A(IN0[17]), .B(IN1[17]), .S(n1), .Z(OUT1[17]) );
  MUX2_X1 U26 ( .A(IN0[15]), .B(IN1[15]), .S(CTRL), .Z(OUT1[15]) );
  MUX2_X1 U27 ( .A(IN0[14]), .B(IN1[14]), .S(CTRL), .Z(OUT1[14]) );
  MUX2_X1 U28 ( .A(IN0[13]), .B(IN1[13]), .S(CTRL), .Z(OUT1[13]) );
  MUX2_X1 U30 ( .A(IN0[11]), .B(IN1[11]), .S(CTRL), .Z(OUT1[11]) );
  MUX2_X1 U31 ( .A(IN0[10]), .B(IN1[10]), .S(CTRL), .Z(OUT1[10]) );
  MUX2_X1 U25 ( .A(IN0[0]), .B(IN1[0]), .S(CTRL), .Z(OUT1[0]) );
  MUX2_X1 U29 ( .A(IN0[12]), .B(IN1[12]), .S(CTRL), .Z(OUT1[12]) );
  MUX2_X1 U32 ( .A(IN0[16]), .B(IN1[16]), .S(CTRL), .Z(OUT1[16]) );
  BUF_X1 U33 ( .A(CTRL), .Z(n1) );
endmodule


module p4add_N32_logN5_0 ( A, B, Cin, sign, S, Cout );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input Cin, sign;
  output Cout;

  wire   [31:0] new_B;
  wire   [7:0] carry_pro;
  wire   SYNOPSYS_UNCONNECTED__0;

  xor_gen_N32_0 xor32 ( .A(B), .B(1'b0), .S(new_B) );
  carry_tree_N32_logN5_0 ct ( .A({1'b0, 1'b0, 1'b0, 1'b0, A[27:0]}), .B({1'b0, 
        1'b0, 1'b0, 1'b0, new_B[27:0]}), .Cin(1'b0), .Cout({
        SYNOPSYS_UNCONNECTED__0, carry_pro[7:1]}) );
  sum_gen_N32_0 add ( .A(A), .B(new_B), .Cin({1'b0, carry_pro[7:1], 1'b0}), 
        .S(S) );
endmodule


module extender_32 ( IN1, CTRL, SIGN, OUT1 );
  input [31:0] IN1;
  output [31:0] OUT1;
  input CTRL, SIGN;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, \OUT1[28] ;
  assign OUT1[15] = IN1[15];
  assign OUT1[14] = IN1[14];
  assign OUT1[13] = IN1[13];
  assign OUT1[12] = IN1[12];
  assign OUT1[11] = IN1[11];
  assign OUT1[10] = IN1[10];
  assign OUT1[9] = IN1[9];
  assign OUT1[8] = IN1[8];
  assign OUT1[7] = IN1[7];
  assign OUT1[6] = IN1[6];
  assign OUT1[5] = IN1[5];
  assign OUT1[4] = IN1[4];
  assign OUT1[3] = IN1[3];
  assign OUT1[2] = IN1[2];
  assign OUT1[1] = IN1[1];
  assign OUT1[0] = IN1[0];
  assign OUT1[26] = OUT1[27];
  assign OUT1[25] = OUT1[27];
  assign OUT1[29] = OUT1[27];
  assign OUT1[30] = \OUT1[28] ;
  assign OUT1[31] = \OUT1[28] ;
  assign OUT1[28] = \OUT1[28] ;

  NAND2_X1 U3 ( .A1(CTRL), .A2(IN1[25]), .ZN(n4) );
  NAND2_X1 U5 ( .A1(CTRL), .A2(IN1[24]), .ZN(n5) );
  NAND2_X1 U4 ( .A1(n3), .A2(n5), .ZN(OUT1[24]) );
  NAND2_X1 U7 ( .A1(CTRL), .A2(IN1[23]), .ZN(n6) );
  NAND2_X1 U6 ( .A1(n3), .A2(n6), .ZN(OUT1[23]) );
  NAND2_X1 U9 ( .A1(CTRL), .A2(IN1[22]), .ZN(n7) );
  NAND2_X1 U8 ( .A1(n3), .A2(n7), .ZN(OUT1[22]) );
  NAND2_X1 U11 ( .A1(CTRL), .A2(IN1[21]), .ZN(n8) );
  NAND2_X1 U10 ( .A1(n3), .A2(n8), .ZN(OUT1[21]) );
  NAND2_X1 U13 ( .A1(CTRL), .A2(IN1[20]), .ZN(n9) );
  NAND2_X1 U12 ( .A1(n3), .A2(n9), .ZN(OUT1[20]) );
  NAND2_X1 U15 ( .A1(CTRL), .A2(IN1[19]), .ZN(n10) );
  NAND2_X1 U14 ( .A1(n3), .A2(n10), .ZN(OUT1[19]) );
  NAND2_X1 U17 ( .A1(CTRL), .A2(IN1[18]), .ZN(n11) );
  NAND2_X1 U16 ( .A1(n3), .A2(n11), .ZN(OUT1[18]) );
  NAND2_X1 U19 ( .A1(CTRL), .A2(IN1[17]), .ZN(n12) );
  NAND2_X1 U18 ( .A1(n3), .A2(n12), .ZN(OUT1[17]) );
  NAND2_X1 U21 ( .A1(CTRL), .A2(IN1[16]), .ZN(n13) );
  NAND2_X1 U20 ( .A1(n3), .A2(n13), .ZN(OUT1[16]) );
  INV_X1 U22 ( .A(CTRL), .ZN(n14) );
  BUF_X1 U2 ( .A(OUT1[27]), .Z(\OUT1[28] ) );
  NAND2_X2 U23 ( .A1(n3), .A2(n4), .ZN(OUT1[27]) );
  NAND3_X1 U24 ( .A1(SIGN), .A2(IN1[15]), .A3(n14), .ZN(n3) );
endmodule


module ff32_en_IR ( D, en, clk, rst, Q );
  input [31:0] D;
  output [31:0] Q;
  input en, clk, rst;
  wire   net338242, n32;

  DFFR_X1 \Q_reg[31]  ( .D(D[31]), .CK(net338242), .RN(n32), .Q(Q[31]) );
  DFFS_X1 \Q_reg[30]  ( .D(D[30]), .CK(net338242), .SN(n32), .Q(Q[30]) );
  DFFR_X1 \Q_reg[29]  ( .D(D[29]), .CK(net338242), .RN(n32), .Q(Q[29]) );
  DFFS_X1 \Q_reg[28]  ( .D(D[28]), .CK(net338242), .SN(n32), .Q(Q[28]) );
  DFFR_X1 \Q_reg[27]  ( .D(D[27]), .CK(net338242), .RN(n32), .Q(Q[27]) );
  DFFS_X1 \Q_reg[26]  ( .D(D[26]), .CK(net338242), .SN(n32), .Q(Q[26]) );
  DFFR_X1 \Q_reg[25]  ( .D(D[25]), .CK(net338242), .RN(n32), .Q(Q[25]) );
  DFFR_X1 \Q_reg[24]  ( .D(D[24]), .CK(net338242), .RN(n32), .Q(Q[24]) );
  DFFR_X1 \Q_reg[23]  ( .D(D[23]), .CK(net338242), .RN(n32), .Q(Q[23]) );
  DFFR_X1 \Q_reg[22]  ( .D(D[22]), .CK(net338242), .RN(n32), .Q(Q[22]) );
  DFFR_X1 \Q_reg[21]  ( .D(D[21]), .CK(net338242), .RN(n32), .Q(Q[21]) );
  DFFR_X1 \Q_reg[20]  ( .D(D[20]), .CK(net338242), .RN(n32), .Q(Q[20]) );
  DFFR_X1 \Q_reg[19]  ( .D(D[19]), .CK(net338242), .RN(n32), .Q(Q[19]) );
  DFFR_X1 \Q_reg[18]  ( .D(D[18]), .CK(net338242), .RN(n32), .Q(Q[18]) );
  DFFR_X1 \Q_reg[17]  ( .D(D[17]), .CK(net338242), .RN(n32), .Q(Q[17]) );
  DFFR_X1 \Q_reg[16]  ( .D(D[16]), .CK(net338242), .RN(n32), .Q(Q[16]) );
  DFFR_X1 \Q_reg[15]  ( .D(D[15]), .CK(net338242), .RN(n32), .Q(Q[15]) );
  DFFR_X1 \Q_reg[14]  ( .D(D[14]), .CK(net338242), .RN(n32), .Q(Q[14]) );
  DFFR_X1 \Q_reg[13]  ( .D(D[13]), .CK(net338242), .RN(n32), .Q(Q[13]) );
  DFFR_X1 \Q_reg[12]  ( .D(D[12]), .CK(net338242), .RN(n32), .Q(Q[12]) );
  DFFR_X1 \Q_reg[11]  ( .D(D[11]), .CK(net338242), .RN(n32), .Q(Q[11]) );
  DFFR_X1 \Q_reg[10]  ( .D(D[10]), .CK(net338242), .RN(n32), .Q(Q[10]) );
  DFFR_X1 \Q_reg[9]  ( .D(D[9]), .CK(net338242), .RN(n32), .Q(Q[9]) );
  DFFR_X1 \Q_reg[8]  ( .D(D[8]), .CK(net338242), .RN(n32), .Q(Q[8]) );
  DFFR_X1 \Q_reg[7]  ( .D(D[7]), .CK(net338242), .RN(n32), .Q(Q[7]) );
  DFFR_X1 \Q_reg[6]  ( .D(D[6]), .CK(net338242), .RN(n32), .Q(Q[6]) );
  DFFR_X1 \Q_reg[5]  ( .D(D[5]), .CK(net338242), .RN(n32), .Q(Q[5]) );
  DFFR_X1 \Q_reg[4]  ( .D(D[4]), .CK(net338242), .RN(n32), .Q(Q[4]) );
  DFFR_X1 \Q_reg[3]  ( .D(D[3]), .CK(net338242), .RN(n32), .Q(Q[3]) );
  DFFR_X1 \Q_reg[2]  ( .D(D[2]), .CK(net338242), .RN(n32), .Q(Q[2]) );
  DFFR_X1 \Q_reg[1]  ( .D(D[1]), .CK(net338242), .RN(n32), .Q(Q[1]) );
  DFFR_X1 \Q_reg[0]  ( .D(D[0]), .CK(net338242), .RN(n32), .Q(Q[0]) );
  SNPS_CLOCK_GATE_HIGH_ff32_en_IR clk_gate_Q_reg ( .CLK(clk), .EN(en), .ENCLK(
        net338242) );
  INV_X2 U2 ( .A(rst), .ZN(n32) );
endmodule


module SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_0 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net338260, net338262, net338263, net338266;
  assign net338260 = CLK;
  assign ENCLK = net338262;
  assign net338263 = EN;

  DLL_X1 latch ( .D(net338263), .GN(net338260), .Q(net338266) );
  AND2_X1 main_gate ( .A1(net338266), .A2(net338260), .ZN(net338262) );
endmodule


module predictor_2_0 ( clock, reset, enable, taken_i, prediction_o );
  input clock, reset, enable, taken_i;
  output prediction_o;
  wire   N11, N12, n3, n4, n6, n8, n9, n1, n2;
  wire   [1:0] next_STATE;

  DLH_X1 \next_STATE_reg[0]  ( .G(enable), .D(N11), .Q(next_STATE[0]) );
  DFFR_X1 \STATE_reg[0]  ( .D(n8), .CK(clock), .RN(n2), .Q(n1), .QN(n9) );
  DLH_X1 \next_STATE_reg[1]  ( .G(enable), .D(N12), .Q(next_STATE[1]) );
  DFFR_X1 \STATE_reg[1]  ( .D(n6), .CK(clock), .RN(n2), .Q(prediction_o) );
  MUX2_X1 U2 ( .A(prediction_o), .B(next_STATE[1]), .S(enable), .Z(n6) );
  MUX2_X1 U4 ( .A(n1), .B(next_STATE[0]), .S(enable), .Z(n8) );
  NOR2_X1 U9 ( .A1(prediction_o), .A2(taken_i), .ZN(n3) );
  NAND2_X1 U7 ( .A1(prediction_o), .A2(taken_i), .ZN(n4) );
  OAI21_X1 U5 ( .B1(n9), .B2(n3), .A(n4), .ZN(N12) );
  OAI21_X1 U6 ( .B1(n3), .B2(n1), .A(n4), .ZN(N11) );
  INV_X1 U3 ( .A(reset), .ZN(n2) );
endmodule


module mux41_0 ( IN0, IN1, IN2, IN3, CTRL, OUT1 );
  input [31:0] IN0;
  input [31:0] IN1;
  input [31:0] IN2;
  input [31:0] IN3;
  input [1:0] CTRL;
  output [31:0] OUT1;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n57, n58, n59, n60, n61,
         n62, n65, n66, n67, n68, n71, n1, n2, n55, n56, n63, n64, n69, n70,
         n72, n73;

  AOI22_X1 U33 ( .A1(n69), .A2(IN1[29]), .B1(n73), .B2(IN0[29]), .ZN(n27) );
  AOI22_X1 U32 ( .A1(n72), .A2(IN3[29]), .B1(n70), .B2(IN2[29]), .ZN(n28) );
  AOI22_X1 U36 ( .A1(n69), .A2(IN1[28]), .B1(n73), .B2(IN0[28]), .ZN(n29) );
  AOI22_X1 U35 ( .A1(n72), .A2(IN3[28]), .B1(n70), .B2(IN2[28]), .ZN(n30) );
  AOI22_X1 U66 ( .A1(n7), .A2(IN1[19]), .B1(n73), .B2(IN0[19]), .ZN(n49) );
  AOI22_X1 U65 ( .A1(n5), .A2(IN3[19]), .B1(n70), .B2(IN2[19]), .ZN(n50) );
  AOI22_X1 U69 ( .A1(n7), .A2(IN1[18]), .B1(n73), .B2(IN0[18]), .ZN(n51) );
  AOI22_X1 U68 ( .A1(n5), .A2(IN3[18]), .B1(n70), .B2(IN2[18]), .ZN(n52) );
  AOI22_X1 U72 ( .A1(n7), .A2(IN1[17]), .B1(n73), .B2(IN0[17]), .ZN(n53) );
  AOI22_X1 U71 ( .A1(n5), .A2(IN3[17]), .B1(n70), .B2(IN2[17]), .ZN(n54) );
  AOI22_X1 U90 ( .A1(n7), .A2(IN1[11]), .B1(n73), .B2(IN0[11]), .ZN(n65) );
  AOI22_X1 U89 ( .A1(n5), .A2(IN3[11]), .B1(n70), .B2(IN2[11]), .ZN(n66) );
  AOI22_X1 U93 ( .A1(n7), .A2(IN1[10]), .B1(n73), .B2(IN0[10]), .ZN(n67) );
  AOI22_X1 U92 ( .A1(n5), .A2(IN3[10]), .B1(n70), .B2(IN2[10]), .ZN(n68) );
  AOI22_X1 U3 ( .A1(n69), .A2(IN1[9]), .B1(n8), .B2(IN0[9]), .ZN(n3) );
  AOI22_X1 U2 ( .A1(n72), .A2(IN3[9]), .B1(n6), .B2(IN2[9]), .ZN(n4) );
  AOI22_X1 U6 ( .A1(n69), .A2(IN1[8]), .B1(n8), .B2(IN0[8]), .ZN(n9) );
  AOI22_X1 U5 ( .A1(n72), .A2(IN3[8]), .B1(n6), .B2(IN2[8]), .ZN(n10) );
  AOI22_X1 U78 ( .A1(n69), .A2(IN1[15]), .B1(n73), .B2(IN0[15]), .ZN(n57) );
  AOI22_X1 U77 ( .A1(n72), .A2(IN3[15]), .B1(n70), .B2(IN2[15]), .ZN(n58) );
  AOI22_X1 U81 ( .A1(n69), .A2(IN1[14]), .B1(n73), .B2(IN0[14]), .ZN(n59) );
  AOI22_X1 U80 ( .A1(n72), .A2(IN3[14]), .B1(n70), .B2(IN2[14]), .ZN(n60) );
  AOI22_X1 U84 ( .A1(n69), .A2(IN1[13]), .B1(n73), .B2(IN0[13]), .ZN(n61) );
  AOI22_X1 U83 ( .A1(n72), .A2(IN3[13]), .B1(n70), .B2(IN2[13]), .ZN(n62) );
  AOI22_X1 U21 ( .A1(n69), .A2(IN1[3]), .B1(n8), .B2(IN0[3]), .ZN(n19) );
  AOI22_X1 U20 ( .A1(n72), .A2(IN3[3]), .B1(n6), .B2(IN2[3]), .ZN(n20) );
  AOI22_X1 U30 ( .A1(n69), .A2(IN1[2]), .B1(n73), .B2(IN0[2]), .ZN(n25) );
  AOI22_X1 U29 ( .A1(n72), .A2(IN3[2]), .B1(n70), .B2(IN2[2]), .ZN(n26) );
  AOI22_X1 U63 ( .A1(n69), .A2(IN1[1]), .B1(n73), .B2(IN0[1]), .ZN(n47) );
  AOI22_X1 U62 ( .A1(n72), .A2(IN3[1]), .B1(n70), .B2(IN2[1]), .ZN(n48) );
  AOI22_X1 U9 ( .A1(n69), .A2(IN1[7]), .B1(n73), .B2(IN0[7]), .ZN(n11) );
  AOI22_X1 U8 ( .A1(n72), .A2(IN3[7]), .B1(n70), .B2(IN2[7]), .ZN(n12) );
  AOI22_X1 U12 ( .A1(n69), .A2(IN1[6]), .B1(n73), .B2(IN0[6]), .ZN(n13) );
  AOI22_X1 U11 ( .A1(n72), .A2(IN3[6]), .B1(n70), .B2(IN2[6]), .ZN(n14) );
  AOI22_X1 U15 ( .A1(n69), .A2(IN1[5]), .B1(n73), .B2(IN0[5]), .ZN(n15) );
  AOI22_X1 U14 ( .A1(n72), .A2(IN3[5]), .B1(n70), .B2(IN2[5]), .ZN(n16) );
  AOI22_X1 U18 ( .A1(n69), .A2(IN1[4]), .B1(n73), .B2(IN0[4]), .ZN(n17) );
  AOI22_X1 U17 ( .A1(n72), .A2(IN3[4]), .B1(n70), .B2(IN2[4]), .ZN(n18) );
  AOI22_X1 U51 ( .A1(n69), .A2(IN1[23]), .B1(n73), .B2(IN0[23]), .ZN(n39) );
  AOI22_X1 U50 ( .A1(n72), .A2(IN3[23]), .B1(n70), .B2(IN2[23]), .ZN(n40) );
  AOI22_X1 U54 ( .A1(n69), .A2(IN1[22]), .B1(n73), .B2(IN0[22]), .ZN(n41) );
  AOI22_X1 U53 ( .A1(n72), .A2(IN3[22]), .B1(n70), .B2(IN2[22]), .ZN(n42) );
  AOI22_X1 U24 ( .A1(n69), .A2(IN1[31]), .B1(n8), .B2(IN0[31]), .ZN(n21) );
  AOI22_X1 U23 ( .A1(n72), .A2(IN3[31]), .B1(n70), .B2(IN2[31]), .ZN(n22) );
  AOI22_X1 U27 ( .A1(n69), .A2(IN1[30]), .B1(n73), .B2(IN0[30]), .ZN(n23) );
  AOI22_X1 U26 ( .A1(n72), .A2(IN3[30]), .B1(n70), .B2(IN2[30]), .ZN(n24) );
  AOI22_X1 U39 ( .A1(n69), .A2(IN1[27]), .B1(n73), .B2(IN0[27]), .ZN(n31) );
  AOI22_X1 U38 ( .A1(n72), .A2(IN3[27]), .B1(n70), .B2(IN2[27]), .ZN(n32) );
  AOI22_X1 U42 ( .A1(n69), .A2(IN1[26]), .B1(n73), .B2(IN0[26]), .ZN(n33) );
  AOI22_X1 U41 ( .A1(n72), .A2(IN3[26]), .B1(n70), .B2(IN2[26]), .ZN(n34) );
  AOI22_X1 U45 ( .A1(n69), .A2(IN1[25]), .B1(n73), .B2(IN0[25]), .ZN(n35) );
  AOI22_X1 U44 ( .A1(n72), .A2(IN3[25]), .B1(n70), .B2(IN2[25]), .ZN(n36) );
  AOI22_X1 U48 ( .A1(n69), .A2(IN1[24]), .B1(n73), .B2(IN0[24]), .ZN(n37) );
  AOI22_X1 U47 ( .A1(n72), .A2(IN3[24]), .B1(n70), .B2(IN2[24]), .ZN(n38) );
  AOI22_X1 U57 ( .A1(n69), .A2(IN1[21]), .B1(n73), .B2(IN0[21]), .ZN(n43) );
  AOI22_X1 U56 ( .A1(n72), .A2(IN3[21]), .B1(n70), .B2(IN2[21]), .ZN(n44) );
  AOI22_X1 U60 ( .A1(n69), .A2(IN1[20]), .B1(n73), .B2(IN0[20]), .ZN(n45) );
  AOI22_X1 U59 ( .A1(n72), .A2(IN3[20]), .B1(n70), .B2(IN2[20]), .ZN(n46) );
  NAND2_X1 U88 ( .A1(n65), .A2(n66), .ZN(OUT1[11]) );
  NAND2_X1 U91 ( .A1(n67), .A2(n68), .ZN(OUT1[10]) );
  NAND2_X1 U76 ( .A1(n57), .A2(n58), .ZN(OUT1[15]) );
  NAND2_X1 U79 ( .A1(n59), .A2(n60), .ZN(OUT1[14]) );
  NAND2_X1 U82 ( .A1(n61), .A2(n62), .ZN(OUT1[13]) );
  NAND2_X1 U13 ( .A1(n15), .A2(n16), .ZN(OUT1[5]) );
  NAND2_X1 U52 ( .A1(n41), .A2(n42), .ZN(OUT1[22]) );
  NAND2_X1 U31 ( .A1(n27), .A2(n28), .ZN(OUT1[29]) );
  NAND2_X1 U34 ( .A1(n29), .A2(n30), .ZN(OUT1[28]) );
  NAND2_X1 U64 ( .A1(n49), .A2(n50), .ZN(OUT1[19]) );
  NAND2_X1 U67 ( .A1(n51), .A2(n52), .ZN(OUT1[18]) );
  NAND2_X1 U70 ( .A1(n53), .A2(n54), .ZN(OUT1[17]) );
  NAND2_X1 U1 ( .A1(n3), .A2(n4), .ZN(OUT1[9]) );
  NAND2_X1 U4 ( .A1(n9), .A2(n10), .ZN(OUT1[8]) );
  NAND2_X1 U19 ( .A1(n19), .A2(n20), .ZN(OUT1[3]) );
  NAND2_X1 U28 ( .A1(n25), .A2(n26), .ZN(OUT1[2]) );
  NAND2_X1 U61 ( .A1(n47), .A2(n48), .ZN(OUT1[1]) );
  NAND2_X1 U7 ( .A1(n11), .A2(n12), .ZN(OUT1[7]) );
  NAND2_X1 U10 ( .A1(n13), .A2(n14), .ZN(OUT1[6]) );
  NAND2_X1 U16 ( .A1(n17), .A2(n18), .ZN(OUT1[4]) );
  NAND2_X1 U49 ( .A1(n39), .A2(n40), .ZN(OUT1[23]) );
  NAND2_X1 U22 ( .A1(n21), .A2(n22), .ZN(OUT1[31]) );
  NAND2_X1 U25 ( .A1(n23), .A2(n24), .ZN(OUT1[30]) );
  NAND2_X1 U37 ( .A1(n31), .A2(n32), .ZN(OUT1[27]) );
  NAND2_X1 U40 ( .A1(n33), .A2(n34), .ZN(OUT1[26]) );
  NAND2_X1 U43 ( .A1(n35), .A2(n36), .ZN(OUT1[25]) );
  NAND2_X1 U46 ( .A1(n37), .A2(n38), .ZN(OUT1[24]) );
  NAND2_X1 U55 ( .A1(n43), .A2(n44), .ZN(OUT1[21]) );
  NAND2_X1 U58 ( .A1(n45), .A2(n46), .ZN(OUT1[20]) );
  INV_X1 U101 ( .A(CTRL[1]), .ZN(n71) );
  AOI22_X1 U73 ( .A1(IN2[0]), .A2(n70), .B1(IN3[0]), .B2(n72), .ZN(n1) );
  AOI22_X1 U74 ( .A1(IN0[0]), .A2(n73), .B1(IN1[0]), .B2(n69), .ZN(n2) );
  NAND2_X1 U75 ( .A1(n1), .A2(n2), .ZN(OUT1[0]) );
  AOI22_X1 U85 ( .A1(IN2[12]), .A2(n70), .B1(IN3[12]), .B2(n72), .ZN(n55) );
  AOI22_X1 U86 ( .A1(IN0[12]), .A2(n73), .B1(IN1[12]), .B2(n69), .ZN(n56) );
  NAND2_X1 U87 ( .A1(n55), .A2(n56), .ZN(OUT1[12]) );
  AOI22_X1 U94 ( .A1(IN2[16]), .A2(n70), .B1(IN3[16]), .B2(n5), .ZN(n63) );
  AOI22_X1 U95 ( .A1(IN0[16]), .A2(n73), .B1(IN1[16]), .B2(n7), .ZN(n64) );
  NAND2_X1 U96 ( .A1(n63), .A2(n64), .ZN(OUT1[16]) );
  BUF_X2 U97 ( .A(n7), .Z(n69) );
  BUF_X2 U98 ( .A(n6), .Z(n70) );
  BUF_X2 U99 ( .A(n5), .Z(n72) );
  BUF_X2 U100 ( .A(n8), .Z(n73) );
  AND2_X1 U102 ( .A1(CTRL[0]), .A2(CTRL[1]), .ZN(n5) );
  AND2_X1 U103 ( .A1(n71), .A2(CTRL[0]), .ZN(n7) );
  NOR2_X1 U104 ( .A1(CTRL[0]), .A2(n71), .ZN(n6) );
  NOR2_X1 U105 ( .A1(CTRL[0]), .A2(CTRL[1]), .ZN(n8) );
endmodule


module add4 ( IN1, OUT1 );
  input [31:0] IN1;
  output [31:0] OUT1;
  wire   \IN1[1] , \IN1[0] , \add_27/carry[4] , \add_27/carry[5] ,
         \add_27/carry[6] , \add_27/carry[7] , \add_27/carry[8] ,
         \add_27/carry[9] , \add_27/carry[10] , \add_27/carry[11] ,
         \add_27/carry[12] , \add_27/carry[13] , \add_27/carry[14] ,
         \add_27/carry[15] , \add_27/carry[16] , \add_27/carry[17] ,
         \add_27/carry[18] , \add_27/carry[19] , \add_27/carry[20] ,
         \add_27/carry[21] , \add_27/carry[22] , \add_27/carry[23] ,
         \add_27/carry[24] , \add_27/carry[25] , \add_27/carry[26] ,
         \add_27/carry[27] , \add_27/carry[28] , \add_27/carry[29] ,
         \add_27/carry[30] , n1;
  assign OUT1[1] = \IN1[1] ;
  assign \IN1[1]  = IN1[1];
  assign OUT1[0] = \IN1[0] ;
  assign \IN1[0]  = IN1[0];

  NAND2_X1 U3 ( .A1(\add_27/carry[30] ), .A2(IN1[30]), .ZN(n1) );
  XNOR2_X1 U4 ( .A(n1), .B(IN1[31]), .ZN(OUT1[31]) );
  INV_X1 U5 ( .A(IN1[2]), .ZN(OUT1[2]) );
  XOR2_X1 U6 ( .A(IN1[3]), .B(IN1[2]), .Z(OUT1[3]) );
  XOR2_X1 U7 ( .A(IN1[4]), .B(\add_27/carry[4] ), .Z(OUT1[4]) );
  XOR2_X1 U8 ( .A(IN1[5]), .B(\add_27/carry[5] ), .Z(OUT1[5]) );
  XOR2_X1 U9 ( .A(IN1[6]), .B(\add_27/carry[6] ), .Z(OUT1[6]) );
  XOR2_X1 U10 ( .A(IN1[7]), .B(\add_27/carry[7] ), .Z(OUT1[7]) );
  XOR2_X1 U11 ( .A(IN1[8]), .B(\add_27/carry[8] ), .Z(OUT1[8]) );
  XOR2_X1 U12 ( .A(IN1[9]), .B(\add_27/carry[9] ), .Z(OUT1[9]) );
  XOR2_X1 U13 ( .A(IN1[10]), .B(\add_27/carry[10] ), .Z(OUT1[10]) );
  XOR2_X1 U14 ( .A(IN1[11]), .B(\add_27/carry[11] ), .Z(OUT1[11]) );
  XOR2_X1 U15 ( .A(IN1[12]), .B(\add_27/carry[12] ), .Z(OUT1[12]) );
  XOR2_X1 U16 ( .A(IN1[13]), .B(\add_27/carry[13] ), .Z(OUT1[13]) );
  XOR2_X1 U17 ( .A(IN1[14]), .B(\add_27/carry[14] ), .Z(OUT1[14]) );
  XOR2_X1 U18 ( .A(IN1[15]), .B(\add_27/carry[15] ), .Z(OUT1[15]) );
  XOR2_X1 U19 ( .A(IN1[16]), .B(\add_27/carry[16] ), .Z(OUT1[16]) );
  XOR2_X1 U20 ( .A(IN1[17]), .B(\add_27/carry[17] ), .Z(OUT1[17]) );
  XOR2_X1 U21 ( .A(IN1[18]), .B(\add_27/carry[18] ), .Z(OUT1[18]) );
  XOR2_X1 U22 ( .A(IN1[19]), .B(\add_27/carry[19] ), .Z(OUT1[19]) );
  XOR2_X1 U23 ( .A(IN1[20]), .B(\add_27/carry[20] ), .Z(OUT1[20]) );
  XOR2_X1 U24 ( .A(IN1[21]), .B(\add_27/carry[21] ), .Z(OUT1[21]) );
  XOR2_X1 U25 ( .A(IN1[22]), .B(\add_27/carry[22] ), .Z(OUT1[22]) );
  XOR2_X1 U26 ( .A(IN1[23]), .B(\add_27/carry[23] ), .Z(OUT1[23]) );
  XOR2_X1 U27 ( .A(IN1[24]), .B(\add_27/carry[24] ), .Z(OUT1[24]) );
  XOR2_X1 U28 ( .A(IN1[25]), .B(\add_27/carry[25] ), .Z(OUT1[25]) );
  XOR2_X1 U29 ( .A(IN1[26]), .B(\add_27/carry[26] ), .Z(OUT1[26]) );
  XOR2_X1 U30 ( .A(IN1[27]), .B(\add_27/carry[27] ), .Z(OUT1[27]) );
  XOR2_X1 U31 ( .A(IN1[28]), .B(\add_27/carry[28] ), .Z(OUT1[28]) );
  XOR2_X1 U32 ( .A(IN1[29]), .B(\add_27/carry[29] ), .Z(OUT1[29]) );
  XOR2_X1 U33 ( .A(IN1[30]), .B(\add_27/carry[30] ), .Z(OUT1[30]) );
  AND2_X1 U34 ( .A1(IN1[2]), .A2(IN1[3]), .ZN(\add_27/carry[4] ) );
  AND2_X1 U35 ( .A1(\add_27/carry[4] ), .A2(IN1[4]), .ZN(\add_27/carry[5] ) );
  AND2_X1 U36 ( .A1(\add_27/carry[5] ), .A2(IN1[5]), .ZN(\add_27/carry[6] ) );
  AND2_X1 U37 ( .A1(\add_27/carry[6] ), .A2(IN1[6]), .ZN(\add_27/carry[7] ) );
  AND2_X1 U38 ( .A1(\add_27/carry[7] ), .A2(IN1[7]), .ZN(\add_27/carry[8] ) );
  AND2_X1 U39 ( .A1(\add_27/carry[8] ), .A2(IN1[8]), .ZN(\add_27/carry[9] ) );
  AND2_X1 U40 ( .A1(\add_27/carry[9] ), .A2(IN1[9]), .ZN(\add_27/carry[10] )
         );
  AND2_X1 U41 ( .A1(\add_27/carry[10] ), .A2(IN1[10]), .ZN(\add_27/carry[11] )
         );
  AND2_X1 U42 ( .A1(\add_27/carry[11] ), .A2(IN1[11]), .ZN(\add_27/carry[12] )
         );
  AND2_X1 U43 ( .A1(\add_27/carry[12] ), .A2(IN1[12]), .ZN(\add_27/carry[13] )
         );
  AND2_X1 U44 ( .A1(\add_27/carry[13] ), .A2(IN1[13]), .ZN(\add_27/carry[14] )
         );
  AND2_X1 U45 ( .A1(\add_27/carry[14] ), .A2(IN1[14]), .ZN(\add_27/carry[15] )
         );
  AND2_X1 U46 ( .A1(\add_27/carry[15] ), .A2(IN1[15]), .ZN(\add_27/carry[16] )
         );
  AND2_X1 U47 ( .A1(\add_27/carry[16] ), .A2(IN1[16]), .ZN(\add_27/carry[17] )
         );
  AND2_X1 U48 ( .A1(\add_27/carry[17] ), .A2(IN1[17]), .ZN(\add_27/carry[18] )
         );
  AND2_X1 U49 ( .A1(\add_27/carry[18] ), .A2(IN1[18]), .ZN(\add_27/carry[19] )
         );
  AND2_X1 U50 ( .A1(\add_27/carry[19] ), .A2(IN1[19]), .ZN(\add_27/carry[20] )
         );
  AND2_X1 U51 ( .A1(\add_27/carry[20] ), .A2(IN1[20]), .ZN(\add_27/carry[21] )
         );
  AND2_X1 U52 ( .A1(\add_27/carry[21] ), .A2(IN1[21]), .ZN(\add_27/carry[22] )
         );
  AND2_X1 U53 ( .A1(\add_27/carry[22] ), .A2(IN1[22]), .ZN(\add_27/carry[23] )
         );
  AND2_X1 U54 ( .A1(\add_27/carry[23] ), .A2(IN1[23]), .ZN(\add_27/carry[24] )
         );
  AND2_X1 U55 ( .A1(\add_27/carry[24] ), .A2(IN1[24]), .ZN(\add_27/carry[25] )
         );
  AND2_X1 U56 ( .A1(\add_27/carry[25] ), .A2(IN1[25]), .ZN(\add_27/carry[26] )
         );
  AND2_X1 U57 ( .A1(\add_27/carry[26] ), .A2(IN1[26]), .ZN(\add_27/carry[27] )
         );
  AND2_X1 U58 ( .A1(\add_27/carry[27] ), .A2(IN1[27]), .ZN(\add_27/carry[28] )
         );
  AND2_X1 U59 ( .A1(\add_27/carry[28] ), .A2(IN1[28]), .ZN(\add_27/carry[29] )
         );
  AND2_X1 U60 ( .A1(\add_27/carry[29] ), .A2(IN1[29]), .ZN(\add_27/carry[30] )
         );
endmodule


module ff32_en_0 ( D, en, clk, rst, Q );
  input [31:0] D;
  output [31:0] Q;
  input en, clk, rst;
  wire   net338257, n32;

  DFFR_X1 \Q_reg[31]  ( .D(D[31]), .CK(net338257), .RN(n32), .Q(Q[31]) );
  DFFR_X1 \Q_reg[30]  ( .D(D[30]), .CK(net338257), .RN(n32), .Q(Q[30]) );
  DFFR_X1 \Q_reg[29]  ( .D(D[29]), .CK(net338257), .RN(n32), .Q(Q[29]) );
  DFFR_X1 \Q_reg[28]  ( .D(D[28]), .CK(net338257), .RN(n32), .Q(Q[28]) );
  DFFR_X1 \Q_reg[27]  ( .D(D[27]), .CK(net338257), .RN(n32), .Q(Q[27]) );
  DFFR_X1 \Q_reg[26]  ( .D(D[26]), .CK(net338257), .RN(n32), .Q(Q[26]) );
  DFFR_X1 \Q_reg[25]  ( .D(D[25]), .CK(net338257), .RN(n32), .Q(Q[25]) );
  DFFR_X1 \Q_reg[24]  ( .D(D[24]), .CK(net338257), .RN(n32), .Q(Q[24]) );
  DFFR_X1 \Q_reg[23]  ( .D(D[23]), .CK(net338257), .RN(n32), .Q(Q[23]) );
  DFFR_X1 \Q_reg[22]  ( .D(D[22]), .CK(net338257), .RN(n32), .Q(Q[22]) );
  DFFR_X1 \Q_reg[21]  ( .D(D[21]), .CK(net338257), .RN(n32), .Q(Q[21]) );
  DFFR_X1 \Q_reg[20]  ( .D(D[20]), .CK(net338257), .RN(n32), .Q(Q[20]) );
  DFFR_X1 \Q_reg[19]  ( .D(D[19]), .CK(net338257), .RN(n32), .Q(Q[19]) );
  DFFR_X1 \Q_reg[18]  ( .D(D[18]), .CK(net338257), .RN(n32), .Q(Q[18]) );
  DFFR_X1 \Q_reg[17]  ( .D(D[17]), .CK(net338257), .RN(n32), .Q(Q[17]) );
  DFFR_X1 \Q_reg[16]  ( .D(D[16]), .CK(net338257), .RN(n32), .Q(Q[16]) );
  DFFR_X1 \Q_reg[15]  ( .D(D[15]), .CK(net338257), .RN(n32), .Q(Q[15]) );
  DFFR_X1 \Q_reg[14]  ( .D(D[14]), .CK(net338257), .RN(n32), .Q(Q[14]) );
  DFFR_X1 \Q_reg[13]  ( .D(D[13]), .CK(net338257), .RN(n32), .Q(Q[13]) );
  DFFR_X1 \Q_reg[12]  ( .D(D[12]), .CK(net338257), .RN(n32), .Q(Q[12]) );
  DFFR_X1 \Q_reg[11]  ( .D(D[11]), .CK(net338257), .RN(n32), .Q(Q[11]) );
  DFFR_X1 \Q_reg[10]  ( .D(D[10]), .CK(net338257), .RN(n32), .Q(Q[10]) );
  DFFR_X1 \Q_reg[9]  ( .D(D[9]), .CK(net338257), .RN(n32), .Q(Q[9]) );
  DFFR_X1 \Q_reg[8]  ( .D(D[8]), .CK(net338257), .RN(n32), .Q(Q[8]) );
  DFFR_X1 \Q_reg[7]  ( .D(D[7]), .CK(net338257), .RN(n32), .Q(Q[7]) );
  DFFR_X1 \Q_reg[6]  ( .D(D[6]), .CK(net338257), .RN(n32), .Q(Q[6]) );
  DFFR_X1 \Q_reg[5]  ( .D(D[5]), .CK(net338257), .RN(n32), .Q(Q[5]) );
  DFFR_X1 \Q_reg[4]  ( .D(D[4]), .CK(net338257), .RN(n32), .Q(Q[4]) );
  DFFR_X1 \Q_reg[3]  ( .D(D[3]), .CK(net338257), .RN(n32), .Q(Q[3]) );
  DFFR_X1 \Q_reg[2]  ( .D(D[2]), .CK(net338257), .RN(n32), .Q(Q[2]) );
  DFFR_X1 \Q_reg[1]  ( .D(D[1]), .CK(net338257), .RN(n32), .Q(Q[1]) );
  DFFR_X1 \Q_reg[0]  ( .D(D[0]), .CK(net338257), .RN(n32), .Q(Q[0]) );
  SNPS_CLOCK_GATE_HIGH_ff32_en_0 clk_gate_Q_reg ( .CLK(clk), .EN(en), .ENCLK(
        net338257) );
  INV_X2 U2 ( .A(rst), .ZN(n32) );
endmodule


module fw_logic ( D1_i, rAdec_i, D2_i, D3_i, rA_i, rB_i, S_mem_W, S_mem_LOAD, 
        S_wb_W, S_exe_W, S_FWAdec, S_FWA, S_FWB );
  input [4:0] D1_i;
  input [4:0] rAdec_i;
  input [4:0] D2_i;
  input [4:0] D3_i;
  input [4:0] rA_i;
  input [4:0] rB_i;
  output [1:0] S_FWAdec;
  output [1:0] S_FWA;
  output [1:0] S_FWB;
  input S_mem_W, S_mem_LOAD, S_wb_W, S_exe_W;
  wire   n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n1;

  XOR2_X1 U53 ( .A(D2_i[4]), .B(rB_i[4]), .Z(n30) );
  XOR2_X1 U54 ( .A(D2_i[4]), .B(rAdec_i[4]), .Z(n46) );
  XOR2_X1 U55 ( .A(D2_i[4]), .B(rA_i[4]), .Z(n61) );
  AOI22_X1 U13 ( .A1(n37), .A2(rB_i[3]), .B1(rB_i[1]), .B2(n38), .ZN(n39) );
  OAI221_X1 U12 ( .B1(n37), .B2(rB_i[3]), .C1(n38), .C2(rB_i[1]), .A(n39), 
        .ZN(n32) );
  AOI22_X1 U11 ( .A1(n34), .A2(rB_i[0]), .B1(rB_i[2]), .B2(n35), .ZN(n36) );
  OAI221_X1 U10 ( .B1(n34), .B2(rB_i[0]), .C1(n35), .C2(rB_i[2]), .A(n36), 
        .ZN(n33) );
  OAI221_X1 U7 ( .B1(D3_i[4]), .B2(n28), .C1(n29), .C2(rB_i[4]), .A(S_wb_W), 
        .ZN(n19) );
  AOI22_X1 U6 ( .A1(n25), .A2(rB_i[3]), .B1(rB_i[1]), .B2(n26), .ZN(n27) );
  OAI221_X1 U5 ( .B1(n25), .B2(rB_i[3]), .C1(n26), .C2(rB_i[1]), .A(n27), .ZN(
        n20) );
  AOI22_X1 U4 ( .A1(n22), .A2(rB_i[0]), .B1(rB_i[2]), .B2(n23), .ZN(n24) );
  OAI221_X1 U3 ( .B1(n22), .B2(rB_i[0]), .C1(n23), .C2(rB_i[2]), .A(n24), .ZN(
        n21) );
  AOI22_X1 U48 ( .A1(n37), .A2(rA_i[3]), .B1(rA_i[1]), .B2(n38), .ZN(n65) );
  OAI221_X1 U47 ( .B1(n37), .B2(rA_i[3]), .C1(n38), .C2(rA_i[1]), .A(n65), 
        .ZN(n62) );
  AOI22_X1 U44 ( .A1(n34), .A2(rA_i[0]), .B1(rA_i[2]), .B2(n35), .ZN(n64) );
  OAI221_X1 U43 ( .B1(n34), .B2(rA_i[0]), .C1(n35), .C2(rA_i[2]), .A(n64), 
        .ZN(n63) );
  OAI221_X1 U39 ( .B1(rA_i[4]), .B2(n29), .C1(n60), .C2(D3_i[4]), .A(S_wb_W), 
        .ZN(n51) );
  AOI22_X1 U36 ( .A1(n57), .A2(D3_i[3]), .B1(D3_i[1]), .B2(n58), .ZN(n59) );
  OAI221_X1 U35 ( .B1(n57), .B2(D3_i[3]), .C1(n58), .C2(D3_i[1]), .A(n59), 
        .ZN(n52) );
  AOI22_X1 U32 ( .A1(n54), .A2(D3_i[0]), .B1(D3_i[2]), .B2(n55), .ZN(n56) );
  OAI221_X1 U31 ( .B1(n54), .B2(D3_i[0]), .C1(n55), .C2(D3_i[2]), .A(n56), 
        .ZN(n53) );
  AOI22_X1 U29 ( .A1(n37), .A2(rAdec_i[3]), .B1(rAdec_i[1]), .B2(n38), .ZN(n50) );
  OAI221_X1 U28 ( .B1(n37), .B2(rAdec_i[3]), .C1(n38), .C2(rAdec_i[1]), .A(n50), .ZN(n47) );
  AOI22_X1 U27 ( .A1(n34), .A2(rAdec_i[0]), .B1(rAdec_i[2]), .B2(n35), .ZN(n49) );
  OAI221_X1 U26 ( .B1(n34), .B2(rAdec_i[0]), .C1(n35), .C2(rAdec_i[2]), .A(n49), .ZN(n48) );
  OAI221_X1 U23 ( .B1(D3_i[4]), .B2(n45), .C1(n29), .C2(rAdec_i[4]), .A(S_wb_W), .ZN(n40) );
  AOI22_X1 U20 ( .A1(n25), .A2(rAdec_i[3]), .B1(rAdec_i[1]), .B2(n26), .ZN(n44) );
  OAI221_X1 U19 ( .B1(n25), .B2(rAdec_i[3]), .C1(n26), .C2(rAdec_i[1]), .A(n44), .ZN(n41) );
  AOI22_X1 U16 ( .A1(n22), .A2(rAdec_i[0]), .B1(rAdec_i[2]), .B2(n23), .ZN(n43) );
  OAI221_X1 U15 ( .B1(n22), .B2(rAdec_i[0]), .C1(n23), .C2(rAdec_i[2]), .A(n43), .ZN(n42) );
  NOR4_X1 U14 ( .A1(S_FWAdec[0]), .A2(n40), .A3(n41), .A4(n42), .ZN(
        S_FWAdec[1]) );
  NAND2_X1 U51 ( .A1(S_mem_W), .A2(n1), .ZN(n31) );
  INV_X1 U50 ( .A(D2_i[3]), .ZN(n37) );
  INV_X1 U49 ( .A(D2_i[1]), .ZN(n38) );
  NOR4_X1 U30 ( .A1(S_FWA[0]), .A2(n51), .A3(n52), .A4(n53), .ZN(S_FWA[1]) );
  INV_X1 U46 ( .A(D2_i[0]), .ZN(n34) );
  INV_X1 U45 ( .A(D2_i[2]), .ZN(n35) );
  NOR4_X1 U2 ( .A1(S_FWB[0]), .A2(n19), .A3(n20), .A4(n21), .ZN(S_FWB[1]) );
  NOR4_X1 U42 ( .A1(n61), .A2(n31), .A3(n62), .A4(n63), .ZN(S_FWA[0]) );
  NOR4_X1 U25 ( .A1(n46), .A2(n31), .A3(n47), .A4(n48), .ZN(S_FWAdec[0]) );
  INV_X1 U8 ( .A(rB_i[4]), .ZN(n28) );
  INV_X1 U41 ( .A(D3_i[4]), .ZN(n29) );
  INV_X1 U22 ( .A(D3_i[3]), .ZN(n25) );
  INV_X1 U21 ( .A(D3_i[1]), .ZN(n26) );
  INV_X1 U18 ( .A(D3_i[0]), .ZN(n22) );
  INV_X1 U17 ( .A(D3_i[2]), .ZN(n23) );
  INV_X1 U40 ( .A(rA_i[4]), .ZN(n60) );
  INV_X1 U38 ( .A(rA_i[3]), .ZN(n57) );
  INV_X1 U37 ( .A(rA_i[1]), .ZN(n58) );
  INV_X1 U34 ( .A(rA_i[0]), .ZN(n54) );
  INV_X1 U33 ( .A(rA_i[2]), .ZN(n55) );
  INV_X1 U24 ( .A(rAdec_i[4]), .ZN(n45) );
  NOR4_X1 U9 ( .A1(n30), .A2(n31), .A3(n32), .A4(n33), .ZN(S_FWB[0]) );
  INV_X1 U52 ( .A(S_mem_LOAD), .ZN(n1) );
endmodule


module mem_block ( X_i, LOAD_i, S_MUX_MEM_i, W_o );
  input [31:0] X_i;
  input [31:0] LOAD_i;
  output [31:0] W_o;
  input S_MUX_MEM_i;


  mux21_2 MUXMEM ( .IN0(X_i), .IN1(LOAD_i), .CTRL(S_MUX_MEM_i), .OUT1(W_o) );
endmodule


module mem_regs ( W_i, D3_i, W_o, D3_o, clk, rst );
  input [31:0] W_i;
  input [4:0] D3_i;
  output [31:0] W_o;
  output [4:0] D3_o;
  input clk, rst;


  ff32_SIZE32 W ( .D(W_i), .clk(clk), .rst(rst), .Q(W_o) );
  ff32_SIZE5 D3 ( .D(D3_i), .clk(clk), .rst(rst), .Q(D3_o) );
endmodule


module execute_block ( IMM_i, A_i, rB_i, rC_i, MUXED_B_i, S_MUX_ALUIN_i, 
        FW_X_i, FW_W_i, S_FW_A_i, S_FW_B_i, muxed_dest, muxed_B, S_MUX_DEST_i, 
    .OP({\OP[4] , \OP[3] , \OP[2] , \OP[1] , \OP[0] }), ALUW_i, DOUT, stall_o, 
        Clock, Reset );
  input [31:0] IMM_i;
  input [31:0] A_i;
  input [4:0] rB_i;
  input [4:0] rC_i;
  input [31:0] MUXED_B_i;
  input [31:0] FW_X_i;
  input [31:0] FW_W_i;
  input [1:0] S_FW_A_i;
  input [1:0] S_FW_B_i;
  output [4:0] muxed_dest;
  output [31:0] muxed_B;
  input [1:0] S_MUX_DEST_i;
  input [12:0] ALUW_i;
  output [31:0] DOUT;
  input S_MUX_ALUIN_i, \OP[4] , \OP[3] , \OP[2] , \OP[1] , \OP[0] , Clock,
         Reset;
  output stall_o;

  wire   [31:0] FWB2alu;
  wire   [31:0] FWA2alu;

  mux21_3 ALUIN_MUX ( .IN0(muxed_B), .IN1(IMM_i), .CTRL(S_MUX_ALUIN_i), .OUT1(
        FWB2alu) );
  real_alu_DATA_SIZE32 ALU ( .IN1(FWA2alu), .IN2(FWB2alu), .ALUW_i(ALUW_i), 
        .DOUT(DOUT), .stall_o(stall_o), .Clock(Clock), .Reset(Reset) );
  mux41_MUX_SIZE5 MUXDEST ( .IN0({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .IN1(rC_i), 
        .IN2(rB_i), .IN3({1'b1, 1'b1, 1'b1, 1'b1, 1'b1}), .CTRL(S_MUX_DEST_i), 
        .OUT1(muxed_dest) );
  mux41_MUX_SIZE32_2 MUX_FWA ( .IN0(A_i), .IN1(FW_X_i), .IN2(FW_W_i), .IN3({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CTRL(S_FW_A_i), 
        .OUT1(FWA2alu) );
  mux41_MUX_SIZE32_1 MUX_FWB ( .IN0(MUXED_B_i), .IN1(FW_X_i), .IN2(FW_W_i), 
        .IN3({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CTRL(S_FW_B_i), .OUT1(muxed_B) );
endmodule


module execute_regs ( X_i, S_i, D2_i, X_o, S_o, D2_o, stall_i, clk, rst );
  input [31:0] X_i;
  input [31:0] S_i;
  input [4:0] D2_i;
  output [31:0] X_o;
  output [31:0] S_o;
  output [4:0] D2_o;
  input stall_i, clk, rst;


  ff32_en_SIZE32_3 X ( .D(X_i), .en(1'b1), .clk(clk), .rst(rst), .Q(X_o) );
  ff32_en_SIZE32_2 S ( .D(S_i), .en(1'b1), .clk(clk), .rst(rst), .Q(S_o) );
  ff32_en_SIZE5_1 D2 ( .D(D2_i), .en(1'b1), .clk(clk), .rst(rst), .Q(D2_o) );
endmodule


module decode_regs ( A_i, B_i, rA_i, rB_i, rC_i, IMM_i, ALUW_i, A_o, B_o, rA_o, 
        rB_o, rC_o, IMM_o, ALUW_o, stall_i, clk, rst );
  input [31:0] A_i;
  input [31:0] B_i;
  input [4:0] rA_i;
  input [4:0] rB_i;
  input [4:0] rC_i;
  input [31:0] IMM_i;
  input [12:0] ALUW_i;
  output [31:0] A_o;
  output [31:0] B_o;
  output [4:0] rA_o;
  output [4:0] rB_o;
  output [4:0] rC_o;
  output [31:0] IMM_o;
  output [12:0] ALUW_o;
  input stall_i, clk, rst;
  wire   enable;

  ff32_en_SIZE32_0 A ( .D(A_i), .en(enable), .clk(clk), .rst(rst), .Q(A_o) );
  ff32_en_SIZE32_5 B ( .D(B_i), .en(enable), .clk(clk), .rst(rst), .Q(B_o) );
  ff32_en_SIZE5_0 rA ( .D(rA_i), .en(enable), .clk(clk), .rst(rst), .Q(rA_o)
         );
  ff32_en_SIZE5_3 rB ( .D(rB_i), .en(enable), .clk(clk), .rst(rst), .Q(rB_o)
         );
  ff32_en_SIZE5_2 rC ( .D(rC_i), .en(enable), .clk(clk), .rst(rst), .Q(rC_o)
         );
  ff32_en_SIZE32_4 IMM ( .D(IMM_i), .en(enable), .clk(clk), .rst(rst), .Q(
        IMM_o) );
  ff32_en_SIZE13 ALUW ( .D(ALUW_i), .en(enable), .clk(clk), .rst(rst), .Q(
        ALUW_o) );
  INV_X1 U1 ( .A(stall_i), .ZN(enable) );
endmodule


module dlx_regfile ( Clk, Rst, ENABLE, RD1, RD2, WR, ADD_WR, ADD_RD1, ADD_RD2, 
        DATAIN, OUT1, OUT2 );
  input [4:0] ADD_WR;
  input [4:0] ADD_RD1;
  input [4:0] ADD_RD2;
  input [31:0] DATAIN;
  output [31:0] OUT1;
  output [31:0] OUT2;
  input Clk, Rst, ENABLE, RD1, RD2, WR;
  wire   N2503, N2567, N2631, N2695, N2759, N2823, N2887, N2951, N3015, N3079,
         N3143, N3207, N3271, N3335, N3399, N3463, N3527, N3591, N3655, N3719,
         N3783, N3847, N3911, N3975, N4039, N4103, N4167, N4231, N4295, N4359,
         N4423, N4487, N4490, N4492, N4494, N4496, N4498, N4500, N4502, N4504,
         N4506, N4508, N4510, N4512, N4514, N4516, N4518, N4520, N4522, N4524,
         N4526, N4528, N4530, N4532, N4534, N4536, N4538, N4540, N4542, N4544,
         N4546, N4548, N4550, N4552, N4554, N4556, N4558, N4560, N4562, N4564,
         N4566, N4568, N4570, N4572, N4574, N4576, N4578, N4580, N4582, N4584,
         N4586, N4588, N4590, N4592, N4594, N4596, N4598, N4600, N4602, N4604,
         N4606, N4608, N4610, N4612, N4614, N4615, N4616, net338042, net338047,
         net338052, net338057, net338062, net338067, net338072, net338077,
         net338082, net338087, net338092, net338097, net338102, net338107,
         net338112, net338117, net338122, net338127, net338132, net338137,
         net338142, net338147, net338152, net338157, net338162, net338167,
         net338172, net338177, net338182, net338187, net338192, net338197,
         net338202, net338207, n1094, n1150, n1172, n1194, n1216, n1238, n1260,
         n1282, n1304, n1326, n1348, n1370, n1392, n1414, n1436, n1458, n1480,
         n1502, n1524, n1546, n1568, n1590, n1612, n1634, n1656, n1678, n1700,
         n1722, n1744, n1766, n1788, n1810, n1, n2, n3, n37, n39, n41, n43,
         n45, n47, n49, n51, n53, n55, n57, n59, n61, n63, n65, n67, n69, n71,
         n73, n75, n77, n79, n81, n83, n85, n87, n89, n91, n93, n95, n97, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
         n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
         n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
         n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
         n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
         n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
         n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
         n1092, n1093, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1195,
         n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
         n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
         n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
         n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
         n1237, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
         n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
         n1258, n1259, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
         n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
         n1279, n1280, n1281, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
         n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
         n1300, n1301, n1302, n1303, n1305, n1306, n1307, n1308, n1309, n1310,
         n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
         n1321, n1322, n1323, n1324, n1325, n1327, n1328, n1329, n1330, n1331,
         n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
         n1342, n1343, n1344, n1345, n1346, n1347, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1371, n1372, n1373,
         n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
         n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1393, n1394,
         n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
         n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1415,
         n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425,
         n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435,
         n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446,
         n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456,
         n1457, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467,
         n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477,
         n1478, n1479, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488,
         n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498,
         n1499, n1500, n1501, n1503, n1504, n1505, n1506, n1507, n1508, n1509,
         n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519,
         n1520, n1521, n1522, n1523, n1525, n1526, n1527, n1528, n1529, n1530,
         n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540,
         n1541, n1542, n1543, n1544, n1545, n1547, n1548, n1549, n1550, n1551,
         n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561,
         n1562, n1563, n1564, n1565, n1566, n1567, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1591, n1592, n1593,
         n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603,
         n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1613, n1614,
         n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
         n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1635,
         n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645,
         n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655,
         n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666,
         n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676,
         n1677, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687,
         n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697,
         n1698, n1699, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708,
         n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718,
         n1719, n1720, n1721, n1723, n1724, n1725, n1726, n1727, n1728, n1729,
         n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739,
         n1740, n1741, n1742, n1743, n1745, n1746, n1747, n1748, n1749, n1750,
         n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760,
         n1761, n1762, n1763, n1764, n1765, n1767, n1768, n1769, n1770, n1771,
         n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781,
         n1782, n1783, n1784, n1785, n1786, n1787, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1811, n1812, n1813,
         n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823,
         n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833,
         n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843,
         n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853,
         n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863,
         n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873,
         n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883,
         n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893,
         n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903,
         n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913,
         n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923,
         n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933,
         n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943,
         n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953,
         n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963,
         n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973,
         n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983,
         n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993,
         n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003,
         n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013,
         n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023,
         n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033,
         n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043,
         n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053,
         n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063,
         n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073,
         n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083,
         n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093,
         n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103,
         n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113,
         n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123,
         n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133,
         n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143,
         n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153,
         n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163,
         n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173,
         n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183,
         n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193,
         n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203,
         n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213,
         n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223,
         n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233,
         n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243,
         n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253,
         n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263,
         n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273,
         n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283,
         n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293,
         n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303,
         n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313,
         n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323,
         n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333,
         n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343,
         n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353,
         n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363,
         n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373,
         n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383,
         n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393,
         n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403,
         n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413,
         n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423,
         n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433,
         n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443,
         n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453,
         n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463,
         n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473,
         n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483,
         n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493,
         n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503,
         n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513,
         n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523,
         n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533,
         n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543,
         n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553,
         n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563,
         n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573,
         n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583,
         n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593,
         n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603,
         n2604, n2605, n2606, n2607, n2608, n2609;
  assign N4487 = Rst;

  DFF_X1 \REGISTERS_reg[0][31]  ( .D(n1094), .CK(net338047), .Q(n177) );
  DFF_X1 \REGISTERS_reg[0][30]  ( .D(n1150), .CK(net338047), .Q(n176) );
  DFF_X1 \REGISTERS_reg[0][29]  ( .D(n1172), .CK(net338047), .Q(n174) );
  DFF_X1 \REGISTERS_reg[0][28]  ( .D(n1194), .CK(net338047), .Q(n173) );
  DFF_X1 \REGISTERS_reg[0][27]  ( .D(n1216), .CK(net338047), .Q(n172) );
  DFF_X1 \REGISTERS_reg[0][26]  ( .D(n1238), .CK(net338047), .Q(n171) );
  DFF_X1 \REGISTERS_reg[0][25]  ( .D(n1260), .CK(net338047), .Q(n170) );
  DFF_X1 \REGISTERS_reg[0][24]  ( .D(n1282), .CK(net338047), .Q(n169) );
  DFF_X1 \REGISTERS_reg[0][23]  ( .D(n1304), .CK(net338047), .Q(n168) );
  DFF_X1 \REGISTERS_reg[0][22]  ( .D(n1326), .CK(net338047), .Q(n167) );
  DFF_X1 \REGISTERS_reg[0][21]  ( .D(n1348), .CK(net338047), .Q(n166) );
  DFF_X1 \REGISTERS_reg[0][20]  ( .D(n1370), .CK(net338047), .Q(n165) );
  DFF_X1 \REGISTERS_reg[0][19]  ( .D(n1392), .CK(net338047), .Q(n163) );
  DFF_X1 \REGISTERS_reg[0][18]  ( .D(n1414), .CK(net338047), .Q(n162) );
  DFF_X1 \REGISTERS_reg[0][17]  ( .D(n1436), .CK(net338047), .Q(n161) );
  DFF_X1 \REGISTERS_reg[0][16]  ( .D(n1458), .CK(net338047), .Q(n160) );
  DFF_X1 \REGISTERS_reg[0][15]  ( .D(n1480), .CK(net338047), .Q(n159) );
  DFF_X1 \REGISTERS_reg[0][14]  ( .D(n1502), .CK(net338047), .Q(n158) );
  DFF_X1 \REGISTERS_reg[0][13]  ( .D(n1524), .CK(net338047), .Q(n157) );
  DFF_X1 \REGISTERS_reg[0][12]  ( .D(n1546), .CK(net338047), .Q(n156) );
  DFF_X1 \REGISTERS_reg[0][11]  ( .D(n1568), .CK(net338047), .Q(n155) );
  DFF_X1 \REGISTERS_reg[0][10]  ( .D(n1590), .CK(net338047), .Q(n154) );
  DFF_X1 \REGISTERS_reg[0][9]  ( .D(n1612), .CK(net338047), .Q(n152) );
  DFF_X1 \REGISTERS_reg[0][8]  ( .D(n1634), .CK(net338047), .Q(n151) );
  DFF_X1 \REGISTERS_reg[0][7]  ( .D(n1656), .CK(net338047), .Q(n150) );
  DFF_X1 \REGISTERS_reg[0][6]  ( .D(n1678), .CK(net338047), .Q(n149) );
  DFF_X1 \REGISTERS_reg[0][5]  ( .D(n1700), .CK(net338047), .Q(n148) );
  DFF_X1 \REGISTERS_reg[0][4]  ( .D(n1722), .CK(net338047), .Q(n147) );
  DFF_X1 \REGISTERS_reg[0][3]  ( .D(n1744), .CK(net338047), .Q(n146) );
  DFF_X1 \REGISTERS_reg[0][2]  ( .D(n1766), .CK(net338047), .Q(n145) );
  DFF_X1 \REGISTERS_reg[0][1]  ( .D(n1788), .CK(net338047), .Q(n144) );
  DFF_X1 \REGISTERS_reg[0][0]  ( .D(n1810), .CK(net338047), .Q(n143) );
  DFF_X1 \REGISTERS_reg[1][31]  ( .D(n1094), .CK(net338052), .Q(n141) );
  DFF_X1 \REGISTERS_reg[1][30]  ( .D(n1150), .CK(net338052), .Q(n140) );
  DFF_X1 \REGISTERS_reg[1][29]  ( .D(n1172), .CK(net338052), .Q(n139) );
  DFF_X1 \REGISTERS_reg[1][28]  ( .D(n1194), .CK(net338052), .Q(n138) );
  DFF_X1 \REGISTERS_reg[1][27]  ( .D(n1216), .CK(net338052), .Q(n137) );
  DFF_X1 \REGISTERS_reg[1][26]  ( .D(n1238), .CK(net338052), .Q(n136) );
  DFF_X1 \REGISTERS_reg[1][25]  ( .D(n1260), .CK(net338052), .Q(n135) );
  DFF_X1 \REGISTERS_reg[1][24]  ( .D(n1282), .CK(net338052), .Q(n134) );
  DFF_X1 \REGISTERS_reg[1][23]  ( .D(n1304), .CK(net338052), .Q(n133) );
  DFF_X1 \REGISTERS_reg[1][22]  ( .D(n1326), .CK(net338052), .Q(n132) );
  DFF_X1 \REGISTERS_reg[1][21]  ( .D(n1348), .CK(net338052), .Q(n130) );
  DFF_X1 \REGISTERS_reg[1][20]  ( .D(n1370), .CK(net338052), .Q(n129) );
  DFF_X1 \REGISTERS_reg[1][19]  ( .D(n1392), .CK(net338052), .Q(n128) );
  DFF_X1 \REGISTERS_reg[1][18]  ( .D(n1414), .CK(net338052), .Q(n127) );
  DFF_X1 \REGISTERS_reg[1][17]  ( .D(n1436), .CK(net338052), .Q(n126) );
  DFF_X1 \REGISTERS_reg[1][16]  ( .D(n1458), .CK(net338052), .Q(n125) );
  DFF_X1 \REGISTERS_reg[1][15]  ( .D(n1480), .CK(net338052), .Q(n124) );
  DFF_X1 \REGISTERS_reg[1][14]  ( .D(n1502), .CK(net338052), .Q(n123) );
  DFF_X1 \REGISTERS_reg[1][13]  ( .D(n1524), .CK(net338052), .Q(n122) );
  DFF_X1 \REGISTERS_reg[1][12]  ( .D(n1546), .CK(net338052), .Q(n121) );
  DFF_X1 \REGISTERS_reg[1][11]  ( .D(n1568), .CK(net338052), .Q(n119) );
  DFF_X1 \REGISTERS_reg[1][10]  ( .D(n1590), .CK(net338052), .Q(n118) );
  DFF_X1 \REGISTERS_reg[1][9]  ( .D(n1612), .CK(net338052), .Q(n117) );
  DFF_X1 \REGISTERS_reg[1][8]  ( .D(n1634), .CK(net338052), .Q(n116) );
  DFF_X1 \REGISTERS_reg[1][7]  ( .D(n1656), .CK(net338052), .Q(n115) );
  DFF_X1 \REGISTERS_reg[1][6]  ( .D(n1678), .CK(net338052), .Q(n114) );
  DFF_X1 \REGISTERS_reg[1][5]  ( .D(n1700), .CK(net338052), .Q(n113) );
  DFF_X1 \REGISTERS_reg[1][4]  ( .D(n1722), .CK(net338052), .Q(n112) );
  DFF_X1 \REGISTERS_reg[1][3]  ( .D(n1744), .CK(net338052), .Q(n111) );
  DFF_X1 \REGISTERS_reg[1][2]  ( .D(n1766), .CK(net338052), .Q(n110) );
  DFF_X1 \REGISTERS_reg[1][1]  ( .D(n1788), .CK(net338052), .Q(n108) );
  DFF_X1 \REGISTERS_reg[1][0]  ( .D(n1810), .CK(net338052), .Q(n107) );
  DFF_X1 \REGISTERS_reg[2][31]  ( .D(n1094), .CK(net338057), .Q(n106) );
  DFF_X1 \REGISTERS_reg[2][30]  ( .D(n1150), .CK(net338057), .Q(n105) );
  DFF_X1 \REGISTERS_reg[2][29]  ( .D(n1172), .CK(net338057), .Q(n104) );
  DFF_X1 \REGISTERS_reg[2][28]  ( .D(n1194), .CK(net338057), .Q(n103) );
  DFF_X1 \REGISTERS_reg[2][27]  ( .D(n1216), .CK(net338057), .Q(n102) );
  DFF_X1 \REGISTERS_reg[2][26]  ( .D(n1238), .CK(net338057), .Q(n101) );
  DFF_X1 \REGISTERS_reg[2][25]  ( .D(n1260), .CK(net338057), .Q(n100) );
  DFF_X1 \REGISTERS_reg[2][24]  ( .D(n1282), .CK(net338057), .Q(n99) );
  DFF_X1 \REGISTERS_reg[2][23]  ( .D(n1304), .CK(net338057), .Q(n95) );
  DFF_X1 \REGISTERS_reg[2][22]  ( .D(n1326), .CK(net338057), .Q(n93) );
  DFF_X1 \REGISTERS_reg[2][21]  ( .D(n1348), .CK(net338057), .Q(n91) );
  DFF_X1 \REGISTERS_reg[2][20]  ( .D(n1370), .CK(net338057), .Q(n89) );
  DFF_X1 \REGISTERS_reg[2][19]  ( .D(n1392), .CK(net338057), .Q(n87) );
  DFF_X1 \REGISTERS_reg[2][18]  ( .D(n1414), .CK(net338057), .Q(n85) );
  DFF_X1 \REGISTERS_reg[2][17]  ( .D(n1436), .CK(net338057), .Q(n83) );
  DFF_X1 \REGISTERS_reg[2][16]  ( .D(n1458), .CK(net338057), .Q(n81) );
  DFF_X1 \REGISTERS_reg[2][15]  ( .D(n1480), .CK(net338057), .Q(n79) );
  DFF_X1 \REGISTERS_reg[2][14]  ( .D(n1502), .CK(net338057), .Q(n77) );
  DFF_X1 \REGISTERS_reg[2][13]  ( .D(n1524), .CK(net338057), .Q(n73) );
  DFF_X1 \REGISTERS_reg[2][12]  ( .D(n1546), .CK(net338057), .Q(n71) );
  DFF_X1 \REGISTERS_reg[2][11]  ( .D(n1568), .CK(net338057), .Q(n69) );
  DFF_X1 \REGISTERS_reg[2][10]  ( .D(n1590), .CK(net338057), .Q(n67) );
  DFF_X1 \REGISTERS_reg[2][9]  ( .D(n1612), .CK(net338057), .Q(n65) );
  DFF_X1 \REGISTERS_reg[2][8]  ( .D(n1634), .CK(net338057), .Q(n63) );
  DFF_X1 \REGISTERS_reg[2][7]  ( .D(n1656), .CK(net338057), .Q(n61) );
  DFF_X1 \REGISTERS_reg[2][6]  ( .D(n1678), .CK(net338057), .Q(n59) );
  DFF_X1 \REGISTERS_reg[2][5]  ( .D(n1700), .CK(net338057), .Q(n57) );
  DFF_X1 \REGISTERS_reg[2][4]  ( .D(n1722), .CK(net338057), .Q(n55) );
  DFF_X1 \REGISTERS_reg[2][3]  ( .D(n1744), .CK(net338057), .Q(n1100) );
  DFF_X1 \REGISTERS_reg[2][2]  ( .D(n1766), .CK(net338057), .Q(n1099) );
  DFF_X1 \REGISTERS_reg[2][1]  ( .D(n1788), .CK(net338057), .Q(n1098) );
  DFF_X1 \REGISTERS_reg[2][0]  ( .D(n1810), .CK(net338057), .Q(n1097) );
  DFF_X1 \REGISTERS_reg[3][31]  ( .D(n1094), .CK(net338062), .Q(n1096) );
  DFF_X1 \REGISTERS_reg[3][30]  ( .D(n1150), .CK(net338062), .Q(n1095) );
  DFF_X1 \REGISTERS_reg[3][29]  ( .D(n1172), .CK(net338062), .Q(n1093) );
  DFF_X1 \REGISTERS_reg[3][28]  ( .D(n1194), .CK(net338062), .Q(n1092) );
  DFF_X1 \REGISTERS_reg[3][27]  ( .D(n1216), .CK(net338062), .Q(n1091) );
  DFF_X1 \REGISTERS_reg[3][26]  ( .D(n1238), .CK(net338062), .Q(n1090) );
  DFF_X1 \REGISTERS_reg[3][25]  ( .D(n1260), .CK(net338062), .Q(n1088) );
  DFF_X1 \REGISTERS_reg[3][24]  ( .D(n1282), .CK(net338062), .Q(n1087) );
  DFF_X1 \REGISTERS_reg[3][23]  ( .D(n1304), .CK(net338062), .Q(n1086) );
  DFF_X1 \REGISTERS_reg[3][22]  ( .D(n1326), .CK(net338062), .Q(n1085) );
  DFF_X1 \REGISTERS_reg[3][21]  ( .D(n1348), .CK(net338062), .Q(n1084) );
  DFF_X1 \REGISTERS_reg[3][20]  ( .D(n1370), .CK(net338062), .Q(n1083) );
  DFF_X1 \REGISTERS_reg[3][19]  ( .D(n1392), .CK(net338062), .Q(n1082) );
  DFF_X1 \REGISTERS_reg[3][18]  ( .D(n1414), .CK(net338062), .Q(n1081) );
  DFF_X1 \REGISTERS_reg[3][17]  ( .D(n1436), .CK(net338062), .Q(n1080) );
  DFF_X1 \REGISTERS_reg[3][16]  ( .D(n1458), .CK(net338062), .Q(n1079) );
  DFF_X1 \REGISTERS_reg[3][15]  ( .D(n1480), .CK(net338062), .Q(n1078) );
  DFF_X1 \REGISTERS_reg[3][14]  ( .D(n1502), .CK(net338062), .Q(n1077) );
  DFF_X1 \REGISTERS_reg[3][13]  ( .D(n1524), .CK(net338062), .Q(n1076) );
  DFF_X1 \REGISTERS_reg[3][12]  ( .D(n1546), .CK(net338062), .Q(n1075) );
  DFF_X1 \REGISTERS_reg[3][11]  ( .D(n1568), .CK(net338062), .Q(n1074) );
  DFF_X1 \REGISTERS_reg[3][10]  ( .D(n1590), .CK(net338062), .Q(n1073) );
  DFF_X1 \REGISTERS_reg[3][9]  ( .D(n1612), .CK(net338062), .Q(n1072) );
  DFF_X1 \REGISTERS_reg[3][8]  ( .D(n1634), .CK(net338062), .Q(n1071) );
  DFF_X1 \REGISTERS_reg[3][7]  ( .D(n1656), .CK(net338062), .Q(n1070) );
  DFF_X1 \REGISTERS_reg[3][6]  ( .D(n1678), .CK(net338062), .Q(n1069) );
  DFF_X1 \REGISTERS_reg[3][5]  ( .D(n1700), .CK(net338062), .Q(n1067) );
  DFF_X1 \REGISTERS_reg[3][4]  ( .D(n1722), .CK(net338062), .Q(n1066) );
  DFF_X1 \REGISTERS_reg[3][3]  ( .D(n1744), .CK(net338062), .Q(n1065) );
  DFF_X1 \REGISTERS_reg[3][2]  ( .D(n1766), .CK(net338062), .Q(n1064) );
  DFF_X1 \REGISTERS_reg[3][1]  ( .D(n1788), .CK(net338062), .Q(n1063) );
  DFF_X1 \REGISTERS_reg[3][0]  ( .D(n1810), .CK(net338062), .Q(n1062) );
  DFF_X1 \REGISTERS_reg[4][31]  ( .D(n1094), .CK(net338067), .Q(n1061) );
  DFF_X1 \REGISTERS_reg[4][30]  ( .D(n1150), .CK(net338067), .Q(n1060) );
  DFF_X1 \REGISTERS_reg[4][29]  ( .D(n1172), .CK(net338067), .Q(n1059) );
  DFF_X1 \REGISTERS_reg[4][28]  ( .D(n1194), .CK(net338067), .Q(n1058) );
  DFF_X1 \REGISTERS_reg[4][27]  ( .D(n1216), .CK(net338067), .Q(n1057) );
  DFF_X1 \REGISTERS_reg[4][26]  ( .D(n1238), .CK(net338067), .Q(n1056) );
  DFF_X1 \REGISTERS_reg[4][25]  ( .D(n1260), .CK(net338067), .Q(n1055) );
  DFF_X1 \REGISTERS_reg[4][24]  ( .D(n1282), .CK(net338067), .Q(n1054) );
  DFF_X1 \REGISTERS_reg[4][23]  ( .D(n1304), .CK(net338067), .Q(n1053) );
  DFF_X1 \REGISTERS_reg[4][22]  ( .D(n1326), .CK(net338067), .Q(n1052) );
  DFF_X1 \REGISTERS_reg[4][21]  ( .D(n1348), .CK(net338067), .Q(n1051) );
  DFF_X1 \REGISTERS_reg[4][20]  ( .D(n1370), .CK(net338067), .Q(n1050) );
  DFF_X1 \REGISTERS_reg[4][19]  ( .D(n1392), .CK(net338067), .Q(n1049) );
  DFF_X1 \REGISTERS_reg[4][18]  ( .D(n1414), .CK(net338067), .Q(n1048) );
  DFF_X1 \REGISTERS_reg[4][17]  ( .D(n1436), .CK(net338067), .Q(n1046) );
  DFF_X1 \REGISTERS_reg[4][16]  ( .D(n1458), .CK(net338067), .Q(n1045) );
  DFF_X1 \REGISTERS_reg[4][15]  ( .D(n1480), .CK(net338067), .Q(n1044) );
  DFF_X1 \REGISTERS_reg[4][14]  ( .D(n1502), .CK(net338067), .Q(n1043) );
  DFF_X1 \REGISTERS_reg[4][13]  ( .D(n1524), .CK(net338067), .Q(n1042) );
  DFF_X1 \REGISTERS_reg[4][12]  ( .D(n1546), .CK(net338067), .Q(n1041) );
  DFF_X1 \REGISTERS_reg[4][11]  ( .D(n1568), .CK(net338067), .Q(n1040) );
  DFF_X1 \REGISTERS_reg[4][10]  ( .D(n1590), .CK(net338067), .Q(n1039) );
  DFF_X1 \REGISTERS_reg[4][9]  ( .D(n1612), .CK(net338067), .Q(n1038) );
  DFF_X1 \REGISTERS_reg[4][8]  ( .D(n1634), .CK(net338067), .Q(n1037) );
  DFF_X1 \REGISTERS_reg[4][7]  ( .D(n1656), .CK(net338067), .Q(n1036) );
  DFF_X1 \REGISTERS_reg[4][6]  ( .D(n1678), .CK(net338067), .Q(n1035) );
  DFF_X1 \REGISTERS_reg[4][5]  ( .D(n1700), .CK(net338067), .Q(n1034) );
  DFF_X1 \REGISTERS_reg[4][4]  ( .D(n1722), .CK(net338067), .Q(n1033) );
  DFF_X1 \REGISTERS_reg[4][3]  ( .D(n1744), .CK(net338067), .Q(n1032) );
  DFF_X1 \REGISTERS_reg[4][2]  ( .D(n1766), .CK(net338067), .Q(n1031) );
  DFF_X1 \REGISTERS_reg[4][1]  ( .D(n1788), .CK(net338067), .Q(n1030) );
  DFF_X1 \REGISTERS_reg[4][0]  ( .D(n1810), .CK(net338067), .Q(n1029) );
  DFF_X1 \REGISTERS_reg[5][31]  ( .D(n1094), .CK(net338072), .Q(n1028) );
  DFF_X1 \REGISTERS_reg[5][30]  ( .D(n1150), .CK(net338072), .Q(n1027) );
  DFF_X1 \REGISTERS_reg[5][29]  ( .D(n1172), .CK(net338072), .Q(n1025) );
  DFF_X1 \REGISTERS_reg[5][28]  ( .D(n1194), .CK(net338072), .Q(n1024) );
  DFF_X1 \REGISTERS_reg[5][27]  ( .D(n1216), .CK(net338072), .Q(n1023) );
  DFF_X1 \REGISTERS_reg[5][26]  ( .D(n1238), .CK(net338072), .Q(n1022) );
  DFF_X1 \REGISTERS_reg[5][25]  ( .D(n1260), .CK(net338072), .Q(n1021) );
  DFF_X1 \REGISTERS_reg[5][24]  ( .D(n1282), .CK(net338072), .Q(n1020) );
  DFF_X1 \REGISTERS_reg[5][23]  ( .D(n1304), .CK(net338072), .Q(n1019) );
  DFF_X1 \REGISTERS_reg[5][22]  ( .D(n1326), .CK(net338072), .Q(n1018) );
  DFF_X1 \REGISTERS_reg[5][21]  ( .D(n1348), .CK(net338072), .Q(n1017) );
  DFF_X1 \REGISTERS_reg[5][20]  ( .D(n1370), .CK(net338072), .Q(n1016) );
  DFF_X1 \REGISTERS_reg[5][19]  ( .D(n1392), .CK(net338072), .Q(n1015) );
  DFF_X1 \REGISTERS_reg[5][18]  ( .D(n1414), .CK(net338072), .Q(n1014) );
  DFF_X1 \REGISTERS_reg[5][17]  ( .D(n1436), .CK(net338072), .Q(n1013) );
  DFF_X1 \REGISTERS_reg[5][16]  ( .D(n1458), .CK(net338072), .Q(n1012) );
  DFF_X1 \REGISTERS_reg[5][15]  ( .D(n1480), .CK(net338072), .Q(n1011) );
  DFF_X1 \REGISTERS_reg[5][14]  ( .D(n1502), .CK(net338072), .Q(n1010) );
  DFF_X1 \REGISTERS_reg[5][13]  ( .D(n1524), .CK(net338072), .Q(n1009) );
  DFF_X1 \REGISTERS_reg[5][12]  ( .D(n1546), .CK(net338072), .Q(n1008) );
  DFF_X1 \REGISTERS_reg[5][11]  ( .D(n1568), .CK(net338072), .Q(n1007) );
  DFF_X1 \REGISTERS_reg[5][10]  ( .D(n1590), .CK(net338072), .Q(n1006) );
  DFF_X1 \REGISTERS_reg[5][9]  ( .D(n1612), .CK(net338072), .Q(n1004) );
  DFF_X1 \REGISTERS_reg[5][8]  ( .D(n1634), .CK(net338072), .Q(n1003) );
  DFF_X1 \REGISTERS_reg[5][7]  ( .D(n1656), .CK(net338072), .Q(n1002) );
  DFF_X1 \REGISTERS_reg[5][6]  ( .D(n1678), .CK(net338072), .Q(n1001) );
  DFF_X1 \REGISTERS_reg[5][5]  ( .D(n1700), .CK(net338072), .Q(n1000) );
  DFF_X1 \REGISTERS_reg[5][4]  ( .D(n1722), .CK(net338072), .Q(n999) );
  DFF_X1 \REGISTERS_reg[5][3]  ( .D(n1744), .CK(net338072), .Q(n998) );
  DFF_X1 \REGISTERS_reg[5][2]  ( .D(n1766), .CK(net338072), .Q(n997) );
  DFF_X1 \REGISTERS_reg[5][1]  ( .D(n1788), .CK(net338072), .Q(n996) );
  DFF_X1 \REGISTERS_reg[5][0]  ( .D(n1810), .CK(net338072), .Q(n995) );
  DFF_X1 \REGISTERS_reg[6][31]  ( .D(n1094), .CK(net338077), .Q(n994) );
  DFF_X1 \REGISTERS_reg[6][30]  ( .D(n1150), .CK(net338077), .Q(n993) );
  DFF_X1 \REGISTERS_reg[6][29]  ( .D(n1172), .CK(net338077), .Q(n992) );
  DFF_X1 \REGISTERS_reg[6][28]  ( .D(n1194), .CK(net338077), .Q(n991) );
  DFF_X1 \REGISTERS_reg[6][27]  ( .D(n1216), .CK(net338077), .Q(n990) );
  DFF_X1 \REGISTERS_reg[6][26]  ( .D(n1238), .CK(net338077), .Q(n989) );
  DFF_X1 \REGISTERS_reg[6][25]  ( .D(n1260), .CK(net338077), .Q(n988) );
  DFF_X1 \REGISTERS_reg[6][24]  ( .D(n1282), .CK(net338077), .Q(n987) );
  DFF_X1 \REGISTERS_reg[6][23]  ( .D(n1304), .CK(net338077), .Q(n986) );
  DFF_X1 \REGISTERS_reg[6][22]  ( .D(n1326), .CK(net338077), .Q(n985) );
  DFF_X1 \REGISTERS_reg[6][21]  ( .D(n1348), .CK(net338077), .Q(n983) );
  DFF_X1 \REGISTERS_reg[6][20]  ( .D(n1370), .CK(net338077), .Q(n982) );
  DFF_X1 \REGISTERS_reg[6][19]  ( .D(n1392), .CK(net338077), .Q(n981) );
  DFF_X1 \REGISTERS_reg[6][18]  ( .D(n1414), .CK(net338077), .Q(n980) );
  DFF_X1 \REGISTERS_reg[6][17]  ( .D(n1436), .CK(net338077), .Q(n979) );
  DFF_X1 \REGISTERS_reg[6][16]  ( .D(n1458), .CK(net338077), .Q(n978) );
  DFF_X1 \REGISTERS_reg[6][15]  ( .D(n1480), .CK(net338077), .Q(n977) );
  DFF_X1 \REGISTERS_reg[6][14]  ( .D(n1502), .CK(net338077), .Q(n976) );
  DFF_X1 \REGISTERS_reg[6][13]  ( .D(n1524), .CK(net338077), .Q(n975) );
  DFF_X1 \REGISTERS_reg[6][12]  ( .D(n1546), .CK(net338077), .Q(n974) );
  DFF_X1 \REGISTERS_reg[6][11]  ( .D(n1568), .CK(net338077), .Q(n973) );
  DFF_X1 \REGISTERS_reg[6][10]  ( .D(n1590), .CK(net338077), .Q(n972) );
  DFF_X1 \REGISTERS_reg[6][9]  ( .D(n1612), .CK(net338077), .Q(n971) );
  DFF_X1 \REGISTERS_reg[6][8]  ( .D(n1634), .CK(net338077), .Q(n970) );
  DFF_X1 \REGISTERS_reg[6][7]  ( .D(n1656), .CK(net338077), .Q(n969) );
  DFF_X1 \REGISTERS_reg[6][6]  ( .D(n1678), .CK(net338077), .Q(n968) );
  DFF_X1 \REGISTERS_reg[6][5]  ( .D(n1700), .CK(net338077), .Q(n967) );
  DFF_X1 \REGISTERS_reg[6][4]  ( .D(n1722), .CK(net338077), .Q(n966) );
  DFF_X1 \REGISTERS_reg[6][3]  ( .D(n1744), .CK(net338077), .Q(n965) );
  DFF_X1 \REGISTERS_reg[6][2]  ( .D(n1766), .CK(net338077), .Q(n964) );
  DFF_X1 \REGISTERS_reg[6][1]  ( .D(n1788), .CK(net338077), .Q(n962) );
  DFF_X1 \REGISTERS_reg[6][0]  ( .D(n1810), .CK(net338077), .Q(n961) );
  DFF_X1 \REGISTERS_reg[7][31]  ( .D(n1094), .CK(net338082), .Q(n960) );
  DFF_X1 \REGISTERS_reg[7][30]  ( .D(n1150), .CK(net338082), .Q(n959) );
  DFF_X1 \REGISTERS_reg[7][29]  ( .D(n1172), .CK(net338082), .Q(n958) );
  DFF_X1 \REGISTERS_reg[7][28]  ( .D(n1194), .CK(net338082), .Q(n957) );
  DFF_X1 \REGISTERS_reg[7][27]  ( .D(n1216), .CK(net338082), .Q(n956) );
  DFF_X1 \REGISTERS_reg[7][26]  ( .D(n1238), .CK(net338082), .Q(n955) );
  DFF_X1 \REGISTERS_reg[7][25]  ( .D(n1260), .CK(net338082), .Q(n954) );
  DFF_X1 \REGISTERS_reg[7][24]  ( .D(n1282), .CK(net338082), .Q(n953) );
  DFF_X1 \REGISTERS_reg[7][23]  ( .D(n1304), .CK(net338082), .Q(n952) );
  DFF_X1 \REGISTERS_reg[7][22]  ( .D(n1326), .CK(net338082), .Q(n951) );
  DFF_X1 \REGISTERS_reg[7][21]  ( .D(n1348), .CK(net338082), .Q(n950) );
  DFF_X1 \REGISTERS_reg[7][20]  ( .D(n1370), .CK(net338082), .Q(n949) );
  DFF_X1 \REGISTERS_reg[7][19]  ( .D(n1392), .CK(net338082), .Q(n948) );
  DFF_X1 \REGISTERS_reg[7][18]  ( .D(n1414), .CK(net338082), .Q(n947) );
  DFF_X1 \REGISTERS_reg[7][17]  ( .D(n1436), .CK(net338082), .Q(n946) );
  DFF_X1 \REGISTERS_reg[7][16]  ( .D(n1458), .CK(net338082), .Q(n945) );
  DFF_X1 \REGISTERS_reg[7][15]  ( .D(n1480), .CK(net338082), .Q(n944) );
  DFF_X1 \REGISTERS_reg[7][14]  ( .D(n1502), .CK(net338082), .Q(n943) );
  DFF_X1 \REGISTERS_reg[7][13]  ( .D(n1524), .CK(net338082), .Q(n941) );
  DFF_X1 \REGISTERS_reg[7][12]  ( .D(n1546), .CK(net338082), .Q(n940) );
  DFF_X1 \REGISTERS_reg[7][11]  ( .D(n1568), .CK(net338082), .Q(n939) );
  DFF_X1 \REGISTERS_reg[7][10]  ( .D(n1590), .CK(net338082), .Q(n938) );
  DFF_X1 \REGISTERS_reg[7][9]  ( .D(n1612), .CK(net338082), .Q(n937) );
  DFF_X1 \REGISTERS_reg[7][8]  ( .D(n1634), .CK(net338082), .Q(n936) );
  DFF_X1 \REGISTERS_reg[7][7]  ( .D(n1656), .CK(net338082), .Q(n935) );
  DFF_X1 \REGISTERS_reg[7][6]  ( .D(n1678), .CK(net338082), .Q(n934) );
  DFF_X1 \REGISTERS_reg[7][5]  ( .D(n1700), .CK(net338082), .Q(n933) );
  DFF_X1 \REGISTERS_reg[7][4]  ( .D(n1722), .CK(net338082), .Q(n932) );
  DFF_X1 \REGISTERS_reg[7][3]  ( .D(n1744), .CK(net338082), .Q(n931) );
  DFF_X1 \REGISTERS_reg[7][2]  ( .D(n1766), .CK(net338082), .Q(n930) );
  DFF_X1 \REGISTERS_reg[7][1]  ( .D(n1788), .CK(net338082), .Q(n929) );
  DFF_X1 \REGISTERS_reg[7][0]  ( .D(n1810), .CK(net338082), .Q(n928) );
  DFF_X1 \REGISTERS_reg[8][31]  ( .D(n1094), .CK(net338087), .Q(n927) );
  DFF_X1 \REGISTERS_reg[8][30]  ( .D(n1150), .CK(net338087), .Q(n926) );
  DFF_X1 \REGISTERS_reg[8][29]  ( .D(n1172), .CK(net338087), .Q(n925) );
  DFF_X1 \REGISTERS_reg[8][28]  ( .D(n1194), .CK(net338087), .Q(n924) );
  DFF_X1 \REGISTERS_reg[8][27]  ( .D(n1216), .CK(net338087), .Q(n923) );
  DFF_X1 \REGISTERS_reg[8][26]  ( .D(n1238), .CK(net338087), .Q(n922) );
  DFF_X1 \REGISTERS_reg[8][25]  ( .D(n1260), .CK(net338087), .Q(n920) );
  DFF_X1 \REGISTERS_reg[8][24]  ( .D(n1282), .CK(net338087), .Q(n919) );
  DFF_X1 \REGISTERS_reg[8][23]  ( .D(n1304), .CK(net338087), .Q(n918) );
  DFF_X1 \REGISTERS_reg[8][22]  ( .D(n1326), .CK(net338087), .Q(n917) );
  DFF_X1 \REGISTERS_reg[8][21]  ( .D(n1348), .CK(net338087), .Q(n916) );
  DFF_X1 \REGISTERS_reg[8][20]  ( .D(n1370), .CK(net338087), .Q(n915) );
  DFF_X1 \REGISTERS_reg[8][19]  ( .D(n1392), .CK(net338087), .Q(n914) );
  DFF_X1 \REGISTERS_reg[8][18]  ( .D(n1414), .CK(net338087), .Q(n913) );
  DFF_X1 \REGISTERS_reg[8][17]  ( .D(n1436), .CK(net338087), .Q(n912) );
  DFF_X1 \REGISTERS_reg[8][16]  ( .D(n1458), .CK(net338087), .Q(n911) );
  DFF_X1 \REGISTERS_reg[8][15]  ( .D(n1480), .CK(net338087), .Q(n910) );
  DFF_X1 \REGISTERS_reg[8][14]  ( .D(n1502), .CK(net338087), .Q(n909) );
  DFF_X1 \REGISTERS_reg[8][13]  ( .D(n1524), .CK(net338087), .Q(n908) );
  DFF_X1 \REGISTERS_reg[8][12]  ( .D(n1546), .CK(net338087), .Q(n907) );
  DFF_X1 \REGISTERS_reg[8][11]  ( .D(n1568), .CK(net338087), .Q(n906) );
  DFF_X1 \REGISTERS_reg[8][10]  ( .D(n1590), .CK(net338087), .Q(n905) );
  DFF_X1 \REGISTERS_reg[8][9]  ( .D(n1612), .CK(net338087), .Q(n904) );
  DFF_X1 \REGISTERS_reg[8][8]  ( .D(n1634), .CK(net338087), .Q(n903) );
  DFF_X1 \REGISTERS_reg[8][7]  ( .D(n1656), .CK(net338087), .Q(n902) );
  DFF_X1 \REGISTERS_reg[8][6]  ( .D(n1678), .CK(net338087), .Q(n901) );
  DFF_X1 \REGISTERS_reg[8][5]  ( .D(n1700), .CK(net338087), .Q(n899) );
  DFF_X1 \REGISTERS_reg[8][4]  ( .D(n1722), .CK(net338087), .Q(n898) );
  DFF_X1 \REGISTERS_reg[8][3]  ( .D(n1744), .CK(net338087), .Q(n897) );
  DFF_X1 \REGISTERS_reg[8][2]  ( .D(n1766), .CK(net338087), .Q(n896) );
  DFF_X1 \REGISTERS_reg[8][1]  ( .D(n1788), .CK(net338087), .Q(n895) );
  DFF_X1 \REGISTERS_reg[8][0]  ( .D(n1810), .CK(net338087), .Q(n894) );
  DFF_X1 \REGISTERS_reg[9][31]  ( .D(n1094), .CK(net338092), .Q(n893) );
  DFF_X1 \REGISTERS_reg[9][30]  ( .D(n1150), .CK(net338092), .Q(n892) );
  DFF_X1 \REGISTERS_reg[9][29]  ( .D(n1172), .CK(net338092), .Q(n891) );
  DFF_X1 \REGISTERS_reg[9][28]  ( .D(n1194), .CK(net338092), .Q(n890) );
  DFF_X1 \REGISTERS_reg[9][27]  ( .D(n1216), .CK(net338092), .Q(n889) );
  DFF_X1 \REGISTERS_reg[9][26]  ( .D(n1238), .CK(net338092), .Q(n888) );
  DFF_X1 \REGISTERS_reg[9][25]  ( .D(n1260), .CK(net338092), .Q(n887) );
  DFF_X1 \REGISTERS_reg[9][24]  ( .D(n1282), .CK(net338092), .Q(n886) );
  DFF_X1 \REGISTERS_reg[9][23]  ( .D(n1304), .CK(net338092), .Q(n885) );
  DFF_X1 \REGISTERS_reg[9][22]  ( .D(n1326), .CK(net338092), .Q(n884) );
  DFF_X1 \REGISTERS_reg[9][21]  ( .D(n1348), .CK(net338092), .Q(n883) );
  DFF_X1 \REGISTERS_reg[9][20]  ( .D(n1370), .CK(net338092), .Q(n882) );
  DFF_X1 \REGISTERS_reg[9][19]  ( .D(n1392), .CK(net338092), .Q(n881) );
  DFF_X1 \REGISTERS_reg[9][18]  ( .D(n1414), .CK(net338092), .Q(n880) );
  DFF_X1 \REGISTERS_reg[9][17]  ( .D(n1436), .CK(net338092), .Q(n878) );
  DFF_X1 \REGISTERS_reg[9][16]  ( .D(n1458), .CK(net338092), .Q(n877) );
  DFF_X1 \REGISTERS_reg[9][15]  ( .D(n1480), .CK(net338092), .Q(n876) );
  DFF_X1 \REGISTERS_reg[9][14]  ( .D(n1502), .CK(net338092), .Q(n875) );
  DFF_X1 \REGISTERS_reg[9][13]  ( .D(n1524), .CK(net338092), .Q(n874) );
  DFF_X1 \REGISTERS_reg[9][12]  ( .D(n1546), .CK(net338092), .Q(n873) );
  DFF_X1 \REGISTERS_reg[9][11]  ( .D(n1568), .CK(net338092), .Q(n872) );
  DFF_X1 \REGISTERS_reg[9][10]  ( .D(n1590), .CK(net338092), .Q(n871) );
  DFF_X1 \REGISTERS_reg[9][9]  ( .D(n1612), .CK(net338092), .Q(n870) );
  DFF_X1 \REGISTERS_reg[9][8]  ( .D(n1634), .CK(net338092), .Q(n869) );
  DFF_X1 \REGISTERS_reg[9][7]  ( .D(n1656), .CK(net338092), .Q(n868) );
  DFF_X1 \REGISTERS_reg[9][6]  ( .D(n1678), .CK(net338092), .Q(n867) );
  DFF_X1 \REGISTERS_reg[9][5]  ( .D(n1700), .CK(net338092), .Q(n866) );
  DFF_X1 \REGISTERS_reg[9][4]  ( .D(n1722), .CK(net338092), .Q(n865) );
  DFF_X1 \REGISTERS_reg[9][3]  ( .D(n1744), .CK(net338092), .Q(n864) );
  DFF_X1 \REGISTERS_reg[9][2]  ( .D(n1766), .CK(net338092), .Q(n863) );
  DFF_X1 \REGISTERS_reg[9][1]  ( .D(n1788), .CK(net338092), .Q(n862) );
  DFF_X1 \REGISTERS_reg[9][0]  ( .D(n1810), .CK(net338092), .Q(n861) );
  DFF_X1 \REGISTERS_reg[10][31]  ( .D(n1094), .CK(net338097), .Q(n860) );
  DFF_X1 \REGISTERS_reg[10][30]  ( .D(n1150), .CK(net338097), .Q(n859) );
  DFF_X1 \REGISTERS_reg[10][29]  ( .D(n1172), .CK(net338097), .Q(n857) );
  DFF_X1 \REGISTERS_reg[10][28]  ( .D(n1194), .CK(net338097), .Q(n856) );
  DFF_X1 \REGISTERS_reg[10][27]  ( .D(n1216), .CK(net338097), .Q(n855) );
  DFF_X1 \REGISTERS_reg[10][26]  ( .D(n1238), .CK(net338097), .Q(n854) );
  DFF_X1 \REGISTERS_reg[10][25]  ( .D(n1260), .CK(net338097), .Q(n853) );
  DFF_X1 \REGISTERS_reg[10][24]  ( .D(n1282), .CK(net338097), .Q(n852) );
  DFF_X1 \REGISTERS_reg[10][23]  ( .D(n1304), .CK(net338097), .Q(n851) );
  DFF_X1 \REGISTERS_reg[10][22]  ( .D(n1326), .CK(net338097), .Q(n850) );
  DFF_X1 \REGISTERS_reg[10][21]  ( .D(n1348), .CK(net338097), .Q(n849) );
  DFF_X1 \REGISTERS_reg[10][20]  ( .D(n1370), .CK(net338097), .Q(n848) );
  DFF_X1 \REGISTERS_reg[10][19]  ( .D(n1392), .CK(net338097), .Q(n847) );
  DFF_X1 \REGISTERS_reg[10][18]  ( .D(n1414), .CK(net338097), .Q(n846) );
  DFF_X1 \REGISTERS_reg[10][17]  ( .D(n1436), .CK(net338097), .Q(n845) );
  DFF_X1 \REGISTERS_reg[10][16]  ( .D(n1458), .CK(net338097), .Q(n844) );
  DFF_X1 \REGISTERS_reg[10][15]  ( .D(n1480), .CK(net338097), .Q(n843) );
  DFF_X1 \REGISTERS_reg[10][14]  ( .D(n1502), .CK(net338097), .Q(n842) );
  DFF_X1 \REGISTERS_reg[10][13]  ( .D(n1524), .CK(net338097), .Q(n841) );
  DFF_X1 \REGISTERS_reg[10][12]  ( .D(n1546), .CK(net338097), .Q(n840) );
  DFF_X1 \REGISTERS_reg[10][11]  ( .D(n1568), .CK(net338097), .Q(n839) );
  DFF_X1 \REGISTERS_reg[10][10]  ( .D(n1590), .CK(net338097), .Q(n838) );
  DFF_X1 \REGISTERS_reg[10][9]  ( .D(n1612), .CK(net338097), .Q(n836) );
  DFF_X1 \REGISTERS_reg[10][8]  ( .D(n1634), .CK(net338097), .Q(n835) );
  DFF_X1 \REGISTERS_reg[10][7]  ( .D(n1656), .CK(net338097), .Q(n834) );
  DFF_X1 \REGISTERS_reg[10][6]  ( .D(n1678), .CK(net338097), .Q(n833) );
  DFF_X1 \REGISTERS_reg[10][5]  ( .D(n1700), .CK(net338097), .Q(n832) );
  DFF_X1 \REGISTERS_reg[10][4]  ( .D(n1722), .CK(net338097), .Q(n831) );
  DFF_X1 \REGISTERS_reg[10][3]  ( .D(n1744), .CK(net338097), .Q(n830) );
  DFF_X1 \REGISTERS_reg[10][2]  ( .D(n1766), .CK(net338097), .Q(n829) );
  DFF_X1 \REGISTERS_reg[10][1]  ( .D(n1788), .CK(net338097), .Q(n828) );
  DFF_X1 \REGISTERS_reg[10][0]  ( .D(n1810), .CK(net338097), .Q(n827) );
  DFF_X1 \REGISTERS_reg[11][31]  ( .D(n1094), .CK(net338102), .Q(n826) );
  DFF_X1 \REGISTERS_reg[11][30]  ( .D(n1150), .CK(net338102), .Q(n825) );
  DFF_X1 \REGISTERS_reg[11][29]  ( .D(n1172), .CK(net338102), .Q(n824) );
  DFF_X1 \REGISTERS_reg[11][28]  ( .D(n1194), .CK(net338102), .Q(n823) );
  DFF_X1 \REGISTERS_reg[11][27]  ( .D(n1216), .CK(net338102), .Q(n822) );
  DFF_X1 \REGISTERS_reg[11][26]  ( .D(n1238), .CK(net338102), .Q(n821) );
  DFF_X1 \REGISTERS_reg[11][25]  ( .D(n1260), .CK(net338102), .Q(n820) );
  DFF_X1 \REGISTERS_reg[11][24]  ( .D(n1282), .CK(net338102), .Q(n819) );
  DFF_X1 \REGISTERS_reg[11][23]  ( .D(n1304), .CK(net338102), .Q(n818) );
  DFF_X1 \REGISTERS_reg[11][22]  ( .D(n1326), .CK(net338102), .Q(n817) );
  DFF_X1 \REGISTERS_reg[11][21]  ( .D(n1348), .CK(net338102), .Q(n815) );
  DFF_X1 \REGISTERS_reg[11][20]  ( .D(n1370), .CK(net338102), .Q(n814) );
  DFF_X1 \REGISTERS_reg[11][19]  ( .D(n1392), .CK(net338102), .Q(n813) );
  DFF_X1 \REGISTERS_reg[11][18]  ( .D(n1414), .CK(net338102), .Q(n812) );
  DFF_X1 \REGISTERS_reg[11][17]  ( .D(n1436), .CK(net338102), .Q(n811) );
  DFF_X1 \REGISTERS_reg[11][16]  ( .D(n1458), .CK(net338102), .Q(n810) );
  DFF_X1 \REGISTERS_reg[11][15]  ( .D(n1480), .CK(net338102), .Q(n809) );
  DFF_X1 \REGISTERS_reg[11][14]  ( .D(n1502), .CK(net338102), .Q(n808) );
  DFF_X1 \REGISTERS_reg[11][13]  ( .D(n1524), .CK(net338102), .Q(n807) );
  DFF_X1 \REGISTERS_reg[11][12]  ( .D(n1546), .CK(net338102), .Q(n806) );
  DFF_X1 \REGISTERS_reg[11][11]  ( .D(n1568), .CK(net338102), .Q(n805) );
  DFF_X1 \REGISTERS_reg[11][10]  ( .D(n1590), .CK(net338102), .Q(n804) );
  DFF_X1 \REGISTERS_reg[11][9]  ( .D(n1612), .CK(net338102), .Q(n803) );
  DFF_X1 \REGISTERS_reg[11][8]  ( .D(n1634), .CK(net338102), .Q(n802) );
  DFF_X1 \REGISTERS_reg[11][7]  ( .D(n1656), .CK(net338102), .Q(n801) );
  DFF_X1 \REGISTERS_reg[11][6]  ( .D(n1678), .CK(net338102), .Q(n800) );
  DFF_X1 \REGISTERS_reg[11][5]  ( .D(n1700), .CK(net338102), .Q(n799) );
  DFF_X1 \REGISTERS_reg[11][4]  ( .D(n1722), .CK(net338102), .Q(n798) );
  DFF_X1 \REGISTERS_reg[11][3]  ( .D(n1744), .CK(net338102), .Q(n797) );
  DFF_X1 \REGISTERS_reg[11][2]  ( .D(n1766), .CK(net338102), .Q(n796) );
  DFF_X1 \REGISTERS_reg[11][1]  ( .D(n1788), .CK(net338102), .Q(n794) );
  DFF_X1 \REGISTERS_reg[11][0]  ( .D(n1810), .CK(net338102), .Q(n793) );
  DFF_X1 \REGISTERS_reg[12][31]  ( .D(n1094), .CK(net338107), .Q(n792) );
  DFF_X1 \REGISTERS_reg[12][30]  ( .D(n1150), .CK(net338107), .Q(n791) );
  DFF_X1 \REGISTERS_reg[12][29]  ( .D(n1172), .CK(net338107), .Q(n790) );
  DFF_X1 \REGISTERS_reg[12][28]  ( .D(n1194), .CK(net338107), .Q(n789) );
  DFF_X1 \REGISTERS_reg[12][27]  ( .D(n1216), .CK(net338107), .Q(n788) );
  DFF_X1 \REGISTERS_reg[12][26]  ( .D(n1238), .CK(net338107), .Q(n787) );
  DFF_X1 \REGISTERS_reg[12][25]  ( .D(n1260), .CK(net338107), .Q(n786) );
  DFF_X1 \REGISTERS_reg[12][24]  ( .D(n1282), .CK(net338107), .Q(n785) );
  DFF_X1 \REGISTERS_reg[12][23]  ( .D(n1304), .CK(net338107), .Q(n784) );
  DFF_X1 \REGISTERS_reg[12][22]  ( .D(n1326), .CK(net338107), .Q(n783) );
  DFF_X1 \REGISTERS_reg[12][21]  ( .D(n1348), .CK(net338107), .Q(n782) );
  DFF_X1 \REGISTERS_reg[12][20]  ( .D(n1370), .CK(net338107), .Q(n781) );
  DFF_X1 \REGISTERS_reg[12][19]  ( .D(n1392), .CK(net338107), .Q(n780) );
  DFF_X1 \REGISTERS_reg[12][18]  ( .D(n1414), .CK(net338107), .Q(n779) );
  DFF_X1 \REGISTERS_reg[12][17]  ( .D(n1436), .CK(net338107), .Q(n778) );
  DFF_X1 \REGISTERS_reg[12][16]  ( .D(n1458), .CK(net338107), .Q(n777) );
  DFF_X1 \REGISTERS_reg[12][15]  ( .D(n1480), .CK(net338107), .Q(n776) );
  DFF_X1 \REGISTERS_reg[12][14]  ( .D(n1502), .CK(net338107), .Q(n775) );
  DFF_X1 \REGISTERS_reg[12][13]  ( .D(n1524), .CK(net338107), .Q(n773) );
  DFF_X1 \REGISTERS_reg[12][12]  ( .D(n1546), .CK(net338107), .Q(n772) );
  DFF_X1 \REGISTERS_reg[12][11]  ( .D(n1568), .CK(net338107), .Q(n771) );
  DFF_X1 \REGISTERS_reg[12][10]  ( .D(n1590), .CK(net338107), .Q(n770) );
  DFF_X1 \REGISTERS_reg[12][9]  ( .D(n1612), .CK(net338107), .Q(n769) );
  DFF_X1 \REGISTERS_reg[12][8]  ( .D(n1634), .CK(net338107), .Q(n768) );
  DFF_X1 \REGISTERS_reg[12][7]  ( .D(n1656), .CK(net338107), .Q(n767) );
  DFF_X1 \REGISTERS_reg[12][6]  ( .D(n1678), .CK(net338107), .Q(n766) );
  DFF_X1 \REGISTERS_reg[12][5]  ( .D(n1700), .CK(net338107), .Q(n765) );
  DFF_X1 \REGISTERS_reg[12][4]  ( .D(n1722), .CK(net338107), .Q(n764) );
  DFF_X1 \REGISTERS_reg[12][3]  ( .D(n1744), .CK(net338107), .Q(n763) );
  DFF_X1 \REGISTERS_reg[12][2]  ( .D(n1766), .CK(net338107), .Q(n762) );
  DFF_X1 \REGISTERS_reg[12][1]  ( .D(n1788), .CK(net338107), .Q(n761) );
  DFF_X1 \REGISTERS_reg[12][0]  ( .D(n1810), .CK(net338107), .Q(n760) );
  DFF_X1 \REGISTERS_reg[13][31]  ( .D(n1094), .CK(net338112), .Q(n759) );
  DFF_X1 \REGISTERS_reg[13][30]  ( .D(n1150), .CK(net338112), .Q(n758) );
  DFF_X1 \REGISTERS_reg[13][29]  ( .D(n1172), .CK(net338112), .Q(n757) );
  DFF_X1 \REGISTERS_reg[13][28]  ( .D(n1194), .CK(net338112), .Q(n756) );
  DFF_X1 \REGISTERS_reg[13][27]  ( .D(n1216), .CK(net338112), .Q(n755) );
  DFF_X1 \REGISTERS_reg[13][26]  ( .D(n1238), .CK(net338112), .Q(n754) );
  DFF_X1 \REGISTERS_reg[13][25]  ( .D(n1260), .CK(net338112), .Q(n752) );
  DFF_X1 \REGISTERS_reg[13][24]  ( .D(n1282), .CK(net338112), .Q(n751) );
  DFF_X1 \REGISTERS_reg[13][23]  ( .D(n1304), .CK(net338112), .Q(n750) );
  DFF_X1 \REGISTERS_reg[13][22]  ( .D(n1326), .CK(net338112), .Q(n749) );
  DFF_X1 \REGISTERS_reg[13][21]  ( .D(n1348), .CK(net338112), .Q(n748) );
  DFF_X1 \REGISTERS_reg[13][20]  ( .D(n1370), .CK(net338112), .Q(n747) );
  DFF_X1 \REGISTERS_reg[13][19]  ( .D(n1392), .CK(net338112), .Q(n746) );
  DFF_X1 \REGISTERS_reg[13][18]  ( .D(n1414), .CK(net338112), .Q(n745) );
  DFF_X1 \REGISTERS_reg[13][17]  ( .D(n1436), .CK(net338112), .Q(n744) );
  DFF_X1 \REGISTERS_reg[13][16]  ( .D(n1458), .CK(net338112), .Q(n743) );
  DFF_X1 \REGISTERS_reg[13][15]  ( .D(n1480), .CK(net338112), .Q(n742) );
  DFF_X1 \REGISTERS_reg[13][14]  ( .D(n1502), .CK(net338112), .Q(n741) );
  DFF_X1 \REGISTERS_reg[13][13]  ( .D(n1524), .CK(net338112), .Q(n740) );
  DFF_X1 \REGISTERS_reg[13][12]  ( .D(n1546), .CK(net338112), .Q(n739) );
  DFF_X1 \REGISTERS_reg[13][11]  ( .D(n1568), .CK(net338112), .Q(n738) );
  DFF_X1 \REGISTERS_reg[13][10]  ( .D(n1590), .CK(net338112), .Q(n737) );
  DFF_X1 \REGISTERS_reg[13][9]  ( .D(n1612), .CK(net338112), .Q(n736) );
  DFF_X1 \REGISTERS_reg[13][8]  ( .D(n1634), .CK(net338112), .Q(n735) );
  DFF_X1 \REGISTERS_reg[13][7]  ( .D(n1656), .CK(net338112), .Q(n734) );
  DFF_X1 \REGISTERS_reg[13][6]  ( .D(n1678), .CK(net338112), .Q(n733) );
  DFF_X1 \REGISTERS_reg[13][5]  ( .D(n1700), .CK(net338112), .Q(n731) );
  DFF_X1 \REGISTERS_reg[13][4]  ( .D(n1722), .CK(net338112), .Q(n730) );
  DFF_X1 \REGISTERS_reg[13][3]  ( .D(n1744), .CK(net338112), .Q(n729) );
  DFF_X1 \REGISTERS_reg[13][2]  ( .D(n1766), .CK(net338112), .Q(n728) );
  DFF_X1 \REGISTERS_reg[13][1]  ( .D(n1788), .CK(net338112), .Q(n727) );
  DFF_X1 \REGISTERS_reg[13][0]  ( .D(n1810), .CK(net338112), .Q(n726) );
  DFF_X1 \REGISTERS_reg[14][31]  ( .D(n1094), .CK(net338117), .Q(n725) );
  DFF_X1 \REGISTERS_reg[14][30]  ( .D(n1150), .CK(net338117), .Q(n724) );
  DFF_X1 \REGISTERS_reg[14][29]  ( .D(n1172), .CK(net338117), .Q(n723) );
  DFF_X1 \REGISTERS_reg[14][28]  ( .D(n1194), .CK(net338117), .Q(n722) );
  DFF_X1 \REGISTERS_reg[14][27]  ( .D(n1216), .CK(net338117), .Q(n721) );
  DFF_X1 \REGISTERS_reg[14][26]  ( .D(n1238), .CK(net338117), .Q(n720) );
  DFF_X1 \REGISTERS_reg[14][25]  ( .D(n1260), .CK(net338117), .Q(n719) );
  DFF_X1 \REGISTERS_reg[14][24]  ( .D(n1282), .CK(net338117), .Q(n718) );
  DFF_X1 \REGISTERS_reg[14][23]  ( .D(n1304), .CK(net338117), .Q(n717) );
  DFF_X1 \REGISTERS_reg[14][22]  ( .D(n1326), .CK(net338117), .Q(n716) );
  DFF_X1 \REGISTERS_reg[14][21]  ( .D(n1348), .CK(net338117), .Q(n715) );
  DFF_X1 \REGISTERS_reg[14][20]  ( .D(n1370), .CK(net338117), .Q(n714) );
  DFF_X1 \REGISTERS_reg[14][19]  ( .D(n1392), .CK(net338117), .Q(n713) );
  DFF_X1 \REGISTERS_reg[14][18]  ( .D(n1414), .CK(net338117), .Q(n712) );
  DFF_X1 \REGISTERS_reg[14][17]  ( .D(n1436), .CK(net338117), .Q(n710) );
  DFF_X1 \REGISTERS_reg[14][16]  ( .D(n1458), .CK(net338117), .Q(n709) );
  DFF_X1 \REGISTERS_reg[14][15]  ( .D(n1480), .CK(net338117), .Q(n708) );
  DFF_X1 \REGISTERS_reg[14][14]  ( .D(n1502), .CK(net338117), .Q(n707) );
  DFF_X1 \REGISTERS_reg[14][13]  ( .D(n1524), .CK(net338117), .Q(n706) );
  DFF_X1 \REGISTERS_reg[14][12]  ( .D(n1546), .CK(net338117), .Q(n705) );
  DFF_X1 \REGISTERS_reg[14][11]  ( .D(n1568), .CK(net338117), .Q(n704) );
  DFF_X1 \REGISTERS_reg[14][10]  ( .D(n1590), .CK(net338117), .Q(n703) );
  DFF_X1 \REGISTERS_reg[14][9]  ( .D(n1612), .CK(net338117), .Q(n702) );
  DFF_X1 \REGISTERS_reg[14][8]  ( .D(n1634), .CK(net338117), .Q(n701) );
  DFF_X1 \REGISTERS_reg[14][7]  ( .D(n1656), .CK(net338117), .Q(n700) );
  DFF_X1 \REGISTERS_reg[14][6]  ( .D(n1678), .CK(net338117), .Q(n699) );
  DFF_X1 \REGISTERS_reg[14][5]  ( .D(n1700), .CK(net338117), .Q(n698) );
  DFF_X1 \REGISTERS_reg[14][4]  ( .D(n1722), .CK(net338117), .Q(n697) );
  DFF_X1 \REGISTERS_reg[14][3]  ( .D(n1744), .CK(net338117), .Q(n696) );
  DFF_X1 \REGISTERS_reg[14][2]  ( .D(n1766), .CK(net338117), .Q(n695) );
  DFF_X1 \REGISTERS_reg[14][1]  ( .D(n1788), .CK(net338117), .Q(n694) );
  DFF_X1 \REGISTERS_reg[14][0]  ( .D(n1810), .CK(net338117), .Q(n693) );
  DFF_X1 \REGISTERS_reg[15][31]  ( .D(n1094), .CK(net338122), .Q(n692) );
  DFF_X1 \REGISTERS_reg[15][30]  ( .D(n1150), .CK(net338122), .Q(n691) );
  DFF_X1 \REGISTERS_reg[15][29]  ( .D(n1172), .CK(net338122), .Q(n689) );
  DFF_X1 \REGISTERS_reg[15][28]  ( .D(n1194), .CK(net338122), .Q(n688) );
  DFF_X1 \REGISTERS_reg[15][27]  ( .D(n1216), .CK(net338122), .Q(n687) );
  DFF_X1 \REGISTERS_reg[15][26]  ( .D(n1238), .CK(net338122), .Q(n686) );
  DFF_X1 \REGISTERS_reg[15][25]  ( .D(n1260), .CK(net338122), .Q(n685) );
  DFF_X1 \REGISTERS_reg[15][24]  ( .D(n1282), .CK(net338122), .Q(n684) );
  DFF_X1 \REGISTERS_reg[15][23]  ( .D(n1304), .CK(net338122), .Q(n683) );
  DFF_X1 \REGISTERS_reg[15][22]  ( .D(n1326), .CK(net338122), .Q(n682) );
  DFF_X1 \REGISTERS_reg[15][21]  ( .D(n1348), .CK(net338122), .Q(n681) );
  DFF_X1 \REGISTERS_reg[15][20]  ( .D(n1370), .CK(net338122), .Q(n680) );
  DFF_X1 \REGISTERS_reg[15][19]  ( .D(n1392), .CK(net338122), .Q(n679) );
  DFF_X1 \REGISTERS_reg[15][18]  ( .D(n1414), .CK(net338122), .Q(n678) );
  DFF_X1 \REGISTERS_reg[15][17]  ( .D(n1436), .CK(net338122), .Q(n677) );
  DFF_X1 \REGISTERS_reg[15][16]  ( .D(n1458), .CK(net338122), .Q(n676) );
  DFF_X1 \REGISTERS_reg[15][15]  ( .D(n1480), .CK(net338122), .Q(n675) );
  DFF_X1 \REGISTERS_reg[15][14]  ( .D(n1502), .CK(net338122), .Q(n674) );
  DFF_X1 \REGISTERS_reg[15][13]  ( .D(n1524), .CK(net338122), .Q(n673) );
  DFF_X1 \REGISTERS_reg[15][12]  ( .D(n1546), .CK(net338122), .Q(n672) );
  DFF_X1 \REGISTERS_reg[15][11]  ( .D(n1568), .CK(net338122), .Q(n671) );
  DFF_X1 \REGISTERS_reg[15][10]  ( .D(n1590), .CK(net338122), .Q(n670) );
  DFF_X1 \REGISTERS_reg[15][9]  ( .D(n1612), .CK(net338122), .Q(n668) );
  DFF_X1 \REGISTERS_reg[15][8]  ( .D(n1634), .CK(net338122), .Q(n667) );
  DFF_X1 \REGISTERS_reg[15][7]  ( .D(n1656), .CK(net338122), .Q(n666) );
  DFF_X1 \REGISTERS_reg[15][6]  ( .D(n1678), .CK(net338122), .Q(n665) );
  DFF_X1 \REGISTERS_reg[15][5]  ( .D(n1700), .CK(net338122), .Q(n664) );
  DFF_X1 \REGISTERS_reg[15][4]  ( .D(n1722), .CK(net338122), .Q(n663) );
  DFF_X1 \REGISTERS_reg[15][3]  ( .D(n1744), .CK(net338122), .Q(n662) );
  DFF_X1 \REGISTERS_reg[15][2]  ( .D(n1766), .CK(net338122), .Q(n661) );
  DFF_X1 \REGISTERS_reg[15][1]  ( .D(n1788), .CK(net338122), .Q(n660) );
  DFF_X1 \REGISTERS_reg[15][0]  ( .D(n1810), .CK(net338122), .Q(n659) );
  DFF_X1 \REGISTERS_reg[16][31]  ( .D(n1094), .CK(net338127), .Q(n658) );
  DFF_X1 \REGISTERS_reg[16][30]  ( .D(n1150), .CK(net338127), .Q(n657) );
  DFF_X1 \REGISTERS_reg[16][29]  ( .D(n1172), .CK(net338127), .Q(n656) );
  DFF_X1 \REGISTERS_reg[16][28]  ( .D(n1194), .CK(net338127), .Q(n655) );
  DFF_X1 \REGISTERS_reg[16][27]  ( .D(n1216), .CK(net338127), .Q(n654) );
  DFF_X1 \REGISTERS_reg[16][26]  ( .D(n1238), .CK(net338127), .Q(n653) );
  DFF_X1 \REGISTERS_reg[16][25]  ( .D(n1260), .CK(net338127), .Q(n652) );
  DFF_X1 \REGISTERS_reg[16][24]  ( .D(n1282), .CK(net338127), .Q(n651) );
  DFF_X1 \REGISTERS_reg[16][23]  ( .D(n1304), .CK(net338127), .Q(n650) );
  DFF_X1 \REGISTERS_reg[16][22]  ( .D(n1326), .CK(net338127), .Q(n649) );
  DFF_X1 \REGISTERS_reg[16][21]  ( .D(n1348), .CK(net338127), .Q(n647) );
  DFF_X1 \REGISTERS_reg[16][20]  ( .D(n1370), .CK(net338127), .Q(n646) );
  DFF_X1 \REGISTERS_reg[16][19]  ( .D(n1392), .CK(net338127), .Q(n645) );
  DFF_X1 \REGISTERS_reg[16][18]  ( .D(n1414), .CK(net338127), .Q(n644) );
  DFF_X1 \REGISTERS_reg[16][17]  ( .D(n1436), .CK(net338127), .Q(n643) );
  DFF_X1 \REGISTERS_reg[16][16]  ( .D(n1458), .CK(net338127), .Q(n642) );
  DFF_X1 \REGISTERS_reg[16][15]  ( .D(n1480), .CK(net338127), .Q(n641) );
  DFF_X1 \REGISTERS_reg[16][14]  ( .D(n1502), .CK(net338127), .Q(n640) );
  DFF_X1 \REGISTERS_reg[16][13]  ( .D(n1524), .CK(net338127), .Q(n639) );
  DFF_X1 \REGISTERS_reg[16][12]  ( .D(n1546), .CK(net338127), .Q(n638) );
  DFF_X1 \REGISTERS_reg[16][11]  ( .D(n1568), .CK(net338127), .Q(n637) );
  DFF_X1 \REGISTERS_reg[16][10]  ( .D(n1590), .CK(net338127), .Q(n636) );
  DFF_X1 \REGISTERS_reg[16][9]  ( .D(n1612), .CK(net338127), .Q(n635) );
  DFF_X1 \REGISTERS_reg[16][8]  ( .D(n1634), .CK(net338127), .Q(n634) );
  DFF_X1 \REGISTERS_reg[16][7]  ( .D(n1656), .CK(net338127), .Q(n633) );
  DFF_X1 \REGISTERS_reg[16][6]  ( .D(n1678), .CK(net338127), .Q(n632) );
  DFF_X1 \REGISTERS_reg[16][5]  ( .D(n1700), .CK(net338127), .Q(n631) );
  DFF_X1 \REGISTERS_reg[16][4]  ( .D(n1722), .CK(net338127), .Q(n630) );
  DFF_X1 \REGISTERS_reg[16][3]  ( .D(n1744), .CK(net338127), .Q(n629) );
  DFF_X1 \REGISTERS_reg[16][2]  ( .D(n1766), .CK(net338127), .Q(n628) );
  DFF_X1 \REGISTERS_reg[16][1]  ( .D(n1788), .CK(net338127), .Q(n626) );
  DFF_X1 \REGISTERS_reg[16][0]  ( .D(n1810), .CK(net338127), .Q(n625) );
  DFF_X1 \REGISTERS_reg[17][31]  ( .D(n1094), .CK(net338132), .Q(n624) );
  DFF_X1 \REGISTERS_reg[17][30]  ( .D(n1150), .CK(net338132), .Q(n623) );
  DFF_X1 \REGISTERS_reg[17][29]  ( .D(n1172), .CK(net338132), .Q(n622) );
  DFF_X1 \REGISTERS_reg[17][28]  ( .D(n1194), .CK(net338132), .Q(n621) );
  DFF_X1 \REGISTERS_reg[17][27]  ( .D(n1216), .CK(net338132), .Q(n620) );
  DFF_X1 \REGISTERS_reg[17][26]  ( .D(n1238), .CK(net338132), .Q(n619) );
  DFF_X1 \REGISTERS_reg[17][25]  ( .D(n1260), .CK(net338132), .Q(n618) );
  DFF_X1 \REGISTERS_reg[17][24]  ( .D(n1282), .CK(net338132), .Q(n617) );
  DFF_X1 \REGISTERS_reg[17][23]  ( .D(n1304), .CK(net338132), .Q(n616) );
  DFF_X1 \REGISTERS_reg[17][22]  ( .D(n1326), .CK(net338132), .Q(n615) );
  DFF_X1 \REGISTERS_reg[17][21]  ( .D(n1348), .CK(net338132), .Q(n614) );
  DFF_X1 \REGISTERS_reg[17][20]  ( .D(n1370), .CK(net338132), .Q(n613) );
  DFF_X1 \REGISTERS_reg[17][19]  ( .D(n1392), .CK(net338132), .Q(n612) );
  DFF_X1 \REGISTERS_reg[17][18]  ( .D(n1414), .CK(net338132), .Q(n611) );
  DFF_X1 \REGISTERS_reg[17][17]  ( .D(n1436), .CK(net338132), .Q(n610) );
  DFF_X1 \REGISTERS_reg[17][16]  ( .D(n1458), .CK(net338132), .Q(n609) );
  DFF_X1 \REGISTERS_reg[17][15]  ( .D(n1480), .CK(net338132), .Q(n608) );
  DFF_X1 \REGISTERS_reg[17][14]  ( .D(n1502), .CK(net338132), .Q(n607) );
  DFF_X1 \REGISTERS_reg[17][13]  ( .D(n1524), .CK(net338132), .Q(n605) );
  DFF_X1 \REGISTERS_reg[17][12]  ( .D(n1546), .CK(net338132), .Q(n604) );
  DFF_X1 \REGISTERS_reg[17][11]  ( .D(n1568), .CK(net338132), .Q(n603) );
  DFF_X1 \REGISTERS_reg[17][10]  ( .D(n1590), .CK(net338132), .Q(n602) );
  DFF_X1 \REGISTERS_reg[17][9]  ( .D(n1612), .CK(net338132), .Q(n601) );
  DFF_X1 \REGISTERS_reg[17][8]  ( .D(n1634), .CK(net338132), .Q(n600) );
  DFF_X1 \REGISTERS_reg[17][7]  ( .D(n1656), .CK(net338132), .Q(n599) );
  DFF_X1 \REGISTERS_reg[17][6]  ( .D(n1678), .CK(net338132), .Q(n598) );
  DFF_X1 \REGISTERS_reg[17][5]  ( .D(n1700), .CK(net338132), .Q(n597) );
  DFF_X1 \REGISTERS_reg[17][4]  ( .D(n1722), .CK(net338132), .Q(n596) );
  DFF_X1 \REGISTERS_reg[17][3]  ( .D(n1744), .CK(net338132), .Q(n595) );
  DFF_X1 \REGISTERS_reg[17][2]  ( .D(n1766), .CK(net338132), .Q(n594) );
  DFF_X1 \REGISTERS_reg[17][1]  ( .D(n1788), .CK(net338132), .Q(n593) );
  DFF_X1 \REGISTERS_reg[17][0]  ( .D(n1810), .CK(net338132), .Q(n592) );
  DFF_X1 \REGISTERS_reg[18][31]  ( .D(n1094), .CK(net338137), .Q(n591) );
  DFF_X1 \REGISTERS_reg[18][30]  ( .D(n1150), .CK(net338137), .Q(n590) );
  DFF_X1 \REGISTERS_reg[18][29]  ( .D(n1172), .CK(net338137), .Q(n589) );
  DFF_X1 \REGISTERS_reg[18][28]  ( .D(n1194), .CK(net338137), .Q(n588) );
  DFF_X1 \REGISTERS_reg[18][27]  ( .D(n1216), .CK(net338137), .Q(n587) );
  DFF_X1 \REGISTERS_reg[18][26]  ( .D(n1238), .CK(net338137), .Q(n586) );
  DFF_X1 \REGISTERS_reg[18][25]  ( .D(n1260), .CK(net338137), .Q(n584) );
  DFF_X1 \REGISTERS_reg[18][24]  ( .D(n1282), .CK(net338137), .Q(n583) );
  DFF_X1 \REGISTERS_reg[18][23]  ( .D(n1304), .CK(net338137), .Q(n582) );
  DFF_X1 \REGISTERS_reg[18][22]  ( .D(n1326), .CK(net338137), .Q(n581) );
  DFF_X1 \REGISTERS_reg[18][21]  ( .D(n1348), .CK(net338137), .Q(n580) );
  DFF_X1 \REGISTERS_reg[18][20]  ( .D(n1370), .CK(net338137), .Q(n579) );
  DFF_X1 \REGISTERS_reg[18][19]  ( .D(n1392), .CK(net338137), .Q(n578) );
  DFF_X1 \REGISTERS_reg[18][18]  ( .D(n1414), .CK(net338137), .Q(n577) );
  DFF_X1 \REGISTERS_reg[18][17]  ( .D(n1436), .CK(net338137), .Q(n576) );
  DFF_X1 \REGISTERS_reg[18][16]  ( .D(n1458), .CK(net338137), .Q(n575) );
  DFF_X1 \REGISTERS_reg[18][15]  ( .D(n1480), .CK(net338137), .Q(n574) );
  DFF_X1 \REGISTERS_reg[18][14]  ( .D(n1502), .CK(net338137), .Q(n573) );
  DFF_X1 \REGISTERS_reg[18][13]  ( .D(n1524), .CK(net338137), .Q(n572) );
  DFF_X1 \REGISTERS_reg[18][12]  ( .D(n1546), .CK(net338137), .Q(n571) );
  DFF_X1 \REGISTERS_reg[18][11]  ( .D(n1568), .CK(net338137), .Q(n570) );
  DFF_X1 \REGISTERS_reg[18][10]  ( .D(n1590), .CK(net338137), .Q(n569) );
  DFF_X1 \REGISTERS_reg[18][9]  ( .D(n1612), .CK(net338137), .Q(n568) );
  DFF_X1 \REGISTERS_reg[18][8]  ( .D(n1634), .CK(net338137), .Q(n567) );
  DFF_X1 \REGISTERS_reg[18][7]  ( .D(n1656), .CK(net338137), .Q(n566) );
  DFF_X1 \REGISTERS_reg[18][6]  ( .D(n1678), .CK(net338137), .Q(n565) );
  DFF_X1 \REGISTERS_reg[18][5]  ( .D(n1700), .CK(net338137), .Q(n563) );
  DFF_X1 \REGISTERS_reg[18][4]  ( .D(n1722), .CK(net338137), .Q(n562) );
  DFF_X1 \REGISTERS_reg[18][3]  ( .D(n1744), .CK(net338137), .Q(n561) );
  DFF_X1 \REGISTERS_reg[18][2]  ( .D(n1766), .CK(net338137), .Q(n560) );
  DFF_X1 \REGISTERS_reg[18][1]  ( .D(n1788), .CK(net338137), .Q(n559) );
  DFF_X1 \REGISTERS_reg[18][0]  ( .D(n1810), .CK(net338137), .Q(n558) );
  DFF_X1 \REGISTERS_reg[19][31]  ( .D(n1094), .CK(net338142), .Q(n557) );
  DFF_X1 \REGISTERS_reg[19][30]  ( .D(n1150), .CK(net338142), .Q(n556) );
  DFF_X1 \REGISTERS_reg[19][29]  ( .D(n1172), .CK(net338142), .Q(n555) );
  DFF_X1 \REGISTERS_reg[19][28]  ( .D(n1194), .CK(net338142), .Q(n554) );
  DFF_X1 \REGISTERS_reg[19][27]  ( .D(n1216), .CK(net338142), .Q(n553) );
  DFF_X1 \REGISTERS_reg[19][26]  ( .D(n1238), .CK(net338142), .Q(n552) );
  DFF_X1 \REGISTERS_reg[19][25]  ( .D(n1260), .CK(net338142), .Q(n551) );
  DFF_X1 \REGISTERS_reg[19][24]  ( .D(n1282), .CK(net338142), .Q(n550) );
  DFF_X1 \REGISTERS_reg[19][23]  ( .D(n1304), .CK(net338142), .Q(n549) );
  DFF_X1 \REGISTERS_reg[19][22]  ( .D(n1326), .CK(net338142), .Q(n548) );
  DFF_X1 \REGISTERS_reg[19][21]  ( .D(n1348), .CK(net338142), .Q(n547) );
  DFF_X1 \REGISTERS_reg[19][20]  ( .D(n1370), .CK(net338142), .Q(n546) );
  DFF_X1 \REGISTERS_reg[19][19]  ( .D(n1392), .CK(net338142), .Q(n545) );
  DFF_X1 \REGISTERS_reg[19][18]  ( .D(n1414), .CK(net338142), .Q(n544) );
  DFF_X1 \REGISTERS_reg[19][17]  ( .D(n1436), .CK(net338142), .Q(n542) );
  DFF_X1 \REGISTERS_reg[19][16]  ( .D(n1458), .CK(net338142), .Q(n541) );
  DFF_X1 \REGISTERS_reg[19][15]  ( .D(n1480), .CK(net338142), .Q(n540) );
  DFF_X1 \REGISTERS_reg[19][14]  ( .D(n1502), .CK(net338142), .Q(n539) );
  DFF_X1 \REGISTERS_reg[19][13]  ( .D(n1524), .CK(net338142), .Q(n538) );
  DFF_X1 \REGISTERS_reg[19][12]  ( .D(n1546), .CK(net338142), .Q(n537) );
  DFF_X1 \REGISTERS_reg[19][11]  ( .D(n1568), .CK(net338142), .Q(n536) );
  DFF_X1 \REGISTERS_reg[19][10]  ( .D(n1590), .CK(net338142), .Q(n535) );
  DFF_X1 \REGISTERS_reg[19][9]  ( .D(n1612), .CK(net338142), .Q(n534) );
  DFF_X1 \REGISTERS_reg[19][8]  ( .D(n1634), .CK(net338142), .Q(n533) );
  DFF_X1 \REGISTERS_reg[19][7]  ( .D(n1656), .CK(net338142), .Q(n532) );
  DFF_X1 \REGISTERS_reg[19][6]  ( .D(n1678), .CK(net338142), .Q(n531) );
  DFF_X1 \REGISTERS_reg[19][5]  ( .D(n1700), .CK(net338142), .Q(n530) );
  DFF_X1 \REGISTERS_reg[19][4]  ( .D(n1722), .CK(net338142), .Q(n529) );
  DFF_X1 \REGISTERS_reg[19][3]  ( .D(n1744), .CK(net338142), .Q(n528) );
  DFF_X1 \REGISTERS_reg[19][2]  ( .D(n1766), .CK(net338142), .Q(n527) );
  DFF_X1 \REGISTERS_reg[19][1]  ( .D(n1788), .CK(net338142), .Q(n526) );
  DFF_X1 \REGISTERS_reg[19][0]  ( .D(n1810), .CK(net338142), .Q(n525) );
  DFF_X1 \REGISTERS_reg[20][31]  ( .D(n1094), .CK(net338147), .Q(n524) );
  DFF_X1 \REGISTERS_reg[20][30]  ( .D(n1150), .CK(net338147), .Q(n523) );
  DFF_X1 \REGISTERS_reg[20][29]  ( .D(n1172), .CK(net338147), .Q(n521) );
  DFF_X1 \REGISTERS_reg[20][28]  ( .D(n1194), .CK(net338147), .Q(n520) );
  DFF_X1 \REGISTERS_reg[20][27]  ( .D(n1216), .CK(net338147), .Q(n519) );
  DFF_X1 \REGISTERS_reg[20][26]  ( .D(n1238), .CK(net338147), .Q(n518) );
  DFF_X1 \REGISTERS_reg[20][25]  ( .D(n1260), .CK(net338147), .Q(n517) );
  DFF_X1 \REGISTERS_reg[20][24]  ( .D(n1282), .CK(net338147), .Q(n516) );
  DFF_X1 \REGISTERS_reg[20][23]  ( .D(n1304), .CK(net338147), .Q(n515) );
  DFF_X1 \REGISTERS_reg[20][22]  ( .D(n1326), .CK(net338147), .Q(n514) );
  DFF_X1 \REGISTERS_reg[20][21]  ( .D(n1348), .CK(net338147), .Q(n513) );
  DFF_X1 \REGISTERS_reg[20][20]  ( .D(n1370), .CK(net338147), .Q(n512) );
  DFF_X1 \REGISTERS_reg[20][19]  ( .D(n1392), .CK(net338147), .Q(n511) );
  DFF_X1 \REGISTERS_reg[20][18]  ( .D(n1414), .CK(net338147), .Q(n510) );
  DFF_X1 \REGISTERS_reg[20][17]  ( .D(n1436), .CK(net338147), .Q(n509) );
  DFF_X1 \REGISTERS_reg[20][16]  ( .D(n1458), .CK(net338147), .Q(n508) );
  DFF_X1 \REGISTERS_reg[20][15]  ( .D(n1480), .CK(net338147), .Q(n507) );
  DFF_X1 \REGISTERS_reg[20][14]  ( .D(n1502), .CK(net338147), .Q(n506) );
  DFF_X1 \REGISTERS_reg[20][13]  ( .D(n1524), .CK(net338147), .Q(n505) );
  DFF_X1 \REGISTERS_reg[20][12]  ( .D(n1546), .CK(net338147), .Q(n504) );
  DFF_X1 \REGISTERS_reg[20][11]  ( .D(n1568), .CK(net338147), .Q(n503) );
  DFF_X1 \REGISTERS_reg[20][10]  ( .D(n1590), .CK(net338147), .Q(n502) );
  DFF_X1 \REGISTERS_reg[20][9]  ( .D(n1612), .CK(net338147), .Q(n500) );
  DFF_X1 \REGISTERS_reg[20][8]  ( .D(n1634), .CK(net338147), .Q(n499) );
  DFF_X1 \REGISTERS_reg[20][7]  ( .D(n1656), .CK(net338147), .Q(n498) );
  DFF_X1 \REGISTERS_reg[20][6]  ( .D(n1678), .CK(net338147), .Q(n497) );
  DFF_X1 \REGISTERS_reg[20][5]  ( .D(n1700), .CK(net338147), .Q(n496) );
  DFF_X1 \REGISTERS_reg[20][4]  ( .D(n1722), .CK(net338147), .Q(n495) );
  DFF_X1 \REGISTERS_reg[20][3]  ( .D(n1744), .CK(net338147), .Q(n494) );
  DFF_X1 \REGISTERS_reg[20][2]  ( .D(n1766), .CK(net338147), .Q(n493) );
  DFF_X1 \REGISTERS_reg[20][1]  ( .D(n1788), .CK(net338147), .Q(n492) );
  DFF_X1 \REGISTERS_reg[20][0]  ( .D(n1810), .CK(net338147), .Q(n491) );
  DFF_X1 \REGISTERS_reg[21][31]  ( .D(n1094), .CK(net338152), .Q(n490) );
  DFF_X1 \REGISTERS_reg[21][30]  ( .D(n1150), .CK(net338152), .Q(n489) );
  DFF_X1 \REGISTERS_reg[21][29]  ( .D(n1172), .CK(net338152), .Q(n488) );
  DFF_X1 \REGISTERS_reg[21][28]  ( .D(n1194), .CK(net338152), .Q(n487) );
  DFF_X1 \REGISTERS_reg[21][27]  ( .D(n1216), .CK(net338152), .Q(n486) );
  DFF_X1 \REGISTERS_reg[21][26]  ( .D(n1238), .CK(net338152), .Q(n485) );
  DFF_X1 \REGISTERS_reg[21][25]  ( .D(n1260), .CK(net338152), .Q(n484) );
  DFF_X1 \REGISTERS_reg[21][24]  ( .D(n1282), .CK(net338152), .Q(n483) );
  DFF_X1 \REGISTERS_reg[21][23]  ( .D(n1304), .CK(net338152), .Q(n482) );
  DFF_X1 \REGISTERS_reg[21][22]  ( .D(n1326), .CK(net338152), .Q(n481) );
  DFF_X1 \REGISTERS_reg[21][21]  ( .D(n1348), .CK(net338152), .Q(n479) );
  DFF_X1 \REGISTERS_reg[21][20]  ( .D(n1370), .CK(net338152), .Q(n478) );
  DFF_X1 \REGISTERS_reg[21][19]  ( .D(n1392), .CK(net338152), .Q(n477) );
  DFF_X1 \REGISTERS_reg[21][18]  ( .D(n1414), .CK(net338152), .Q(n476) );
  DFF_X1 \REGISTERS_reg[21][17]  ( .D(n1436), .CK(net338152), .Q(n475) );
  DFF_X1 \REGISTERS_reg[21][16]  ( .D(n1458), .CK(net338152), .Q(n474) );
  DFF_X1 \REGISTERS_reg[21][15]  ( .D(n1480), .CK(net338152), .Q(n473) );
  DFF_X1 \REGISTERS_reg[21][14]  ( .D(n1502), .CK(net338152), .Q(n472) );
  DFF_X1 \REGISTERS_reg[21][13]  ( .D(n1524), .CK(net338152), .Q(n471) );
  DFF_X1 \REGISTERS_reg[21][12]  ( .D(n1546), .CK(net338152), .Q(n470) );
  DFF_X1 \REGISTERS_reg[21][11]  ( .D(n1568), .CK(net338152), .Q(n469) );
  DFF_X1 \REGISTERS_reg[21][10]  ( .D(n1590), .CK(net338152), .Q(n468) );
  DFF_X1 \REGISTERS_reg[21][9]  ( .D(n1612), .CK(net338152), .Q(n467) );
  DFF_X1 \REGISTERS_reg[21][8]  ( .D(n1634), .CK(net338152), .Q(n466) );
  DFF_X1 \REGISTERS_reg[21][7]  ( .D(n1656), .CK(net338152), .Q(n465) );
  DFF_X1 \REGISTERS_reg[21][6]  ( .D(n1678), .CK(net338152), .Q(n464) );
  DFF_X1 \REGISTERS_reg[21][5]  ( .D(n1700), .CK(net338152), .Q(n463) );
  DFF_X1 \REGISTERS_reg[21][4]  ( .D(n1722), .CK(net338152), .Q(n462) );
  DFF_X1 \REGISTERS_reg[21][3]  ( .D(n1744), .CK(net338152), .Q(n461) );
  DFF_X1 \REGISTERS_reg[21][2]  ( .D(n1766), .CK(net338152), .Q(n460) );
  DFF_X1 \REGISTERS_reg[21][1]  ( .D(n1788), .CK(net338152), .Q(n458) );
  DFF_X1 \REGISTERS_reg[21][0]  ( .D(n1810), .CK(net338152), .Q(n457) );
  DFF_X1 \REGISTERS_reg[22][31]  ( .D(n1094), .CK(net338157), .Q(n456) );
  DFF_X1 \REGISTERS_reg[22][30]  ( .D(n1150), .CK(net338157), .Q(n455) );
  DFF_X1 \REGISTERS_reg[22][29]  ( .D(n1172), .CK(net338157), .Q(n454) );
  DFF_X1 \REGISTERS_reg[22][28]  ( .D(n1194), .CK(net338157), .Q(n453) );
  DFF_X1 \REGISTERS_reg[22][27]  ( .D(n1216), .CK(net338157), .Q(n452) );
  DFF_X1 \REGISTERS_reg[22][26]  ( .D(n1238), .CK(net338157), .Q(n451) );
  DFF_X1 \REGISTERS_reg[22][25]  ( .D(n1260), .CK(net338157), .Q(n450) );
  DFF_X1 \REGISTERS_reg[22][24]  ( .D(n1282), .CK(net338157), .Q(n449) );
  DFF_X1 \REGISTERS_reg[22][23]  ( .D(n1304), .CK(net338157), .Q(n448) );
  DFF_X1 \REGISTERS_reg[22][22]  ( .D(n1326), .CK(net338157), .Q(n447) );
  DFF_X1 \REGISTERS_reg[22][21]  ( .D(n1348), .CK(net338157), .Q(n446) );
  DFF_X1 \REGISTERS_reg[22][20]  ( .D(n1370), .CK(net338157), .Q(n445) );
  DFF_X1 \REGISTERS_reg[22][19]  ( .D(n1392), .CK(net338157), .Q(n444) );
  DFF_X1 \REGISTERS_reg[22][18]  ( .D(n1414), .CK(net338157), .Q(n443) );
  DFF_X1 \REGISTERS_reg[22][17]  ( .D(n1436), .CK(net338157), .Q(n442) );
  DFF_X1 \REGISTERS_reg[22][16]  ( .D(n1458), .CK(net338157), .Q(n441) );
  DFF_X1 \REGISTERS_reg[22][15]  ( .D(n1480), .CK(net338157), .Q(n440) );
  DFF_X1 \REGISTERS_reg[22][14]  ( .D(n1502), .CK(net338157), .Q(n439) );
  DFF_X1 \REGISTERS_reg[22][13]  ( .D(n1524), .CK(net338157), .Q(n437) );
  DFF_X1 \REGISTERS_reg[22][12]  ( .D(n1546), .CK(net338157), .Q(n436) );
  DFF_X1 \REGISTERS_reg[22][11]  ( .D(n1568), .CK(net338157), .Q(n435) );
  DFF_X1 \REGISTERS_reg[22][10]  ( .D(n1590), .CK(net338157), .Q(n434) );
  DFF_X1 \REGISTERS_reg[22][9]  ( .D(n1612), .CK(net338157), .Q(n433) );
  DFF_X1 \REGISTERS_reg[22][8]  ( .D(n1634), .CK(net338157), .Q(n432) );
  DFF_X1 \REGISTERS_reg[22][7]  ( .D(n1656), .CK(net338157), .Q(n431) );
  DFF_X1 \REGISTERS_reg[22][6]  ( .D(n1678), .CK(net338157), .Q(n430) );
  DFF_X1 \REGISTERS_reg[22][5]  ( .D(n1700), .CK(net338157), .Q(n429) );
  DFF_X1 \REGISTERS_reg[22][4]  ( .D(n1722), .CK(net338157), .Q(n428) );
  DFF_X1 \REGISTERS_reg[22][3]  ( .D(n1744), .CK(net338157), .Q(n427) );
  DFF_X1 \REGISTERS_reg[22][2]  ( .D(n1766), .CK(net338157), .Q(n426) );
  DFF_X1 \REGISTERS_reg[22][1]  ( .D(n1788), .CK(net338157), .Q(n425) );
  DFF_X1 \REGISTERS_reg[22][0]  ( .D(n1810), .CK(net338157), .Q(n424) );
  DFF_X1 \REGISTERS_reg[23][31]  ( .D(n1094), .CK(net338162), .Q(n423) );
  DFF_X1 \REGISTERS_reg[23][30]  ( .D(n1150), .CK(net338162), .Q(n422) );
  DFF_X1 \REGISTERS_reg[23][29]  ( .D(n1172), .CK(net338162), .Q(n421) );
  DFF_X1 \REGISTERS_reg[23][28]  ( .D(n1194), .CK(net338162), .Q(n420) );
  DFF_X1 \REGISTERS_reg[23][27]  ( .D(n1216), .CK(net338162), .Q(n419) );
  DFF_X1 \REGISTERS_reg[23][26]  ( .D(n1238), .CK(net338162), .Q(n418) );
  DFF_X1 \REGISTERS_reg[23][25]  ( .D(n1260), .CK(net338162), .Q(n417) );
  DFF_X1 \REGISTERS_reg[23][24]  ( .D(n1282), .CK(net338162), .Q(n416) );
  DFF_X1 \REGISTERS_reg[23][23]  ( .D(n1304), .CK(net338162), .Q(n415) );
  DFF_X1 \REGISTERS_reg[23][22]  ( .D(n1326), .CK(net338162), .Q(n414) );
  DFF_X1 \REGISTERS_reg[23][21]  ( .D(n1348), .CK(net338162), .Q(n413) );
  DFF_X1 \REGISTERS_reg[23][20]  ( .D(n1370), .CK(net338162), .Q(n412) );
  DFF_X1 \REGISTERS_reg[23][19]  ( .D(n1392), .CK(net338162), .Q(n411) );
  DFF_X1 \REGISTERS_reg[23][18]  ( .D(n1414), .CK(net338162), .Q(n410) );
  DFF_X1 \REGISTERS_reg[23][17]  ( .D(n1436), .CK(net338162), .Q(n409) );
  DFF_X1 \REGISTERS_reg[23][16]  ( .D(n1458), .CK(net338162), .Q(n408) );
  DFF_X1 \REGISTERS_reg[23][15]  ( .D(n1480), .CK(net338162), .Q(n407) );
  DFF_X1 \REGISTERS_reg[23][14]  ( .D(n1502), .CK(net338162), .Q(n406) );
  DFF_X1 \REGISTERS_reg[23][13]  ( .D(n1524), .CK(net338162), .Q(n405) );
  DFF_X1 \REGISTERS_reg[23][12]  ( .D(n1546), .CK(net338162), .Q(n404) );
  DFF_X1 \REGISTERS_reg[23][11]  ( .D(n1568), .CK(net338162), .Q(n403) );
  DFF_X1 \REGISTERS_reg[23][10]  ( .D(n1590), .CK(net338162), .Q(n402) );
  DFF_X1 \REGISTERS_reg[23][9]  ( .D(n1612), .CK(net338162), .Q(n401) );
  DFF_X1 \REGISTERS_reg[23][8]  ( .D(n1634), .CK(net338162), .Q(n400) );
  DFF_X1 \REGISTERS_reg[23][7]  ( .D(n1656), .CK(net338162), .Q(n399) );
  DFF_X1 \REGISTERS_reg[23][6]  ( .D(n1678), .CK(net338162), .Q(n398) );
  DFF_X1 \REGISTERS_reg[23][5]  ( .D(n1700), .CK(net338162), .Q(n397) );
  DFF_X1 \REGISTERS_reg[23][4]  ( .D(n1722), .CK(net338162), .Q(n396) );
  DFF_X1 \REGISTERS_reg[23][3]  ( .D(n1744), .CK(net338162), .Q(n395) );
  DFF_X1 \REGISTERS_reg[23][2]  ( .D(n1766), .CK(net338162), .Q(n394) );
  DFF_X1 \REGISTERS_reg[23][1]  ( .D(n1788), .CK(net338162), .Q(n393) );
  DFF_X1 \REGISTERS_reg[23][0]  ( .D(n1810), .CK(net338162), .Q(n392) );
  DFF_X1 \REGISTERS_reg[24][31]  ( .D(n1094), .CK(net338167), .Q(n391) );
  DFF_X1 \REGISTERS_reg[24][30]  ( .D(n1150), .CK(net338167), .Q(n390) );
  DFF_X1 \REGISTERS_reg[24][29]  ( .D(n1172), .CK(net338167), .Q(n389) );
  DFF_X1 \REGISTERS_reg[24][28]  ( .D(n1194), .CK(net338167), .Q(n388) );
  DFF_X1 \REGISTERS_reg[24][27]  ( .D(n1216), .CK(net338167), .Q(n387) );
  DFF_X1 \REGISTERS_reg[24][26]  ( .D(n1238), .CK(net338167), .Q(n386) );
  DFF_X1 \REGISTERS_reg[24][25]  ( .D(n1260), .CK(net338167), .Q(n385) );
  DFF_X1 \REGISTERS_reg[24][24]  ( .D(n1282), .CK(net338167), .Q(n384) );
  DFF_X1 \REGISTERS_reg[24][23]  ( .D(n1304), .CK(net338167), .Q(n383) );
  DFF_X1 \REGISTERS_reg[24][22]  ( .D(n1326), .CK(net338167), .Q(n382) );
  DFF_X1 \REGISTERS_reg[24][21]  ( .D(n1348), .CK(net338167), .Q(n381) );
  DFF_X1 \REGISTERS_reg[24][20]  ( .D(n1370), .CK(net338167), .Q(n380) );
  DFF_X1 \REGISTERS_reg[24][19]  ( .D(n1392), .CK(net338167), .Q(n379) );
  DFF_X1 \REGISTERS_reg[24][18]  ( .D(n1414), .CK(net338167), .Q(n378) );
  DFF_X1 \REGISTERS_reg[24][17]  ( .D(n1436), .CK(net338167), .Q(n377) );
  DFF_X1 \REGISTERS_reg[24][16]  ( .D(n1458), .CK(net338167), .Q(n376) );
  DFF_X1 \REGISTERS_reg[24][15]  ( .D(n1480), .CK(net338167), .Q(n375) );
  DFF_X1 \REGISTERS_reg[24][14]  ( .D(n1502), .CK(net338167), .Q(n374) );
  DFF_X1 \REGISTERS_reg[24][13]  ( .D(n1524), .CK(net338167), .Q(n373) );
  DFF_X1 \REGISTERS_reg[24][12]  ( .D(n1546), .CK(net338167), .Q(n372) );
  DFF_X1 \REGISTERS_reg[24][11]  ( .D(n1568), .CK(net338167), .Q(n371) );
  DFF_X1 \REGISTERS_reg[24][10]  ( .D(n1590), .CK(net338167), .Q(n370) );
  DFF_X1 \REGISTERS_reg[24][9]  ( .D(n1612), .CK(net338167), .Q(n369) );
  DFF_X1 \REGISTERS_reg[24][8]  ( .D(n1634), .CK(net338167), .Q(n368) );
  DFF_X1 \REGISTERS_reg[24][7]  ( .D(n1656), .CK(net338167), .Q(n367) );
  DFF_X1 \REGISTERS_reg[24][6]  ( .D(n1678), .CK(net338167), .Q(n366) );
  DFF_X1 \REGISTERS_reg[24][5]  ( .D(n1700), .CK(net338167), .Q(n365) );
  DFF_X1 \REGISTERS_reg[24][4]  ( .D(n1722), .CK(net338167), .Q(n364) );
  DFF_X1 \REGISTERS_reg[24][3]  ( .D(n1744), .CK(net338167), .Q(n363) );
  DFF_X1 \REGISTERS_reg[24][2]  ( .D(n1766), .CK(net338167), .Q(n362) );
  DFF_X1 \REGISTERS_reg[24][1]  ( .D(n1788), .CK(net338167), .Q(n361) );
  DFF_X1 \REGISTERS_reg[24][0]  ( .D(n1810), .CK(net338167), .Q(n360) );
  DFF_X1 \REGISTERS_reg[25][31]  ( .D(n1094), .CK(net338172), .Q(n359) );
  DFF_X1 \REGISTERS_reg[25][30]  ( .D(n1150), .CK(net338172), .Q(n358) );
  DFF_X1 \REGISTERS_reg[25][29]  ( .D(n1172), .CK(net338172), .Q(n357) );
  DFF_X1 \REGISTERS_reg[25][28]  ( .D(n1194), .CK(net338172), .Q(n356) );
  DFF_X1 \REGISTERS_reg[25][27]  ( .D(n1216), .CK(net338172), .Q(n355) );
  DFF_X1 \REGISTERS_reg[25][26]  ( .D(n1238), .CK(net338172), .Q(n354) );
  DFF_X1 \REGISTERS_reg[25][25]  ( .D(n1260), .CK(net338172), .Q(n353) );
  DFF_X1 \REGISTERS_reg[25][24]  ( .D(n1282), .CK(net338172), .Q(n352) );
  DFF_X1 \REGISTERS_reg[25][23]  ( .D(n1304), .CK(net338172), .Q(n351) );
  DFF_X1 \REGISTERS_reg[25][22]  ( .D(n1326), .CK(net338172), .Q(n350) );
  DFF_X1 \REGISTERS_reg[25][21]  ( .D(n1348), .CK(net338172), .Q(n349) );
  DFF_X1 \REGISTERS_reg[25][20]  ( .D(n1370), .CK(net338172), .Q(n348) );
  DFF_X1 \REGISTERS_reg[25][19]  ( .D(n1392), .CK(net338172), .Q(n347) );
  DFF_X1 \REGISTERS_reg[25][18]  ( .D(n1414), .CK(net338172), .Q(n346) );
  DFF_X1 \REGISTERS_reg[25][17]  ( .D(n1436), .CK(net338172), .Q(n345) );
  DFF_X1 \REGISTERS_reg[25][16]  ( .D(n1458), .CK(net338172), .Q(n344) );
  DFF_X1 \REGISTERS_reg[25][15]  ( .D(n1480), .CK(net338172), .Q(n343) );
  DFF_X1 \REGISTERS_reg[25][14]  ( .D(n1502), .CK(net338172), .Q(n342) );
  DFF_X1 \REGISTERS_reg[25][13]  ( .D(n1524), .CK(net338172), .Q(n341) );
  DFF_X1 \REGISTERS_reg[25][12]  ( .D(n1546), .CK(net338172), .Q(n340) );
  DFF_X1 \REGISTERS_reg[25][11]  ( .D(n1568), .CK(net338172), .Q(n339) );
  DFF_X1 \REGISTERS_reg[25][10]  ( .D(n1590), .CK(net338172), .Q(n338) );
  DFF_X1 \REGISTERS_reg[25][9]  ( .D(n1612), .CK(net338172), .Q(n337) );
  DFF_X1 \REGISTERS_reg[25][8]  ( .D(n1634), .CK(net338172), .Q(n336) );
  DFF_X1 \REGISTERS_reg[25][7]  ( .D(n1656), .CK(net338172), .Q(n335) );
  DFF_X1 \REGISTERS_reg[25][6]  ( .D(n1678), .CK(net338172), .Q(n334) );
  DFF_X1 \REGISTERS_reg[25][5]  ( .D(n1700), .CK(net338172), .Q(n333) );
  DFF_X1 \REGISTERS_reg[25][4]  ( .D(n1722), .CK(net338172), .Q(n332) );
  DFF_X1 \REGISTERS_reg[25][3]  ( .D(n1744), .CK(net338172), .Q(n331) );
  DFF_X1 \REGISTERS_reg[25][2]  ( .D(n1766), .CK(net338172), .Q(n330) );
  DFF_X1 \REGISTERS_reg[25][1]  ( .D(n1788), .CK(net338172), .Q(n329) );
  DFF_X1 \REGISTERS_reg[25][0]  ( .D(n1810), .CK(net338172), .Q(n328) );
  DFF_X1 \REGISTERS_reg[26][31]  ( .D(n1094), .CK(net338177), .Q(n327) );
  DFF_X1 \REGISTERS_reg[26][30]  ( .D(n1150), .CK(net338177), .Q(n326) );
  DFF_X1 \REGISTERS_reg[26][29]  ( .D(n1172), .CK(net338177), .Q(n325) );
  DFF_X1 \REGISTERS_reg[26][28]  ( .D(n1194), .CK(net338177), .Q(n324) );
  DFF_X1 \REGISTERS_reg[26][27]  ( .D(n1216), .CK(net338177), .Q(n323) );
  DFF_X1 \REGISTERS_reg[26][26]  ( .D(n1238), .CK(net338177), .Q(n322) );
  DFF_X1 \REGISTERS_reg[26][25]  ( .D(n1260), .CK(net338177), .Q(n321) );
  DFF_X1 \REGISTERS_reg[26][24]  ( .D(n1282), .CK(net338177), .Q(n320) );
  DFF_X1 \REGISTERS_reg[26][23]  ( .D(n1304), .CK(net338177), .Q(n319) );
  DFF_X1 \REGISTERS_reg[26][22]  ( .D(n1326), .CK(net338177), .Q(n318) );
  DFF_X1 \REGISTERS_reg[26][21]  ( .D(n1348), .CK(net338177), .Q(n317) );
  DFF_X1 \REGISTERS_reg[26][20]  ( .D(n1370), .CK(net338177), .Q(n316) );
  DFF_X1 \REGISTERS_reg[26][19]  ( .D(n1392), .CK(net338177), .Q(n315) );
  DFF_X1 \REGISTERS_reg[26][18]  ( .D(n1414), .CK(net338177), .Q(n314) );
  DFF_X1 \REGISTERS_reg[26][17]  ( .D(n1436), .CK(net338177), .Q(n313) );
  DFF_X1 \REGISTERS_reg[26][16]  ( .D(n1458), .CK(net338177), .Q(n312) );
  DFF_X1 \REGISTERS_reg[26][15]  ( .D(n1480), .CK(net338177), .Q(n311) );
  DFF_X1 \REGISTERS_reg[26][14]  ( .D(n1502), .CK(net338177), .Q(n310) );
  DFF_X1 \REGISTERS_reg[26][13]  ( .D(n1524), .CK(net338177), .Q(n309) );
  DFF_X1 \REGISTERS_reg[26][12]  ( .D(n1546), .CK(net338177), .Q(n308) );
  DFF_X1 \REGISTERS_reg[26][11]  ( .D(n1568), .CK(net338177), .Q(n307) );
  DFF_X1 \REGISTERS_reg[26][10]  ( .D(n1590), .CK(net338177), .Q(n306) );
  DFF_X1 \REGISTERS_reg[26][9]  ( .D(n1612), .CK(net338177), .Q(n305) );
  DFF_X1 \REGISTERS_reg[26][8]  ( .D(n1634), .CK(net338177), .Q(n304) );
  DFF_X1 \REGISTERS_reg[26][7]  ( .D(n1656), .CK(net338177), .Q(n303) );
  DFF_X1 \REGISTERS_reg[26][6]  ( .D(n1678), .CK(net338177), .Q(n302) );
  DFF_X1 \REGISTERS_reg[26][5]  ( .D(n1700), .CK(net338177), .Q(n301) );
  DFF_X1 \REGISTERS_reg[26][4]  ( .D(n1722), .CK(net338177), .Q(n300) );
  DFF_X1 \REGISTERS_reg[26][3]  ( .D(n1744), .CK(net338177), .Q(n299) );
  DFF_X1 \REGISTERS_reg[26][2]  ( .D(n1766), .CK(net338177), .Q(n298) );
  DFF_X1 \REGISTERS_reg[26][1]  ( .D(n1788), .CK(net338177), .Q(n297) );
  DFF_X1 \REGISTERS_reg[26][0]  ( .D(n1810), .CK(net338177), .Q(n296) );
  DFF_X1 \REGISTERS_reg[27][31]  ( .D(n1094), .CK(net338182), .Q(n295) );
  DFF_X1 \REGISTERS_reg[27][30]  ( .D(n1150), .CK(net338182), .Q(n294) );
  DFF_X1 \REGISTERS_reg[27][29]  ( .D(n1172), .CK(net338182), .Q(n293) );
  DFF_X1 \REGISTERS_reg[27][28]  ( .D(n1194), .CK(net338182), .Q(n292) );
  DFF_X1 \REGISTERS_reg[27][27]  ( .D(n1216), .CK(net338182), .Q(n291) );
  DFF_X1 \REGISTERS_reg[27][26]  ( .D(n1238), .CK(net338182), .Q(n290) );
  DFF_X1 \REGISTERS_reg[27][25]  ( .D(n1260), .CK(net338182), .Q(n289) );
  DFF_X1 \REGISTERS_reg[27][24]  ( .D(n1282), .CK(net338182), .Q(n288) );
  DFF_X1 \REGISTERS_reg[27][23]  ( .D(n1304), .CK(net338182), .Q(n287) );
  DFF_X1 \REGISTERS_reg[27][22]  ( .D(n1326), .CK(net338182), .Q(n286) );
  DFF_X1 \REGISTERS_reg[27][21]  ( .D(n1348), .CK(net338182), .Q(n285) );
  DFF_X1 \REGISTERS_reg[27][20]  ( .D(n1370), .CK(net338182), .Q(n284) );
  DFF_X1 \REGISTERS_reg[27][19]  ( .D(n1392), .CK(net338182), .Q(n283) );
  DFF_X1 \REGISTERS_reg[27][18]  ( .D(n1414), .CK(net338182), .Q(n282) );
  DFF_X1 \REGISTERS_reg[27][17]  ( .D(n1436), .CK(net338182), .Q(n281) );
  DFF_X1 \REGISTERS_reg[27][16]  ( .D(n1458), .CK(net338182), .Q(n280) );
  DFF_X1 \REGISTERS_reg[27][15]  ( .D(n1480), .CK(net338182), .Q(n279) );
  DFF_X1 \REGISTERS_reg[27][14]  ( .D(n1502), .CK(net338182), .Q(n278) );
  DFF_X1 \REGISTERS_reg[27][13]  ( .D(n1524), .CK(net338182), .Q(n277) );
  DFF_X1 \REGISTERS_reg[27][12]  ( .D(n1546), .CK(net338182), .Q(n276) );
  DFF_X1 \REGISTERS_reg[27][11]  ( .D(n1568), .CK(net338182), .Q(n275) );
  DFF_X1 \REGISTERS_reg[27][10]  ( .D(n1590), .CK(net338182), .Q(n274) );
  DFF_X1 \REGISTERS_reg[27][9]  ( .D(n1612), .CK(net338182), .Q(n273) );
  DFF_X1 \REGISTERS_reg[27][8]  ( .D(n1634), .CK(net338182), .Q(n272) );
  DFF_X1 \REGISTERS_reg[27][7]  ( .D(n1656), .CK(net338182), .Q(n271) );
  DFF_X1 \REGISTERS_reg[27][6]  ( .D(n1678), .CK(net338182), .Q(n270) );
  DFF_X1 \REGISTERS_reg[27][5]  ( .D(n1700), .CK(net338182), .Q(n269) );
  DFF_X1 \REGISTERS_reg[27][4]  ( .D(n1722), .CK(net338182), .Q(n268) );
  DFF_X1 \REGISTERS_reg[27][3]  ( .D(n1744), .CK(net338182), .Q(n267) );
  DFF_X1 \REGISTERS_reg[27][2]  ( .D(n1766), .CK(net338182), .Q(n266) );
  DFF_X1 \REGISTERS_reg[27][1]  ( .D(n1788), .CK(net338182), .Q(n265) );
  DFF_X1 \REGISTERS_reg[27][0]  ( .D(n1810), .CK(net338182), .Q(n264) );
  DFF_X1 \REGISTERS_reg[28][31]  ( .D(n1094), .CK(net338187), .Q(n263) );
  DFF_X1 \REGISTERS_reg[28][30]  ( .D(n1150), .CK(net338187), .Q(n262) );
  DFF_X1 \REGISTERS_reg[28][29]  ( .D(n1172), .CK(net338187), .Q(n261) );
  DFF_X1 \REGISTERS_reg[28][28]  ( .D(n1194), .CK(net338187), .Q(n260) );
  DFF_X1 \REGISTERS_reg[28][27]  ( .D(n1216), .CK(net338187), .Q(n259) );
  DFF_X1 \REGISTERS_reg[28][26]  ( .D(n1238), .CK(net338187), .Q(n258) );
  DFF_X1 \REGISTERS_reg[28][25]  ( .D(n1260), .CK(net338187), .Q(n257) );
  DFF_X1 \REGISTERS_reg[28][24]  ( .D(n1282), .CK(net338187), .Q(n256) );
  DFF_X1 \REGISTERS_reg[28][23]  ( .D(n1304), .CK(net338187), .Q(n255) );
  DFF_X1 \REGISTERS_reg[28][22]  ( .D(n1326), .CK(net338187), .Q(n254) );
  DFF_X1 \REGISTERS_reg[28][21]  ( .D(n1348), .CK(net338187), .Q(n253) );
  DFF_X1 \REGISTERS_reg[28][20]  ( .D(n1370), .CK(net338187), .Q(n252) );
  DFF_X1 \REGISTERS_reg[28][19]  ( .D(n1392), .CK(net338187), .Q(n251) );
  DFF_X1 \REGISTERS_reg[28][18]  ( .D(n1414), .CK(net338187), .Q(n250) );
  DFF_X1 \REGISTERS_reg[28][17]  ( .D(n1436), .CK(net338187), .Q(n249) );
  DFF_X1 \REGISTERS_reg[28][16]  ( .D(n1458), .CK(net338187), .Q(n248) );
  DFF_X1 \REGISTERS_reg[28][15]  ( .D(n1480), .CK(net338187), .Q(n247) );
  DFF_X1 \REGISTERS_reg[28][14]  ( .D(n1502), .CK(net338187), .Q(n246) );
  DFF_X1 \REGISTERS_reg[28][13]  ( .D(n1524), .CK(net338187), .Q(n245) );
  DFF_X1 \REGISTERS_reg[28][12]  ( .D(n1546), .CK(net338187), .Q(n244) );
  DFF_X1 \REGISTERS_reg[28][11]  ( .D(n1568), .CK(net338187), .Q(n243) );
  DFF_X1 \REGISTERS_reg[28][10]  ( .D(n1590), .CK(net338187), .Q(n242) );
  DFF_X1 \REGISTERS_reg[28][9]  ( .D(n1612), .CK(net338187), .Q(n241) );
  DFF_X1 \REGISTERS_reg[28][8]  ( .D(n1634), .CK(net338187), .Q(n240) );
  DFF_X1 \REGISTERS_reg[28][7]  ( .D(n1656), .CK(net338187), .Q(n239) );
  DFF_X1 \REGISTERS_reg[28][6]  ( .D(n1678), .CK(net338187), .Q(n238) );
  DFF_X1 \REGISTERS_reg[28][5]  ( .D(n1700), .CK(net338187), .Q(n237) );
  DFF_X1 \REGISTERS_reg[28][4]  ( .D(n1722), .CK(net338187), .Q(n236) );
  DFF_X1 \REGISTERS_reg[28][3]  ( .D(n1744), .CK(net338187), .Q(n235) );
  DFF_X1 \REGISTERS_reg[28][2]  ( .D(n1766), .CK(net338187), .Q(n234) );
  DFF_X1 \REGISTERS_reg[28][1]  ( .D(n1788), .CK(net338187), .Q(n233) );
  DFF_X1 \REGISTERS_reg[28][0]  ( .D(n1810), .CK(net338187), .Q(n232) );
  DFF_X1 \REGISTERS_reg[29][31]  ( .D(n1094), .CK(net338192), .Q(n231) );
  DFF_X1 \REGISTERS_reg[29][30]  ( .D(n1150), .CK(net338192), .Q(n230) );
  DFF_X1 \REGISTERS_reg[29][29]  ( .D(n1172), .CK(net338192), .Q(n229) );
  DFF_X1 \REGISTERS_reg[29][28]  ( .D(n1194), .CK(net338192), .Q(n228) );
  DFF_X1 \REGISTERS_reg[29][27]  ( .D(n1216), .CK(net338192), .Q(n227) );
  DFF_X1 \REGISTERS_reg[29][26]  ( .D(n1238), .CK(net338192), .Q(n226) );
  DFF_X1 \REGISTERS_reg[29][25]  ( .D(n1260), .CK(net338192), .Q(n225) );
  DFF_X1 \REGISTERS_reg[29][24]  ( .D(n1282), .CK(net338192), .Q(n224) );
  DFF_X1 \REGISTERS_reg[29][23]  ( .D(n1304), .CK(net338192), .Q(n223) );
  DFF_X1 \REGISTERS_reg[29][22]  ( .D(n1326), .CK(net338192), .Q(n222) );
  DFF_X1 \REGISTERS_reg[29][21]  ( .D(n1348), .CK(net338192), .Q(n221) );
  DFF_X1 \REGISTERS_reg[29][20]  ( .D(n1370), .CK(net338192), .Q(n220) );
  DFF_X1 \REGISTERS_reg[29][19]  ( .D(n1392), .CK(net338192), .Q(n219) );
  DFF_X1 \REGISTERS_reg[29][18]  ( .D(n1414), .CK(net338192), .Q(n218) );
  DFF_X1 \REGISTERS_reg[29][17]  ( .D(n1436), .CK(net338192), .Q(n217) );
  DFF_X1 \REGISTERS_reg[29][16]  ( .D(n1458), .CK(net338192), .Q(n216) );
  DFF_X1 \REGISTERS_reg[29][15]  ( .D(n1480), .CK(net338192), .Q(n215) );
  DFF_X1 \REGISTERS_reg[29][14]  ( .D(n1502), .CK(net338192), .Q(n214) );
  DFF_X1 \REGISTERS_reg[29][13]  ( .D(n1524), .CK(net338192), .Q(n213) );
  DFF_X1 \REGISTERS_reg[29][12]  ( .D(n1546), .CK(net338192), .Q(n212) );
  DFF_X1 \REGISTERS_reg[29][11]  ( .D(n1568), .CK(net338192), .Q(n211) );
  DFF_X1 \REGISTERS_reg[29][10]  ( .D(n1590), .CK(net338192), .Q(n210) );
  DFF_X1 \REGISTERS_reg[29][9]  ( .D(n1612), .CK(net338192), .Q(n209) );
  DFF_X1 \REGISTERS_reg[29][8]  ( .D(n1634), .CK(net338192), .Q(n208) );
  DFF_X1 \REGISTERS_reg[29][7]  ( .D(n1656), .CK(net338192), .Q(n207) );
  DFF_X1 \REGISTERS_reg[29][6]  ( .D(n1678), .CK(net338192), .Q(n206) );
  DFF_X1 \REGISTERS_reg[29][5]  ( .D(n1700), .CK(net338192), .Q(n205) );
  DFF_X1 \REGISTERS_reg[29][4]  ( .D(n1722), .CK(net338192), .Q(n204) );
  DFF_X1 \REGISTERS_reg[29][3]  ( .D(n1744), .CK(net338192), .Q(n203) );
  DFF_X1 \REGISTERS_reg[29][2]  ( .D(n1766), .CK(net338192), .Q(n202) );
  DFF_X1 \REGISTERS_reg[29][1]  ( .D(n1788), .CK(net338192), .Q(n201) );
  DFF_X1 \REGISTERS_reg[29][0]  ( .D(n1810), .CK(net338192), .Q(n200) );
  DFF_X1 \REGISTERS_reg[30][31]  ( .D(n1094), .CK(net338197), .Q(n199) );
  DFF_X1 \REGISTERS_reg[30][30]  ( .D(n1150), .CK(net338197), .Q(n198) );
  DFF_X1 \REGISTERS_reg[30][29]  ( .D(n1172), .CK(net338197), .Q(n197) );
  DFF_X1 \REGISTERS_reg[30][28]  ( .D(n1194), .CK(net338197), .Q(n196) );
  DFF_X1 \REGISTERS_reg[30][27]  ( .D(n1216), .CK(net338197), .Q(n195) );
  DFF_X1 \REGISTERS_reg[30][26]  ( .D(n1238), .CK(net338197), .Q(n194) );
  DFF_X1 \REGISTERS_reg[30][25]  ( .D(n1260), .CK(net338197), .Q(n193) );
  DFF_X1 \REGISTERS_reg[30][24]  ( .D(n1282), .CK(net338197), .Q(n192) );
  DFF_X1 \REGISTERS_reg[30][23]  ( .D(n1304), .CK(net338197), .Q(n191) );
  DFF_X1 \REGISTERS_reg[30][22]  ( .D(n1326), .CK(net338197), .Q(n190) );
  DFF_X1 \REGISTERS_reg[30][21]  ( .D(n1348), .CK(net338197), .Q(n189) );
  DFF_X1 \REGISTERS_reg[30][20]  ( .D(n1370), .CK(net338197), .Q(n188) );
  DFF_X1 \REGISTERS_reg[30][19]  ( .D(n1392), .CK(net338197), .Q(n187) );
  DFF_X1 \REGISTERS_reg[30][18]  ( .D(n1414), .CK(net338197), .Q(n186) );
  DFF_X1 \REGISTERS_reg[30][17]  ( .D(n1436), .CK(net338197), .Q(n185) );
  DFF_X1 \REGISTERS_reg[30][16]  ( .D(n1458), .CK(net338197), .Q(n184) );
  DFF_X1 \REGISTERS_reg[30][15]  ( .D(n1480), .CK(net338197), .Q(n183) );
  DFF_X1 \REGISTERS_reg[30][14]  ( .D(n1502), .CK(net338197), .Q(n182) );
  DFF_X1 \REGISTERS_reg[30][13]  ( .D(n1524), .CK(net338197), .Q(n181) );
  DFF_X1 \REGISTERS_reg[30][12]  ( .D(n1546), .CK(net338197), .Q(n180) );
  DFF_X1 \REGISTERS_reg[30][11]  ( .D(n1568), .CK(net338197), .Q(n179) );
  DFF_X1 \REGISTERS_reg[30][10]  ( .D(n1590), .CK(net338197), .Q(n178) );
  DFF_X1 \REGISTERS_reg[30][9]  ( .D(n1612), .CK(net338197), .Q(n175) );
  DFF_X1 \REGISTERS_reg[30][8]  ( .D(n1634), .CK(net338197), .Q(n164) );
  DFF_X1 \REGISTERS_reg[30][7]  ( .D(n1656), .CK(net338197), .Q(n153) );
  DFF_X1 \REGISTERS_reg[30][6]  ( .D(n1678), .CK(net338197), .Q(n142) );
  DFF_X1 \REGISTERS_reg[30][5]  ( .D(n1700), .CK(net338197), .Q(n131) );
  DFF_X1 \REGISTERS_reg[30][4]  ( .D(n1722), .CK(net338197), .Q(n120) );
  DFF_X1 \REGISTERS_reg[30][3]  ( .D(n1744), .CK(net338197), .Q(n109) );
  DFF_X1 \REGISTERS_reg[30][2]  ( .D(n1766), .CK(net338197), .Q(n97) );
  DFF_X1 \REGISTERS_reg[30][1]  ( .D(n1788), .CK(net338197), .Q(n75) );
  DFF_X1 \REGISTERS_reg[30][0]  ( .D(n1810), .CK(net338197), .Q(n53) );
  DFF_X1 \REGISTERS_reg[31][31]  ( .D(n1094), .CK(net338202), .Q(n1089) );
  DFF_X1 \OUT2_reg[31]  ( .D(N4616), .CK(net338042), .Q(OUT2[31]) );
  DFF_X1 \REGISTERS_reg[31][30]  ( .D(n1150), .CK(net338202), .Q(n1068) );
  DFF_X1 \OUT2_reg[30]  ( .D(N4614), .CK(net338042), .Q(OUT2[30]) );
  DFF_X1 \REGISTERS_reg[31][29]  ( .D(n1172), .CK(net338202), .Q(n1047) );
  DFF_X1 \OUT2_reg[29]  ( .D(N4612), .CK(net338042), .Q(OUT2[29]) );
  DFF_X1 \REGISTERS_reg[31][28]  ( .D(n1194), .CK(net338202), .Q(n1026) );
  DFF_X1 \OUT2_reg[28]  ( .D(N4610), .CK(net338042), .Q(OUT2[28]) );
  DFF_X1 \REGISTERS_reg[31][27]  ( .D(n1216), .CK(net338202), .Q(n1005) );
  DFF_X1 \OUT2_reg[27]  ( .D(N4608), .CK(net338042), .Q(OUT2[27]) );
  DFF_X1 \REGISTERS_reg[31][26]  ( .D(n1238), .CK(net338202), .Q(n984) );
  DFF_X1 \OUT2_reg[26]  ( .D(N4606), .CK(net338042), .Q(OUT2[26]) );
  DFF_X1 \REGISTERS_reg[31][25]  ( .D(n1260), .CK(net338202), .Q(n963) );
  DFF_X1 \OUT2_reg[25]  ( .D(N4604), .CK(net338042), .Q(OUT2[25]) );
  DFF_X1 \REGISTERS_reg[31][24]  ( .D(n1282), .CK(net338202), .Q(n942) );
  DFF_X1 \OUT2_reg[24]  ( .D(N4602), .CK(net338042), .Q(OUT2[24]) );
  DFF_X1 \REGISTERS_reg[31][23]  ( .D(n1304), .CK(net338202), .Q(n921) );
  DFF_X1 \OUT2_reg[23]  ( .D(N4600), .CK(net338042), .Q(OUT2[23]) );
  DFF_X1 \REGISTERS_reg[31][22]  ( .D(n1326), .CK(net338202), .Q(n900) );
  DFF_X1 \OUT2_reg[22]  ( .D(N4598), .CK(net338042), .Q(OUT2[22]) );
  DFF_X1 \REGISTERS_reg[31][21]  ( .D(n1348), .CK(net338202), .Q(n879) );
  DFF_X1 \OUT2_reg[21]  ( .D(N4596), .CK(net338042), .Q(OUT2[21]) );
  DFF_X1 \REGISTERS_reg[31][20]  ( .D(n1370), .CK(net338202), .Q(n858) );
  DFF_X1 \OUT2_reg[20]  ( .D(N4594), .CK(net338042), .Q(OUT2[20]) );
  DFF_X1 \REGISTERS_reg[31][19]  ( .D(n1392), .CK(net338202), .Q(n837) );
  DFF_X1 \OUT2_reg[19]  ( .D(N4592), .CK(net338042), .Q(OUT2[19]) );
  DFF_X1 \REGISTERS_reg[31][18]  ( .D(n1414), .CK(net338202), .Q(n816) );
  DFF_X1 \OUT2_reg[18]  ( .D(N4590), .CK(net338042), .Q(OUT2[18]) );
  DFF_X1 \REGISTERS_reg[31][17]  ( .D(n1436), .CK(net338202), .Q(n795) );
  DFF_X1 \OUT2_reg[17]  ( .D(N4588), .CK(net338042), .Q(OUT2[17]) );
  DFF_X1 \REGISTERS_reg[31][16]  ( .D(n1458), .CK(net338202), .Q(n774) );
  DFF_X1 \OUT2_reg[16]  ( .D(N4586), .CK(net338042), .Q(OUT2[16]) );
  DFF_X1 \REGISTERS_reg[31][15]  ( .D(n1480), .CK(net338202), .Q(n753) );
  DFF_X1 \OUT2_reg[15]  ( .D(N4584), .CK(net338042), .Q(OUT2[15]) );
  DFF_X1 \REGISTERS_reg[31][14]  ( .D(n1502), .CK(net338202), .Q(n732) );
  DFF_X1 \OUT2_reg[14]  ( .D(N4582), .CK(net338042), .Q(OUT2[14]) );
  DFF_X1 \REGISTERS_reg[31][13]  ( .D(n1524), .CK(net338202), .Q(n711) );
  DFF_X1 \OUT2_reg[13]  ( .D(N4580), .CK(net338042), .Q(OUT2[13]) );
  DFF_X1 \REGISTERS_reg[31][12]  ( .D(n1546), .CK(net338202), .Q(n690) );
  DFF_X1 \OUT2_reg[12]  ( .D(N4578), .CK(net338042), .Q(OUT2[12]) );
  DFF_X1 \REGISTERS_reg[31][11]  ( .D(n1568), .CK(net338202), .Q(n669) );
  DFF_X1 \OUT2_reg[11]  ( .D(N4576), .CK(net338042), .Q(OUT2[11]) );
  DFF_X1 \REGISTERS_reg[31][10]  ( .D(n1590), .CK(net338202), .Q(n648) );
  DFF_X1 \OUT2_reg[10]  ( .D(N4574), .CK(net338042), .Q(OUT2[10]) );
  DFF_X1 \REGISTERS_reg[31][9]  ( .D(n1612), .CK(net338202), .Q(n627) );
  DFF_X1 \OUT2_reg[9]  ( .D(N4572), .CK(net338042), .Q(OUT2[9]) );
  DFF_X1 \REGISTERS_reg[31][8]  ( .D(n1634), .CK(net338202), .Q(n606) );
  DFF_X1 \OUT2_reg[8]  ( .D(N4570), .CK(net338042), .Q(OUT2[8]) );
  DFF_X1 \REGISTERS_reg[31][7]  ( .D(n1656), .CK(net338202), .Q(n585) );
  DFF_X1 \OUT2_reg[7]  ( .D(N4568), .CK(net338042), .Q(OUT2[7]) );
  DFF_X1 \REGISTERS_reg[31][6]  ( .D(n1678), .CK(net338202), .Q(n564) );
  DFF_X1 \OUT2_reg[6]  ( .D(N4566), .CK(net338042), .Q(OUT2[6]) );
  DFF_X1 \REGISTERS_reg[31][5]  ( .D(n1700), .CK(net338202), .Q(n543) );
  DFF_X1 \OUT2_reg[5]  ( .D(N4564), .CK(net338042), .Q(OUT2[5]) );
  DFF_X1 \REGISTERS_reg[31][4]  ( .D(n1722), .CK(net338202), .Q(n522) );
  DFF_X1 \OUT2_reg[4]  ( .D(N4562), .CK(net338042), .Q(OUT2[4]) );
  DFF_X1 \REGISTERS_reg[31][3]  ( .D(n1744), .CK(net338202), .Q(n501) );
  DFF_X1 \OUT2_reg[3]  ( .D(N4560), .CK(net338042), .Q(OUT2[3]) );
  DFF_X1 \REGISTERS_reg[31][2]  ( .D(n1766), .CK(net338202), .Q(n480) );
  DFF_X1 \OUT2_reg[2]  ( .D(N4558), .CK(net338042), .Q(OUT2[2]) );
  DFF_X1 \REGISTERS_reg[31][1]  ( .D(n1788), .CK(net338202), .Q(n459) );
  DFF_X1 \OUT2_reg[1]  ( .D(N4556), .CK(net338042), .Q(OUT2[1]) );
  DFF_X1 \REGISTERS_reg[31][0]  ( .D(n1810), .CK(net338202), .Q(n438) );
  DFF_X1 \OUT2_reg[0]  ( .D(N4554), .CK(net338042), .Q(OUT2[0]) );
  DFF_X1 \OUT1_reg[31]  ( .D(N4552), .CK(net338207), .Q(OUT1[31]) );
  DFF_X1 \OUT1_reg[30]  ( .D(N4550), .CK(net338207), .Q(OUT1[30]) );
  DFF_X1 \OUT1_reg[29]  ( .D(N4548), .CK(net338207), .Q(OUT1[29]) );
  DFF_X1 \OUT1_reg[28]  ( .D(N4546), .CK(net338207), .Q(OUT1[28]) );
  DFF_X1 \OUT1_reg[27]  ( .D(N4544), .CK(net338207), .Q(OUT1[27]) );
  DFF_X1 \OUT1_reg[26]  ( .D(N4542), .CK(net338207), .Q(OUT1[26]) );
  DFF_X1 \OUT1_reg[25]  ( .D(N4540), .CK(net338207), .Q(OUT1[25]) );
  DFF_X1 \OUT1_reg[24]  ( .D(N4538), .CK(net338207), .Q(OUT1[24]) );
  DFF_X1 \OUT1_reg[23]  ( .D(N4536), .CK(net338207), .Q(OUT1[23]) );
  DFF_X1 \OUT1_reg[22]  ( .D(N4534), .CK(net338207), .Q(OUT1[22]) );
  DFF_X1 \OUT1_reg[21]  ( .D(N4532), .CK(net338207), .Q(OUT1[21]) );
  DFF_X1 \OUT1_reg[20]  ( .D(N4530), .CK(net338207), .Q(OUT1[20]) );
  DFF_X1 \OUT1_reg[19]  ( .D(N4528), .CK(net338207), .Q(OUT1[19]) );
  DFF_X1 \OUT1_reg[18]  ( .D(N4526), .CK(net338207), .Q(OUT1[18]) );
  DFF_X1 \OUT1_reg[17]  ( .D(N4524), .CK(net338207), .Q(OUT1[17]) );
  DFF_X1 \OUT1_reg[16]  ( .D(N4522), .CK(net338207), .Q(OUT1[16]) );
  DFF_X1 \OUT1_reg[15]  ( .D(N4520), .CK(net338207), .Q(OUT1[15]) );
  DFF_X1 \OUT1_reg[14]  ( .D(N4518), .CK(net338207), .Q(OUT1[14]) );
  DFF_X1 \OUT1_reg[13]  ( .D(N4516), .CK(net338207), .Q(OUT1[13]) );
  DFF_X1 \OUT1_reg[12]  ( .D(N4514), .CK(net338207), .Q(OUT1[12]) );
  DFF_X1 \OUT1_reg[11]  ( .D(N4512), .CK(net338207), .Q(OUT1[11]) );
  DFF_X1 \OUT1_reg[10]  ( .D(N4510), .CK(net338207), .Q(OUT1[10]) );
  DFF_X1 \OUT1_reg[9]  ( .D(N4508), .CK(net338207), .Q(OUT1[9]) );
  DFF_X1 \OUT1_reg[8]  ( .D(N4506), .CK(net338207), .Q(OUT1[8]) );
  DFF_X1 \OUT1_reg[7]  ( .D(N4504), .CK(net338207), .Q(OUT1[7]) );
  DFF_X1 \OUT1_reg[6]  ( .D(N4502), .CK(net338207), .Q(OUT1[6]) );
  DFF_X1 \OUT1_reg[5]  ( .D(N4500), .CK(net338207), .Q(OUT1[5]) );
  DFF_X1 \OUT1_reg[4]  ( .D(N4498), .CK(net338207), .Q(OUT1[4]) );
  DFF_X1 \OUT1_reg[3]  ( .D(N4496), .CK(net338207), .Q(OUT1[3]) );
  DFF_X1 \OUT1_reg[2]  ( .D(N4494), .CK(net338207), .Q(OUT1[2]) );
  DFF_X1 \OUT1_reg[1]  ( .D(N4492), .CK(net338207), .Q(OUT1[1]) );
  DFF_X1 \OUT1_reg[0]  ( .D(N4490), .CK(net338207), .Q(OUT1[0]) );
  SNPS_CLOCK_GATE_HIGH_dlx_regfile_0 clk_gate_OUT2_reg ( .CLK(Clk), .EN(N4615), 
        .ENCLK(net338042) );
  SNPS_CLOCK_GATE_HIGH_dlx_regfile_33 \clk_gate_REGISTERS_reg[0]  ( .CLK(Clk), 
        .EN(N4487), .ENCLK(net338047) );
  SNPS_CLOCK_GATE_HIGH_dlx_regfile_32 \clk_gate_REGISTERS_reg[1]  ( .CLK(Clk), 
        .EN(N4423), .ENCLK(net338052) );
  SNPS_CLOCK_GATE_HIGH_dlx_regfile_31 \clk_gate_REGISTERS_reg[2]  ( .CLK(Clk), 
        .EN(N4359), .ENCLK(net338057) );
  SNPS_CLOCK_GATE_HIGH_dlx_regfile_30 \clk_gate_REGISTERS_reg[3]  ( .CLK(Clk), 
        .EN(N4295), .ENCLK(net338062) );
  SNPS_CLOCK_GATE_HIGH_dlx_regfile_29 \clk_gate_REGISTERS_reg[4]  ( .CLK(Clk), 
        .EN(N4231), .ENCLK(net338067) );
  SNPS_CLOCK_GATE_HIGH_dlx_regfile_28 \clk_gate_REGISTERS_reg[5]  ( .CLK(Clk), 
        .EN(N4167), .ENCLK(net338072) );
  SNPS_CLOCK_GATE_HIGH_dlx_regfile_27 \clk_gate_REGISTERS_reg[6]  ( .CLK(Clk), 
        .EN(N4103), .ENCLK(net338077) );
  SNPS_CLOCK_GATE_HIGH_dlx_regfile_26 \clk_gate_REGISTERS_reg[7]  ( .CLK(Clk), 
        .EN(N4039), .ENCLK(net338082) );
  SNPS_CLOCK_GATE_HIGH_dlx_regfile_25 \clk_gate_REGISTERS_reg[8]  ( .CLK(Clk), 
        .EN(N3975), .ENCLK(net338087) );
  SNPS_CLOCK_GATE_HIGH_dlx_regfile_24 \clk_gate_REGISTERS_reg[9]  ( .CLK(Clk), 
        .EN(N3911), .ENCLK(net338092) );
  SNPS_CLOCK_GATE_HIGH_dlx_regfile_23 \clk_gate_REGISTERS_reg[10]  ( .CLK(Clk), 
        .EN(N3847), .ENCLK(net338097) );
  SNPS_CLOCK_GATE_HIGH_dlx_regfile_22 \clk_gate_REGISTERS_reg[11]  ( .CLK(Clk), 
        .EN(N3783), .ENCLK(net338102) );
  SNPS_CLOCK_GATE_HIGH_dlx_regfile_21 \clk_gate_REGISTERS_reg[12]  ( .CLK(Clk), 
        .EN(N3719), .ENCLK(net338107) );
  SNPS_CLOCK_GATE_HIGH_dlx_regfile_20 \clk_gate_REGISTERS_reg[13]  ( .CLK(Clk), 
        .EN(N3655), .ENCLK(net338112) );
  SNPS_CLOCK_GATE_HIGH_dlx_regfile_19 \clk_gate_REGISTERS_reg[14]  ( .CLK(Clk), 
        .EN(N3591), .ENCLK(net338117) );
  SNPS_CLOCK_GATE_HIGH_dlx_regfile_18 \clk_gate_REGISTERS_reg[15]  ( .CLK(Clk), 
        .EN(N3527), .ENCLK(net338122) );
  SNPS_CLOCK_GATE_HIGH_dlx_regfile_17 \clk_gate_REGISTERS_reg[16]  ( .CLK(Clk), 
        .EN(N3463), .ENCLK(net338127) );
  SNPS_CLOCK_GATE_HIGH_dlx_regfile_16 \clk_gate_REGISTERS_reg[17]  ( .CLK(Clk), 
        .EN(N3399), .ENCLK(net338132) );
  SNPS_CLOCK_GATE_HIGH_dlx_regfile_15 \clk_gate_REGISTERS_reg[18]  ( .CLK(Clk), 
        .EN(N3335), .ENCLK(net338137) );
  SNPS_CLOCK_GATE_HIGH_dlx_regfile_14 \clk_gate_REGISTERS_reg[19]  ( .CLK(Clk), 
        .EN(N3271), .ENCLK(net338142) );
  SNPS_CLOCK_GATE_HIGH_dlx_regfile_13 \clk_gate_REGISTERS_reg[20]  ( .CLK(Clk), 
        .EN(N3207), .ENCLK(net338147) );
  SNPS_CLOCK_GATE_HIGH_dlx_regfile_12 \clk_gate_REGISTERS_reg[21]  ( .CLK(Clk), 
        .EN(N3143), .ENCLK(net338152) );
  SNPS_CLOCK_GATE_HIGH_dlx_regfile_11 \clk_gate_REGISTERS_reg[22]  ( .CLK(Clk), 
        .EN(N3079), .ENCLK(net338157) );
  SNPS_CLOCK_GATE_HIGH_dlx_regfile_10 \clk_gate_REGISTERS_reg[23]  ( .CLK(Clk), 
        .EN(N3015), .ENCLK(net338162) );
  SNPS_CLOCK_GATE_HIGH_dlx_regfile_9 \clk_gate_REGISTERS_reg[24]  ( .CLK(Clk), 
        .EN(N2951), .ENCLK(net338167) );
  SNPS_CLOCK_GATE_HIGH_dlx_regfile_8 \clk_gate_REGISTERS_reg[25]  ( .CLK(Clk), 
        .EN(N2887), .ENCLK(net338172) );
  SNPS_CLOCK_GATE_HIGH_dlx_regfile_7 \clk_gate_REGISTERS_reg[26]  ( .CLK(Clk), 
        .EN(N2823), .ENCLK(net338177) );
  SNPS_CLOCK_GATE_HIGH_dlx_regfile_6 \clk_gate_REGISTERS_reg[27]  ( .CLK(Clk), 
        .EN(N2759), .ENCLK(net338182) );
  SNPS_CLOCK_GATE_HIGH_dlx_regfile_5 \clk_gate_REGISTERS_reg[28]  ( .CLK(Clk), 
        .EN(N2695), .ENCLK(net338187) );
  SNPS_CLOCK_GATE_HIGH_dlx_regfile_4 \clk_gate_REGISTERS_reg[29]  ( .CLK(Clk), 
        .EN(N2631), .ENCLK(net338192) );
  SNPS_CLOCK_GATE_HIGH_dlx_regfile_3 \clk_gate_REGISTERS_reg[30]  ( .CLK(Clk), 
        .EN(N2567), .ENCLK(net338197) );
  SNPS_CLOCK_GATE_HIGH_dlx_regfile_2 \clk_gate_REGISTERS_reg[31]  ( .CLK(Clk), 
        .EN(N2503), .ENCLK(net338202) );
  SNPS_CLOCK_GATE_HIGH_dlx_regfile_1 clk_gate_OUT1_reg ( .CLK(Clk), .EN(N4615), 
        .ENCLK(net338207) );
  INV_X1 U3 ( .A(N4487), .ZN(n51) );
  NAND2_X2 U4 ( .A1(n2575), .A2(n2597), .ZN(n1916) );
  NAND2_X2 U5 ( .A1(n1842), .A2(n1859), .ZN(n1138) );
  NAND2_X2 U6 ( .A1(n1842), .A2(n1864), .ZN(n1152) );
  NAND2_X2 U7 ( .A1(n1839), .A2(n1840), .ZN(n1113) );
  NAND2_X2 U8 ( .A1(n2572), .A2(n2573), .ZN(n1878) );
  NAND2_X2 U9 ( .A1(n2575), .A2(n2592), .ZN(n1903) );
  INV_X2 U10 ( .A(N4487), .ZN(n49) );
  INV_X1 U11 ( .A(N4487), .ZN(n47) );
  NAND2_X2 U12 ( .A1(n47), .A2(n1103), .ZN(n1102) );
  NAND2_X2 U13 ( .A1(n49), .A2(n1868), .ZN(n1867) );
  NAND3_X2 U14 ( .A1(n1819), .A2(n1820), .A3(n1821), .ZN(n1103) );
  NAND3_X2 U15 ( .A1(n1819), .A2(n2553), .A3(n2554), .ZN(n1868) );
  BUF_X1 U16 ( .A(n1154), .Z(n2) );
  BUF_X1 U17 ( .A(n1153), .Z(n1) );
  BUF_X1 U18 ( .A(n1156), .Z(n37) );
  BUF_X1 U19 ( .A(n1917), .Z(n41) );
  BUF_X1 U20 ( .A(n1883), .Z(n39) );
  BUF_X1 U21 ( .A(n1918), .Z(n43) );
  NAND2_X2 U22 ( .A1(DATAIN[12]), .A2(n51), .ZN(n1546) );
  NAND2_X2 U23 ( .A1(DATAIN[13]), .A2(n51), .ZN(n1524) );
  NAND2_X2 U24 ( .A1(DATAIN[14]), .A2(n51), .ZN(n1502) );
  NAND2_X2 U25 ( .A1(DATAIN[15]), .A2(n49), .ZN(n1480) );
  NAND2_X2 U26 ( .A1(DATAIN[16]), .A2(n49), .ZN(n1458) );
  NAND2_X2 U27 ( .A1(DATAIN[17]), .A2(n49), .ZN(n1436) );
  NAND2_X2 U28 ( .A1(DATAIN[18]), .A2(n49), .ZN(n1414) );
  NAND2_X2 U29 ( .A1(DATAIN[19]), .A2(n49), .ZN(n1392) );
  NAND2_X2 U30 ( .A1(DATAIN[20]), .A2(n49), .ZN(n1370) );
  NAND2_X2 U31 ( .A1(DATAIN[21]), .A2(n49), .ZN(n1348) );
  NAND2_X2 U32 ( .A1(DATAIN[22]), .A2(n49), .ZN(n1326) );
  NAND2_X2 U33 ( .A1(DATAIN[23]), .A2(n49), .ZN(n1304) );
  NAND2_X2 U34 ( .A1(DATAIN[24]), .A2(n49), .ZN(n1282) );
  NAND2_X2 U35 ( .A1(DATAIN[25]), .A2(n49), .ZN(n1260) );
  NAND2_X2 U36 ( .A1(DATAIN[26]), .A2(n49), .ZN(n1238) );
  NAND2_X2 U37 ( .A1(DATAIN[27]), .A2(n47), .ZN(n1216) );
  NAND2_X2 U38 ( .A1(DATAIN[28]), .A2(n47), .ZN(n1194) );
  NAND2_X2 U39 ( .A1(DATAIN[29]), .A2(n47), .ZN(n1172) );
  NAND2_X2 U40 ( .A1(DATAIN[30]), .A2(n47), .ZN(n1150) );
  NAND2_X2 U41 ( .A1(DATAIN[31]), .A2(n47), .ZN(n1094) );
  NAND2_X2 U42 ( .A1(DATAIN[0]), .A2(n49), .ZN(n1810) );
  NAND2_X2 U43 ( .A1(DATAIN[1]), .A2(n49), .ZN(n1788) );
  NAND2_X2 U44 ( .A1(DATAIN[2]), .A2(n47), .ZN(n1766) );
  NAND2_X2 U45 ( .A1(DATAIN[3]), .A2(n51), .ZN(n1744) );
  NAND2_X2 U46 ( .A1(DATAIN[4]), .A2(n51), .ZN(n1722) );
  NAND2_X2 U47 ( .A1(DATAIN[5]), .A2(n51), .ZN(n1700) );
  NAND2_X2 U48 ( .A1(DATAIN[6]), .A2(n51), .ZN(n1678) );
  NAND2_X2 U49 ( .A1(DATAIN[7]), .A2(n51), .ZN(n1656) );
  NAND2_X2 U50 ( .A1(DATAIN[8]), .A2(n51), .ZN(n1634) );
  NAND2_X2 U51 ( .A1(DATAIN[9]), .A2(n51), .ZN(n1612) );
  NAND2_X2 U52 ( .A1(DATAIN[10]), .A2(n51), .ZN(n1590) );
  NAND2_X2 U53 ( .A1(DATAIN[11]), .A2(n51), .ZN(n1568) );
  NAND2_X2 U54 ( .A1(n2572), .A2(n2585), .ZN(n1890) );
  NAND2_X2 U55 ( .A1(n2577), .A2(n2573), .ZN(n1884) );
  NAND2_X2 U56 ( .A1(n2576), .A2(n2574), .ZN(n1881) );
  NAND2_X2 U57 ( .A1(n2576), .A2(n2573), .ZN(n1882) );
  NAND2_X2 U58 ( .A1(n2575), .A2(n2574), .ZN(n1879) );
  NAND2_X2 U59 ( .A1(n2575), .A2(n2573), .ZN(n1880) );
  NAND2_X2 U60 ( .A1(n2572), .A2(n2574), .ZN(n1877) );
  NAND2_X2 U61 ( .A1(n2572), .A2(n2586), .ZN(n1889) );
  BUF_X1 U62 ( .A(n1919), .Z(n45) );
  NAND2_X2 U63 ( .A1(n2577), .A2(n2597), .ZN(n1920) );
  NAND2_X2 U64 ( .A1(n2598), .A2(n2575), .ZN(n1915) );
  NAND2_X2 U65 ( .A1(n2572), .A2(n2597), .ZN(n1914) );
  NAND2_X2 U66 ( .A1(n2577), .A2(n2592), .ZN(n1907) );
  NAND2_X2 U67 ( .A1(n2591), .A2(n2577), .ZN(n1908) );
  NAND2_X2 U68 ( .A1(n2576), .A2(n2592), .ZN(n1905) );
  NAND2_X2 U69 ( .A1(n2576), .A2(n2591), .ZN(n1906) );
  NAND2_X2 U70 ( .A1(n2591), .A2(n2575), .ZN(n1904) );
  NAND2_X2 U71 ( .A1(n2572), .A2(n2592), .ZN(n1901) );
  NAND2_X2 U72 ( .A1(n2572), .A2(n2591), .ZN(n1902) );
  NAND2_X2 U73 ( .A1(n2577), .A2(n2586), .ZN(n1895) );
  NAND2_X2 U74 ( .A1(n2577), .A2(n2585), .ZN(n1896) );
  NAND2_X2 U75 ( .A1(n2576), .A2(n2586), .ZN(n1893) );
  NAND2_X2 U76 ( .A1(n2576), .A2(n2585), .ZN(n1894) );
  NAND2_X2 U77 ( .A1(n2586), .A2(n2575), .ZN(n1891) );
  NAND2_X2 U78 ( .A1(n2585), .A2(n2575), .ZN(n1892) );
  NAND2_X2 U79 ( .A1(n1842), .A2(n1841), .ZN(n1114) );
  NAND2_X2 U80 ( .A1(n1843), .A2(n1840), .ZN(n1117) );
  NAND2_X2 U81 ( .A1(n1843), .A2(n1841), .ZN(n1116) );
  NAND2_X2 U82 ( .A1(n1844), .A2(n1840), .ZN(n1119) );
  NAND2_X2 U83 ( .A1(n1844), .A2(n1841), .ZN(n1118) );
  NAND2_X2 U84 ( .A1(n1839), .A2(n1852), .ZN(n1125) );
  NAND2_X2 U85 ( .A1(n1839), .A2(n1853), .ZN(n1124) );
  NAND2_X2 U86 ( .A1(n1852), .A2(n1842), .ZN(n1127) );
  NAND2_X2 U87 ( .A1(n1853), .A2(n1842), .ZN(n1126) );
  NAND2_X2 U88 ( .A1(n1843), .A2(n1852), .ZN(n1129) );
  NAND2_X2 U89 ( .A1(n1843), .A2(n1853), .ZN(n1128) );
  NAND2_X2 U90 ( .A1(n1844), .A2(n1852), .ZN(n1131) );
  NAND2_X2 U91 ( .A1(n1844), .A2(n1853), .ZN(n1130) );
  NAND2_X2 U92 ( .A1(n1839), .A2(n1858), .ZN(n1137) );
  NAND2_X2 U93 ( .A1(n1839), .A2(n1859), .ZN(n1136) );
  NAND2_X2 U94 ( .A1(n1858), .A2(n1842), .ZN(n1139) );
  NAND2_X2 U95 ( .A1(n1843), .A2(n1858), .ZN(n1141) );
  NAND2_X2 U96 ( .A1(n1843), .A2(n1859), .ZN(n1140) );
  NAND2_X2 U97 ( .A1(n1858), .A2(n1844), .ZN(n1143) );
  NAND2_X2 U98 ( .A1(n1839), .A2(n1841), .ZN(n1112) );
  NAND2_X2 U99 ( .A1(n1842), .A2(n1840), .ZN(n1115) );
  NAND2_X2 U100 ( .A1(n1839), .A2(n1864), .ZN(n1149) );
  NAND2_X2 U101 ( .A1(n1865), .A2(n1842), .ZN(n1151) );
  NAND2_X2 U102 ( .A1(n1844), .A2(n1859), .ZN(n1142) );
  BUF_X1 U103 ( .A(n1155), .Z(n3) );
  INV_X1 U104 ( .A(ADD_WR[0]), .ZN(n1826) );
  INV_X1 U105 ( .A(ADD_WR[3]), .ZN(n1829) );
  INV_X1 U106 ( .A(ADD_WR[2]), .ZN(n1825) );
  INV_X1 U107 ( .A(ADD_WR[1]), .ZN(n1823) );
  NAND2_X2 U108 ( .A1(n2598), .A2(n2572), .ZN(n1913) );
  NAND2_X2 U109 ( .A1(n1865), .A2(n1839), .ZN(n1148) );
  AND4_X1 U110 ( .A1(n1488), .A2(n1489), .A3(n1490), .A4(n1491), .ZN(n1487) );
  AND4_X1 U111 ( .A1(n1400), .A2(n1401), .A3(n1402), .A4(n1403), .ZN(n1399) );
  AND4_X1 U112 ( .A1(n1356), .A2(n1357), .A3(n1358), .A4(n1359), .ZN(n1355) );
  AND4_X1 U113 ( .A1(n1378), .A2(n1379), .A3(n1380), .A4(n1381), .ZN(n1377) );
  AND4_X1 U114 ( .A1(n1444), .A2(n1445), .A3(n1446), .A4(n1447), .ZN(n1443) );
  AND4_X1 U115 ( .A1(n1422), .A2(n1423), .A3(n1424), .A4(n1425), .ZN(n1421) );
  AND4_X1 U116 ( .A1(n1104), .A2(n1105), .A3(n1106), .A4(n1107), .ZN(n1101) );
  AND4_X1 U117 ( .A1(n1180), .A2(n1181), .A3(n1182), .A4(n1183), .ZN(n1179) );
  AND4_X1 U118 ( .A1(n1312), .A2(n1313), .A3(n1314), .A4(n1315), .ZN(n1311) );
  AND4_X1 U119 ( .A1(n1334), .A2(n1335), .A3(n1336), .A4(n1337), .ZN(n1333) );
  AND4_X1 U120 ( .A1(n1532), .A2(n1533), .A3(n1534), .A4(n1535), .ZN(n1531) );
  AND4_X1 U121 ( .A1(n1554), .A2(n1555), .A3(n1556), .A4(n1557), .ZN(n1553) );
  AND4_X1 U122 ( .A1(n1268), .A2(n1269), .A3(n1270), .A4(n1271), .ZN(n1267) );
  AND4_X1 U123 ( .A1(n1202), .A2(n1203), .A3(n1204), .A4(n1205), .ZN(n1201) );
  AND4_X1 U124 ( .A1(n1510), .A2(n1511), .A3(n1512), .A4(n1513), .ZN(n1509) );
  AND4_X1 U125 ( .A1(n1290), .A2(n1291), .A3(n1292), .A4(n1293), .ZN(n1289) );
  AND4_X1 U126 ( .A1(n1158), .A2(n1159), .A3(n1160), .A4(n1161), .ZN(n1157) );
  AND4_X1 U127 ( .A1(n1224), .A2(n1225), .A3(n1226), .A4(n1227), .ZN(n1223) );
  AND4_X1 U128 ( .A1(n1466), .A2(n1467), .A3(n1468), .A4(n1469), .ZN(n1465) );
  AND4_X1 U129 ( .A1(n2237), .A2(n2238), .A3(n2239), .A4(n2240), .ZN(n2236) );
  AND4_X1 U130 ( .A1(n2300), .A2(n2301), .A3(n2302), .A4(n2303), .ZN(n2299) );
  AND4_X1 U131 ( .A1(n1985), .A2(n1986), .A3(n1987), .A4(n1988), .ZN(n1984) );
  AND4_X1 U132 ( .A1(n2153), .A2(n2154), .A3(n2155), .A4(n2156), .ZN(n2152) );
  AND4_X1 U133 ( .A1(n1964), .A2(n1965), .A3(n1966), .A4(n1967), .ZN(n1963) );
  AND4_X1 U134 ( .A1(n1869), .A2(n1870), .A3(n1871), .A4(n1872), .ZN(n1866) );
  AND4_X1 U135 ( .A1(n2258), .A2(n2259), .A3(n2260), .A4(n2261), .ZN(n2257) );
  AND4_X1 U136 ( .A1(n2279), .A2(n2280), .A3(n2281), .A4(n2282), .ZN(n2278) );
  AND4_X1 U137 ( .A1(n2069), .A2(n2070), .A3(n2071), .A4(n2072), .ZN(n2068) );
  AND4_X1 U138 ( .A1(n2132), .A2(n2133), .A3(n2134), .A4(n2135), .ZN(n2131) );
  AND4_X1 U139 ( .A1(n2048), .A2(n2049), .A3(n2050), .A4(n2051), .ZN(n2047) );
  AND4_X1 U140 ( .A1(n2111), .A2(n2112), .A3(n2113), .A4(n2114), .ZN(n2110) );
  AND4_X1 U141 ( .A1(n2216), .A2(n2217), .A3(n2218), .A4(n2219), .ZN(n2215) );
  AND4_X1 U142 ( .A1(n2174), .A2(n2175), .A3(n2176), .A4(n2177), .ZN(n2173) );
  AND4_X1 U143 ( .A1(n2027), .A2(n2028), .A3(n2029), .A4(n2030), .ZN(n2026) );
  AND4_X1 U144 ( .A1(n2195), .A2(n2196), .A3(n2197), .A4(n2198), .ZN(n2194) );
  AND4_X1 U145 ( .A1(n1922), .A2(n1923), .A3(n1924), .A4(n1925), .ZN(n1921) );
  AND4_X1 U146 ( .A1(n2090), .A2(n2091), .A3(n2092), .A4(n2093), .ZN(n2089) );
  AND4_X1 U147 ( .A1(n1943), .A2(n1944), .A3(n1945), .A4(n1946), .ZN(n1942) );
  AND4_X1 U148 ( .A1(n1664), .A2(n1665), .A3(n1666), .A4(n1667), .ZN(n1663) );
  AND4_X1 U149 ( .A1(n1797), .A2(n1798), .A3(n1799), .A4(n1800), .ZN(n1796) );
  INV_X1 U150 ( .A(n1773), .ZN(n1767) );
  AND4_X1 U151 ( .A1(n1686), .A2(n1687), .A3(n1688), .A4(n1689), .ZN(n1685) );
  AND4_X1 U152 ( .A1(n1708), .A2(n1709), .A3(n1710), .A4(n1711), .ZN(n1707) );
  AND4_X1 U153 ( .A1(n1831), .A2(n1832), .A3(n1833), .A4(n1834), .ZN(n1818) );
  AND4_X1 U154 ( .A1(n1730), .A2(n1731), .A3(n1732), .A4(n1733), .ZN(n1729) );
  AND4_X1 U155 ( .A1(n1775), .A2(n1776), .A3(n1777), .A4(n1778), .ZN(n1774) );
  AND4_X1 U156 ( .A1(n2532), .A2(n2533), .A3(n2534), .A4(n2535), .ZN(n2531) );
  INV_X1 U157 ( .A(n2509), .ZN(n2503) );
  AND4_X1 U158 ( .A1(n2426), .A2(n2427), .A3(n2428), .A4(n2429), .ZN(n2425) );
  AND4_X1 U159 ( .A1(n2564), .A2(n2565), .A3(n2566), .A4(n2567), .ZN(n2552) );
  AND4_X1 U160 ( .A1(n2447), .A2(n2448), .A3(n2449), .A4(n2450), .ZN(n2446) );
  AND4_X1 U161 ( .A1(n2405), .A2(n2406), .A3(n2407), .A4(n2408), .ZN(n2404) );
  AND4_X1 U162 ( .A1(n2511), .A2(n2512), .A3(n2513), .A4(n2514), .ZN(n2510) );
  AND4_X1 U163 ( .A1(n2468), .A2(n2469), .A3(n2470), .A4(n2471), .ZN(n2467) );
  AND4_X1 U164 ( .A1(n1246), .A2(n1247), .A3(n1248), .A4(n1249), .ZN(n1245) );
  AND4_X1 U165 ( .A1(n1598), .A2(n1599), .A3(n1600), .A4(n1601), .ZN(n1597) );
  AND4_X1 U166 ( .A1(n1620), .A2(n1621), .A3(n1622), .A4(n1623), .ZN(n1619) );
  AND4_X1 U167 ( .A1(n1576), .A2(n1577), .A3(n1578), .A4(n1579), .ZN(n1575) );
  AND4_X1 U168 ( .A1(n1642), .A2(n1643), .A3(n1644), .A4(n1645), .ZN(n1641) );
  INV_X1 U169 ( .A(ADD_RD2[4]), .ZN(n1828) );
  INV_X1 U170 ( .A(ADD_RD2[3]), .ZN(n1845) );
  AND2_X1 U171 ( .A1(ADD_RD2[1]), .A2(ADD_RD2[2]), .ZN(n1839) );
  AND2_X1 U172 ( .A1(n1822), .A2(ADD_RD2[2]), .ZN(n1842) );
  INV_X1 U173 ( .A(ADD_RD2[1]), .ZN(n1822) );
  INV_X1 U174 ( .A(ADD_RD2[0]), .ZN(n1846) );
  AND4_X1 U175 ( .A1(n2363), .A2(n2364), .A3(n2365), .A4(n2366), .ZN(n2362) );
  AND4_X1 U176 ( .A1(n2384), .A2(n2385), .A3(n2386), .A4(n2387), .ZN(n2383) );
  AND4_X1 U177 ( .A1(n2006), .A2(n2007), .A3(n2008), .A4(n2009), .ZN(n2005) );
  AND4_X1 U178 ( .A1(n2321), .A2(n2322), .A3(n2323), .A4(n2324), .ZN(n2320) );
  INV_X1 U179 ( .A(n2563), .ZN(n2560) );
  AND4_X1 U180 ( .A1(n2342), .A2(n2343), .A3(n2344), .A4(n2345), .ZN(n2341) );
  INV_X1 U181 ( .A(ADD_RD1[4]), .ZN(n2558) );
  INV_X1 U182 ( .A(ADD_RD1[3]), .ZN(n2578) );
  AND2_X1 U183 ( .A1(ADD_RD1[1]), .A2(ADD_RD1[2]), .ZN(n2572) );
  AND2_X1 U184 ( .A1(n2555), .A2(ADD_RD1[2]), .ZN(n2575) );
  INV_X1 U185 ( .A(ADD_RD1[1]), .ZN(n2555) );
  INV_X1 U186 ( .A(ADD_RD1[0]), .ZN(n2579) );
  OR2_X1 U187 ( .A1(N4487), .A2(ENABLE), .ZN(N4615) );
  OR3_X1 U188 ( .A1(n1829), .A2(n2562), .A3(ADD_WR[4]), .ZN(n2607) );
  NOR2_X1 U189 ( .A1(ADD_RD2[0]), .A2(n1847), .ZN(n1841) );
  NOR2_X1 U190 ( .A1(ADD_RD2[2]), .A2(n1822), .ZN(n1843) );
  NOR2_X1 U191 ( .A1(ADD_RD2[1]), .A2(ADD_RD2[2]), .ZN(n1844) );
  AOI21_X1 U192 ( .B1(n2560), .B2(n2561), .A(n2562), .ZN(n1819) );
  NOR2_X1 U193 ( .A1(ADD_RD1[0]), .A2(n2580), .ZN(n2574) );
  NOR2_X1 U194 ( .A1(ADD_RD1[2]), .A2(n2555), .ZN(n2576) );
  NOR2_X1 U195 ( .A1(ADD_RD1[1]), .A2(ADD_RD1[2]), .ZN(n2577) );
  NAND2_X1 U196 ( .A1(n2577), .A2(n2574), .ZN(n1883) );
  OAI22_X1 U197 ( .A1(n1101), .A2(n1102), .B1(n1103), .B2(n1094), .ZN(N4616)
         );
  NOR4_X1 U198 ( .A1(n1108), .A2(n1109), .A3(n1110), .A4(n1111), .ZN(n1107) );
  OAI22_X1 U199 ( .A1(n199), .A2(n1112), .B1(n1089), .B2(n1113), .ZN(n1111) );
  OAI22_X1 U200 ( .A1(n263), .A2(n1114), .B1(n231), .B2(n1115), .ZN(n1110) );
  OAI22_X1 U201 ( .A1(n327), .A2(n1116), .B1(n295), .B2(n1117), .ZN(n1109) );
  OAI22_X1 U202 ( .A1(n391), .A2(n1118), .B1(n359), .B2(n1119), .ZN(n1108) );
  NOR4_X1 U203 ( .A1(n1120), .A2(n1121), .A3(n1122), .A4(n1123), .ZN(n1106) );
  OAI22_X1 U204 ( .A1(n456), .A2(n1124), .B1(n423), .B2(n1125), .ZN(n1123) );
  OAI22_X1 U205 ( .A1(n524), .A2(n1126), .B1(n490), .B2(n1127), .ZN(n1122) );
  OAI22_X1 U206 ( .A1(n591), .A2(n1128), .B1(n557), .B2(n1129), .ZN(n1121) );
  OAI22_X1 U207 ( .A1(n658), .A2(n1130), .B1(n624), .B2(n1131), .ZN(n1120) );
  NOR4_X1 U208 ( .A1(n1132), .A2(n1133), .A3(n1134), .A4(n1135), .ZN(n1105) );
  OAI22_X1 U209 ( .A1(n725), .A2(n1136), .B1(n692), .B2(n1137), .ZN(n1135) );
  OAI22_X1 U210 ( .A1(n792), .A2(n1138), .B1(n759), .B2(n1139), .ZN(n1134) );
  OAI22_X1 U211 ( .A1(n860), .A2(n1140), .B1(n826), .B2(n1141), .ZN(n1133) );
  OAI22_X1 U212 ( .A1(n927), .A2(n1142), .B1(n893), .B2(n1143), .ZN(n1132) );
  NOR4_X1 U213 ( .A1(n1144), .A2(n1145), .A3(n1146), .A4(n1147), .ZN(n1104) );
  OAI22_X1 U214 ( .A1(n994), .A2(n1148), .B1(n960), .B2(n1149), .ZN(n1147) );
  OAI22_X1 U215 ( .A1(n1061), .A2(n1151), .B1(n1028), .B2(n1152), .ZN(n1146)
         );
  OAI22_X1 U216 ( .A1(n106), .A2(n1), .B1(n1096), .B2(n1154), .ZN(n1145) );
  OAI22_X1 U217 ( .A1(n177), .A2(n1155), .B1(n141), .B2(n1156), .ZN(n1144) );
  OAI22_X1 U218 ( .A1(n1157), .A2(n1102), .B1(n1103), .B2(n1150), .ZN(N4614)
         );
  NOR4_X1 U219 ( .A1(n1162), .A2(n1163), .A3(n1164), .A4(n1165), .ZN(n1161) );
  OAI22_X1 U220 ( .A1(n198), .A2(n1112), .B1(n1068), .B2(n1113), .ZN(n1165) );
  OAI22_X1 U221 ( .A1(n262), .A2(n1114), .B1(n230), .B2(n1115), .ZN(n1164) );
  OAI22_X1 U222 ( .A1(n326), .A2(n1116), .B1(n294), .B2(n1117), .ZN(n1163) );
  OAI22_X1 U223 ( .A1(n390), .A2(n1118), .B1(n358), .B2(n1119), .ZN(n1162) );
  NOR4_X1 U224 ( .A1(n1166), .A2(n1167), .A3(n1168), .A4(n1169), .ZN(n1160) );
  OAI22_X1 U225 ( .A1(n455), .A2(n1124), .B1(n422), .B2(n1125), .ZN(n1169) );
  OAI22_X1 U226 ( .A1(n523), .A2(n1126), .B1(n489), .B2(n1127), .ZN(n1168) );
  OAI22_X1 U227 ( .A1(n590), .A2(n1128), .B1(n556), .B2(n1129), .ZN(n1167) );
  OAI22_X1 U228 ( .A1(n657), .A2(n1130), .B1(n623), .B2(n1131), .ZN(n1166) );
  NOR4_X1 U229 ( .A1(n1170), .A2(n1171), .A3(n1173), .A4(n1174), .ZN(n1159) );
  OAI22_X1 U230 ( .A1(n724), .A2(n1136), .B1(n691), .B2(n1137), .ZN(n1174) );
  OAI22_X1 U231 ( .A1(n791), .A2(n1138), .B1(n758), .B2(n1139), .ZN(n1173) );
  OAI22_X1 U232 ( .A1(n859), .A2(n1140), .B1(n825), .B2(n1141), .ZN(n1171) );
  OAI22_X1 U233 ( .A1(n926), .A2(n1142), .B1(n892), .B2(n1143), .ZN(n1170) );
  NOR4_X1 U234 ( .A1(n1175), .A2(n1176), .A3(n1177), .A4(n1178), .ZN(n1158) );
  OAI22_X1 U235 ( .A1(n993), .A2(n1148), .B1(n959), .B2(n1149), .ZN(n1178) );
  OAI22_X1 U236 ( .A1(n1060), .A2(n1151), .B1(n1027), .B2(n1152), .ZN(n1177)
         );
  OAI22_X1 U237 ( .A1(n105), .A2(n1153), .B1(n1095), .B2(n1154), .ZN(n1176) );
  OAI22_X1 U238 ( .A1(n176), .A2(n3), .B1(n140), .B2(n37), .ZN(n1175) );
  OAI22_X1 U239 ( .A1(n1179), .A2(n1102), .B1(n1103), .B2(n1172), .ZN(N4612)
         );
  NOR4_X1 U240 ( .A1(n1184), .A2(n1185), .A3(n1186), .A4(n1187), .ZN(n1183) );
  OAI22_X1 U241 ( .A1(n197), .A2(n1112), .B1(n1047), .B2(n1113), .ZN(n1187) );
  OAI22_X1 U242 ( .A1(n261), .A2(n1114), .B1(n229), .B2(n1115), .ZN(n1186) );
  OAI22_X1 U243 ( .A1(n325), .A2(n1116), .B1(n293), .B2(n1117), .ZN(n1185) );
  OAI22_X1 U244 ( .A1(n389), .A2(n1118), .B1(n357), .B2(n1119), .ZN(n1184) );
  NOR4_X1 U245 ( .A1(n1188), .A2(n1189), .A3(n1190), .A4(n1191), .ZN(n1182) );
  OAI22_X1 U246 ( .A1(n454), .A2(n1124), .B1(n421), .B2(n1125), .ZN(n1191) );
  OAI22_X1 U247 ( .A1(n521), .A2(n1126), .B1(n488), .B2(n1127), .ZN(n1190) );
  OAI22_X1 U248 ( .A1(n589), .A2(n1128), .B1(n555), .B2(n1129), .ZN(n1189) );
  OAI22_X1 U249 ( .A1(n656), .A2(n1130), .B1(n622), .B2(n1131), .ZN(n1188) );
  NOR4_X1 U250 ( .A1(n1192), .A2(n1193), .A3(n1195), .A4(n1196), .ZN(n1181) );
  OAI22_X1 U251 ( .A1(n723), .A2(n1136), .B1(n689), .B2(n1137), .ZN(n1196) );
  OAI22_X1 U252 ( .A1(n790), .A2(n1138), .B1(n757), .B2(n1139), .ZN(n1195) );
  OAI22_X1 U253 ( .A1(n857), .A2(n1140), .B1(n824), .B2(n1141), .ZN(n1193) );
  OAI22_X1 U254 ( .A1(n925), .A2(n1142), .B1(n891), .B2(n1143), .ZN(n1192) );
  NOR4_X1 U255 ( .A1(n1197), .A2(n1198), .A3(n1199), .A4(n1200), .ZN(n1180) );
  OAI22_X1 U256 ( .A1(n992), .A2(n1148), .B1(n958), .B2(n1149), .ZN(n1200) );
  OAI22_X1 U257 ( .A1(n1059), .A2(n1151), .B1(n1025), .B2(n1152), .ZN(n1199)
         );
  OAI22_X1 U258 ( .A1(n104), .A2(n1153), .B1(n1093), .B2(n1154), .ZN(n1198) );
  OAI22_X1 U259 ( .A1(n174), .A2(n3), .B1(n139), .B2(n37), .ZN(n1197) );
  OAI22_X1 U260 ( .A1(n1201), .A2(n1102), .B1(n1103), .B2(n1194), .ZN(N4610)
         );
  NOR4_X1 U261 ( .A1(n1206), .A2(n1207), .A3(n1208), .A4(n1209), .ZN(n1205) );
  OAI22_X1 U262 ( .A1(n196), .A2(n1112), .B1(n1026), .B2(n1113), .ZN(n1209) );
  OAI22_X1 U263 ( .A1(n260), .A2(n1114), .B1(n228), .B2(n1115), .ZN(n1208) );
  OAI22_X1 U264 ( .A1(n324), .A2(n1116), .B1(n292), .B2(n1117), .ZN(n1207) );
  OAI22_X1 U265 ( .A1(n388), .A2(n1118), .B1(n356), .B2(n1119), .ZN(n1206) );
  NOR4_X1 U266 ( .A1(n1210), .A2(n1211), .A3(n1212), .A4(n1213), .ZN(n1204) );
  OAI22_X1 U267 ( .A1(n453), .A2(n1124), .B1(n420), .B2(n1125), .ZN(n1213) );
  OAI22_X1 U268 ( .A1(n520), .A2(n1126), .B1(n487), .B2(n1127), .ZN(n1212) );
  OAI22_X1 U269 ( .A1(n588), .A2(n1128), .B1(n554), .B2(n1129), .ZN(n1211) );
  OAI22_X1 U270 ( .A1(n655), .A2(n1130), .B1(n621), .B2(n1131), .ZN(n1210) );
  NOR4_X1 U271 ( .A1(n1214), .A2(n1215), .A3(n1217), .A4(n1218), .ZN(n1203) );
  OAI22_X1 U272 ( .A1(n722), .A2(n1136), .B1(n688), .B2(n1137), .ZN(n1218) );
  OAI22_X1 U273 ( .A1(n789), .A2(n1138), .B1(n756), .B2(n1139), .ZN(n1217) );
  OAI22_X1 U274 ( .A1(n856), .A2(n1140), .B1(n823), .B2(n1141), .ZN(n1215) );
  OAI22_X1 U275 ( .A1(n924), .A2(n1142), .B1(n890), .B2(n1143), .ZN(n1214) );
  NOR4_X1 U276 ( .A1(n1219), .A2(n1220), .A3(n1221), .A4(n1222), .ZN(n1202) );
  OAI22_X1 U277 ( .A1(n991), .A2(n1148), .B1(n957), .B2(n1149), .ZN(n1222) );
  OAI22_X1 U278 ( .A1(n1058), .A2(n1151), .B1(n1024), .B2(n1152), .ZN(n1221)
         );
  OAI22_X1 U279 ( .A1(n103), .A2(n1153), .B1(n1092), .B2(n2), .ZN(n1220) );
  OAI22_X1 U280 ( .A1(n173), .A2(n3), .B1(n138), .B2(n37), .ZN(n1219) );
  OAI22_X1 U281 ( .A1(n1223), .A2(n1102), .B1(n1103), .B2(n1216), .ZN(N4608)
         );
  NOR4_X1 U282 ( .A1(n1228), .A2(n1229), .A3(n1230), .A4(n1231), .ZN(n1227) );
  OAI22_X1 U283 ( .A1(n195), .A2(n1112), .B1(n1005), .B2(n1113), .ZN(n1231) );
  OAI22_X1 U284 ( .A1(n259), .A2(n1114), .B1(n227), .B2(n1115), .ZN(n1230) );
  OAI22_X1 U285 ( .A1(n323), .A2(n1116), .B1(n291), .B2(n1117), .ZN(n1229) );
  OAI22_X1 U286 ( .A1(n387), .A2(n1118), .B1(n355), .B2(n1119), .ZN(n1228) );
  NOR4_X1 U287 ( .A1(n1232), .A2(n1233), .A3(n1234), .A4(n1235), .ZN(n1226) );
  OAI22_X1 U288 ( .A1(n452), .A2(n1124), .B1(n419), .B2(n1125), .ZN(n1235) );
  OAI22_X1 U289 ( .A1(n519), .A2(n1126), .B1(n486), .B2(n1127), .ZN(n1234) );
  OAI22_X1 U290 ( .A1(n587), .A2(n1128), .B1(n553), .B2(n1129), .ZN(n1233) );
  OAI22_X1 U291 ( .A1(n654), .A2(n1130), .B1(n620), .B2(n1131), .ZN(n1232) );
  NOR4_X1 U292 ( .A1(n1236), .A2(n1237), .A3(n1239), .A4(n1240), .ZN(n1225) );
  OAI22_X1 U293 ( .A1(n721), .A2(n1136), .B1(n687), .B2(n1137), .ZN(n1240) );
  OAI22_X1 U294 ( .A1(n788), .A2(n1138), .B1(n755), .B2(n1139), .ZN(n1239) );
  OAI22_X1 U295 ( .A1(n855), .A2(n1140), .B1(n822), .B2(n1141), .ZN(n1237) );
  OAI22_X1 U296 ( .A1(n923), .A2(n1142), .B1(n889), .B2(n1143), .ZN(n1236) );
  NOR4_X1 U297 ( .A1(n1241), .A2(n1242), .A3(n1243), .A4(n1244), .ZN(n1224) );
  OAI22_X1 U298 ( .A1(n990), .A2(n1148), .B1(n956), .B2(n1149), .ZN(n1244) );
  OAI22_X1 U299 ( .A1(n1057), .A2(n1151), .B1(n1023), .B2(n1152), .ZN(n1243)
         );
  OAI22_X1 U300 ( .A1(n102), .A2(n1153), .B1(n1091), .B2(n2), .ZN(n1242) );
  OAI22_X1 U301 ( .A1(n172), .A2(n3), .B1(n137), .B2(n37), .ZN(n1241) );
  OAI22_X1 U302 ( .A1(n1245), .A2(n1102), .B1(n1103), .B2(n1238), .ZN(N4606)
         );
  NOR4_X1 U303 ( .A1(n1250), .A2(n1251), .A3(n1252), .A4(n1253), .ZN(n1249) );
  OAI22_X1 U304 ( .A1(n194), .A2(n1112), .B1(n984), .B2(n1113), .ZN(n1253) );
  OAI22_X1 U305 ( .A1(n258), .A2(n1114), .B1(n226), .B2(n1115), .ZN(n1252) );
  OAI22_X1 U306 ( .A1(n322), .A2(n1116), .B1(n290), .B2(n1117), .ZN(n1251) );
  OAI22_X1 U307 ( .A1(n386), .A2(n1118), .B1(n354), .B2(n1119), .ZN(n1250) );
  NOR4_X1 U308 ( .A1(n1254), .A2(n1255), .A3(n1256), .A4(n1257), .ZN(n1248) );
  OAI22_X1 U309 ( .A1(n451), .A2(n1124), .B1(n418), .B2(n1125), .ZN(n1257) );
  OAI22_X1 U310 ( .A1(n518), .A2(n1126), .B1(n485), .B2(n1127), .ZN(n1256) );
  OAI22_X1 U311 ( .A1(n586), .A2(n1128), .B1(n552), .B2(n1129), .ZN(n1255) );
  OAI22_X1 U312 ( .A1(n653), .A2(n1130), .B1(n619), .B2(n1131), .ZN(n1254) );
  NOR4_X1 U313 ( .A1(n1258), .A2(n1259), .A3(n1261), .A4(n1262), .ZN(n1247) );
  OAI22_X1 U314 ( .A1(n720), .A2(n1136), .B1(n686), .B2(n1137), .ZN(n1262) );
  OAI22_X1 U315 ( .A1(n787), .A2(n1138), .B1(n754), .B2(n1139), .ZN(n1261) );
  OAI22_X1 U316 ( .A1(n854), .A2(n1140), .B1(n821), .B2(n1141), .ZN(n1259) );
  OAI22_X1 U317 ( .A1(n922), .A2(n1142), .B1(n888), .B2(n1143), .ZN(n1258) );
  NOR4_X1 U318 ( .A1(n1263), .A2(n1264), .A3(n1265), .A4(n1266), .ZN(n1246) );
  OAI22_X1 U319 ( .A1(n989), .A2(n1148), .B1(n955), .B2(n1149), .ZN(n1266) );
  OAI22_X1 U320 ( .A1(n1056), .A2(n1151), .B1(n1022), .B2(n1152), .ZN(n1265)
         );
  OAI22_X1 U321 ( .A1(n101), .A2(n1153), .B1(n1090), .B2(n1154), .ZN(n1264) );
  OAI22_X1 U322 ( .A1(n171), .A2(n3), .B1(n136), .B2(n37), .ZN(n1263) );
  OAI22_X1 U323 ( .A1(n1267), .A2(n1102), .B1(n1103), .B2(n1260), .ZN(N4604)
         );
  NOR4_X1 U324 ( .A1(n1272), .A2(n1273), .A3(n1274), .A4(n1275), .ZN(n1271) );
  OAI22_X1 U325 ( .A1(n193), .A2(n1112), .B1(n963), .B2(n1113), .ZN(n1275) );
  OAI22_X1 U326 ( .A1(n257), .A2(n1114), .B1(n225), .B2(n1115), .ZN(n1274) );
  OAI22_X1 U327 ( .A1(n321), .A2(n1116), .B1(n289), .B2(n1117), .ZN(n1273) );
  OAI22_X1 U328 ( .A1(n385), .A2(n1118), .B1(n353), .B2(n1119), .ZN(n1272) );
  NOR4_X1 U329 ( .A1(n1276), .A2(n1277), .A3(n1278), .A4(n1279), .ZN(n1270) );
  OAI22_X1 U330 ( .A1(n450), .A2(n1124), .B1(n417), .B2(n1125), .ZN(n1279) );
  OAI22_X1 U331 ( .A1(n517), .A2(n1126), .B1(n484), .B2(n1127), .ZN(n1278) );
  OAI22_X1 U332 ( .A1(n584), .A2(n1128), .B1(n551), .B2(n1129), .ZN(n1277) );
  OAI22_X1 U333 ( .A1(n652), .A2(n1130), .B1(n618), .B2(n1131), .ZN(n1276) );
  NOR4_X1 U334 ( .A1(n1280), .A2(n1281), .A3(n1283), .A4(n1284), .ZN(n1269) );
  OAI22_X1 U335 ( .A1(n719), .A2(n1136), .B1(n685), .B2(n1137), .ZN(n1284) );
  OAI22_X1 U336 ( .A1(n786), .A2(n1138), .B1(n752), .B2(n1139), .ZN(n1283) );
  OAI22_X1 U337 ( .A1(n853), .A2(n1140), .B1(n820), .B2(n1141), .ZN(n1281) );
  OAI22_X1 U338 ( .A1(n920), .A2(n1142), .B1(n887), .B2(n1143), .ZN(n1280) );
  NOR4_X1 U339 ( .A1(n1285), .A2(n1286), .A3(n1287), .A4(n1288), .ZN(n1268) );
  OAI22_X1 U340 ( .A1(n988), .A2(n1148), .B1(n954), .B2(n1149), .ZN(n1288) );
  OAI22_X1 U341 ( .A1(n1055), .A2(n1151), .B1(n1021), .B2(n1152), .ZN(n1287)
         );
  OAI22_X1 U342 ( .A1(n100), .A2(n1153), .B1(n1088), .B2(n2), .ZN(n1286) );
  OAI22_X1 U343 ( .A1(n170), .A2(n3), .B1(n135), .B2(n37), .ZN(n1285) );
  OAI22_X1 U344 ( .A1(n1289), .A2(n1102), .B1(n1103), .B2(n1282), .ZN(N4602)
         );
  NOR4_X1 U345 ( .A1(n1294), .A2(n1295), .A3(n1296), .A4(n1297), .ZN(n1293) );
  OAI22_X1 U346 ( .A1(n192), .A2(n1112), .B1(n942), .B2(n1113), .ZN(n1297) );
  OAI22_X1 U347 ( .A1(n256), .A2(n1114), .B1(n224), .B2(n1115), .ZN(n1296) );
  OAI22_X1 U348 ( .A1(n320), .A2(n1116), .B1(n288), .B2(n1117), .ZN(n1295) );
  OAI22_X1 U349 ( .A1(n384), .A2(n1118), .B1(n352), .B2(n1119), .ZN(n1294) );
  NOR4_X1 U350 ( .A1(n1298), .A2(n1299), .A3(n1300), .A4(n1301), .ZN(n1292) );
  OAI22_X1 U351 ( .A1(n449), .A2(n1124), .B1(n416), .B2(n1125), .ZN(n1301) );
  OAI22_X1 U352 ( .A1(n516), .A2(n1126), .B1(n483), .B2(n1127), .ZN(n1300) );
  OAI22_X1 U353 ( .A1(n583), .A2(n1128), .B1(n550), .B2(n1129), .ZN(n1299) );
  OAI22_X1 U354 ( .A1(n651), .A2(n1130), .B1(n617), .B2(n1131), .ZN(n1298) );
  NOR4_X1 U355 ( .A1(n1302), .A2(n1303), .A3(n1305), .A4(n1306), .ZN(n1291) );
  OAI22_X1 U356 ( .A1(n718), .A2(n1136), .B1(n684), .B2(n1137), .ZN(n1306) );
  OAI22_X1 U357 ( .A1(n785), .A2(n1138), .B1(n751), .B2(n1139), .ZN(n1305) );
  OAI22_X1 U358 ( .A1(n852), .A2(n1140), .B1(n819), .B2(n1141), .ZN(n1303) );
  OAI22_X1 U359 ( .A1(n919), .A2(n1142), .B1(n886), .B2(n1143), .ZN(n1302) );
  NOR4_X1 U360 ( .A1(n1307), .A2(n1308), .A3(n1309), .A4(n1310), .ZN(n1290) );
  OAI22_X1 U361 ( .A1(n987), .A2(n1148), .B1(n953), .B2(n1149), .ZN(n1310) );
  OAI22_X1 U362 ( .A1(n1054), .A2(n1151), .B1(n1020), .B2(n1152), .ZN(n1309)
         );
  OAI22_X1 U363 ( .A1(n99), .A2(n1153), .B1(n1087), .B2(n1154), .ZN(n1308) );
  OAI22_X1 U364 ( .A1(n169), .A2(n3), .B1(n134), .B2(n37), .ZN(n1307) );
  OAI22_X1 U365 ( .A1(n1311), .A2(n1102), .B1(n1103), .B2(n1304), .ZN(N4600)
         );
  NOR4_X1 U366 ( .A1(n1316), .A2(n1317), .A3(n1318), .A4(n1319), .ZN(n1315) );
  OAI22_X1 U367 ( .A1(n191), .A2(n1112), .B1(n921), .B2(n1113), .ZN(n1319) );
  OAI22_X1 U368 ( .A1(n255), .A2(n1114), .B1(n223), .B2(n1115), .ZN(n1318) );
  OAI22_X1 U369 ( .A1(n319), .A2(n1116), .B1(n287), .B2(n1117), .ZN(n1317) );
  OAI22_X1 U370 ( .A1(n383), .A2(n1118), .B1(n351), .B2(n1119), .ZN(n1316) );
  NOR4_X1 U371 ( .A1(n1320), .A2(n1321), .A3(n1322), .A4(n1323), .ZN(n1314) );
  OAI22_X1 U372 ( .A1(n448), .A2(n1124), .B1(n415), .B2(n1125), .ZN(n1323) );
  OAI22_X1 U373 ( .A1(n515), .A2(n1126), .B1(n482), .B2(n1127), .ZN(n1322) );
  OAI22_X1 U374 ( .A1(n582), .A2(n1128), .B1(n549), .B2(n1129), .ZN(n1321) );
  OAI22_X1 U375 ( .A1(n650), .A2(n1130), .B1(n616), .B2(n1131), .ZN(n1320) );
  NOR4_X1 U376 ( .A1(n1324), .A2(n1325), .A3(n1327), .A4(n1328), .ZN(n1313) );
  OAI22_X1 U377 ( .A1(n717), .A2(n1136), .B1(n683), .B2(n1137), .ZN(n1328) );
  OAI22_X1 U378 ( .A1(n784), .A2(n1138), .B1(n750), .B2(n1139), .ZN(n1327) );
  OAI22_X1 U379 ( .A1(n851), .A2(n1140), .B1(n818), .B2(n1141), .ZN(n1325) );
  OAI22_X1 U380 ( .A1(n918), .A2(n1142), .B1(n885), .B2(n1143), .ZN(n1324) );
  NOR4_X1 U381 ( .A1(n1329), .A2(n1330), .A3(n1331), .A4(n1332), .ZN(n1312) );
  OAI22_X1 U382 ( .A1(n986), .A2(n1148), .B1(n952), .B2(n1149), .ZN(n1332) );
  OAI22_X1 U383 ( .A1(n1053), .A2(n1151), .B1(n1019), .B2(n1152), .ZN(n1331)
         );
  OAI22_X1 U384 ( .A1(n95), .A2(n1153), .B1(n1086), .B2(n2), .ZN(n1330) );
  OAI22_X1 U385 ( .A1(n168), .A2(n3), .B1(n133), .B2(n37), .ZN(n1329) );
  OAI22_X1 U386 ( .A1(n1333), .A2(n1102), .B1(n1103), .B2(n1326), .ZN(N4598)
         );
  NOR4_X1 U387 ( .A1(n1338), .A2(n1339), .A3(n1340), .A4(n1341), .ZN(n1337) );
  OAI22_X1 U388 ( .A1(n190), .A2(n1112), .B1(n900), .B2(n1113), .ZN(n1341) );
  OAI22_X1 U389 ( .A1(n254), .A2(n1114), .B1(n222), .B2(n1115), .ZN(n1340) );
  OAI22_X1 U390 ( .A1(n318), .A2(n1116), .B1(n286), .B2(n1117), .ZN(n1339) );
  OAI22_X1 U391 ( .A1(n382), .A2(n1118), .B1(n350), .B2(n1119), .ZN(n1338) );
  NOR4_X1 U392 ( .A1(n1342), .A2(n1343), .A3(n1344), .A4(n1345), .ZN(n1336) );
  OAI22_X1 U393 ( .A1(n447), .A2(n1124), .B1(n414), .B2(n1125), .ZN(n1345) );
  OAI22_X1 U394 ( .A1(n514), .A2(n1126), .B1(n481), .B2(n1127), .ZN(n1344) );
  OAI22_X1 U395 ( .A1(n581), .A2(n1128), .B1(n548), .B2(n1129), .ZN(n1343) );
  OAI22_X1 U396 ( .A1(n649), .A2(n1130), .B1(n615), .B2(n1131), .ZN(n1342) );
  NOR4_X1 U397 ( .A1(n1346), .A2(n1347), .A3(n1349), .A4(n1350), .ZN(n1335) );
  OAI22_X1 U398 ( .A1(n716), .A2(n1136), .B1(n682), .B2(n1137), .ZN(n1350) );
  OAI22_X1 U399 ( .A1(n783), .A2(n1138), .B1(n749), .B2(n1139), .ZN(n1349) );
  OAI22_X1 U400 ( .A1(n850), .A2(n1140), .B1(n817), .B2(n1141), .ZN(n1347) );
  OAI22_X1 U401 ( .A1(n917), .A2(n1142), .B1(n884), .B2(n1143), .ZN(n1346) );
  NOR4_X1 U402 ( .A1(n1351), .A2(n1352), .A3(n1353), .A4(n1354), .ZN(n1334) );
  OAI22_X1 U403 ( .A1(n985), .A2(n1148), .B1(n951), .B2(n1149), .ZN(n1354) );
  OAI22_X1 U404 ( .A1(n1052), .A2(n1151), .B1(n1018), .B2(n1152), .ZN(n1353)
         );
  OAI22_X1 U405 ( .A1(n93), .A2(n1153), .B1(n1085), .B2(n2), .ZN(n1352) );
  OAI22_X1 U406 ( .A1(n167), .A2(n3), .B1(n132), .B2(n37), .ZN(n1351) );
  OAI22_X1 U407 ( .A1(n1355), .A2(n1102), .B1(n1103), .B2(n1348), .ZN(N4596)
         );
  NOR4_X1 U408 ( .A1(n1360), .A2(n1361), .A3(n1362), .A4(n1363), .ZN(n1359) );
  OAI22_X1 U409 ( .A1(n189), .A2(n1112), .B1(n879), .B2(n1113), .ZN(n1363) );
  OAI22_X1 U410 ( .A1(n253), .A2(n1114), .B1(n221), .B2(n1115), .ZN(n1362) );
  OAI22_X1 U411 ( .A1(n317), .A2(n1116), .B1(n285), .B2(n1117), .ZN(n1361) );
  OAI22_X1 U412 ( .A1(n381), .A2(n1118), .B1(n349), .B2(n1119), .ZN(n1360) );
  NOR4_X1 U413 ( .A1(n1364), .A2(n1365), .A3(n1366), .A4(n1367), .ZN(n1358) );
  OAI22_X1 U414 ( .A1(n446), .A2(n1124), .B1(n413), .B2(n1125), .ZN(n1367) );
  OAI22_X1 U415 ( .A1(n513), .A2(n1126), .B1(n479), .B2(n1127), .ZN(n1366) );
  OAI22_X1 U416 ( .A1(n580), .A2(n1128), .B1(n547), .B2(n1129), .ZN(n1365) );
  OAI22_X1 U417 ( .A1(n647), .A2(n1130), .B1(n614), .B2(n1131), .ZN(n1364) );
  NOR4_X1 U418 ( .A1(n1368), .A2(n1369), .A3(n1371), .A4(n1372), .ZN(n1357) );
  OAI22_X1 U419 ( .A1(n715), .A2(n1136), .B1(n681), .B2(n1137), .ZN(n1372) );
  OAI22_X1 U420 ( .A1(n782), .A2(n1138), .B1(n748), .B2(n1139), .ZN(n1371) );
  OAI22_X1 U421 ( .A1(n849), .A2(n1140), .B1(n815), .B2(n1141), .ZN(n1369) );
  OAI22_X1 U422 ( .A1(n916), .A2(n1142), .B1(n883), .B2(n1143), .ZN(n1368) );
  NOR4_X1 U423 ( .A1(n1373), .A2(n1374), .A3(n1375), .A4(n1376), .ZN(n1356) );
  OAI22_X1 U424 ( .A1(n983), .A2(n1148), .B1(n950), .B2(n1149), .ZN(n1376) );
  OAI22_X1 U425 ( .A1(n1051), .A2(n1151), .B1(n1017), .B2(n1152), .ZN(n1375)
         );
  OAI22_X1 U426 ( .A1(n91), .A2(n1153), .B1(n1084), .B2(n2), .ZN(n1374) );
  OAI22_X1 U427 ( .A1(n166), .A2(n3), .B1(n130), .B2(n37), .ZN(n1373) );
  OAI22_X1 U428 ( .A1(n1377), .A2(n1102), .B1(n1103), .B2(n1370), .ZN(N4594)
         );
  NOR4_X1 U429 ( .A1(n1382), .A2(n1383), .A3(n1384), .A4(n1385), .ZN(n1381) );
  OAI22_X1 U430 ( .A1(n188), .A2(n1112), .B1(n858), .B2(n1113), .ZN(n1385) );
  OAI22_X1 U431 ( .A1(n252), .A2(n1114), .B1(n220), .B2(n1115), .ZN(n1384) );
  OAI22_X1 U432 ( .A1(n316), .A2(n1116), .B1(n284), .B2(n1117), .ZN(n1383) );
  OAI22_X1 U433 ( .A1(n380), .A2(n1118), .B1(n348), .B2(n1119), .ZN(n1382) );
  NOR4_X1 U434 ( .A1(n1386), .A2(n1387), .A3(n1388), .A4(n1389), .ZN(n1380) );
  OAI22_X1 U435 ( .A1(n445), .A2(n1124), .B1(n412), .B2(n1125), .ZN(n1389) );
  OAI22_X1 U436 ( .A1(n512), .A2(n1126), .B1(n478), .B2(n1127), .ZN(n1388) );
  OAI22_X1 U437 ( .A1(n579), .A2(n1128), .B1(n546), .B2(n1129), .ZN(n1387) );
  OAI22_X1 U438 ( .A1(n646), .A2(n1130), .B1(n613), .B2(n1131), .ZN(n1386) );
  NOR4_X1 U439 ( .A1(n1390), .A2(n1391), .A3(n1393), .A4(n1394), .ZN(n1379) );
  OAI22_X1 U440 ( .A1(n714), .A2(n1136), .B1(n680), .B2(n1137), .ZN(n1394) );
  OAI22_X1 U441 ( .A1(n781), .A2(n1138), .B1(n747), .B2(n1139), .ZN(n1393) );
  OAI22_X1 U442 ( .A1(n848), .A2(n1140), .B1(n814), .B2(n1141), .ZN(n1391) );
  OAI22_X1 U443 ( .A1(n915), .A2(n1142), .B1(n882), .B2(n1143), .ZN(n1390) );
  NOR4_X1 U444 ( .A1(n1395), .A2(n1396), .A3(n1397), .A4(n1398), .ZN(n1378) );
  OAI22_X1 U445 ( .A1(n982), .A2(n1148), .B1(n949), .B2(n1149), .ZN(n1398) );
  OAI22_X1 U446 ( .A1(n1050), .A2(n1151), .B1(n1016), .B2(n1152), .ZN(n1397)
         );
  OAI22_X1 U447 ( .A1(n89), .A2(n1153), .B1(n1083), .B2(n2), .ZN(n1396) );
  OAI22_X1 U448 ( .A1(n165), .A2(n3), .B1(n129), .B2(n1156), .ZN(n1395) );
  OAI22_X1 U449 ( .A1(n1399), .A2(n1102), .B1(n1103), .B2(n1392), .ZN(N4592)
         );
  NOR4_X1 U450 ( .A1(n1404), .A2(n1405), .A3(n1406), .A4(n1407), .ZN(n1403) );
  OAI22_X1 U451 ( .A1(n187), .A2(n1112), .B1(n837), .B2(n1113), .ZN(n1407) );
  OAI22_X1 U452 ( .A1(n251), .A2(n1114), .B1(n219), .B2(n1115), .ZN(n1406) );
  OAI22_X1 U453 ( .A1(n315), .A2(n1116), .B1(n283), .B2(n1117), .ZN(n1405) );
  OAI22_X1 U454 ( .A1(n379), .A2(n1118), .B1(n347), .B2(n1119), .ZN(n1404) );
  NOR4_X1 U455 ( .A1(n1408), .A2(n1409), .A3(n1410), .A4(n1411), .ZN(n1402) );
  OAI22_X1 U456 ( .A1(n444), .A2(n1124), .B1(n411), .B2(n1125), .ZN(n1411) );
  OAI22_X1 U457 ( .A1(n511), .A2(n1126), .B1(n477), .B2(n1127), .ZN(n1410) );
  OAI22_X1 U458 ( .A1(n578), .A2(n1128), .B1(n545), .B2(n1129), .ZN(n1409) );
  OAI22_X1 U459 ( .A1(n645), .A2(n1130), .B1(n612), .B2(n1131), .ZN(n1408) );
  NOR4_X1 U460 ( .A1(n1412), .A2(n1413), .A3(n1415), .A4(n1416), .ZN(n1401) );
  OAI22_X1 U461 ( .A1(n713), .A2(n1136), .B1(n679), .B2(n1137), .ZN(n1416) );
  OAI22_X1 U462 ( .A1(n780), .A2(n1138), .B1(n746), .B2(n1139), .ZN(n1415) );
  OAI22_X1 U463 ( .A1(n847), .A2(n1140), .B1(n813), .B2(n1141), .ZN(n1413) );
  OAI22_X1 U464 ( .A1(n914), .A2(n1142), .B1(n881), .B2(n1143), .ZN(n1412) );
  NOR4_X1 U465 ( .A1(n1417), .A2(n1418), .A3(n1419), .A4(n1420), .ZN(n1400) );
  OAI22_X1 U466 ( .A1(n981), .A2(n1148), .B1(n948), .B2(n1149), .ZN(n1420) );
  OAI22_X1 U467 ( .A1(n1049), .A2(n1151), .B1(n1015), .B2(n1152), .ZN(n1419)
         );
  OAI22_X1 U468 ( .A1(n87), .A2(n1), .B1(n1082), .B2(n2), .ZN(n1418) );
  OAI22_X1 U469 ( .A1(n163), .A2(n1155), .B1(n128), .B2(n1156), .ZN(n1417) );
  OAI22_X1 U470 ( .A1(n1421), .A2(n1102), .B1(n1103), .B2(n1414), .ZN(N4590)
         );
  NOR4_X1 U471 ( .A1(n1426), .A2(n1427), .A3(n1428), .A4(n1429), .ZN(n1425) );
  OAI22_X1 U472 ( .A1(n186), .A2(n1112), .B1(n816), .B2(n1113), .ZN(n1429) );
  OAI22_X1 U473 ( .A1(n250), .A2(n1114), .B1(n218), .B2(n1115), .ZN(n1428) );
  OAI22_X1 U474 ( .A1(n314), .A2(n1116), .B1(n282), .B2(n1117), .ZN(n1427) );
  OAI22_X1 U475 ( .A1(n378), .A2(n1118), .B1(n346), .B2(n1119), .ZN(n1426) );
  NOR4_X1 U476 ( .A1(n1430), .A2(n1431), .A3(n1432), .A4(n1433), .ZN(n1424) );
  OAI22_X1 U477 ( .A1(n443), .A2(n1124), .B1(n410), .B2(n1125), .ZN(n1433) );
  OAI22_X1 U478 ( .A1(n510), .A2(n1126), .B1(n476), .B2(n1127), .ZN(n1432) );
  OAI22_X1 U479 ( .A1(n577), .A2(n1128), .B1(n544), .B2(n1129), .ZN(n1431) );
  OAI22_X1 U480 ( .A1(n644), .A2(n1130), .B1(n611), .B2(n1131), .ZN(n1430) );
  NOR4_X1 U481 ( .A1(n1434), .A2(n1435), .A3(n1437), .A4(n1438), .ZN(n1423) );
  OAI22_X1 U482 ( .A1(n712), .A2(n1136), .B1(n678), .B2(n1137), .ZN(n1438) );
  OAI22_X1 U483 ( .A1(n779), .A2(n1138), .B1(n745), .B2(n1139), .ZN(n1437) );
  OAI22_X1 U484 ( .A1(n846), .A2(n1140), .B1(n812), .B2(n1141), .ZN(n1435) );
  OAI22_X1 U485 ( .A1(n913), .A2(n1142), .B1(n880), .B2(n1143), .ZN(n1434) );
  NOR4_X1 U486 ( .A1(n1439), .A2(n1440), .A3(n1441), .A4(n1442), .ZN(n1422) );
  OAI22_X1 U487 ( .A1(n980), .A2(n1148), .B1(n947), .B2(n1149), .ZN(n1442) );
  OAI22_X1 U488 ( .A1(n1048), .A2(n1151), .B1(n1014), .B2(n1152), .ZN(n1441)
         );
  OAI22_X1 U489 ( .A1(n85), .A2(n1), .B1(n1081), .B2(n2), .ZN(n1440) );
  OAI22_X1 U490 ( .A1(n162), .A2(n1155), .B1(n127), .B2(n1156), .ZN(n1439) );
  OAI22_X1 U491 ( .A1(n1443), .A2(n1102), .B1(n1103), .B2(n1436), .ZN(N4588)
         );
  NOR4_X1 U492 ( .A1(n1448), .A2(n1449), .A3(n1450), .A4(n1451), .ZN(n1447) );
  OAI22_X1 U493 ( .A1(n185), .A2(n1112), .B1(n795), .B2(n1113), .ZN(n1451) );
  OAI22_X1 U494 ( .A1(n249), .A2(n1114), .B1(n217), .B2(n1115), .ZN(n1450) );
  OAI22_X1 U495 ( .A1(n313), .A2(n1116), .B1(n281), .B2(n1117), .ZN(n1449) );
  OAI22_X1 U496 ( .A1(n377), .A2(n1118), .B1(n345), .B2(n1119), .ZN(n1448) );
  NOR4_X1 U497 ( .A1(n1452), .A2(n1453), .A3(n1454), .A4(n1455), .ZN(n1446) );
  OAI22_X1 U498 ( .A1(n442), .A2(n1124), .B1(n409), .B2(n1125), .ZN(n1455) );
  OAI22_X1 U499 ( .A1(n509), .A2(n1126), .B1(n475), .B2(n1127), .ZN(n1454) );
  OAI22_X1 U500 ( .A1(n576), .A2(n1128), .B1(n542), .B2(n1129), .ZN(n1453) );
  OAI22_X1 U501 ( .A1(n643), .A2(n1130), .B1(n610), .B2(n1131), .ZN(n1452) );
  NOR4_X1 U502 ( .A1(n1456), .A2(n1457), .A3(n1459), .A4(n1460), .ZN(n1445) );
  OAI22_X1 U503 ( .A1(n710), .A2(n1136), .B1(n677), .B2(n1137), .ZN(n1460) );
  OAI22_X1 U504 ( .A1(n778), .A2(n1138), .B1(n744), .B2(n1139), .ZN(n1459) );
  OAI22_X1 U505 ( .A1(n845), .A2(n1140), .B1(n811), .B2(n1141), .ZN(n1457) );
  OAI22_X1 U506 ( .A1(n912), .A2(n1142), .B1(n878), .B2(n1143), .ZN(n1456) );
  NOR4_X1 U507 ( .A1(n1461), .A2(n1462), .A3(n1463), .A4(n1464), .ZN(n1444) );
  OAI22_X1 U508 ( .A1(n979), .A2(n1148), .B1(n946), .B2(n1149), .ZN(n1464) );
  OAI22_X1 U509 ( .A1(n1046), .A2(n1151), .B1(n1013), .B2(n1152), .ZN(n1463)
         );
  OAI22_X1 U510 ( .A1(n83), .A2(n1), .B1(n1080), .B2(n2), .ZN(n1462) );
  OAI22_X1 U511 ( .A1(n161), .A2(n1155), .B1(n126), .B2(n1156), .ZN(n1461) );
  OAI22_X1 U512 ( .A1(n1465), .A2(n1102), .B1(n1103), .B2(n1458), .ZN(N4586)
         );
  NOR4_X1 U513 ( .A1(n1470), .A2(n1471), .A3(n1472), .A4(n1473), .ZN(n1469) );
  OAI22_X1 U514 ( .A1(n184), .A2(n1112), .B1(n774), .B2(n1113), .ZN(n1473) );
  OAI22_X1 U515 ( .A1(n248), .A2(n1114), .B1(n216), .B2(n1115), .ZN(n1472) );
  OAI22_X1 U516 ( .A1(n312), .A2(n1116), .B1(n280), .B2(n1117), .ZN(n1471) );
  OAI22_X1 U517 ( .A1(n376), .A2(n1118), .B1(n344), .B2(n1119), .ZN(n1470) );
  NOR4_X1 U518 ( .A1(n1474), .A2(n1475), .A3(n1476), .A4(n1477), .ZN(n1468) );
  OAI22_X1 U519 ( .A1(n441), .A2(n1124), .B1(n408), .B2(n1125), .ZN(n1477) );
  OAI22_X1 U520 ( .A1(n508), .A2(n1126), .B1(n474), .B2(n1127), .ZN(n1476) );
  OAI22_X1 U521 ( .A1(n575), .A2(n1128), .B1(n541), .B2(n1129), .ZN(n1475) );
  OAI22_X1 U522 ( .A1(n642), .A2(n1130), .B1(n609), .B2(n1131), .ZN(n1474) );
  NOR4_X1 U523 ( .A1(n1478), .A2(n1479), .A3(n1481), .A4(n1482), .ZN(n1467) );
  OAI22_X1 U524 ( .A1(n709), .A2(n1136), .B1(n676), .B2(n1137), .ZN(n1482) );
  OAI22_X1 U525 ( .A1(n777), .A2(n1138), .B1(n743), .B2(n1139), .ZN(n1481) );
  OAI22_X1 U526 ( .A1(n844), .A2(n1140), .B1(n810), .B2(n1141), .ZN(n1479) );
  OAI22_X1 U527 ( .A1(n911), .A2(n1142), .B1(n877), .B2(n1143), .ZN(n1478) );
  NOR4_X1 U528 ( .A1(n1483), .A2(n1484), .A3(n1485), .A4(n1486), .ZN(n1466) );
  OAI22_X1 U529 ( .A1(n978), .A2(n1148), .B1(n945), .B2(n1149), .ZN(n1486) );
  OAI22_X1 U530 ( .A1(n1045), .A2(n1151), .B1(n1012), .B2(n1152), .ZN(n1485)
         );
  OAI22_X1 U531 ( .A1(n81), .A2(n1), .B1(n1079), .B2(n2), .ZN(n1484) );
  OAI22_X1 U532 ( .A1(n160), .A2(n1155), .B1(n125), .B2(n1156), .ZN(n1483) );
  OAI22_X1 U533 ( .A1(n1487), .A2(n1102), .B1(n1103), .B2(n1480), .ZN(N4584)
         );
  NOR4_X1 U534 ( .A1(n1492), .A2(n1493), .A3(n1494), .A4(n1495), .ZN(n1491) );
  OAI22_X1 U535 ( .A1(n183), .A2(n1112), .B1(n753), .B2(n1113), .ZN(n1495) );
  OAI22_X1 U536 ( .A1(n247), .A2(n1114), .B1(n215), .B2(n1115), .ZN(n1494) );
  OAI22_X1 U537 ( .A1(n311), .A2(n1116), .B1(n279), .B2(n1117), .ZN(n1493) );
  OAI22_X1 U538 ( .A1(n375), .A2(n1118), .B1(n343), .B2(n1119), .ZN(n1492) );
  NOR4_X1 U539 ( .A1(n1496), .A2(n1497), .A3(n1498), .A4(n1499), .ZN(n1490) );
  OAI22_X1 U540 ( .A1(n440), .A2(n1124), .B1(n407), .B2(n1125), .ZN(n1499) );
  OAI22_X1 U541 ( .A1(n507), .A2(n1126), .B1(n473), .B2(n1127), .ZN(n1498) );
  OAI22_X1 U542 ( .A1(n574), .A2(n1128), .B1(n540), .B2(n1129), .ZN(n1497) );
  OAI22_X1 U543 ( .A1(n641), .A2(n1130), .B1(n608), .B2(n1131), .ZN(n1496) );
  NOR4_X1 U544 ( .A1(n1500), .A2(n1501), .A3(n1503), .A4(n1504), .ZN(n1489) );
  OAI22_X1 U545 ( .A1(n708), .A2(n1136), .B1(n675), .B2(n1137), .ZN(n1504) );
  OAI22_X1 U546 ( .A1(n776), .A2(n1138), .B1(n742), .B2(n1139), .ZN(n1503) );
  OAI22_X1 U547 ( .A1(n843), .A2(n1140), .B1(n809), .B2(n1141), .ZN(n1501) );
  OAI22_X1 U548 ( .A1(n910), .A2(n1142), .B1(n876), .B2(n1143), .ZN(n1500) );
  NOR4_X1 U549 ( .A1(n1505), .A2(n1506), .A3(n1507), .A4(n1508), .ZN(n1488) );
  OAI22_X1 U550 ( .A1(n977), .A2(n1148), .B1(n944), .B2(n1149), .ZN(n1508) );
  OAI22_X1 U551 ( .A1(n1044), .A2(n1151), .B1(n1011), .B2(n1152), .ZN(n1507)
         );
  OAI22_X1 U552 ( .A1(n79), .A2(n1), .B1(n1078), .B2(n2), .ZN(n1506) );
  OAI22_X1 U553 ( .A1(n159), .A2(n1155), .B1(n124), .B2(n1156), .ZN(n1505) );
  OAI22_X1 U554 ( .A1(n1509), .A2(n1102), .B1(n1103), .B2(n1502), .ZN(N4582)
         );
  NOR4_X1 U555 ( .A1(n1514), .A2(n1515), .A3(n1516), .A4(n1517), .ZN(n1513) );
  OAI22_X1 U556 ( .A1(n182), .A2(n1112), .B1(n732), .B2(n1113), .ZN(n1517) );
  OAI22_X1 U557 ( .A1(n246), .A2(n1114), .B1(n214), .B2(n1115), .ZN(n1516) );
  OAI22_X1 U558 ( .A1(n310), .A2(n1116), .B1(n278), .B2(n1117), .ZN(n1515) );
  OAI22_X1 U559 ( .A1(n374), .A2(n1118), .B1(n342), .B2(n1119), .ZN(n1514) );
  NOR4_X1 U560 ( .A1(n1518), .A2(n1519), .A3(n1520), .A4(n1521), .ZN(n1512) );
  OAI22_X1 U561 ( .A1(n439), .A2(n1124), .B1(n406), .B2(n1125), .ZN(n1521) );
  OAI22_X1 U562 ( .A1(n506), .A2(n1126), .B1(n472), .B2(n1127), .ZN(n1520) );
  OAI22_X1 U563 ( .A1(n573), .A2(n1128), .B1(n539), .B2(n1129), .ZN(n1519) );
  OAI22_X1 U564 ( .A1(n640), .A2(n1130), .B1(n607), .B2(n1131), .ZN(n1518) );
  NOR4_X1 U565 ( .A1(n1522), .A2(n1523), .A3(n1525), .A4(n1526), .ZN(n1511) );
  OAI22_X1 U566 ( .A1(n707), .A2(n1136), .B1(n674), .B2(n1137), .ZN(n1526) );
  OAI22_X1 U567 ( .A1(n775), .A2(n1138), .B1(n741), .B2(n1139), .ZN(n1525) );
  OAI22_X1 U568 ( .A1(n842), .A2(n1140), .B1(n808), .B2(n1141), .ZN(n1523) );
  OAI22_X1 U569 ( .A1(n909), .A2(n1142), .B1(n875), .B2(n1143), .ZN(n1522) );
  NOR4_X1 U570 ( .A1(n1527), .A2(n1528), .A3(n1529), .A4(n1530), .ZN(n1510) );
  OAI22_X1 U571 ( .A1(n976), .A2(n1148), .B1(n943), .B2(n1149), .ZN(n1530) );
  OAI22_X1 U572 ( .A1(n1043), .A2(n1151), .B1(n1010), .B2(n1152), .ZN(n1529)
         );
  OAI22_X1 U573 ( .A1(n77), .A2(n1), .B1(n1077), .B2(n2), .ZN(n1528) );
  OAI22_X1 U574 ( .A1(n158), .A2(n1155), .B1(n123), .B2(n1156), .ZN(n1527) );
  OAI22_X1 U575 ( .A1(n1531), .A2(n1102), .B1(n1103), .B2(n1524), .ZN(N4580)
         );
  NOR4_X1 U576 ( .A1(n1536), .A2(n1537), .A3(n1538), .A4(n1539), .ZN(n1535) );
  OAI22_X1 U577 ( .A1(n181), .A2(n1112), .B1(n711), .B2(n1113), .ZN(n1539) );
  OAI22_X1 U578 ( .A1(n245), .A2(n1114), .B1(n213), .B2(n1115), .ZN(n1538) );
  OAI22_X1 U579 ( .A1(n309), .A2(n1116), .B1(n277), .B2(n1117), .ZN(n1537) );
  OAI22_X1 U580 ( .A1(n373), .A2(n1118), .B1(n341), .B2(n1119), .ZN(n1536) );
  NOR4_X1 U581 ( .A1(n1540), .A2(n1541), .A3(n1542), .A4(n1543), .ZN(n1534) );
  OAI22_X1 U582 ( .A1(n437), .A2(n1124), .B1(n405), .B2(n1125), .ZN(n1543) );
  OAI22_X1 U583 ( .A1(n505), .A2(n1126), .B1(n471), .B2(n1127), .ZN(n1542) );
  OAI22_X1 U584 ( .A1(n572), .A2(n1128), .B1(n538), .B2(n1129), .ZN(n1541) );
  OAI22_X1 U585 ( .A1(n639), .A2(n1130), .B1(n605), .B2(n1131), .ZN(n1540) );
  NOR4_X1 U586 ( .A1(n1544), .A2(n1545), .A3(n1547), .A4(n1548), .ZN(n1533) );
  OAI22_X1 U587 ( .A1(n706), .A2(n1136), .B1(n673), .B2(n1137), .ZN(n1548) );
  OAI22_X1 U588 ( .A1(n773), .A2(n1138), .B1(n740), .B2(n1139), .ZN(n1547) );
  OAI22_X1 U589 ( .A1(n841), .A2(n1140), .B1(n807), .B2(n1141), .ZN(n1545) );
  OAI22_X1 U590 ( .A1(n908), .A2(n1142), .B1(n874), .B2(n1143), .ZN(n1544) );
  NOR4_X1 U591 ( .A1(n1549), .A2(n1550), .A3(n1551), .A4(n1552), .ZN(n1532) );
  OAI22_X1 U592 ( .A1(n975), .A2(n1148), .B1(n941), .B2(n1149), .ZN(n1552) );
  OAI22_X1 U593 ( .A1(n1042), .A2(n1151), .B1(n1009), .B2(n1152), .ZN(n1551)
         );
  OAI22_X1 U594 ( .A1(n73), .A2(n1), .B1(n1076), .B2(n2), .ZN(n1550) );
  OAI22_X1 U595 ( .A1(n157), .A2(n1155), .B1(n122), .B2(n1156), .ZN(n1549) );
  OAI22_X1 U596 ( .A1(n1553), .A2(n1102), .B1(n1103), .B2(n1546), .ZN(N4578)
         );
  NOR4_X1 U597 ( .A1(n1558), .A2(n1559), .A3(n1560), .A4(n1561), .ZN(n1557) );
  OAI22_X1 U598 ( .A1(n180), .A2(n1112), .B1(n690), .B2(n1113), .ZN(n1561) );
  OAI22_X1 U599 ( .A1(n244), .A2(n1114), .B1(n212), .B2(n1115), .ZN(n1560) );
  OAI22_X1 U600 ( .A1(n308), .A2(n1116), .B1(n276), .B2(n1117), .ZN(n1559) );
  OAI22_X1 U601 ( .A1(n372), .A2(n1118), .B1(n340), .B2(n1119), .ZN(n1558) );
  NOR4_X1 U602 ( .A1(n1562), .A2(n1563), .A3(n1564), .A4(n1565), .ZN(n1556) );
  OAI22_X1 U603 ( .A1(n436), .A2(n1124), .B1(n404), .B2(n1125), .ZN(n1565) );
  OAI22_X1 U604 ( .A1(n504), .A2(n1126), .B1(n470), .B2(n1127), .ZN(n1564) );
  OAI22_X1 U605 ( .A1(n571), .A2(n1128), .B1(n537), .B2(n1129), .ZN(n1563) );
  OAI22_X1 U606 ( .A1(n638), .A2(n1130), .B1(n604), .B2(n1131), .ZN(n1562) );
  NOR4_X1 U607 ( .A1(n1566), .A2(n1567), .A3(n1569), .A4(n1570), .ZN(n1555) );
  OAI22_X1 U608 ( .A1(n705), .A2(n1136), .B1(n672), .B2(n1137), .ZN(n1570) );
  OAI22_X1 U609 ( .A1(n772), .A2(n1138), .B1(n739), .B2(n1139), .ZN(n1569) );
  OAI22_X1 U610 ( .A1(n840), .A2(n1140), .B1(n806), .B2(n1141), .ZN(n1567) );
  OAI22_X1 U611 ( .A1(n907), .A2(n1142), .B1(n873), .B2(n1143), .ZN(n1566) );
  NOR4_X1 U612 ( .A1(n1571), .A2(n1572), .A3(n1573), .A4(n1574), .ZN(n1554) );
  OAI22_X1 U613 ( .A1(n974), .A2(n1148), .B1(n940), .B2(n1149), .ZN(n1574) );
  OAI22_X1 U614 ( .A1(n1041), .A2(n1151), .B1(n1008), .B2(n1152), .ZN(n1573)
         );
  OAI22_X1 U615 ( .A1(n71), .A2(n1), .B1(n1075), .B2(n2), .ZN(n1572) );
  OAI22_X1 U616 ( .A1(n156), .A2(n1155), .B1(n121), .B2(n1156), .ZN(n1571) );
  OAI22_X1 U617 ( .A1(n1575), .A2(n1102), .B1(n1103), .B2(n1568), .ZN(N4576)
         );
  NOR4_X1 U618 ( .A1(n1580), .A2(n1581), .A3(n1582), .A4(n1583), .ZN(n1579) );
  OAI22_X1 U619 ( .A1(n179), .A2(n1112), .B1(n669), .B2(n1113), .ZN(n1583) );
  OAI22_X1 U620 ( .A1(n243), .A2(n1114), .B1(n211), .B2(n1115), .ZN(n1582) );
  OAI22_X1 U621 ( .A1(n307), .A2(n1116), .B1(n275), .B2(n1117), .ZN(n1581) );
  OAI22_X1 U622 ( .A1(n371), .A2(n1118), .B1(n339), .B2(n1119), .ZN(n1580) );
  NOR4_X1 U623 ( .A1(n1584), .A2(n1585), .A3(n1586), .A4(n1587), .ZN(n1578) );
  OAI22_X1 U624 ( .A1(n435), .A2(n1124), .B1(n403), .B2(n1125), .ZN(n1587) );
  OAI22_X1 U625 ( .A1(n503), .A2(n1126), .B1(n469), .B2(n1127), .ZN(n1586) );
  OAI22_X1 U626 ( .A1(n570), .A2(n1128), .B1(n536), .B2(n1129), .ZN(n1585) );
  OAI22_X1 U627 ( .A1(n637), .A2(n1130), .B1(n603), .B2(n1131), .ZN(n1584) );
  NOR4_X1 U628 ( .A1(n1588), .A2(n1589), .A3(n1591), .A4(n1592), .ZN(n1577) );
  OAI22_X1 U629 ( .A1(n704), .A2(n1136), .B1(n671), .B2(n1137), .ZN(n1592) );
  OAI22_X1 U630 ( .A1(n771), .A2(n1138), .B1(n738), .B2(n1139), .ZN(n1591) );
  OAI22_X1 U631 ( .A1(n839), .A2(n1140), .B1(n805), .B2(n1141), .ZN(n1589) );
  OAI22_X1 U632 ( .A1(n906), .A2(n1142), .B1(n872), .B2(n1143), .ZN(n1588) );
  NOR4_X1 U633 ( .A1(n1593), .A2(n1594), .A3(n1595), .A4(n1596), .ZN(n1576) );
  OAI22_X1 U634 ( .A1(n973), .A2(n1148), .B1(n939), .B2(n1149), .ZN(n1596) );
  OAI22_X1 U635 ( .A1(n1040), .A2(n1151), .B1(n1007), .B2(n1152), .ZN(n1595)
         );
  OAI22_X1 U636 ( .A1(n69), .A2(n1), .B1(n1074), .B2(n1154), .ZN(n1594) );
  OAI22_X1 U637 ( .A1(n155), .A2(n1155), .B1(n119), .B2(n1156), .ZN(n1593) );
  OAI22_X1 U638 ( .A1(n1597), .A2(n1102), .B1(n1103), .B2(n1590), .ZN(N4574)
         );
  NOR4_X1 U639 ( .A1(n1602), .A2(n1603), .A3(n1604), .A4(n1605), .ZN(n1601) );
  OAI22_X1 U640 ( .A1(n178), .A2(n1112), .B1(n648), .B2(n1113), .ZN(n1605) );
  OAI22_X1 U641 ( .A1(n242), .A2(n1114), .B1(n210), .B2(n1115), .ZN(n1604) );
  OAI22_X1 U642 ( .A1(n306), .A2(n1116), .B1(n274), .B2(n1117), .ZN(n1603) );
  OAI22_X1 U643 ( .A1(n370), .A2(n1118), .B1(n338), .B2(n1119), .ZN(n1602) );
  NOR4_X1 U644 ( .A1(n1606), .A2(n1607), .A3(n1608), .A4(n1609), .ZN(n1600) );
  OAI22_X1 U645 ( .A1(n434), .A2(n1124), .B1(n402), .B2(n1125), .ZN(n1609) );
  OAI22_X1 U646 ( .A1(n502), .A2(n1126), .B1(n468), .B2(n1127), .ZN(n1608) );
  OAI22_X1 U647 ( .A1(n569), .A2(n1128), .B1(n535), .B2(n1129), .ZN(n1607) );
  OAI22_X1 U648 ( .A1(n636), .A2(n1130), .B1(n602), .B2(n1131), .ZN(n1606) );
  NOR4_X1 U649 ( .A1(n1610), .A2(n1611), .A3(n1613), .A4(n1614), .ZN(n1599) );
  OAI22_X1 U650 ( .A1(n703), .A2(n1136), .B1(n670), .B2(n1137), .ZN(n1614) );
  OAI22_X1 U651 ( .A1(n770), .A2(n1138), .B1(n737), .B2(n1139), .ZN(n1613) );
  OAI22_X1 U652 ( .A1(n838), .A2(n1140), .B1(n804), .B2(n1141), .ZN(n1611) );
  OAI22_X1 U653 ( .A1(n905), .A2(n1142), .B1(n871), .B2(n1143), .ZN(n1610) );
  NOR4_X1 U654 ( .A1(n1615), .A2(n1616), .A3(n1617), .A4(n1618), .ZN(n1598) );
  OAI22_X1 U655 ( .A1(n972), .A2(n1148), .B1(n938), .B2(n1149), .ZN(n1618) );
  OAI22_X1 U656 ( .A1(n1039), .A2(n1151), .B1(n1006), .B2(n1152), .ZN(n1617)
         );
  OAI22_X1 U657 ( .A1(n67), .A2(n1), .B1(n1073), .B2(n1154), .ZN(n1616) );
  OAI22_X1 U658 ( .A1(n154), .A2(n1155), .B1(n118), .B2(n1156), .ZN(n1615) );
  OAI22_X1 U659 ( .A1(n1619), .A2(n1102), .B1(n1103), .B2(n1612), .ZN(N4572)
         );
  NOR4_X1 U660 ( .A1(n1624), .A2(n1625), .A3(n1626), .A4(n1627), .ZN(n1623) );
  OAI22_X1 U661 ( .A1(n175), .A2(n1112), .B1(n627), .B2(n1113), .ZN(n1627) );
  OAI22_X1 U662 ( .A1(n241), .A2(n1114), .B1(n209), .B2(n1115), .ZN(n1626) );
  OAI22_X1 U663 ( .A1(n305), .A2(n1116), .B1(n273), .B2(n1117), .ZN(n1625) );
  OAI22_X1 U664 ( .A1(n369), .A2(n1118), .B1(n337), .B2(n1119), .ZN(n1624) );
  NOR4_X1 U665 ( .A1(n1628), .A2(n1629), .A3(n1630), .A4(n1631), .ZN(n1622) );
  OAI22_X1 U666 ( .A1(n433), .A2(n1124), .B1(n401), .B2(n1125), .ZN(n1631) );
  OAI22_X1 U667 ( .A1(n500), .A2(n1126), .B1(n467), .B2(n1127), .ZN(n1630) );
  OAI22_X1 U668 ( .A1(n568), .A2(n1128), .B1(n534), .B2(n1129), .ZN(n1629) );
  OAI22_X1 U669 ( .A1(n635), .A2(n1130), .B1(n601), .B2(n1131), .ZN(n1628) );
  NOR4_X1 U670 ( .A1(n1632), .A2(n1633), .A3(n1635), .A4(n1636), .ZN(n1621) );
  OAI22_X1 U671 ( .A1(n702), .A2(n1136), .B1(n668), .B2(n1137), .ZN(n1636) );
  OAI22_X1 U672 ( .A1(n769), .A2(n1138), .B1(n736), .B2(n1139), .ZN(n1635) );
  OAI22_X1 U673 ( .A1(n836), .A2(n1140), .B1(n803), .B2(n1141), .ZN(n1633) );
  OAI22_X1 U674 ( .A1(n904), .A2(n1142), .B1(n870), .B2(n1143), .ZN(n1632) );
  NOR4_X1 U675 ( .A1(n1637), .A2(n1638), .A3(n1639), .A4(n1640), .ZN(n1620) );
  OAI22_X1 U676 ( .A1(n971), .A2(n1148), .B1(n937), .B2(n1149), .ZN(n1640) );
  OAI22_X1 U677 ( .A1(n1038), .A2(n1151), .B1(n1004), .B2(n1152), .ZN(n1639)
         );
  OAI22_X1 U678 ( .A1(n65), .A2(n1), .B1(n1072), .B2(n1154), .ZN(n1638) );
  OAI22_X1 U679 ( .A1(n152), .A2(n1155), .B1(n117), .B2(n1156), .ZN(n1637) );
  OAI22_X1 U680 ( .A1(n1641), .A2(n1102), .B1(n1103), .B2(n1634), .ZN(N4570)
         );
  NOR4_X1 U681 ( .A1(n1646), .A2(n1647), .A3(n1648), .A4(n1649), .ZN(n1645) );
  OAI22_X1 U682 ( .A1(n164), .A2(n1112), .B1(n606), .B2(n1113), .ZN(n1649) );
  OAI22_X1 U683 ( .A1(n240), .A2(n1114), .B1(n208), .B2(n1115), .ZN(n1648) );
  OAI22_X1 U684 ( .A1(n304), .A2(n1116), .B1(n272), .B2(n1117), .ZN(n1647) );
  OAI22_X1 U685 ( .A1(n368), .A2(n1118), .B1(n336), .B2(n1119), .ZN(n1646) );
  NOR4_X1 U686 ( .A1(n1650), .A2(n1651), .A3(n1652), .A4(n1653), .ZN(n1644) );
  OAI22_X1 U687 ( .A1(n432), .A2(n1124), .B1(n400), .B2(n1125), .ZN(n1653) );
  OAI22_X1 U688 ( .A1(n499), .A2(n1126), .B1(n466), .B2(n1127), .ZN(n1652) );
  OAI22_X1 U689 ( .A1(n567), .A2(n1128), .B1(n533), .B2(n1129), .ZN(n1651) );
  OAI22_X1 U690 ( .A1(n634), .A2(n1130), .B1(n600), .B2(n1131), .ZN(n1650) );
  NOR4_X1 U691 ( .A1(n1654), .A2(n1655), .A3(n1657), .A4(n1658), .ZN(n1643) );
  OAI22_X1 U692 ( .A1(n701), .A2(n1136), .B1(n667), .B2(n1137), .ZN(n1658) );
  OAI22_X1 U693 ( .A1(n768), .A2(n1138), .B1(n735), .B2(n1139), .ZN(n1657) );
  OAI22_X1 U694 ( .A1(n835), .A2(n1140), .B1(n802), .B2(n1141), .ZN(n1655) );
  OAI22_X1 U695 ( .A1(n903), .A2(n1142), .B1(n869), .B2(n1143), .ZN(n1654) );
  NOR4_X1 U696 ( .A1(n1659), .A2(n1660), .A3(n1661), .A4(n1662), .ZN(n1642) );
  OAI22_X1 U697 ( .A1(n970), .A2(n1148), .B1(n936), .B2(n1149), .ZN(n1662) );
  OAI22_X1 U698 ( .A1(n1037), .A2(n1151), .B1(n1003), .B2(n1152), .ZN(n1661)
         );
  OAI22_X1 U699 ( .A1(n63), .A2(n1), .B1(n1071), .B2(n1154), .ZN(n1660) );
  OAI22_X1 U700 ( .A1(n151), .A2(n3), .B1(n116), .B2(n37), .ZN(n1659) );
  OAI22_X1 U701 ( .A1(n1663), .A2(n1102), .B1(n1103), .B2(n1656), .ZN(N4568)
         );
  NOR4_X1 U702 ( .A1(n1668), .A2(n1669), .A3(n1670), .A4(n1671), .ZN(n1667) );
  OAI22_X1 U703 ( .A1(n153), .A2(n1112), .B1(n585), .B2(n1113), .ZN(n1671) );
  OAI22_X1 U704 ( .A1(n239), .A2(n1114), .B1(n207), .B2(n1115), .ZN(n1670) );
  OAI22_X1 U705 ( .A1(n303), .A2(n1116), .B1(n271), .B2(n1117), .ZN(n1669) );
  OAI22_X1 U706 ( .A1(n367), .A2(n1118), .B1(n335), .B2(n1119), .ZN(n1668) );
  NOR4_X1 U707 ( .A1(n1672), .A2(n1673), .A3(n1674), .A4(n1675), .ZN(n1666) );
  OAI22_X1 U708 ( .A1(n431), .A2(n1124), .B1(n399), .B2(n1125), .ZN(n1675) );
  OAI22_X1 U709 ( .A1(n498), .A2(n1126), .B1(n465), .B2(n1127), .ZN(n1674) );
  OAI22_X1 U710 ( .A1(n566), .A2(n1128), .B1(n532), .B2(n1129), .ZN(n1673) );
  OAI22_X1 U711 ( .A1(n633), .A2(n1130), .B1(n599), .B2(n1131), .ZN(n1672) );
  NOR4_X1 U712 ( .A1(n1676), .A2(n1677), .A3(n1679), .A4(n1680), .ZN(n1665) );
  OAI22_X1 U713 ( .A1(n700), .A2(n1136), .B1(n666), .B2(n1137), .ZN(n1680) );
  OAI22_X1 U714 ( .A1(n767), .A2(n1138), .B1(n734), .B2(n1139), .ZN(n1679) );
  OAI22_X1 U715 ( .A1(n834), .A2(n1140), .B1(n801), .B2(n1141), .ZN(n1677) );
  OAI22_X1 U716 ( .A1(n902), .A2(n1142), .B1(n868), .B2(n1143), .ZN(n1676) );
  NOR4_X1 U717 ( .A1(n1681), .A2(n1682), .A3(n1683), .A4(n1684), .ZN(n1664) );
  OAI22_X1 U718 ( .A1(n969), .A2(n1148), .B1(n935), .B2(n1149), .ZN(n1684) );
  OAI22_X1 U719 ( .A1(n1036), .A2(n1151), .B1(n1002), .B2(n1152), .ZN(n1683)
         );
  OAI22_X1 U720 ( .A1(n61), .A2(n1), .B1(n1070), .B2(n1154), .ZN(n1682) );
  OAI22_X1 U721 ( .A1(n150), .A2(n3), .B1(n115), .B2(n1156), .ZN(n1681) );
  OAI22_X1 U722 ( .A1(n1685), .A2(n1102), .B1(n1103), .B2(n1678), .ZN(N4566)
         );
  NOR4_X1 U723 ( .A1(n1690), .A2(n1691), .A3(n1692), .A4(n1693), .ZN(n1689) );
  OAI22_X1 U724 ( .A1(n142), .A2(n1112), .B1(n564), .B2(n1113), .ZN(n1693) );
  OAI22_X1 U725 ( .A1(n238), .A2(n1114), .B1(n206), .B2(n1115), .ZN(n1692) );
  OAI22_X1 U726 ( .A1(n302), .A2(n1116), .B1(n270), .B2(n1117), .ZN(n1691) );
  OAI22_X1 U727 ( .A1(n366), .A2(n1118), .B1(n334), .B2(n1119), .ZN(n1690) );
  NOR4_X1 U728 ( .A1(n1694), .A2(n1695), .A3(n1696), .A4(n1697), .ZN(n1688) );
  OAI22_X1 U729 ( .A1(n430), .A2(n1124), .B1(n398), .B2(n1125), .ZN(n1697) );
  OAI22_X1 U730 ( .A1(n497), .A2(n1126), .B1(n464), .B2(n1127), .ZN(n1696) );
  OAI22_X1 U731 ( .A1(n565), .A2(n1128), .B1(n531), .B2(n1129), .ZN(n1695) );
  OAI22_X1 U732 ( .A1(n632), .A2(n1130), .B1(n598), .B2(n1131), .ZN(n1694) );
  NOR4_X1 U733 ( .A1(n1698), .A2(n1699), .A3(n1701), .A4(n1702), .ZN(n1687) );
  OAI22_X1 U734 ( .A1(n699), .A2(n1136), .B1(n665), .B2(n1137), .ZN(n1702) );
  OAI22_X1 U735 ( .A1(n766), .A2(n1138), .B1(n733), .B2(n1139), .ZN(n1701) );
  OAI22_X1 U736 ( .A1(n833), .A2(n1140), .B1(n800), .B2(n1141), .ZN(n1699) );
  OAI22_X1 U737 ( .A1(n901), .A2(n1142), .B1(n867), .B2(n1143), .ZN(n1698) );
  NOR4_X1 U738 ( .A1(n1703), .A2(n1704), .A3(n1705), .A4(n1706), .ZN(n1686) );
  OAI22_X1 U739 ( .A1(n968), .A2(n1148), .B1(n934), .B2(n1149), .ZN(n1706) );
  OAI22_X1 U740 ( .A1(n1035), .A2(n1151), .B1(n1001), .B2(n1152), .ZN(n1705)
         );
  OAI22_X1 U741 ( .A1(n59), .A2(n1153), .B1(n1069), .B2(n1154), .ZN(n1704) );
  OAI22_X1 U742 ( .A1(n149), .A2(n3), .B1(n114), .B2(n37), .ZN(n1703) );
  OAI22_X1 U743 ( .A1(n1707), .A2(n1102), .B1(n1103), .B2(n1700), .ZN(N4564)
         );
  NOR4_X1 U744 ( .A1(n1712), .A2(n1713), .A3(n1714), .A4(n1715), .ZN(n1711) );
  OAI22_X1 U745 ( .A1(n131), .A2(n1112), .B1(n543), .B2(n1113), .ZN(n1715) );
  OAI22_X1 U746 ( .A1(n237), .A2(n1114), .B1(n205), .B2(n1115), .ZN(n1714) );
  OAI22_X1 U747 ( .A1(n301), .A2(n1116), .B1(n269), .B2(n1117), .ZN(n1713) );
  OAI22_X1 U748 ( .A1(n365), .A2(n1118), .B1(n333), .B2(n1119), .ZN(n1712) );
  NOR4_X1 U749 ( .A1(n1716), .A2(n1717), .A3(n1718), .A4(n1719), .ZN(n1710) );
  OAI22_X1 U750 ( .A1(n429), .A2(n1124), .B1(n397), .B2(n1125), .ZN(n1719) );
  OAI22_X1 U751 ( .A1(n496), .A2(n1126), .B1(n463), .B2(n1127), .ZN(n1718) );
  OAI22_X1 U752 ( .A1(n563), .A2(n1128), .B1(n530), .B2(n1129), .ZN(n1717) );
  OAI22_X1 U753 ( .A1(n631), .A2(n1130), .B1(n597), .B2(n1131), .ZN(n1716) );
  NOR4_X1 U754 ( .A1(n1720), .A2(n1721), .A3(n1723), .A4(n1724), .ZN(n1709) );
  OAI22_X1 U755 ( .A1(n698), .A2(n1136), .B1(n664), .B2(n1137), .ZN(n1724) );
  OAI22_X1 U756 ( .A1(n765), .A2(n1138), .B1(n731), .B2(n1139), .ZN(n1723) );
  OAI22_X1 U757 ( .A1(n832), .A2(n1140), .B1(n799), .B2(n1141), .ZN(n1721) );
  OAI22_X1 U758 ( .A1(n899), .A2(n1142), .B1(n866), .B2(n1143), .ZN(n1720) );
  NOR4_X1 U759 ( .A1(n1725), .A2(n1726), .A3(n1727), .A4(n1728), .ZN(n1708) );
  OAI22_X1 U760 ( .A1(n967), .A2(n1148), .B1(n933), .B2(n1149), .ZN(n1728) );
  OAI22_X1 U761 ( .A1(n1034), .A2(n1151), .B1(n1000), .B2(n1152), .ZN(n1727)
         );
  OAI22_X1 U762 ( .A1(n57), .A2(n1153), .B1(n1067), .B2(n1154), .ZN(n1726) );
  OAI22_X1 U763 ( .A1(n148), .A2(n1155), .B1(n113), .B2(n1156), .ZN(n1725) );
  OAI22_X1 U764 ( .A1(n1729), .A2(n1102), .B1(n1103), .B2(n1722), .ZN(N4562)
         );
  NOR4_X1 U765 ( .A1(n1734), .A2(n1735), .A3(n1736), .A4(n1737), .ZN(n1733) );
  OAI22_X1 U766 ( .A1(n120), .A2(n1112), .B1(n522), .B2(n1113), .ZN(n1737) );
  OAI22_X1 U767 ( .A1(n236), .A2(n1114), .B1(n204), .B2(n1115), .ZN(n1736) );
  OAI22_X1 U768 ( .A1(n300), .A2(n1116), .B1(n268), .B2(n1117), .ZN(n1735) );
  OAI22_X1 U769 ( .A1(n364), .A2(n1118), .B1(n332), .B2(n1119), .ZN(n1734) );
  NOR4_X1 U770 ( .A1(n1738), .A2(n1739), .A3(n1740), .A4(n1741), .ZN(n1732) );
  OAI22_X1 U771 ( .A1(n428), .A2(n1124), .B1(n396), .B2(n1125), .ZN(n1741) );
  OAI22_X1 U772 ( .A1(n495), .A2(n1126), .B1(n462), .B2(n1127), .ZN(n1740) );
  OAI22_X1 U773 ( .A1(n562), .A2(n1128), .B1(n529), .B2(n1129), .ZN(n1739) );
  OAI22_X1 U774 ( .A1(n630), .A2(n1130), .B1(n596), .B2(n1131), .ZN(n1738) );
  NOR4_X1 U775 ( .A1(n1742), .A2(n1743), .A3(n1745), .A4(n1746), .ZN(n1731) );
  OAI22_X1 U776 ( .A1(n697), .A2(n1136), .B1(n663), .B2(n1137), .ZN(n1746) );
  OAI22_X1 U777 ( .A1(n764), .A2(n1138), .B1(n730), .B2(n1139), .ZN(n1745) );
  OAI22_X1 U778 ( .A1(n831), .A2(n1140), .B1(n798), .B2(n1141), .ZN(n1743) );
  OAI22_X1 U779 ( .A1(n898), .A2(n1142), .B1(n865), .B2(n1143), .ZN(n1742) );
  NOR4_X1 U780 ( .A1(n1747), .A2(n1748), .A3(n1749), .A4(n1750), .ZN(n1730) );
  OAI22_X1 U781 ( .A1(n966), .A2(n1148), .B1(n932), .B2(n1149), .ZN(n1750) );
  OAI22_X1 U782 ( .A1(n1033), .A2(n1151), .B1(n999), .B2(n1152), .ZN(n1749) );
  OAI22_X1 U783 ( .A1(n55), .A2(n1153), .B1(n1066), .B2(n1154), .ZN(n1748) );
  OAI22_X1 U784 ( .A1(n147), .A2(n1155), .B1(n112), .B2(n1156), .ZN(n1747) );
  OAI22_X1 U785 ( .A1(n1751), .A2(n1102), .B1(n1744), .B2(n1103), .ZN(N4560)
         );
  NOR4_X1 U786 ( .A1(n1752), .A2(n1753), .A3(n1754), .A4(n1755), .ZN(n1751) );
  OAI211_X1 U787 ( .C1(n1100), .C2(n1153), .A(n1756), .B(n1757), .ZN(n1755) );
  NOR4_X1 U788 ( .A1(n1758), .A2(n1759), .A3(n1760), .A4(n1761), .ZN(n1757) );
  OAI22_X1 U789 ( .A1(n109), .A2(n1112), .B1(n203), .B2(n1115), .ZN(n1761) );
  OAI22_X1 U790 ( .A1(n235), .A2(n1114), .B1(n267), .B2(n1117), .ZN(n1760) );
  OAI22_X1 U791 ( .A1(n299), .A2(n1116), .B1(n331), .B2(n1119), .ZN(n1759) );
  OAI22_X1 U792 ( .A1(n363), .A2(n1118), .B1(n395), .B2(n1125), .ZN(n1758) );
  NOR4_X1 U793 ( .A1(n1762), .A2(n1763), .A3(n1764), .A4(n1765), .ZN(n1756) );
  OAI22_X1 U794 ( .A1(n427), .A2(n1124), .B1(n461), .B2(n1127), .ZN(n1765) );
  OAI22_X1 U795 ( .A1(n494), .A2(n1126), .B1(n528), .B2(n1129), .ZN(n1764) );
  OAI22_X1 U796 ( .A1(n561), .A2(n1128), .B1(n595), .B2(n1131), .ZN(n1763) );
  OAI22_X1 U797 ( .A1(n629), .A2(n1130), .B1(n662), .B2(n1137), .ZN(n1762) );
  OAI211_X1 U798 ( .C1(n146), .C2(n1155), .A(n1767), .B(n1768), .ZN(n1754) );
  NOR4_X1 U799 ( .A1(n1769), .A2(n1770), .A3(n1771), .A4(n1772), .ZN(n1768) );
  OAI22_X1 U800 ( .A1(n763), .A2(n1138), .B1(n797), .B2(n1141), .ZN(n1772) );
  OAI22_X1 U801 ( .A1(n696), .A2(n1136), .B1(n729), .B2(n1139), .ZN(n1771) );
  OAI22_X1 U802 ( .A1(n897), .A2(n1142), .B1(n931), .B2(n1149), .ZN(n1770) );
  OAI22_X1 U803 ( .A1(n830), .A2(n1140), .B1(n864), .B2(n1143), .ZN(n1769) );
  OAI22_X1 U804 ( .A1(n1113), .A2(n501), .B1(n37), .B2(n111), .ZN(n1773) );
  OAI22_X1 U805 ( .A1(n1032), .A2(n1151), .B1(n1065), .B2(n1154), .ZN(n1753)
         );
  OAI22_X1 U806 ( .A1(n965), .A2(n1148), .B1(n998), .B2(n1152), .ZN(n1752) );
  OAI22_X1 U807 ( .A1(n1774), .A2(n1102), .B1(n1103), .B2(n1766), .ZN(N4558)
         );
  NOR4_X1 U808 ( .A1(n1779), .A2(n1780), .A3(n1781), .A4(n1782), .ZN(n1778) );
  OAI22_X1 U809 ( .A1(n97), .A2(n1112), .B1(n480), .B2(n1113), .ZN(n1782) );
  OAI22_X1 U810 ( .A1(n234), .A2(n1114), .B1(n202), .B2(n1115), .ZN(n1781) );
  OAI22_X1 U811 ( .A1(n298), .A2(n1116), .B1(n266), .B2(n1117), .ZN(n1780) );
  OAI22_X1 U812 ( .A1(n362), .A2(n1118), .B1(n330), .B2(n1119), .ZN(n1779) );
  NOR4_X1 U813 ( .A1(n1783), .A2(n1784), .A3(n1785), .A4(n1786), .ZN(n1777) );
  OAI22_X1 U814 ( .A1(n426), .A2(n1124), .B1(n394), .B2(n1125), .ZN(n1786) );
  OAI22_X1 U815 ( .A1(n493), .A2(n1126), .B1(n460), .B2(n1127), .ZN(n1785) );
  OAI22_X1 U816 ( .A1(n560), .A2(n1128), .B1(n527), .B2(n1129), .ZN(n1784) );
  OAI22_X1 U817 ( .A1(n628), .A2(n1130), .B1(n594), .B2(n1131), .ZN(n1783) );
  NOR4_X1 U818 ( .A1(n1787), .A2(n1789), .A3(n1790), .A4(n1791), .ZN(n1776) );
  OAI22_X1 U819 ( .A1(n695), .A2(n1136), .B1(n661), .B2(n1137), .ZN(n1791) );
  OAI22_X1 U820 ( .A1(n762), .A2(n1138), .B1(n728), .B2(n1139), .ZN(n1790) );
  OAI22_X1 U821 ( .A1(n829), .A2(n1140), .B1(n796), .B2(n1141), .ZN(n1789) );
  OAI22_X1 U822 ( .A1(n896), .A2(n1142), .B1(n863), .B2(n1143), .ZN(n1787) );
  NOR4_X1 U823 ( .A1(n1792), .A2(n1793), .A3(n1794), .A4(n1795), .ZN(n1775) );
  OAI22_X1 U824 ( .A1(n964), .A2(n1148), .B1(n930), .B2(n1149), .ZN(n1795) );
  OAI22_X1 U825 ( .A1(n1031), .A2(n1151), .B1(n997), .B2(n1152), .ZN(n1794) );
  OAI22_X1 U826 ( .A1(n1099), .A2(n1153), .B1(n1064), .B2(n1154), .ZN(n1793)
         );
  OAI22_X1 U827 ( .A1(n145), .A2(n1155), .B1(n110), .B2(n1156), .ZN(n1792) );
  OAI22_X1 U828 ( .A1(n1796), .A2(n1102), .B1(n1103), .B2(n1788), .ZN(N4556)
         );
  NOR4_X1 U829 ( .A1(n1801), .A2(n1802), .A3(n1803), .A4(n1804), .ZN(n1800) );
  OAI22_X1 U830 ( .A1(n75), .A2(n1112), .B1(n459), .B2(n1113), .ZN(n1804) );
  OAI22_X1 U831 ( .A1(n233), .A2(n1114), .B1(n201), .B2(n1115), .ZN(n1803) );
  OAI22_X1 U832 ( .A1(n297), .A2(n1116), .B1(n265), .B2(n1117), .ZN(n1802) );
  OAI22_X1 U833 ( .A1(n361), .A2(n1118), .B1(n329), .B2(n1119), .ZN(n1801) );
  NOR4_X1 U834 ( .A1(n1805), .A2(n1806), .A3(n1807), .A4(n1808), .ZN(n1799) );
  OAI22_X1 U835 ( .A1(n425), .A2(n1124), .B1(n393), .B2(n1125), .ZN(n1808) );
  OAI22_X1 U836 ( .A1(n492), .A2(n1126), .B1(n458), .B2(n1127), .ZN(n1807) );
  OAI22_X1 U837 ( .A1(n559), .A2(n1128), .B1(n526), .B2(n1129), .ZN(n1806) );
  OAI22_X1 U838 ( .A1(n626), .A2(n1130), .B1(n593), .B2(n1131), .ZN(n1805) );
  NOR4_X1 U839 ( .A1(n1809), .A2(n1811), .A3(n1812), .A4(n1813), .ZN(n1798) );
  OAI22_X1 U840 ( .A1(n694), .A2(n1136), .B1(n660), .B2(n1137), .ZN(n1813) );
  OAI22_X1 U841 ( .A1(n761), .A2(n1138), .B1(n727), .B2(n1139), .ZN(n1812) );
  OAI22_X1 U842 ( .A1(n828), .A2(n1140), .B1(n794), .B2(n1141), .ZN(n1811) );
  OAI22_X1 U843 ( .A1(n895), .A2(n1142), .B1(n862), .B2(n1143), .ZN(n1809) );
  NOR4_X1 U844 ( .A1(n1814), .A2(n1815), .A3(n1816), .A4(n1817), .ZN(n1797) );
  OAI22_X1 U845 ( .A1(n962), .A2(n1148), .B1(n929), .B2(n1149), .ZN(n1817) );
  OAI22_X1 U846 ( .A1(n1030), .A2(n1151), .B1(n996), .B2(n1152), .ZN(n1816) );
  OAI22_X1 U847 ( .A1(n1098), .A2(n1153), .B1(n1063), .B2(n1154), .ZN(n1815)
         );
  OAI22_X1 U848 ( .A1(n144), .A2(n1155), .B1(n108), .B2(n1156), .ZN(n1814) );
  OAI22_X1 U849 ( .A1(n1818), .A2(n1102), .B1(n1103), .B2(n1810), .ZN(N4554)
         );
  AOI221_X1 U850 ( .B1(ADD_WR[1]), .B2(n1822), .C1(n1823), .C2(ADD_RD2[1]), 
        .A(n1824), .ZN(n1821) );
  OAI221_X1 U851 ( .B1(n1825), .B2(ADD_RD2[2]), .C1(n1826), .C2(ADD_RD2[0]), 
        .A(n1827), .ZN(n1824) );
  AOI22_X1 U852 ( .A1(n1825), .A2(ADD_RD2[2]), .B1(n1826), .B2(ADD_RD2[0]), 
        .ZN(n1827) );
  AOI221_X1 U853 ( .B1(n1828), .B2(ADD_WR[4]), .C1(n1829), .C2(ADD_RD2[3]), 
        .A(n1830), .ZN(n1820) );
  OAI22_X1 U854 ( .A1(ADD_WR[4]), .A2(n1828), .B1(n1829), .B2(ADD_RD2[3]), 
        .ZN(n1830) );
  NOR4_X1 U855 ( .A1(n1835), .A2(n1836), .A3(n1837), .A4(n1838), .ZN(n1834) );
  OAI22_X1 U856 ( .A1(n53), .A2(n1112), .B1(n438), .B2(n1113), .ZN(n1838) );
  OAI22_X1 U857 ( .A1(n232), .A2(n1114), .B1(n200), .B2(n1115), .ZN(n1837) );
  OAI22_X1 U858 ( .A1(n296), .A2(n1116), .B1(n264), .B2(n1117), .ZN(n1836) );
  OAI22_X1 U859 ( .A1(n360), .A2(n1118), .B1(n328), .B2(n1119), .ZN(n1835) );
  NOR3_X1 U860 ( .A1(n1828), .A2(n1845), .A3(n1846), .ZN(n1840) );
  NAND2_X1 U861 ( .A1(ADD_RD2[4]), .A2(ADD_RD2[3]), .ZN(n1847) );
  NOR4_X1 U862 ( .A1(n1848), .A2(n1849), .A3(n1850), .A4(n1851), .ZN(n1833) );
  OAI22_X1 U863 ( .A1(n424), .A2(n1124), .B1(n392), .B2(n1125), .ZN(n1851) );
  OAI22_X1 U864 ( .A1(n491), .A2(n1126), .B1(n457), .B2(n1127), .ZN(n1850) );
  OAI22_X1 U865 ( .A1(n558), .A2(n1128), .B1(n525), .B2(n1129), .ZN(n1849) );
  OAI22_X1 U866 ( .A1(n625), .A2(n1130), .B1(n592), .B2(n1131), .ZN(n1848) );
  NOR3_X1 U867 ( .A1(ADD_RD2[3]), .A2(n1828), .A3(n1846), .ZN(n1852) );
  NOR3_X1 U868 ( .A1(ADD_RD2[3]), .A2(ADD_RD2[0]), .A3(n1828), .ZN(n1853) );
  NOR4_X1 U869 ( .A1(n1854), .A2(n1855), .A3(n1856), .A4(n1857), .ZN(n1832) );
  OAI22_X1 U870 ( .A1(n693), .A2(n1136), .B1(n659), .B2(n1137), .ZN(n1857) );
  OAI22_X1 U871 ( .A1(n760), .A2(n1138), .B1(n726), .B2(n1139), .ZN(n1856) );
  OAI22_X1 U872 ( .A1(n827), .A2(n1140), .B1(n793), .B2(n1141), .ZN(n1855) );
  OAI22_X1 U873 ( .A1(n894), .A2(n1142), .B1(n861), .B2(n1143), .ZN(n1854) );
  NOR3_X1 U874 ( .A1(ADD_RD2[4]), .A2(n1845), .A3(n1846), .ZN(n1858) );
  NOR3_X1 U875 ( .A1(ADD_RD2[4]), .A2(ADD_RD2[0]), .A3(n1845), .ZN(n1859) );
  NOR4_X1 U876 ( .A1(n1860), .A2(n1861), .A3(n1862), .A4(n1863), .ZN(n1831) );
  OAI22_X1 U877 ( .A1(n961), .A2(n1148), .B1(n928), .B2(n1149), .ZN(n1863) );
  OAI22_X1 U878 ( .A1(n1029), .A2(n1151), .B1(n995), .B2(n1152), .ZN(n1862) );
  OAI22_X1 U879 ( .A1(n1097), .A2(n1153), .B1(n1062), .B2(n1154), .ZN(n1861)
         );
  NAND2_X1 U880 ( .A1(n1843), .A2(n1864), .ZN(n1154) );
  NAND2_X1 U881 ( .A1(n1865), .A2(n1843), .ZN(n1153) );
  OAI22_X1 U882 ( .A1(n143), .A2(n3), .B1(n107), .B2(n37), .ZN(n1860) );
  NAND2_X1 U883 ( .A1(n1844), .A2(n1864), .ZN(n1156) );
  NOR3_X1 U884 ( .A1(ADD_RD2[4]), .A2(ADD_RD2[3]), .A3(n1846), .ZN(n1864) );
  NAND2_X1 U885 ( .A1(n1865), .A2(n1844), .ZN(n1155) );
  NOR3_X1 U886 ( .A1(ADD_RD2[4]), .A2(ADD_RD2[3]), .A3(ADD_RD2[0]), .ZN(n1865)
         );
  OAI22_X1 U887 ( .A1(n1866), .A2(n1867), .B1(n1868), .B2(n1094), .ZN(N4552)
         );
  NOR4_X1 U888 ( .A1(n1873), .A2(n1874), .A3(n1875), .A4(n1876), .ZN(n1872) );
  OAI22_X1 U889 ( .A1(n199), .A2(n1877), .B1(n1089), .B2(n1878), .ZN(n1876) );
  OAI22_X1 U890 ( .A1(n263), .A2(n1879), .B1(n231), .B2(n1880), .ZN(n1875) );
  OAI22_X1 U891 ( .A1(n327), .A2(n1881), .B1(n295), .B2(n1882), .ZN(n1874) );
  OAI22_X1 U892 ( .A1(n391), .A2(n1883), .B1(n359), .B2(n1884), .ZN(n1873) );
  NOR4_X1 U893 ( .A1(n1885), .A2(n1886), .A3(n1887), .A4(n1888), .ZN(n1871) );
  OAI22_X1 U894 ( .A1(n456), .A2(n1889), .B1(n423), .B2(n1890), .ZN(n1888) );
  OAI22_X1 U895 ( .A1(n524), .A2(n1891), .B1(n490), .B2(n1892), .ZN(n1887) );
  OAI22_X1 U896 ( .A1(n591), .A2(n1893), .B1(n557), .B2(n1894), .ZN(n1886) );
  OAI22_X1 U897 ( .A1(n658), .A2(n1895), .B1(n624), .B2(n1896), .ZN(n1885) );
  NOR4_X1 U898 ( .A1(n1897), .A2(n1898), .A3(n1899), .A4(n1900), .ZN(n1870) );
  OAI22_X1 U899 ( .A1(n725), .A2(n1901), .B1(n692), .B2(n1902), .ZN(n1900) );
  OAI22_X1 U900 ( .A1(n792), .A2(n1903), .B1(n759), .B2(n1904), .ZN(n1899) );
  OAI22_X1 U901 ( .A1(n860), .A2(n1905), .B1(n826), .B2(n1906), .ZN(n1898) );
  OAI22_X1 U902 ( .A1(n927), .A2(n1907), .B1(n893), .B2(n1908), .ZN(n1897) );
  NOR4_X1 U903 ( .A1(n1909), .A2(n1910), .A3(n1911), .A4(n1912), .ZN(n1869) );
  OAI22_X1 U904 ( .A1(n994), .A2(n1913), .B1(n960), .B2(n1914), .ZN(n1912) );
  OAI22_X1 U905 ( .A1(n1061), .A2(n1915), .B1(n1028), .B2(n1916), .ZN(n1911)
         );
  OAI22_X1 U906 ( .A1(n106), .A2(n41), .B1(n1096), .B2(n1918), .ZN(n1910) );
  OAI22_X1 U907 ( .A1(n177), .A2(n1919), .B1(n141), .B2(n1920), .ZN(n1909) );
  OAI22_X1 U908 ( .A1(n1921), .A2(n1867), .B1(n1868), .B2(n1150), .ZN(N4550)
         );
  NOR4_X1 U909 ( .A1(n1926), .A2(n1927), .A3(n1928), .A4(n1929), .ZN(n1925) );
  OAI22_X1 U910 ( .A1(n198), .A2(n1877), .B1(n1068), .B2(n1878), .ZN(n1929) );
  OAI22_X1 U911 ( .A1(n262), .A2(n1879), .B1(n230), .B2(n1880), .ZN(n1928) );
  OAI22_X1 U912 ( .A1(n326), .A2(n1881), .B1(n294), .B2(n1882), .ZN(n1927) );
  OAI22_X1 U913 ( .A1(n390), .A2(n39), .B1(n358), .B2(n1884), .ZN(n1926) );
  NOR4_X1 U914 ( .A1(n1930), .A2(n1931), .A3(n1932), .A4(n1933), .ZN(n1924) );
  OAI22_X1 U915 ( .A1(n455), .A2(n1889), .B1(n422), .B2(n1890), .ZN(n1933) );
  OAI22_X1 U916 ( .A1(n523), .A2(n1891), .B1(n489), .B2(n1892), .ZN(n1932) );
  OAI22_X1 U917 ( .A1(n590), .A2(n1893), .B1(n556), .B2(n1894), .ZN(n1931) );
  OAI22_X1 U918 ( .A1(n657), .A2(n1895), .B1(n623), .B2(n1896), .ZN(n1930) );
  NOR4_X1 U919 ( .A1(n1934), .A2(n1935), .A3(n1936), .A4(n1937), .ZN(n1923) );
  OAI22_X1 U920 ( .A1(n724), .A2(n1901), .B1(n691), .B2(n1902), .ZN(n1937) );
  OAI22_X1 U921 ( .A1(n791), .A2(n1903), .B1(n758), .B2(n1904), .ZN(n1936) );
  OAI22_X1 U922 ( .A1(n859), .A2(n1905), .B1(n825), .B2(n1906), .ZN(n1935) );
  OAI22_X1 U923 ( .A1(n926), .A2(n1907), .B1(n892), .B2(n1908), .ZN(n1934) );
  NOR4_X1 U924 ( .A1(n1938), .A2(n1939), .A3(n1940), .A4(n1941), .ZN(n1922) );
  OAI22_X1 U925 ( .A1(n993), .A2(n1913), .B1(n959), .B2(n1914), .ZN(n1941) );
  OAI22_X1 U926 ( .A1(n1060), .A2(n1915), .B1(n1027), .B2(n1916), .ZN(n1940)
         );
  OAI22_X1 U927 ( .A1(n105), .A2(n1917), .B1(n1095), .B2(n1918), .ZN(n1939) );
  OAI22_X1 U928 ( .A1(n176), .A2(n45), .B1(n140), .B2(n1920), .ZN(n1938) );
  OAI22_X1 U929 ( .A1(n1942), .A2(n1867), .B1(n1868), .B2(n1172), .ZN(N4548)
         );
  NOR4_X1 U930 ( .A1(n1947), .A2(n1948), .A3(n1949), .A4(n1950), .ZN(n1946) );
  OAI22_X1 U931 ( .A1(n197), .A2(n1877), .B1(n1047), .B2(n1878), .ZN(n1950) );
  OAI22_X1 U932 ( .A1(n261), .A2(n1879), .B1(n229), .B2(n1880), .ZN(n1949) );
  OAI22_X1 U933 ( .A1(n325), .A2(n1881), .B1(n293), .B2(n1882), .ZN(n1948) );
  OAI22_X1 U934 ( .A1(n389), .A2(n1883), .B1(n357), .B2(n1884), .ZN(n1947) );
  NOR4_X1 U935 ( .A1(n1951), .A2(n1952), .A3(n1953), .A4(n1954), .ZN(n1945) );
  OAI22_X1 U936 ( .A1(n454), .A2(n1889), .B1(n421), .B2(n1890), .ZN(n1954) );
  OAI22_X1 U937 ( .A1(n521), .A2(n1891), .B1(n488), .B2(n1892), .ZN(n1953) );
  OAI22_X1 U938 ( .A1(n589), .A2(n1893), .B1(n555), .B2(n1894), .ZN(n1952) );
  OAI22_X1 U939 ( .A1(n656), .A2(n1895), .B1(n622), .B2(n1896), .ZN(n1951) );
  NOR4_X1 U940 ( .A1(n1955), .A2(n1956), .A3(n1957), .A4(n1958), .ZN(n1944) );
  OAI22_X1 U941 ( .A1(n723), .A2(n1901), .B1(n689), .B2(n1902), .ZN(n1958) );
  OAI22_X1 U942 ( .A1(n790), .A2(n1903), .B1(n757), .B2(n1904), .ZN(n1957) );
  OAI22_X1 U943 ( .A1(n857), .A2(n1905), .B1(n824), .B2(n1906), .ZN(n1956) );
  OAI22_X1 U944 ( .A1(n925), .A2(n1907), .B1(n891), .B2(n1908), .ZN(n1955) );
  NOR4_X1 U945 ( .A1(n1959), .A2(n1960), .A3(n1961), .A4(n1962), .ZN(n1943) );
  OAI22_X1 U946 ( .A1(n992), .A2(n1913), .B1(n958), .B2(n1914), .ZN(n1962) );
  OAI22_X1 U947 ( .A1(n1059), .A2(n1915), .B1(n1025), .B2(n1916), .ZN(n1961)
         );
  OAI22_X1 U948 ( .A1(n104), .A2(n1917), .B1(n1093), .B2(n1918), .ZN(n1960) );
  OAI22_X1 U949 ( .A1(n174), .A2(n45), .B1(n139), .B2(n1920), .ZN(n1959) );
  OAI22_X1 U950 ( .A1(n1963), .A2(n1867), .B1(n1868), .B2(n1194), .ZN(N4546)
         );
  NOR4_X1 U951 ( .A1(n1968), .A2(n1969), .A3(n1970), .A4(n1971), .ZN(n1967) );
  OAI22_X1 U952 ( .A1(n196), .A2(n1877), .B1(n1026), .B2(n1878), .ZN(n1971) );
  OAI22_X1 U953 ( .A1(n260), .A2(n1879), .B1(n228), .B2(n1880), .ZN(n1970) );
  OAI22_X1 U954 ( .A1(n324), .A2(n1881), .B1(n292), .B2(n1882), .ZN(n1969) );
  OAI22_X1 U955 ( .A1(n388), .A2(n1883), .B1(n356), .B2(n1884), .ZN(n1968) );
  NOR4_X1 U956 ( .A1(n1972), .A2(n1973), .A3(n1974), .A4(n1975), .ZN(n1966) );
  OAI22_X1 U957 ( .A1(n453), .A2(n1889), .B1(n420), .B2(n1890), .ZN(n1975) );
  OAI22_X1 U958 ( .A1(n520), .A2(n1891), .B1(n487), .B2(n1892), .ZN(n1974) );
  OAI22_X1 U959 ( .A1(n588), .A2(n1893), .B1(n554), .B2(n1894), .ZN(n1973) );
  OAI22_X1 U960 ( .A1(n655), .A2(n1895), .B1(n621), .B2(n1896), .ZN(n1972) );
  NOR4_X1 U961 ( .A1(n1976), .A2(n1977), .A3(n1978), .A4(n1979), .ZN(n1965) );
  OAI22_X1 U962 ( .A1(n722), .A2(n1901), .B1(n688), .B2(n1902), .ZN(n1979) );
  OAI22_X1 U963 ( .A1(n789), .A2(n1903), .B1(n756), .B2(n1904), .ZN(n1978) );
  OAI22_X1 U964 ( .A1(n856), .A2(n1905), .B1(n823), .B2(n1906), .ZN(n1977) );
  OAI22_X1 U965 ( .A1(n924), .A2(n1907), .B1(n890), .B2(n1908), .ZN(n1976) );
  NOR4_X1 U966 ( .A1(n1980), .A2(n1981), .A3(n1982), .A4(n1983), .ZN(n1964) );
  OAI22_X1 U967 ( .A1(n991), .A2(n1913), .B1(n957), .B2(n1914), .ZN(n1983) );
  OAI22_X1 U968 ( .A1(n1058), .A2(n1915), .B1(n1024), .B2(n1916), .ZN(n1982)
         );
  OAI22_X1 U969 ( .A1(n103), .A2(n1917), .B1(n1092), .B2(n43), .ZN(n1981) );
  OAI22_X1 U970 ( .A1(n173), .A2(n45), .B1(n138), .B2(n1920), .ZN(n1980) );
  OAI22_X1 U971 ( .A1(n1984), .A2(n1867), .B1(n1868), .B2(n1216), .ZN(N4544)
         );
  NOR4_X1 U972 ( .A1(n1989), .A2(n1990), .A3(n1991), .A4(n1992), .ZN(n1988) );
  OAI22_X1 U973 ( .A1(n195), .A2(n1877), .B1(n1005), .B2(n1878), .ZN(n1992) );
  OAI22_X1 U974 ( .A1(n259), .A2(n1879), .B1(n227), .B2(n1880), .ZN(n1991) );
  OAI22_X1 U975 ( .A1(n323), .A2(n1881), .B1(n291), .B2(n1882), .ZN(n1990) );
  OAI22_X1 U976 ( .A1(n387), .A2(n1883), .B1(n355), .B2(n1884), .ZN(n1989) );
  NOR4_X1 U977 ( .A1(n1993), .A2(n1994), .A3(n1995), .A4(n1996), .ZN(n1987) );
  OAI22_X1 U978 ( .A1(n452), .A2(n1889), .B1(n419), .B2(n1890), .ZN(n1996) );
  OAI22_X1 U979 ( .A1(n519), .A2(n1891), .B1(n486), .B2(n1892), .ZN(n1995) );
  OAI22_X1 U980 ( .A1(n587), .A2(n1893), .B1(n553), .B2(n1894), .ZN(n1994) );
  OAI22_X1 U981 ( .A1(n654), .A2(n1895), .B1(n620), .B2(n1896), .ZN(n1993) );
  NOR4_X1 U982 ( .A1(n1997), .A2(n1998), .A3(n1999), .A4(n2000), .ZN(n1986) );
  OAI22_X1 U983 ( .A1(n721), .A2(n1901), .B1(n687), .B2(n1902), .ZN(n2000) );
  OAI22_X1 U984 ( .A1(n788), .A2(n1903), .B1(n755), .B2(n1904), .ZN(n1999) );
  OAI22_X1 U985 ( .A1(n855), .A2(n1905), .B1(n822), .B2(n1906), .ZN(n1998) );
  OAI22_X1 U986 ( .A1(n923), .A2(n1907), .B1(n889), .B2(n1908), .ZN(n1997) );
  NOR4_X1 U987 ( .A1(n2001), .A2(n2002), .A3(n2003), .A4(n2004), .ZN(n1985) );
  OAI22_X1 U988 ( .A1(n990), .A2(n1913), .B1(n956), .B2(n1914), .ZN(n2004) );
  OAI22_X1 U989 ( .A1(n1057), .A2(n1915), .B1(n1023), .B2(n1916), .ZN(n2003)
         );
  OAI22_X1 U990 ( .A1(n102), .A2(n1917), .B1(n1091), .B2(n43), .ZN(n2002) );
  OAI22_X1 U991 ( .A1(n172), .A2(n45), .B1(n137), .B2(n1920), .ZN(n2001) );
  OAI22_X1 U992 ( .A1(n2005), .A2(n1867), .B1(n1868), .B2(n1238), .ZN(N4542)
         );
  NOR4_X1 U993 ( .A1(n2010), .A2(n2011), .A3(n2012), .A4(n2013), .ZN(n2009) );
  OAI22_X1 U994 ( .A1(n194), .A2(n1877), .B1(n984), .B2(n1878), .ZN(n2013) );
  OAI22_X1 U995 ( .A1(n258), .A2(n1879), .B1(n226), .B2(n1880), .ZN(n2012) );
  OAI22_X1 U996 ( .A1(n322), .A2(n1881), .B1(n290), .B2(n1882), .ZN(n2011) );
  OAI22_X1 U997 ( .A1(n386), .A2(n1883), .B1(n354), .B2(n1884), .ZN(n2010) );
  NOR4_X1 U998 ( .A1(n2014), .A2(n2015), .A3(n2016), .A4(n2017), .ZN(n2008) );
  OAI22_X1 U999 ( .A1(n451), .A2(n1889), .B1(n418), .B2(n1890), .ZN(n2017) );
  OAI22_X1 U1000 ( .A1(n518), .A2(n1891), .B1(n485), .B2(n1892), .ZN(n2016) );
  OAI22_X1 U1001 ( .A1(n586), .A2(n1893), .B1(n552), .B2(n1894), .ZN(n2015) );
  OAI22_X1 U1002 ( .A1(n653), .A2(n1895), .B1(n619), .B2(n1896), .ZN(n2014) );
  NOR4_X1 U1003 ( .A1(n2018), .A2(n2019), .A3(n2020), .A4(n2021), .ZN(n2007)
         );
  OAI22_X1 U1004 ( .A1(n720), .A2(n1901), .B1(n686), .B2(n1902), .ZN(n2021) );
  OAI22_X1 U1005 ( .A1(n787), .A2(n1903), .B1(n754), .B2(n1904), .ZN(n2020) );
  OAI22_X1 U1006 ( .A1(n854), .A2(n1905), .B1(n821), .B2(n1906), .ZN(n2019) );
  OAI22_X1 U1007 ( .A1(n922), .A2(n1907), .B1(n888), .B2(n1908), .ZN(n2018) );
  NOR4_X1 U1008 ( .A1(n2022), .A2(n2023), .A3(n2024), .A4(n2025), .ZN(n2006)
         );
  OAI22_X1 U1009 ( .A1(n989), .A2(n1913), .B1(n955), .B2(n1914), .ZN(n2025) );
  OAI22_X1 U1010 ( .A1(n1056), .A2(n1915), .B1(n1022), .B2(n1916), .ZN(n2024)
         );
  OAI22_X1 U1011 ( .A1(n101), .A2(n1917), .B1(n1090), .B2(n1918), .ZN(n2023)
         );
  OAI22_X1 U1012 ( .A1(n171), .A2(n45), .B1(n136), .B2(n1920), .ZN(n2022) );
  OAI22_X1 U1013 ( .A1(n2026), .A2(n1867), .B1(n1868), .B2(n1260), .ZN(N4540)
         );
  NOR4_X1 U1014 ( .A1(n2031), .A2(n2032), .A3(n2033), .A4(n2034), .ZN(n2030)
         );
  OAI22_X1 U1015 ( .A1(n193), .A2(n1877), .B1(n963), .B2(n1878), .ZN(n2034) );
  OAI22_X1 U1016 ( .A1(n257), .A2(n1879), .B1(n225), .B2(n1880), .ZN(n2033) );
  OAI22_X1 U1017 ( .A1(n321), .A2(n1881), .B1(n289), .B2(n1882), .ZN(n2032) );
  OAI22_X1 U1018 ( .A1(n385), .A2(n1883), .B1(n353), .B2(n1884), .ZN(n2031) );
  NOR4_X1 U1019 ( .A1(n2035), .A2(n2036), .A3(n2037), .A4(n2038), .ZN(n2029)
         );
  OAI22_X1 U1020 ( .A1(n450), .A2(n1889), .B1(n417), .B2(n1890), .ZN(n2038) );
  OAI22_X1 U1021 ( .A1(n517), .A2(n1891), .B1(n484), .B2(n1892), .ZN(n2037) );
  OAI22_X1 U1022 ( .A1(n584), .A2(n1893), .B1(n551), .B2(n1894), .ZN(n2036) );
  OAI22_X1 U1023 ( .A1(n652), .A2(n1895), .B1(n618), .B2(n1896), .ZN(n2035) );
  NOR4_X1 U1024 ( .A1(n2039), .A2(n2040), .A3(n2041), .A4(n2042), .ZN(n2028)
         );
  OAI22_X1 U1025 ( .A1(n719), .A2(n1901), .B1(n685), .B2(n1902), .ZN(n2042) );
  OAI22_X1 U1026 ( .A1(n786), .A2(n1903), .B1(n752), .B2(n1904), .ZN(n2041) );
  OAI22_X1 U1027 ( .A1(n853), .A2(n1905), .B1(n820), .B2(n1906), .ZN(n2040) );
  OAI22_X1 U1028 ( .A1(n920), .A2(n1907), .B1(n887), .B2(n1908), .ZN(n2039) );
  NOR4_X1 U1029 ( .A1(n2043), .A2(n2044), .A3(n2045), .A4(n2046), .ZN(n2027)
         );
  OAI22_X1 U1030 ( .A1(n988), .A2(n1913), .B1(n954), .B2(n1914), .ZN(n2046) );
  OAI22_X1 U1031 ( .A1(n1055), .A2(n1915), .B1(n1021), .B2(n1916), .ZN(n2045)
         );
  OAI22_X1 U1032 ( .A1(n100), .A2(n1917), .B1(n1088), .B2(n43), .ZN(n2044) );
  OAI22_X1 U1033 ( .A1(n170), .A2(n45), .B1(n135), .B2(n1920), .ZN(n2043) );
  OAI22_X1 U1034 ( .A1(n2047), .A2(n1867), .B1(n1868), .B2(n1282), .ZN(N4538)
         );
  NOR4_X1 U1035 ( .A1(n2052), .A2(n2053), .A3(n2054), .A4(n2055), .ZN(n2051)
         );
  OAI22_X1 U1036 ( .A1(n192), .A2(n1877), .B1(n942), .B2(n1878), .ZN(n2055) );
  OAI22_X1 U1037 ( .A1(n256), .A2(n1879), .B1(n224), .B2(n1880), .ZN(n2054) );
  OAI22_X1 U1038 ( .A1(n320), .A2(n1881), .B1(n288), .B2(n1882), .ZN(n2053) );
  OAI22_X1 U1039 ( .A1(n384), .A2(n1883), .B1(n352), .B2(n1884), .ZN(n2052) );
  NOR4_X1 U1040 ( .A1(n2056), .A2(n2057), .A3(n2058), .A4(n2059), .ZN(n2050)
         );
  OAI22_X1 U1041 ( .A1(n449), .A2(n1889), .B1(n416), .B2(n1890), .ZN(n2059) );
  OAI22_X1 U1042 ( .A1(n516), .A2(n1891), .B1(n483), .B2(n1892), .ZN(n2058) );
  OAI22_X1 U1043 ( .A1(n583), .A2(n1893), .B1(n550), .B2(n1894), .ZN(n2057) );
  OAI22_X1 U1044 ( .A1(n651), .A2(n1895), .B1(n617), .B2(n1896), .ZN(n2056) );
  NOR4_X1 U1045 ( .A1(n2060), .A2(n2061), .A3(n2062), .A4(n2063), .ZN(n2049)
         );
  OAI22_X1 U1046 ( .A1(n718), .A2(n1901), .B1(n684), .B2(n1902), .ZN(n2063) );
  OAI22_X1 U1047 ( .A1(n785), .A2(n1903), .B1(n751), .B2(n1904), .ZN(n2062) );
  OAI22_X1 U1048 ( .A1(n852), .A2(n1905), .B1(n819), .B2(n1906), .ZN(n2061) );
  OAI22_X1 U1049 ( .A1(n919), .A2(n1907), .B1(n886), .B2(n1908), .ZN(n2060) );
  NOR4_X1 U1050 ( .A1(n2064), .A2(n2065), .A3(n2066), .A4(n2067), .ZN(n2048)
         );
  OAI22_X1 U1051 ( .A1(n987), .A2(n1913), .B1(n953), .B2(n1914), .ZN(n2067) );
  OAI22_X1 U1052 ( .A1(n1054), .A2(n1915), .B1(n1020), .B2(n1916), .ZN(n2066)
         );
  OAI22_X1 U1053 ( .A1(n99), .A2(n1917), .B1(n1087), .B2(n1918), .ZN(n2065) );
  OAI22_X1 U1054 ( .A1(n169), .A2(n45), .B1(n134), .B2(n1920), .ZN(n2064) );
  OAI22_X1 U1055 ( .A1(n2068), .A2(n1867), .B1(n1868), .B2(n1304), .ZN(N4536)
         );
  NOR4_X1 U1056 ( .A1(n2073), .A2(n2074), .A3(n2075), .A4(n2076), .ZN(n2072)
         );
  OAI22_X1 U1057 ( .A1(n191), .A2(n1877), .B1(n921), .B2(n1878), .ZN(n2076) );
  OAI22_X1 U1058 ( .A1(n255), .A2(n1879), .B1(n223), .B2(n1880), .ZN(n2075) );
  OAI22_X1 U1059 ( .A1(n319), .A2(n1881), .B1(n287), .B2(n1882), .ZN(n2074) );
  OAI22_X1 U1060 ( .A1(n383), .A2(n1883), .B1(n351), .B2(n1884), .ZN(n2073) );
  NOR4_X1 U1061 ( .A1(n2077), .A2(n2078), .A3(n2079), .A4(n2080), .ZN(n2071)
         );
  OAI22_X1 U1062 ( .A1(n448), .A2(n1889), .B1(n415), .B2(n1890), .ZN(n2080) );
  OAI22_X1 U1063 ( .A1(n515), .A2(n1891), .B1(n482), .B2(n1892), .ZN(n2079) );
  OAI22_X1 U1064 ( .A1(n582), .A2(n1893), .B1(n549), .B2(n1894), .ZN(n2078) );
  OAI22_X1 U1065 ( .A1(n650), .A2(n1895), .B1(n616), .B2(n1896), .ZN(n2077) );
  NOR4_X1 U1066 ( .A1(n2081), .A2(n2082), .A3(n2083), .A4(n2084), .ZN(n2070)
         );
  OAI22_X1 U1067 ( .A1(n717), .A2(n1901), .B1(n683), .B2(n1902), .ZN(n2084) );
  OAI22_X1 U1068 ( .A1(n784), .A2(n1903), .B1(n750), .B2(n1904), .ZN(n2083) );
  OAI22_X1 U1069 ( .A1(n851), .A2(n1905), .B1(n818), .B2(n1906), .ZN(n2082) );
  OAI22_X1 U1070 ( .A1(n918), .A2(n1907), .B1(n885), .B2(n1908), .ZN(n2081) );
  NOR4_X1 U1071 ( .A1(n2085), .A2(n2086), .A3(n2087), .A4(n2088), .ZN(n2069)
         );
  OAI22_X1 U1072 ( .A1(n986), .A2(n1913), .B1(n952), .B2(n1914), .ZN(n2088) );
  OAI22_X1 U1073 ( .A1(n1053), .A2(n1915), .B1(n1019), .B2(n1916), .ZN(n2087)
         );
  OAI22_X1 U1074 ( .A1(n95), .A2(n1917), .B1(n1086), .B2(n43), .ZN(n2086) );
  OAI22_X1 U1075 ( .A1(n168), .A2(n45), .B1(n133), .B2(n1920), .ZN(n2085) );
  OAI22_X1 U1076 ( .A1(n2089), .A2(n1867), .B1(n1868), .B2(n1326), .ZN(N4534)
         );
  NOR4_X1 U1077 ( .A1(n2094), .A2(n2095), .A3(n2096), .A4(n2097), .ZN(n2093)
         );
  OAI22_X1 U1078 ( .A1(n190), .A2(n1877), .B1(n900), .B2(n1878), .ZN(n2097) );
  OAI22_X1 U1079 ( .A1(n254), .A2(n1879), .B1(n222), .B2(n1880), .ZN(n2096) );
  OAI22_X1 U1080 ( .A1(n318), .A2(n1881), .B1(n286), .B2(n1882), .ZN(n2095) );
  OAI22_X1 U1081 ( .A1(n382), .A2(n1883), .B1(n350), .B2(n1884), .ZN(n2094) );
  NOR4_X1 U1082 ( .A1(n2098), .A2(n2099), .A3(n2100), .A4(n2101), .ZN(n2092)
         );
  OAI22_X1 U1083 ( .A1(n447), .A2(n1889), .B1(n414), .B2(n1890), .ZN(n2101) );
  OAI22_X1 U1084 ( .A1(n514), .A2(n1891), .B1(n481), .B2(n1892), .ZN(n2100) );
  OAI22_X1 U1085 ( .A1(n581), .A2(n1893), .B1(n548), .B2(n1894), .ZN(n2099) );
  OAI22_X1 U1086 ( .A1(n649), .A2(n1895), .B1(n615), .B2(n1896), .ZN(n2098) );
  NOR4_X1 U1087 ( .A1(n2102), .A2(n2103), .A3(n2104), .A4(n2105), .ZN(n2091)
         );
  OAI22_X1 U1088 ( .A1(n716), .A2(n1901), .B1(n682), .B2(n1902), .ZN(n2105) );
  OAI22_X1 U1089 ( .A1(n783), .A2(n1903), .B1(n749), .B2(n1904), .ZN(n2104) );
  OAI22_X1 U1090 ( .A1(n850), .A2(n1905), .B1(n817), .B2(n1906), .ZN(n2103) );
  OAI22_X1 U1091 ( .A1(n917), .A2(n1907), .B1(n884), .B2(n1908), .ZN(n2102) );
  NOR4_X1 U1092 ( .A1(n2106), .A2(n2107), .A3(n2108), .A4(n2109), .ZN(n2090)
         );
  OAI22_X1 U1093 ( .A1(n985), .A2(n1913), .B1(n951), .B2(n1914), .ZN(n2109) );
  OAI22_X1 U1094 ( .A1(n1052), .A2(n1915), .B1(n1018), .B2(n1916), .ZN(n2108)
         );
  OAI22_X1 U1095 ( .A1(n93), .A2(n1917), .B1(n1085), .B2(n43), .ZN(n2107) );
  OAI22_X1 U1096 ( .A1(n167), .A2(n45), .B1(n132), .B2(n1920), .ZN(n2106) );
  OAI22_X1 U1097 ( .A1(n2110), .A2(n1867), .B1(n1868), .B2(n1348), .ZN(N4532)
         );
  NOR4_X1 U1098 ( .A1(n2115), .A2(n2116), .A3(n2117), .A4(n2118), .ZN(n2114)
         );
  OAI22_X1 U1099 ( .A1(n189), .A2(n1877), .B1(n879), .B2(n1878), .ZN(n2118) );
  OAI22_X1 U1100 ( .A1(n253), .A2(n1879), .B1(n221), .B2(n1880), .ZN(n2117) );
  OAI22_X1 U1101 ( .A1(n317), .A2(n1881), .B1(n285), .B2(n1882), .ZN(n2116) );
  OAI22_X1 U1102 ( .A1(n381), .A2(n1883), .B1(n349), .B2(n1884), .ZN(n2115) );
  NOR4_X1 U1103 ( .A1(n2119), .A2(n2120), .A3(n2121), .A4(n2122), .ZN(n2113)
         );
  OAI22_X1 U1104 ( .A1(n446), .A2(n1889), .B1(n413), .B2(n1890), .ZN(n2122) );
  OAI22_X1 U1105 ( .A1(n513), .A2(n1891), .B1(n479), .B2(n1892), .ZN(n2121) );
  OAI22_X1 U1106 ( .A1(n580), .A2(n1893), .B1(n547), .B2(n1894), .ZN(n2120) );
  OAI22_X1 U1107 ( .A1(n647), .A2(n1895), .B1(n614), .B2(n1896), .ZN(n2119) );
  NOR4_X1 U1108 ( .A1(n2123), .A2(n2124), .A3(n2125), .A4(n2126), .ZN(n2112)
         );
  OAI22_X1 U1109 ( .A1(n715), .A2(n1901), .B1(n681), .B2(n1902), .ZN(n2126) );
  OAI22_X1 U1110 ( .A1(n782), .A2(n1903), .B1(n748), .B2(n1904), .ZN(n2125) );
  OAI22_X1 U1111 ( .A1(n849), .A2(n1905), .B1(n815), .B2(n1906), .ZN(n2124) );
  OAI22_X1 U1112 ( .A1(n916), .A2(n1907), .B1(n883), .B2(n1908), .ZN(n2123) );
  NOR4_X1 U1113 ( .A1(n2127), .A2(n2128), .A3(n2129), .A4(n2130), .ZN(n2111)
         );
  OAI22_X1 U1114 ( .A1(n983), .A2(n1913), .B1(n950), .B2(n1914), .ZN(n2130) );
  OAI22_X1 U1115 ( .A1(n1051), .A2(n1915), .B1(n1017), .B2(n1916), .ZN(n2129)
         );
  OAI22_X1 U1116 ( .A1(n91), .A2(n1917), .B1(n1084), .B2(n43), .ZN(n2128) );
  OAI22_X1 U1117 ( .A1(n166), .A2(n45), .B1(n130), .B2(n1920), .ZN(n2127) );
  OAI22_X1 U1118 ( .A1(n2131), .A2(n1867), .B1(n1868), .B2(n1370), .ZN(N4530)
         );
  NOR4_X1 U1119 ( .A1(n2136), .A2(n2137), .A3(n2138), .A4(n2139), .ZN(n2135)
         );
  OAI22_X1 U1120 ( .A1(n188), .A2(n1877), .B1(n858), .B2(n1878), .ZN(n2139) );
  OAI22_X1 U1121 ( .A1(n252), .A2(n1879), .B1(n220), .B2(n1880), .ZN(n2138) );
  OAI22_X1 U1122 ( .A1(n316), .A2(n1881), .B1(n284), .B2(n1882), .ZN(n2137) );
  OAI22_X1 U1123 ( .A1(n380), .A2(n1883), .B1(n348), .B2(n1884), .ZN(n2136) );
  NOR4_X1 U1124 ( .A1(n2140), .A2(n2141), .A3(n2142), .A4(n2143), .ZN(n2134)
         );
  OAI22_X1 U1125 ( .A1(n445), .A2(n1889), .B1(n412), .B2(n1890), .ZN(n2143) );
  OAI22_X1 U1126 ( .A1(n512), .A2(n1891), .B1(n478), .B2(n1892), .ZN(n2142) );
  OAI22_X1 U1127 ( .A1(n579), .A2(n1893), .B1(n546), .B2(n1894), .ZN(n2141) );
  OAI22_X1 U1128 ( .A1(n646), .A2(n1895), .B1(n613), .B2(n1896), .ZN(n2140) );
  NOR4_X1 U1129 ( .A1(n2144), .A2(n2145), .A3(n2146), .A4(n2147), .ZN(n2133)
         );
  OAI22_X1 U1130 ( .A1(n714), .A2(n1901), .B1(n680), .B2(n1902), .ZN(n2147) );
  OAI22_X1 U1131 ( .A1(n781), .A2(n1903), .B1(n747), .B2(n1904), .ZN(n2146) );
  OAI22_X1 U1132 ( .A1(n848), .A2(n1905), .B1(n814), .B2(n1906), .ZN(n2145) );
  OAI22_X1 U1133 ( .A1(n915), .A2(n1907), .B1(n882), .B2(n1908), .ZN(n2144) );
  NOR4_X1 U1134 ( .A1(n2148), .A2(n2149), .A3(n2150), .A4(n2151), .ZN(n2132)
         );
  OAI22_X1 U1135 ( .A1(n982), .A2(n1913), .B1(n949), .B2(n1914), .ZN(n2151) );
  OAI22_X1 U1136 ( .A1(n1050), .A2(n1915), .B1(n1016), .B2(n1916), .ZN(n2150)
         );
  OAI22_X1 U1137 ( .A1(n89), .A2(n1917), .B1(n1083), .B2(n43), .ZN(n2149) );
  OAI22_X1 U1138 ( .A1(n165), .A2(n45), .B1(n129), .B2(n1920), .ZN(n2148) );
  OAI22_X1 U1139 ( .A1(n2152), .A2(n1867), .B1(n1868), .B2(n1392), .ZN(N4528)
         );
  NOR4_X1 U1140 ( .A1(n2157), .A2(n2158), .A3(n2159), .A4(n2160), .ZN(n2156)
         );
  OAI22_X1 U1141 ( .A1(n187), .A2(n1877), .B1(n837), .B2(n1878), .ZN(n2160) );
  OAI22_X1 U1142 ( .A1(n251), .A2(n1879), .B1(n219), .B2(n1880), .ZN(n2159) );
  OAI22_X1 U1143 ( .A1(n315), .A2(n1881), .B1(n283), .B2(n1882), .ZN(n2158) );
  OAI22_X1 U1144 ( .A1(n379), .A2(n1883), .B1(n347), .B2(n1884), .ZN(n2157) );
  NOR4_X1 U1145 ( .A1(n2161), .A2(n2162), .A3(n2163), .A4(n2164), .ZN(n2155)
         );
  OAI22_X1 U1146 ( .A1(n444), .A2(n1889), .B1(n411), .B2(n1890), .ZN(n2164) );
  OAI22_X1 U1147 ( .A1(n511), .A2(n1891), .B1(n477), .B2(n1892), .ZN(n2163) );
  OAI22_X1 U1148 ( .A1(n578), .A2(n1893), .B1(n545), .B2(n1894), .ZN(n2162) );
  OAI22_X1 U1149 ( .A1(n645), .A2(n1895), .B1(n612), .B2(n1896), .ZN(n2161) );
  NOR4_X1 U1150 ( .A1(n2165), .A2(n2166), .A3(n2167), .A4(n2168), .ZN(n2154)
         );
  OAI22_X1 U1151 ( .A1(n713), .A2(n1901), .B1(n679), .B2(n1902), .ZN(n2168) );
  OAI22_X1 U1152 ( .A1(n780), .A2(n1903), .B1(n746), .B2(n1904), .ZN(n2167) );
  OAI22_X1 U1153 ( .A1(n847), .A2(n1905), .B1(n813), .B2(n1906), .ZN(n2166) );
  OAI22_X1 U1154 ( .A1(n914), .A2(n1907), .B1(n881), .B2(n1908), .ZN(n2165) );
  NOR4_X1 U1155 ( .A1(n2169), .A2(n2170), .A3(n2171), .A4(n2172), .ZN(n2153)
         );
  OAI22_X1 U1156 ( .A1(n981), .A2(n1913), .B1(n948), .B2(n1914), .ZN(n2172) );
  OAI22_X1 U1157 ( .A1(n1049), .A2(n1915), .B1(n1015), .B2(n1916), .ZN(n2171)
         );
  OAI22_X1 U1158 ( .A1(n87), .A2(n41), .B1(n1082), .B2(n43), .ZN(n2170) );
  OAI22_X1 U1159 ( .A1(n163), .A2(n1919), .B1(n128), .B2(n1920), .ZN(n2169) );
  OAI22_X1 U1160 ( .A1(n2173), .A2(n1867), .B1(n1868), .B2(n1414), .ZN(N4526)
         );
  NOR4_X1 U1161 ( .A1(n2178), .A2(n2179), .A3(n2180), .A4(n2181), .ZN(n2177)
         );
  OAI22_X1 U1162 ( .A1(n186), .A2(n1877), .B1(n816), .B2(n1878), .ZN(n2181) );
  OAI22_X1 U1163 ( .A1(n250), .A2(n1879), .B1(n218), .B2(n1880), .ZN(n2180) );
  OAI22_X1 U1164 ( .A1(n314), .A2(n1881), .B1(n282), .B2(n1882), .ZN(n2179) );
  OAI22_X1 U1165 ( .A1(n378), .A2(n1883), .B1(n346), .B2(n1884), .ZN(n2178) );
  NOR4_X1 U1166 ( .A1(n2182), .A2(n2183), .A3(n2184), .A4(n2185), .ZN(n2176)
         );
  OAI22_X1 U1167 ( .A1(n443), .A2(n1889), .B1(n410), .B2(n1890), .ZN(n2185) );
  OAI22_X1 U1168 ( .A1(n510), .A2(n1891), .B1(n476), .B2(n1892), .ZN(n2184) );
  OAI22_X1 U1169 ( .A1(n577), .A2(n1893), .B1(n544), .B2(n1894), .ZN(n2183) );
  OAI22_X1 U1170 ( .A1(n644), .A2(n1895), .B1(n611), .B2(n1896), .ZN(n2182) );
  NOR4_X1 U1171 ( .A1(n2186), .A2(n2187), .A3(n2188), .A4(n2189), .ZN(n2175)
         );
  OAI22_X1 U1172 ( .A1(n712), .A2(n1901), .B1(n678), .B2(n1902), .ZN(n2189) );
  OAI22_X1 U1173 ( .A1(n779), .A2(n1903), .B1(n745), .B2(n1904), .ZN(n2188) );
  OAI22_X1 U1174 ( .A1(n846), .A2(n1905), .B1(n812), .B2(n1906), .ZN(n2187) );
  OAI22_X1 U1175 ( .A1(n913), .A2(n1907), .B1(n880), .B2(n1908), .ZN(n2186) );
  NOR4_X1 U1176 ( .A1(n2190), .A2(n2191), .A3(n2192), .A4(n2193), .ZN(n2174)
         );
  OAI22_X1 U1177 ( .A1(n980), .A2(n1913), .B1(n947), .B2(n1914), .ZN(n2193) );
  OAI22_X1 U1178 ( .A1(n1048), .A2(n1915), .B1(n1014), .B2(n1916), .ZN(n2192)
         );
  OAI22_X1 U1179 ( .A1(n85), .A2(n41), .B1(n1081), .B2(n43), .ZN(n2191) );
  OAI22_X1 U1180 ( .A1(n162), .A2(n1919), .B1(n127), .B2(n1920), .ZN(n2190) );
  OAI22_X1 U1181 ( .A1(n2194), .A2(n1867), .B1(n1868), .B2(n1436), .ZN(N4524)
         );
  NOR4_X1 U1182 ( .A1(n2199), .A2(n2200), .A3(n2201), .A4(n2202), .ZN(n2198)
         );
  OAI22_X1 U1183 ( .A1(n185), .A2(n1877), .B1(n795), .B2(n1878), .ZN(n2202) );
  OAI22_X1 U1184 ( .A1(n249), .A2(n1879), .B1(n217), .B2(n1880), .ZN(n2201) );
  OAI22_X1 U1185 ( .A1(n313), .A2(n1881), .B1(n281), .B2(n1882), .ZN(n2200) );
  OAI22_X1 U1186 ( .A1(n377), .A2(n1883), .B1(n345), .B2(n1884), .ZN(n2199) );
  NOR4_X1 U1187 ( .A1(n2203), .A2(n2204), .A3(n2205), .A4(n2206), .ZN(n2197)
         );
  OAI22_X1 U1188 ( .A1(n442), .A2(n1889), .B1(n409), .B2(n1890), .ZN(n2206) );
  OAI22_X1 U1189 ( .A1(n509), .A2(n1891), .B1(n475), .B2(n1892), .ZN(n2205) );
  OAI22_X1 U1190 ( .A1(n576), .A2(n1893), .B1(n542), .B2(n1894), .ZN(n2204) );
  OAI22_X1 U1191 ( .A1(n643), .A2(n1895), .B1(n610), .B2(n1896), .ZN(n2203) );
  NOR4_X1 U1192 ( .A1(n2207), .A2(n2208), .A3(n2209), .A4(n2210), .ZN(n2196)
         );
  OAI22_X1 U1193 ( .A1(n710), .A2(n1901), .B1(n677), .B2(n1902), .ZN(n2210) );
  OAI22_X1 U1194 ( .A1(n778), .A2(n1903), .B1(n744), .B2(n1904), .ZN(n2209) );
  OAI22_X1 U1195 ( .A1(n845), .A2(n1905), .B1(n811), .B2(n1906), .ZN(n2208) );
  OAI22_X1 U1196 ( .A1(n912), .A2(n1907), .B1(n878), .B2(n1908), .ZN(n2207) );
  NOR4_X1 U1197 ( .A1(n2211), .A2(n2212), .A3(n2213), .A4(n2214), .ZN(n2195)
         );
  OAI22_X1 U1198 ( .A1(n979), .A2(n1913), .B1(n946), .B2(n1914), .ZN(n2214) );
  OAI22_X1 U1199 ( .A1(n1046), .A2(n1915), .B1(n1013), .B2(n1916), .ZN(n2213)
         );
  OAI22_X1 U1200 ( .A1(n83), .A2(n41), .B1(n1080), .B2(n43), .ZN(n2212) );
  OAI22_X1 U1201 ( .A1(n161), .A2(n1919), .B1(n126), .B2(n1920), .ZN(n2211) );
  OAI22_X1 U1202 ( .A1(n2215), .A2(n1867), .B1(n1868), .B2(n1458), .ZN(N4522)
         );
  NOR4_X1 U1203 ( .A1(n2220), .A2(n2221), .A3(n2222), .A4(n2223), .ZN(n2219)
         );
  OAI22_X1 U1204 ( .A1(n184), .A2(n1877), .B1(n774), .B2(n1878), .ZN(n2223) );
  OAI22_X1 U1205 ( .A1(n248), .A2(n1879), .B1(n216), .B2(n1880), .ZN(n2222) );
  OAI22_X1 U1206 ( .A1(n312), .A2(n1881), .B1(n280), .B2(n1882), .ZN(n2221) );
  OAI22_X1 U1207 ( .A1(n376), .A2(n1883), .B1(n344), .B2(n1884), .ZN(n2220) );
  NOR4_X1 U1208 ( .A1(n2224), .A2(n2225), .A3(n2226), .A4(n2227), .ZN(n2218)
         );
  OAI22_X1 U1209 ( .A1(n441), .A2(n1889), .B1(n408), .B2(n1890), .ZN(n2227) );
  OAI22_X1 U1210 ( .A1(n508), .A2(n1891), .B1(n474), .B2(n1892), .ZN(n2226) );
  OAI22_X1 U1211 ( .A1(n575), .A2(n1893), .B1(n541), .B2(n1894), .ZN(n2225) );
  OAI22_X1 U1212 ( .A1(n642), .A2(n1895), .B1(n609), .B2(n1896), .ZN(n2224) );
  NOR4_X1 U1213 ( .A1(n2228), .A2(n2229), .A3(n2230), .A4(n2231), .ZN(n2217)
         );
  OAI22_X1 U1214 ( .A1(n709), .A2(n1901), .B1(n676), .B2(n1902), .ZN(n2231) );
  OAI22_X1 U1215 ( .A1(n777), .A2(n1903), .B1(n743), .B2(n1904), .ZN(n2230) );
  OAI22_X1 U1216 ( .A1(n844), .A2(n1905), .B1(n810), .B2(n1906), .ZN(n2229) );
  OAI22_X1 U1217 ( .A1(n911), .A2(n1907), .B1(n877), .B2(n1908), .ZN(n2228) );
  NOR4_X1 U1218 ( .A1(n2232), .A2(n2233), .A3(n2234), .A4(n2235), .ZN(n2216)
         );
  OAI22_X1 U1219 ( .A1(n978), .A2(n1913), .B1(n945), .B2(n1914), .ZN(n2235) );
  OAI22_X1 U1220 ( .A1(n1045), .A2(n1915), .B1(n1012), .B2(n1916), .ZN(n2234)
         );
  OAI22_X1 U1221 ( .A1(n81), .A2(n41), .B1(n1079), .B2(n43), .ZN(n2233) );
  OAI22_X1 U1222 ( .A1(n160), .A2(n1919), .B1(n125), .B2(n1920), .ZN(n2232) );
  OAI22_X1 U1223 ( .A1(n2236), .A2(n1867), .B1(n1868), .B2(n1480), .ZN(N4520)
         );
  NOR4_X1 U1224 ( .A1(n2241), .A2(n2242), .A3(n2243), .A4(n2244), .ZN(n2240)
         );
  OAI22_X1 U1225 ( .A1(n183), .A2(n1877), .B1(n753), .B2(n1878), .ZN(n2244) );
  OAI22_X1 U1226 ( .A1(n247), .A2(n1879), .B1(n215), .B2(n1880), .ZN(n2243) );
  OAI22_X1 U1227 ( .A1(n311), .A2(n1881), .B1(n279), .B2(n1882), .ZN(n2242) );
  OAI22_X1 U1228 ( .A1(n375), .A2(n1883), .B1(n343), .B2(n1884), .ZN(n2241) );
  NOR4_X1 U1229 ( .A1(n2245), .A2(n2246), .A3(n2247), .A4(n2248), .ZN(n2239)
         );
  OAI22_X1 U1230 ( .A1(n440), .A2(n1889), .B1(n407), .B2(n1890), .ZN(n2248) );
  OAI22_X1 U1231 ( .A1(n507), .A2(n1891), .B1(n473), .B2(n1892), .ZN(n2247) );
  OAI22_X1 U1232 ( .A1(n574), .A2(n1893), .B1(n540), .B2(n1894), .ZN(n2246) );
  OAI22_X1 U1233 ( .A1(n641), .A2(n1895), .B1(n608), .B2(n1896), .ZN(n2245) );
  NOR4_X1 U1234 ( .A1(n2249), .A2(n2250), .A3(n2251), .A4(n2252), .ZN(n2238)
         );
  OAI22_X1 U1235 ( .A1(n708), .A2(n1901), .B1(n675), .B2(n1902), .ZN(n2252) );
  OAI22_X1 U1236 ( .A1(n776), .A2(n1903), .B1(n742), .B2(n1904), .ZN(n2251) );
  OAI22_X1 U1237 ( .A1(n843), .A2(n1905), .B1(n809), .B2(n1906), .ZN(n2250) );
  OAI22_X1 U1238 ( .A1(n910), .A2(n1907), .B1(n876), .B2(n1908), .ZN(n2249) );
  NOR4_X1 U1239 ( .A1(n2253), .A2(n2254), .A3(n2255), .A4(n2256), .ZN(n2237)
         );
  OAI22_X1 U1240 ( .A1(n977), .A2(n1913), .B1(n944), .B2(n1914), .ZN(n2256) );
  OAI22_X1 U1241 ( .A1(n1044), .A2(n1915), .B1(n1011), .B2(n1916), .ZN(n2255)
         );
  OAI22_X1 U1242 ( .A1(n79), .A2(n41), .B1(n1078), .B2(n43), .ZN(n2254) );
  OAI22_X1 U1243 ( .A1(n159), .A2(n1919), .B1(n124), .B2(n1920), .ZN(n2253) );
  OAI22_X1 U1244 ( .A1(n2257), .A2(n1867), .B1(n1868), .B2(n1502), .ZN(N4518)
         );
  NOR4_X1 U1245 ( .A1(n2262), .A2(n2263), .A3(n2264), .A4(n2265), .ZN(n2261)
         );
  OAI22_X1 U1246 ( .A1(n182), .A2(n1877), .B1(n732), .B2(n1878), .ZN(n2265) );
  OAI22_X1 U1247 ( .A1(n246), .A2(n1879), .B1(n214), .B2(n1880), .ZN(n2264) );
  OAI22_X1 U1248 ( .A1(n310), .A2(n1881), .B1(n278), .B2(n1882), .ZN(n2263) );
  OAI22_X1 U1249 ( .A1(n374), .A2(n1883), .B1(n342), .B2(n1884), .ZN(n2262) );
  NOR4_X1 U1250 ( .A1(n2266), .A2(n2267), .A3(n2268), .A4(n2269), .ZN(n2260)
         );
  OAI22_X1 U1251 ( .A1(n439), .A2(n1889), .B1(n406), .B2(n1890), .ZN(n2269) );
  OAI22_X1 U1252 ( .A1(n506), .A2(n1891), .B1(n472), .B2(n1892), .ZN(n2268) );
  OAI22_X1 U1253 ( .A1(n573), .A2(n1893), .B1(n539), .B2(n1894), .ZN(n2267) );
  OAI22_X1 U1254 ( .A1(n640), .A2(n1895), .B1(n607), .B2(n1896), .ZN(n2266) );
  NOR4_X1 U1255 ( .A1(n2270), .A2(n2271), .A3(n2272), .A4(n2273), .ZN(n2259)
         );
  OAI22_X1 U1256 ( .A1(n707), .A2(n1901), .B1(n674), .B2(n1902), .ZN(n2273) );
  OAI22_X1 U1257 ( .A1(n775), .A2(n1903), .B1(n741), .B2(n1904), .ZN(n2272) );
  OAI22_X1 U1258 ( .A1(n842), .A2(n1905), .B1(n808), .B2(n1906), .ZN(n2271) );
  OAI22_X1 U1259 ( .A1(n909), .A2(n1907), .B1(n875), .B2(n1908), .ZN(n2270) );
  NOR4_X1 U1260 ( .A1(n2274), .A2(n2275), .A3(n2276), .A4(n2277), .ZN(n2258)
         );
  OAI22_X1 U1261 ( .A1(n976), .A2(n1913), .B1(n943), .B2(n1914), .ZN(n2277) );
  OAI22_X1 U1262 ( .A1(n1043), .A2(n1915), .B1(n1010), .B2(n1916), .ZN(n2276)
         );
  OAI22_X1 U1263 ( .A1(n77), .A2(n41), .B1(n1077), .B2(n43), .ZN(n2275) );
  OAI22_X1 U1264 ( .A1(n158), .A2(n1919), .B1(n123), .B2(n1920), .ZN(n2274) );
  OAI22_X1 U1265 ( .A1(n2278), .A2(n1867), .B1(n1868), .B2(n1524), .ZN(N4516)
         );
  NOR4_X1 U1266 ( .A1(n2283), .A2(n2284), .A3(n2285), .A4(n2286), .ZN(n2282)
         );
  OAI22_X1 U1267 ( .A1(n181), .A2(n1877), .B1(n711), .B2(n1878), .ZN(n2286) );
  OAI22_X1 U1268 ( .A1(n245), .A2(n1879), .B1(n213), .B2(n1880), .ZN(n2285) );
  OAI22_X1 U1269 ( .A1(n309), .A2(n1881), .B1(n277), .B2(n1882), .ZN(n2284) );
  OAI22_X1 U1270 ( .A1(n373), .A2(n1883), .B1(n341), .B2(n1884), .ZN(n2283) );
  NOR4_X1 U1271 ( .A1(n2287), .A2(n2288), .A3(n2289), .A4(n2290), .ZN(n2281)
         );
  OAI22_X1 U1272 ( .A1(n437), .A2(n1889), .B1(n405), .B2(n1890), .ZN(n2290) );
  OAI22_X1 U1273 ( .A1(n505), .A2(n1891), .B1(n471), .B2(n1892), .ZN(n2289) );
  OAI22_X1 U1274 ( .A1(n572), .A2(n1893), .B1(n538), .B2(n1894), .ZN(n2288) );
  OAI22_X1 U1275 ( .A1(n639), .A2(n1895), .B1(n605), .B2(n1896), .ZN(n2287) );
  NOR4_X1 U1276 ( .A1(n2291), .A2(n2292), .A3(n2293), .A4(n2294), .ZN(n2280)
         );
  OAI22_X1 U1277 ( .A1(n706), .A2(n1901), .B1(n673), .B2(n1902), .ZN(n2294) );
  OAI22_X1 U1278 ( .A1(n773), .A2(n1903), .B1(n740), .B2(n1904), .ZN(n2293) );
  OAI22_X1 U1279 ( .A1(n841), .A2(n1905), .B1(n807), .B2(n1906), .ZN(n2292) );
  OAI22_X1 U1280 ( .A1(n908), .A2(n1907), .B1(n874), .B2(n1908), .ZN(n2291) );
  NOR4_X1 U1281 ( .A1(n2295), .A2(n2296), .A3(n2297), .A4(n2298), .ZN(n2279)
         );
  OAI22_X1 U1282 ( .A1(n975), .A2(n1913), .B1(n941), .B2(n1914), .ZN(n2298) );
  OAI22_X1 U1283 ( .A1(n1042), .A2(n1915), .B1(n1009), .B2(n1916), .ZN(n2297)
         );
  OAI22_X1 U1284 ( .A1(n73), .A2(n41), .B1(n1076), .B2(n43), .ZN(n2296) );
  OAI22_X1 U1285 ( .A1(n157), .A2(n1919), .B1(n122), .B2(n1920), .ZN(n2295) );
  OAI22_X1 U1286 ( .A1(n2299), .A2(n1867), .B1(n1868), .B2(n1546), .ZN(N4514)
         );
  NOR4_X1 U1287 ( .A1(n2304), .A2(n2305), .A3(n2306), .A4(n2307), .ZN(n2303)
         );
  OAI22_X1 U1288 ( .A1(n180), .A2(n1877), .B1(n690), .B2(n1878), .ZN(n2307) );
  OAI22_X1 U1289 ( .A1(n244), .A2(n1879), .B1(n212), .B2(n1880), .ZN(n2306) );
  OAI22_X1 U1290 ( .A1(n308), .A2(n1881), .B1(n276), .B2(n1882), .ZN(n2305) );
  OAI22_X1 U1291 ( .A1(n372), .A2(n1883), .B1(n340), .B2(n1884), .ZN(n2304) );
  NOR4_X1 U1292 ( .A1(n2308), .A2(n2309), .A3(n2310), .A4(n2311), .ZN(n2302)
         );
  OAI22_X1 U1293 ( .A1(n436), .A2(n1889), .B1(n404), .B2(n1890), .ZN(n2311) );
  OAI22_X1 U1294 ( .A1(n504), .A2(n1891), .B1(n470), .B2(n1892), .ZN(n2310) );
  OAI22_X1 U1295 ( .A1(n571), .A2(n1893), .B1(n537), .B2(n1894), .ZN(n2309) );
  OAI22_X1 U1296 ( .A1(n638), .A2(n1895), .B1(n604), .B2(n1896), .ZN(n2308) );
  NOR4_X1 U1297 ( .A1(n2312), .A2(n2313), .A3(n2314), .A4(n2315), .ZN(n2301)
         );
  OAI22_X1 U1298 ( .A1(n705), .A2(n1901), .B1(n672), .B2(n1902), .ZN(n2315) );
  OAI22_X1 U1299 ( .A1(n772), .A2(n1903), .B1(n739), .B2(n1904), .ZN(n2314) );
  OAI22_X1 U1300 ( .A1(n840), .A2(n1905), .B1(n806), .B2(n1906), .ZN(n2313) );
  OAI22_X1 U1301 ( .A1(n907), .A2(n1907), .B1(n873), .B2(n1908), .ZN(n2312) );
  NOR4_X1 U1302 ( .A1(n2316), .A2(n2317), .A3(n2318), .A4(n2319), .ZN(n2300)
         );
  OAI22_X1 U1303 ( .A1(n974), .A2(n1913), .B1(n940), .B2(n1914), .ZN(n2319) );
  OAI22_X1 U1304 ( .A1(n1041), .A2(n1915), .B1(n1008), .B2(n1916), .ZN(n2318)
         );
  OAI22_X1 U1305 ( .A1(n71), .A2(n41), .B1(n1075), .B2(n43), .ZN(n2317) );
  OAI22_X1 U1306 ( .A1(n156), .A2(n1919), .B1(n121), .B2(n1920), .ZN(n2316) );
  OAI22_X1 U1307 ( .A1(n2320), .A2(n1867), .B1(n1868), .B2(n1568), .ZN(N4512)
         );
  NOR4_X1 U1308 ( .A1(n2325), .A2(n2326), .A3(n2327), .A4(n2328), .ZN(n2324)
         );
  OAI22_X1 U1309 ( .A1(n179), .A2(n1877), .B1(n669), .B2(n1878), .ZN(n2328) );
  OAI22_X1 U1310 ( .A1(n243), .A2(n1879), .B1(n211), .B2(n1880), .ZN(n2327) );
  OAI22_X1 U1311 ( .A1(n307), .A2(n1881), .B1(n275), .B2(n1882), .ZN(n2326) );
  OAI22_X1 U1312 ( .A1(n371), .A2(n39), .B1(n339), .B2(n1884), .ZN(n2325) );
  NOR4_X1 U1313 ( .A1(n2329), .A2(n2330), .A3(n2331), .A4(n2332), .ZN(n2323)
         );
  OAI22_X1 U1314 ( .A1(n435), .A2(n1889), .B1(n403), .B2(n1890), .ZN(n2332) );
  OAI22_X1 U1315 ( .A1(n503), .A2(n1891), .B1(n469), .B2(n1892), .ZN(n2331) );
  OAI22_X1 U1316 ( .A1(n570), .A2(n1893), .B1(n536), .B2(n1894), .ZN(n2330) );
  OAI22_X1 U1317 ( .A1(n637), .A2(n1895), .B1(n603), .B2(n1896), .ZN(n2329) );
  NOR4_X1 U1318 ( .A1(n2333), .A2(n2334), .A3(n2335), .A4(n2336), .ZN(n2322)
         );
  OAI22_X1 U1319 ( .A1(n704), .A2(n1901), .B1(n671), .B2(n1902), .ZN(n2336) );
  OAI22_X1 U1320 ( .A1(n771), .A2(n1903), .B1(n738), .B2(n1904), .ZN(n2335) );
  OAI22_X1 U1321 ( .A1(n839), .A2(n1905), .B1(n805), .B2(n1906), .ZN(n2334) );
  OAI22_X1 U1322 ( .A1(n906), .A2(n1907), .B1(n872), .B2(n1908), .ZN(n2333) );
  NOR4_X1 U1323 ( .A1(n2337), .A2(n2338), .A3(n2339), .A4(n2340), .ZN(n2321)
         );
  OAI22_X1 U1324 ( .A1(n973), .A2(n1913), .B1(n939), .B2(n1914), .ZN(n2340) );
  OAI22_X1 U1325 ( .A1(n1040), .A2(n1915), .B1(n1007), .B2(n1916), .ZN(n2339)
         );
  OAI22_X1 U1326 ( .A1(n69), .A2(n41), .B1(n1074), .B2(n1918), .ZN(n2338) );
  OAI22_X1 U1327 ( .A1(n155), .A2(n1919), .B1(n119), .B2(n1920), .ZN(n2337) );
  OAI22_X1 U1328 ( .A1(n2341), .A2(n1867), .B1(n1868), .B2(n1590), .ZN(N4510)
         );
  NOR4_X1 U1329 ( .A1(n2346), .A2(n2347), .A3(n2348), .A4(n2349), .ZN(n2345)
         );
  OAI22_X1 U1330 ( .A1(n178), .A2(n1877), .B1(n648), .B2(n1878), .ZN(n2349) );
  OAI22_X1 U1331 ( .A1(n242), .A2(n1879), .B1(n210), .B2(n1880), .ZN(n2348) );
  OAI22_X1 U1332 ( .A1(n306), .A2(n1881), .B1(n274), .B2(n1882), .ZN(n2347) );
  OAI22_X1 U1333 ( .A1(n370), .A2(n39), .B1(n338), .B2(n1884), .ZN(n2346) );
  NOR4_X1 U1334 ( .A1(n2350), .A2(n2351), .A3(n2352), .A4(n2353), .ZN(n2344)
         );
  OAI22_X1 U1335 ( .A1(n434), .A2(n1889), .B1(n402), .B2(n1890), .ZN(n2353) );
  OAI22_X1 U1336 ( .A1(n502), .A2(n1891), .B1(n468), .B2(n1892), .ZN(n2352) );
  OAI22_X1 U1337 ( .A1(n569), .A2(n1893), .B1(n535), .B2(n1894), .ZN(n2351) );
  OAI22_X1 U1338 ( .A1(n636), .A2(n1895), .B1(n602), .B2(n1896), .ZN(n2350) );
  NOR4_X1 U1339 ( .A1(n2354), .A2(n2355), .A3(n2356), .A4(n2357), .ZN(n2343)
         );
  OAI22_X1 U1340 ( .A1(n703), .A2(n1901), .B1(n670), .B2(n1902), .ZN(n2357) );
  OAI22_X1 U1341 ( .A1(n770), .A2(n1903), .B1(n737), .B2(n1904), .ZN(n2356) );
  OAI22_X1 U1342 ( .A1(n838), .A2(n1905), .B1(n804), .B2(n1906), .ZN(n2355) );
  OAI22_X1 U1343 ( .A1(n905), .A2(n1907), .B1(n871), .B2(n1908), .ZN(n2354) );
  NOR4_X1 U1344 ( .A1(n2358), .A2(n2359), .A3(n2360), .A4(n2361), .ZN(n2342)
         );
  OAI22_X1 U1345 ( .A1(n972), .A2(n1913), .B1(n938), .B2(n1914), .ZN(n2361) );
  OAI22_X1 U1346 ( .A1(n1039), .A2(n1915), .B1(n1006), .B2(n1916), .ZN(n2360)
         );
  OAI22_X1 U1347 ( .A1(n67), .A2(n41), .B1(n1073), .B2(n1918), .ZN(n2359) );
  OAI22_X1 U1348 ( .A1(n154), .A2(n1919), .B1(n118), .B2(n1920), .ZN(n2358) );
  OAI22_X1 U1349 ( .A1(n2362), .A2(n1867), .B1(n1868), .B2(n1612), .ZN(N4508)
         );
  NOR4_X1 U1350 ( .A1(n2367), .A2(n2368), .A3(n2369), .A4(n2370), .ZN(n2366)
         );
  OAI22_X1 U1351 ( .A1(n175), .A2(n1877), .B1(n627), .B2(n1878), .ZN(n2370) );
  OAI22_X1 U1352 ( .A1(n241), .A2(n1879), .B1(n209), .B2(n1880), .ZN(n2369) );
  OAI22_X1 U1353 ( .A1(n305), .A2(n1881), .B1(n273), .B2(n1882), .ZN(n2368) );
  OAI22_X1 U1354 ( .A1(n369), .A2(n39), .B1(n337), .B2(n1884), .ZN(n2367) );
  NOR4_X1 U1355 ( .A1(n2371), .A2(n2372), .A3(n2373), .A4(n2374), .ZN(n2365)
         );
  OAI22_X1 U1356 ( .A1(n433), .A2(n1889), .B1(n401), .B2(n1890), .ZN(n2374) );
  OAI22_X1 U1357 ( .A1(n500), .A2(n1891), .B1(n467), .B2(n1892), .ZN(n2373) );
  OAI22_X1 U1358 ( .A1(n568), .A2(n1893), .B1(n534), .B2(n1894), .ZN(n2372) );
  OAI22_X1 U1359 ( .A1(n635), .A2(n1895), .B1(n601), .B2(n1896), .ZN(n2371) );
  NOR4_X1 U1360 ( .A1(n2375), .A2(n2376), .A3(n2377), .A4(n2378), .ZN(n2364)
         );
  OAI22_X1 U1361 ( .A1(n702), .A2(n1901), .B1(n668), .B2(n1902), .ZN(n2378) );
  OAI22_X1 U1362 ( .A1(n769), .A2(n1903), .B1(n736), .B2(n1904), .ZN(n2377) );
  OAI22_X1 U1363 ( .A1(n836), .A2(n1905), .B1(n803), .B2(n1906), .ZN(n2376) );
  OAI22_X1 U1364 ( .A1(n904), .A2(n1907), .B1(n870), .B2(n1908), .ZN(n2375) );
  NOR4_X1 U1365 ( .A1(n2379), .A2(n2380), .A3(n2381), .A4(n2382), .ZN(n2363)
         );
  OAI22_X1 U1366 ( .A1(n971), .A2(n1913), .B1(n937), .B2(n1914), .ZN(n2382) );
  OAI22_X1 U1367 ( .A1(n1038), .A2(n1915), .B1(n1004), .B2(n1916), .ZN(n2381)
         );
  OAI22_X1 U1368 ( .A1(n65), .A2(n41), .B1(n1072), .B2(n1918), .ZN(n2380) );
  OAI22_X1 U1369 ( .A1(n152), .A2(n1919), .B1(n117), .B2(n1920), .ZN(n2379) );
  OAI22_X1 U1370 ( .A1(n2383), .A2(n1867), .B1(n1868), .B2(n1634), .ZN(N4506)
         );
  NOR4_X1 U1371 ( .A1(n2388), .A2(n2389), .A3(n2390), .A4(n2391), .ZN(n2387)
         );
  OAI22_X1 U1372 ( .A1(n164), .A2(n1877), .B1(n606), .B2(n1878), .ZN(n2391) );
  OAI22_X1 U1373 ( .A1(n240), .A2(n1879), .B1(n208), .B2(n1880), .ZN(n2390) );
  OAI22_X1 U1374 ( .A1(n304), .A2(n1881), .B1(n272), .B2(n1882), .ZN(n2389) );
  OAI22_X1 U1375 ( .A1(n368), .A2(n39), .B1(n336), .B2(n1884), .ZN(n2388) );
  NOR4_X1 U1376 ( .A1(n2392), .A2(n2393), .A3(n2394), .A4(n2395), .ZN(n2386)
         );
  OAI22_X1 U1377 ( .A1(n432), .A2(n1889), .B1(n400), .B2(n1890), .ZN(n2395) );
  OAI22_X1 U1378 ( .A1(n499), .A2(n1891), .B1(n466), .B2(n1892), .ZN(n2394) );
  OAI22_X1 U1379 ( .A1(n567), .A2(n1893), .B1(n533), .B2(n1894), .ZN(n2393) );
  OAI22_X1 U1380 ( .A1(n634), .A2(n1895), .B1(n600), .B2(n1896), .ZN(n2392) );
  NOR4_X1 U1381 ( .A1(n2396), .A2(n2397), .A3(n2398), .A4(n2399), .ZN(n2385)
         );
  OAI22_X1 U1382 ( .A1(n701), .A2(n1901), .B1(n667), .B2(n1902), .ZN(n2399) );
  OAI22_X1 U1383 ( .A1(n768), .A2(n1903), .B1(n735), .B2(n1904), .ZN(n2398) );
  OAI22_X1 U1384 ( .A1(n835), .A2(n1905), .B1(n802), .B2(n1906), .ZN(n2397) );
  OAI22_X1 U1385 ( .A1(n903), .A2(n1907), .B1(n869), .B2(n1908), .ZN(n2396) );
  NOR4_X1 U1386 ( .A1(n2400), .A2(n2401), .A3(n2402), .A4(n2403), .ZN(n2384)
         );
  OAI22_X1 U1387 ( .A1(n970), .A2(n1913), .B1(n936), .B2(n1914), .ZN(n2403) );
  OAI22_X1 U1388 ( .A1(n1037), .A2(n1915), .B1(n1003), .B2(n1916), .ZN(n2402)
         );
  OAI22_X1 U1389 ( .A1(n63), .A2(n41), .B1(n1071), .B2(n1918), .ZN(n2401) );
  OAI22_X1 U1390 ( .A1(n151), .A2(n45), .B1(n116), .B2(n1920), .ZN(n2400) );
  OAI22_X1 U1391 ( .A1(n2404), .A2(n1867), .B1(n1868), .B2(n1656), .ZN(N4504)
         );
  NOR4_X1 U1392 ( .A1(n2409), .A2(n2410), .A3(n2411), .A4(n2412), .ZN(n2408)
         );
  OAI22_X1 U1393 ( .A1(n153), .A2(n1877), .B1(n585), .B2(n1878), .ZN(n2412) );
  OAI22_X1 U1394 ( .A1(n239), .A2(n1879), .B1(n207), .B2(n1880), .ZN(n2411) );
  OAI22_X1 U1395 ( .A1(n303), .A2(n1881), .B1(n271), .B2(n1882), .ZN(n2410) );
  OAI22_X1 U1396 ( .A1(n367), .A2(n39), .B1(n335), .B2(n1884), .ZN(n2409) );
  NOR4_X1 U1397 ( .A1(n2413), .A2(n2414), .A3(n2415), .A4(n2416), .ZN(n2407)
         );
  OAI22_X1 U1398 ( .A1(n431), .A2(n1889), .B1(n399), .B2(n1890), .ZN(n2416) );
  OAI22_X1 U1399 ( .A1(n498), .A2(n1891), .B1(n465), .B2(n1892), .ZN(n2415) );
  OAI22_X1 U1400 ( .A1(n566), .A2(n1893), .B1(n532), .B2(n1894), .ZN(n2414) );
  OAI22_X1 U1401 ( .A1(n633), .A2(n1895), .B1(n599), .B2(n1896), .ZN(n2413) );
  NOR4_X1 U1402 ( .A1(n2417), .A2(n2418), .A3(n2419), .A4(n2420), .ZN(n2406)
         );
  OAI22_X1 U1403 ( .A1(n700), .A2(n1901), .B1(n666), .B2(n1902), .ZN(n2420) );
  OAI22_X1 U1404 ( .A1(n767), .A2(n1903), .B1(n734), .B2(n1904), .ZN(n2419) );
  OAI22_X1 U1405 ( .A1(n834), .A2(n1905), .B1(n801), .B2(n1906), .ZN(n2418) );
  OAI22_X1 U1406 ( .A1(n902), .A2(n1907), .B1(n868), .B2(n1908), .ZN(n2417) );
  NOR4_X1 U1407 ( .A1(n2421), .A2(n2422), .A3(n2423), .A4(n2424), .ZN(n2405)
         );
  OAI22_X1 U1408 ( .A1(n969), .A2(n1913), .B1(n935), .B2(n1914), .ZN(n2424) );
  OAI22_X1 U1409 ( .A1(n1036), .A2(n1915), .B1(n1002), .B2(n1916), .ZN(n2423)
         );
  OAI22_X1 U1410 ( .A1(n61), .A2(n41), .B1(n1070), .B2(n1918), .ZN(n2422) );
  OAI22_X1 U1411 ( .A1(n150), .A2(n45), .B1(n115), .B2(n1920), .ZN(n2421) );
  OAI22_X1 U1412 ( .A1(n2425), .A2(n1867), .B1(n1868), .B2(n1678), .ZN(N4502)
         );
  NOR4_X1 U1413 ( .A1(n2430), .A2(n2431), .A3(n2432), .A4(n2433), .ZN(n2429)
         );
  OAI22_X1 U1414 ( .A1(n142), .A2(n1877), .B1(n564), .B2(n1878), .ZN(n2433) );
  OAI22_X1 U1415 ( .A1(n238), .A2(n1879), .B1(n206), .B2(n1880), .ZN(n2432) );
  OAI22_X1 U1416 ( .A1(n302), .A2(n1881), .B1(n270), .B2(n1882), .ZN(n2431) );
  OAI22_X1 U1417 ( .A1(n366), .A2(n39), .B1(n334), .B2(n1884), .ZN(n2430) );
  NOR4_X1 U1418 ( .A1(n2434), .A2(n2435), .A3(n2436), .A4(n2437), .ZN(n2428)
         );
  OAI22_X1 U1419 ( .A1(n430), .A2(n1889), .B1(n398), .B2(n1890), .ZN(n2437) );
  OAI22_X1 U1420 ( .A1(n497), .A2(n1891), .B1(n464), .B2(n1892), .ZN(n2436) );
  OAI22_X1 U1421 ( .A1(n565), .A2(n1893), .B1(n531), .B2(n1894), .ZN(n2435) );
  OAI22_X1 U1422 ( .A1(n632), .A2(n1895), .B1(n598), .B2(n1896), .ZN(n2434) );
  NOR4_X1 U1423 ( .A1(n2438), .A2(n2439), .A3(n2440), .A4(n2441), .ZN(n2427)
         );
  OAI22_X1 U1424 ( .A1(n699), .A2(n1901), .B1(n665), .B2(n1902), .ZN(n2441) );
  OAI22_X1 U1425 ( .A1(n766), .A2(n1903), .B1(n733), .B2(n1904), .ZN(n2440) );
  OAI22_X1 U1426 ( .A1(n833), .A2(n1905), .B1(n800), .B2(n1906), .ZN(n2439) );
  OAI22_X1 U1427 ( .A1(n901), .A2(n1907), .B1(n867), .B2(n1908), .ZN(n2438) );
  NOR4_X1 U1428 ( .A1(n2442), .A2(n2443), .A3(n2444), .A4(n2445), .ZN(n2426)
         );
  OAI22_X1 U1429 ( .A1(n968), .A2(n1913), .B1(n934), .B2(n1914), .ZN(n2445) );
  OAI22_X1 U1430 ( .A1(n1035), .A2(n1915), .B1(n1001), .B2(n1916), .ZN(n2444)
         );
  OAI22_X1 U1431 ( .A1(n59), .A2(n1917), .B1(n1069), .B2(n1918), .ZN(n2443) );
  OAI22_X1 U1432 ( .A1(n149), .A2(n45), .B1(n114), .B2(n1920), .ZN(n2442) );
  OAI22_X1 U1433 ( .A1(n2446), .A2(n1867), .B1(n1868), .B2(n1700), .ZN(N4500)
         );
  NOR4_X1 U1434 ( .A1(n2451), .A2(n2452), .A3(n2453), .A4(n2454), .ZN(n2450)
         );
  OAI22_X1 U1435 ( .A1(n131), .A2(n1877), .B1(n543), .B2(n1878), .ZN(n2454) );
  OAI22_X1 U1436 ( .A1(n237), .A2(n1879), .B1(n205), .B2(n1880), .ZN(n2453) );
  OAI22_X1 U1437 ( .A1(n301), .A2(n1881), .B1(n269), .B2(n1882), .ZN(n2452) );
  OAI22_X1 U1438 ( .A1(n365), .A2(n39), .B1(n333), .B2(n1884), .ZN(n2451) );
  NOR4_X1 U1439 ( .A1(n2455), .A2(n2456), .A3(n2457), .A4(n2458), .ZN(n2449)
         );
  OAI22_X1 U1440 ( .A1(n429), .A2(n1889), .B1(n397), .B2(n1890), .ZN(n2458) );
  OAI22_X1 U1441 ( .A1(n496), .A2(n1891), .B1(n463), .B2(n1892), .ZN(n2457) );
  OAI22_X1 U1442 ( .A1(n563), .A2(n1893), .B1(n530), .B2(n1894), .ZN(n2456) );
  OAI22_X1 U1443 ( .A1(n631), .A2(n1895), .B1(n597), .B2(n1896), .ZN(n2455) );
  NOR4_X1 U1444 ( .A1(n2459), .A2(n2460), .A3(n2461), .A4(n2462), .ZN(n2448)
         );
  OAI22_X1 U1445 ( .A1(n698), .A2(n1901), .B1(n664), .B2(n1902), .ZN(n2462) );
  OAI22_X1 U1446 ( .A1(n765), .A2(n1903), .B1(n731), .B2(n1904), .ZN(n2461) );
  OAI22_X1 U1447 ( .A1(n832), .A2(n1905), .B1(n799), .B2(n1906), .ZN(n2460) );
  OAI22_X1 U1448 ( .A1(n899), .A2(n1907), .B1(n866), .B2(n1908), .ZN(n2459) );
  NOR4_X1 U1449 ( .A1(n2463), .A2(n2464), .A3(n2465), .A4(n2466), .ZN(n2447)
         );
  OAI22_X1 U1450 ( .A1(n967), .A2(n1913), .B1(n933), .B2(n1914), .ZN(n2466) );
  OAI22_X1 U1451 ( .A1(n1034), .A2(n1915), .B1(n1000), .B2(n1916), .ZN(n2465)
         );
  OAI22_X1 U1452 ( .A1(n57), .A2(n1917), .B1(n1067), .B2(n1918), .ZN(n2464) );
  OAI22_X1 U1453 ( .A1(n148), .A2(n1919), .B1(n113), .B2(n1920), .ZN(n2463) );
  OAI22_X1 U1454 ( .A1(n2467), .A2(n1867), .B1(n1868), .B2(n1722), .ZN(N4498)
         );
  NOR4_X1 U1455 ( .A1(n2472), .A2(n2473), .A3(n2474), .A4(n2475), .ZN(n2471)
         );
  OAI22_X1 U1456 ( .A1(n120), .A2(n1877), .B1(n522), .B2(n1878), .ZN(n2475) );
  OAI22_X1 U1457 ( .A1(n236), .A2(n1879), .B1(n204), .B2(n1880), .ZN(n2474) );
  OAI22_X1 U1458 ( .A1(n300), .A2(n1881), .B1(n268), .B2(n1882), .ZN(n2473) );
  OAI22_X1 U1459 ( .A1(n364), .A2(n39), .B1(n332), .B2(n1884), .ZN(n2472) );
  NOR4_X1 U1460 ( .A1(n2476), .A2(n2477), .A3(n2478), .A4(n2479), .ZN(n2470)
         );
  OAI22_X1 U1461 ( .A1(n428), .A2(n1889), .B1(n396), .B2(n1890), .ZN(n2479) );
  OAI22_X1 U1462 ( .A1(n495), .A2(n1891), .B1(n462), .B2(n1892), .ZN(n2478) );
  OAI22_X1 U1463 ( .A1(n562), .A2(n1893), .B1(n529), .B2(n1894), .ZN(n2477) );
  OAI22_X1 U1464 ( .A1(n630), .A2(n1895), .B1(n596), .B2(n1896), .ZN(n2476) );
  NOR4_X1 U1465 ( .A1(n2480), .A2(n2481), .A3(n2482), .A4(n2483), .ZN(n2469)
         );
  OAI22_X1 U1466 ( .A1(n697), .A2(n1901), .B1(n663), .B2(n1902), .ZN(n2483) );
  OAI22_X1 U1467 ( .A1(n764), .A2(n1903), .B1(n730), .B2(n1904), .ZN(n2482) );
  OAI22_X1 U1468 ( .A1(n831), .A2(n1905), .B1(n798), .B2(n1906), .ZN(n2481) );
  OAI22_X1 U1469 ( .A1(n898), .A2(n1907), .B1(n865), .B2(n1908), .ZN(n2480) );
  NOR4_X1 U1470 ( .A1(n2484), .A2(n2485), .A3(n2486), .A4(n2487), .ZN(n2468)
         );
  OAI22_X1 U1471 ( .A1(n966), .A2(n1913), .B1(n932), .B2(n1914), .ZN(n2487) );
  OAI22_X1 U1472 ( .A1(n1033), .A2(n1915), .B1(n999), .B2(n1916), .ZN(n2486)
         );
  OAI22_X1 U1473 ( .A1(n55), .A2(n1917), .B1(n1066), .B2(n1918), .ZN(n2485) );
  OAI22_X1 U1474 ( .A1(n147), .A2(n1919), .B1(n112), .B2(n1920), .ZN(n2484) );
  OAI22_X1 U1475 ( .A1(n2488), .A2(n1867), .B1(n1868), .B2(n1744), .ZN(N4496)
         );
  NOR4_X1 U1476 ( .A1(n2489), .A2(n2490), .A3(n2491), .A4(n2492), .ZN(n2488)
         );
  OAI211_X1 U1477 ( .C1(n1100), .C2(n1917), .A(n2493), .B(n2494), .ZN(n2492)
         );
  NOR4_X1 U1478 ( .A1(n2495), .A2(n2496), .A3(n2497), .A4(n2498), .ZN(n2494)
         );
  OAI22_X1 U1479 ( .A1(n109), .A2(n1877), .B1(n203), .B2(n1880), .ZN(n2498) );
  OAI22_X1 U1480 ( .A1(n235), .A2(n1879), .B1(n267), .B2(n1882), .ZN(n2497) );
  OAI22_X1 U1481 ( .A1(n299), .A2(n1881), .B1(n331), .B2(n1884), .ZN(n2496) );
  OAI22_X1 U1482 ( .A1(n363), .A2(n39), .B1(n395), .B2(n1890), .ZN(n2495) );
  NOR4_X1 U1483 ( .A1(n2499), .A2(n2500), .A3(n2501), .A4(n2502), .ZN(n2493)
         );
  OAI22_X1 U1484 ( .A1(n427), .A2(n1889), .B1(n461), .B2(n1892), .ZN(n2502) );
  OAI22_X1 U1485 ( .A1(n494), .A2(n1891), .B1(n528), .B2(n1894), .ZN(n2501) );
  OAI22_X1 U1486 ( .A1(n561), .A2(n1893), .B1(n595), .B2(n1896), .ZN(n2500) );
  OAI22_X1 U1487 ( .A1(n629), .A2(n1895), .B1(n662), .B2(n1902), .ZN(n2499) );
  OAI211_X1 U1488 ( .C1(n146), .C2(n1919), .A(n2503), .B(n2504), .ZN(n2491) );
  NOR4_X1 U1489 ( .A1(n2505), .A2(n2506), .A3(n2507), .A4(n2508), .ZN(n2504)
         );
  OAI22_X1 U1490 ( .A1(n763), .A2(n1903), .B1(n797), .B2(n1906), .ZN(n2508) );
  OAI22_X1 U1491 ( .A1(n696), .A2(n1901), .B1(n729), .B2(n1904), .ZN(n2507) );
  OAI22_X1 U1492 ( .A1(n897), .A2(n1907), .B1(n931), .B2(n1914), .ZN(n2506) );
  OAI22_X1 U1493 ( .A1(n830), .A2(n1905), .B1(n864), .B2(n1908), .ZN(n2505) );
  OAI22_X1 U1494 ( .A1(n1878), .A2(n501), .B1(n1920), .B2(n111), .ZN(n2509) );
  OAI22_X1 U1495 ( .A1(n1032), .A2(n1915), .B1(n1065), .B2(n1918), .ZN(n2490)
         );
  OAI22_X1 U1496 ( .A1(n965), .A2(n1913), .B1(n998), .B2(n1916), .ZN(n2489) );
  OAI22_X1 U1497 ( .A1(n2510), .A2(n1867), .B1(n1868), .B2(n1766), .ZN(N4494)
         );
  NOR4_X1 U1498 ( .A1(n2515), .A2(n2516), .A3(n2517), .A4(n2518), .ZN(n2514)
         );
  OAI22_X1 U1499 ( .A1(n97), .A2(n1877), .B1(n480), .B2(n1878), .ZN(n2518) );
  OAI22_X1 U1500 ( .A1(n234), .A2(n1879), .B1(n202), .B2(n1880), .ZN(n2517) );
  OAI22_X1 U1501 ( .A1(n298), .A2(n1881), .B1(n266), .B2(n1882), .ZN(n2516) );
  OAI22_X1 U1502 ( .A1(n362), .A2(n39), .B1(n330), .B2(n1884), .ZN(n2515) );
  NOR4_X1 U1503 ( .A1(n2519), .A2(n2520), .A3(n2521), .A4(n2522), .ZN(n2513)
         );
  OAI22_X1 U1504 ( .A1(n426), .A2(n1889), .B1(n394), .B2(n1890), .ZN(n2522) );
  OAI22_X1 U1505 ( .A1(n493), .A2(n1891), .B1(n460), .B2(n1892), .ZN(n2521) );
  OAI22_X1 U1506 ( .A1(n560), .A2(n1893), .B1(n527), .B2(n1894), .ZN(n2520) );
  OAI22_X1 U1507 ( .A1(n628), .A2(n1895), .B1(n594), .B2(n1896), .ZN(n2519) );
  NOR4_X1 U1508 ( .A1(n2523), .A2(n2524), .A3(n2525), .A4(n2526), .ZN(n2512)
         );
  OAI22_X1 U1509 ( .A1(n695), .A2(n1901), .B1(n661), .B2(n1902), .ZN(n2526) );
  OAI22_X1 U1510 ( .A1(n762), .A2(n1903), .B1(n728), .B2(n1904), .ZN(n2525) );
  OAI22_X1 U1511 ( .A1(n829), .A2(n1905), .B1(n796), .B2(n1906), .ZN(n2524) );
  OAI22_X1 U1512 ( .A1(n896), .A2(n1907), .B1(n863), .B2(n1908), .ZN(n2523) );
  NOR4_X1 U1513 ( .A1(n2527), .A2(n2528), .A3(n2529), .A4(n2530), .ZN(n2511)
         );
  OAI22_X1 U1514 ( .A1(n964), .A2(n1913), .B1(n930), .B2(n1914), .ZN(n2530) );
  OAI22_X1 U1515 ( .A1(n1031), .A2(n1915), .B1(n997), .B2(n1916), .ZN(n2529)
         );
  OAI22_X1 U1516 ( .A1(n1099), .A2(n1917), .B1(n1064), .B2(n1918), .ZN(n2528)
         );
  OAI22_X1 U1517 ( .A1(n145), .A2(n1919), .B1(n110), .B2(n1920), .ZN(n2527) );
  OAI22_X1 U1518 ( .A1(n2531), .A2(n1867), .B1(n1868), .B2(n1788), .ZN(N4492)
         );
  NOR4_X1 U1519 ( .A1(n2536), .A2(n2537), .A3(n2538), .A4(n2539), .ZN(n2535)
         );
  OAI22_X1 U1520 ( .A1(n75), .A2(n1877), .B1(n459), .B2(n1878), .ZN(n2539) );
  OAI22_X1 U1521 ( .A1(n233), .A2(n1879), .B1(n201), .B2(n1880), .ZN(n2538) );
  OAI22_X1 U1522 ( .A1(n297), .A2(n1881), .B1(n265), .B2(n1882), .ZN(n2537) );
  OAI22_X1 U1523 ( .A1(n361), .A2(n39), .B1(n329), .B2(n1884), .ZN(n2536) );
  NOR4_X1 U1524 ( .A1(n2540), .A2(n2541), .A3(n2542), .A4(n2543), .ZN(n2534)
         );
  OAI22_X1 U1525 ( .A1(n425), .A2(n1889), .B1(n393), .B2(n1890), .ZN(n2543) );
  OAI22_X1 U1526 ( .A1(n492), .A2(n1891), .B1(n458), .B2(n1892), .ZN(n2542) );
  OAI22_X1 U1527 ( .A1(n559), .A2(n1893), .B1(n526), .B2(n1894), .ZN(n2541) );
  OAI22_X1 U1528 ( .A1(n626), .A2(n1895), .B1(n593), .B2(n1896), .ZN(n2540) );
  NOR4_X1 U1529 ( .A1(n2544), .A2(n2545), .A3(n2546), .A4(n2547), .ZN(n2533)
         );
  OAI22_X1 U1530 ( .A1(n694), .A2(n1901), .B1(n660), .B2(n1902), .ZN(n2547) );
  OAI22_X1 U1531 ( .A1(n761), .A2(n1903), .B1(n727), .B2(n1904), .ZN(n2546) );
  OAI22_X1 U1532 ( .A1(n828), .A2(n1905), .B1(n794), .B2(n1906), .ZN(n2545) );
  OAI22_X1 U1533 ( .A1(n895), .A2(n1907), .B1(n862), .B2(n1908), .ZN(n2544) );
  NOR4_X1 U1534 ( .A1(n2548), .A2(n2549), .A3(n2550), .A4(n2551), .ZN(n2532)
         );
  OAI22_X1 U1535 ( .A1(n962), .A2(n1913), .B1(n929), .B2(n1914), .ZN(n2551) );
  OAI22_X1 U1536 ( .A1(n1030), .A2(n1915), .B1(n996), .B2(n1916), .ZN(n2550)
         );
  OAI22_X1 U1537 ( .A1(n1098), .A2(n1917), .B1(n1063), .B2(n1918), .ZN(n2549)
         );
  OAI22_X1 U1538 ( .A1(n144), .A2(n1919), .B1(n108), .B2(n1920), .ZN(n2548) );
  OAI22_X1 U1539 ( .A1(n2552), .A2(n1867), .B1(n1868), .B2(n1810), .ZN(N4490)
         );
  AOI221_X1 U1540 ( .B1(ADD_WR[1]), .B2(n2555), .C1(n1823), .C2(ADD_RD1[1]), 
        .A(n2556), .ZN(n2554) );
  OAI221_X1 U1541 ( .B1(n1825), .B2(ADD_RD1[2]), .C1(n1826), .C2(ADD_RD1[0]), 
        .A(n2557), .ZN(n2556) );
  AOI22_X1 U1542 ( .A1(n1825), .A2(ADD_RD1[2]), .B1(n1826), .B2(ADD_RD1[0]), 
        .ZN(n2557) );
  AOI221_X1 U1543 ( .B1(n2558), .B2(ADD_WR[4]), .C1(n1829), .C2(ADD_RD1[3]), 
        .A(n2559), .ZN(n2553) );
  OAI22_X1 U1544 ( .A1(ADD_WR[4]), .A2(n2558), .B1(n1829), .B2(ADD_RD1[3]), 
        .ZN(n2559) );
  NOR4_X1 U1545 ( .A1(n2568), .A2(n2569), .A3(n2570), .A4(n2571), .ZN(n2567)
         );
  OAI22_X1 U1546 ( .A1(n53), .A2(n1877), .B1(n438), .B2(n1878), .ZN(n2571) );
  OAI22_X1 U1547 ( .A1(n232), .A2(n1879), .B1(n200), .B2(n1880), .ZN(n2570) );
  OAI22_X1 U1548 ( .A1(n296), .A2(n1881), .B1(n264), .B2(n1882), .ZN(n2569) );
  OAI22_X1 U1549 ( .A1(n360), .A2(n39), .B1(n328), .B2(n1884), .ZN(n2568) );
  NOR3_X1 U1550 ( .A1(n2558), .A2(n2578), .A3(n2579), .ZN(n2573) );
  NAND2_X1 U1551 ( .A1(ADD_RD1[4]), .A2(ADD_RD1[3]), .ZN(n2580) );
  NOR4_X1 U1552 ( .A1(n2581), .A2(n2582), .A3(n2583), .A4(n2584), .ZN(n2566)
         );
  OAI22_X1 U1553 ( .A1(n424), .A2(n1889), .B1(n392), .B2(n1890), .ZN(n2584) );
  OAI22_X1 U1554 ( .A1(n491), .A2(n1891), .B1(n457), .B2(n1892), .ZN(n2583) );
  OAI22_X1 U1555 ( .A1(n558), .A2(n1893), .B1(n525), .B2(n1894), .ZN(n2582) );
  OAI22_X1 U1556 ( .A1(n625), .A2(n1895), .B1(n592), .B2(n1896), .ZN(n2581) );
  NOR3_X1 U1557 ( .A1(ADD_RD1[3]), .A2(n2558), .A3(n2579), .ZN(n2585) );
  NOR3_X1 U1558 ( .A1(ADD_RD1[3]), .A2(ADD_RD1[0]), .A3(n2558), .ZN(n2586) );
  NOR4_X1 U1559 ( .A1(n2587), .A2(n2588), .A3(n2589), .A4(n2590), .ZN(n2565)
         );
  OAI22_X1 U1560 ( .A1(n693), .A2(n1901), .B1(n659), .B2(n1902), .ZN(n2590) );
  OAI22_X1 U1561 ( .A1(n760), .A2(n1903), .B1(n726), .B2(n1904), .ZN(n2589) );
  OAI22_X1 U1562 ( .A1(n827), .A2(n1905), .B1(n793), .B2(n1906), .ZN(n2588) );
  OAI22_X1 U1563 ( .A1(n894), .A2(n1907), .B1(n861), .B2(n1908), .ZN(n2587) );
  NOR3_X1 U1564 ( .A1(ADD_RD1[4]), .A2(n2578), .A3(n2579), .ZN(n2591) );
  NOR3_X1 U1565 ( .A1(ADD_RD1[4]), .A2(ADD_RD1[0]), .A3(n2578), .ZN(n2592) );
  NOR4_X1 U1566 ( .A1(n2593), .A2(n2594), .A3(n2595), .A4(n2596), .ZN(n2564)
         );
  OAI22_X1 U1567 ( .A1(n961), .A2(n1913), .B1(n928), .B2(n1914), .ZN(n2596) );
  OAI22_X1 U1568 ( .A1(n1029), .A2(n1915), .B1(n995), .B2(n1916), .ZN(n2595)
         );
  OAI22_X1 U1569 ( .A1(n1097), .A2(n1917), .B1(n1062), .B2(n1918), .ZN(n2594)
         );
  NAND2_X1 U1570 ( .A1(n2576), .A2(n2597), .ZN(n1918) );
  NAND2_X1 U1571 ( .A1(n2598), .A2(n2576), .ZN(n1917) );
  OAI22_X1 U1572 ( .A1(n143), .A2(n45), .B1(n107), .B2(n1920), .ZN(n2593) );
  NOR3_X1 U1573 ( .A1(ADD_RD1[4]), .A2(ADD_RD1[3]), .A3(n2579), .ZN(n2597) );
  NAND2_X1 U1574 ( .A1(n2598), .A2(n2577), .ZN(n1919) );
  NOR3_X1 U1575 ( .A1(ADD_RD1[4]), .A2(ADD_RD1[3]), .A3(ADD_RD1[0]), .ZN(n2598) );
  OAI21_X1 U1576 ( .B1(n2599), .B2(n2600), .A(n47), .ZN(N4423) );
  OAI21_X1 U1577 ( .B1(n2600), .B2(n2601), .A(n47), .ZN(N4359) );
  OAI21_X1 U1578 ( .B1(n2600), .B2(n2602), .A(n47), .ZN(N4295) );
  OAI21_X1 U1579 ( .B1(n2600), .B2(n2603), .A(n47), .ZN(N4231) );
  OAI21_X1 U1580 ( .B1(n2600), .B2(n2604), .A(n47), .ZN(N4167) );
  OAI21_X1 U1581 ( .B1(n2600), .B2(n2605), .A(n47), .ZN(N4103) );
  OAI21_X1 U1582 ( .B1(n2600), .B2(n2606), .A(n47), .ZN(N4039) );
  NAND2_X1 U1583 ( .A1(n2561), .A2(WR), .ZN(n2600) );
  NOR2_X1 U1584 ( .A1(ADD_WR[4]), .A2(ADD_WR[3]), .ZN(n2561) );
  OAI21_X1 U1585 ( .B1(n2563), .B2(n2607), .A(n49), .ZN(N3975) );
  OAI21_X1 U1586 ( .B1(n2599), .B2(n2607), .A(n51), .ZN(N3911) );
  OAI21_X1 U1587 ( .B1(n2607), .B2(n2601), .A(n49), .ZN(N3847) );
  OAI21_X1 U1588 ( .B1(n2607), .B2(n2602), .A(n49), .ZN(N3783) );
  OAI21_X1 U1589 ( .B1(n2607), .B2(n2603), .A(n49), .ZN(N3719) );
  OAI21_X1 U1590 ( .B1(n2607), .B2(n2604), .A(n49), .ZN(N3655) );
  OAI21_X1 U1591 ( .B1(n2607), .B2(n2605), .A(n49), .ZN(N3591) );
  OAI21_X1 U1592 ( .B1(n2607), .B2(n2606), .A(n49), .ZN(N3527) );
  INV_X1 U1593 ( .A(WR), .ZN(n2562) );
  OAI21_X1 U1594 ( .B1(n2563), .B2(n2608), .A(n49), .ZN(N3463) );
  OAI21_X1 U1595 ( .B1(n2599), .B2(n2608), .A(n47), .ZN(N3399) );
  OAI21_X1 U1596 ( .B1(n2608), .B2(n2601), .A(n49), .ZN(N3335) );
  OAI21_X1 U1597 ( .B1(n2608), .B2(n2602), .A(n49), .ZN(N3271) );
  OAI21_X1 U1598 ( .B1(n2608), .B2(n2603), .A(n47), .ZN(N3207) );
  OAI21_X1 U1599 ( .B1(n2608), .B2(n2604), .A(n47), .ZN(N3143) );
  OAI21_X1 U1600 ( .B1(n2608), .B2(n2605), .A(n51), .ZN(N3079) );
  OAI21_X1 U1601 ( .B1(n2608), .B2(n2606), .A(n49), .ZN(N3015) );
  NAND3_X1 U1602 ( .A1(ADD_WR[4]), .A2(WR), .A3(n1829), .ZN(n2608) );
  OAI21_X1 U1603 ( .B1(n2563), .B2(n2609), .A(n51), .ZN(N2951) );
  NAND3_X1 U1604 ( .A1(n1826), .A2(n1825), .A3(n1823), .ZN(n2563) );
  OAI21_X1 U1605 ( .B1(n2599), .B2(n2609), .A(n49), .ZN(N2887) );
  NAND3_X1 U1606 ( .A1(ADD_WR[0]), .A2(n1825), .A3(n1823), .ZN(n2599) );
  OAI21_X1 U1607 ( .B1(n2609), .B2(n2601), .A(n47), .ZN(N2823) );
  NAND3_X1 U1608 ( .A1(ADD_WR[1]), .A2(n1826), .A3(n1825), .ZN(n2601) );
  OAI21_X1 U1609 ( .B1(n2609), .B2(n2602), .A(n47), .ZN(N2759) );
  NAND3_X1 U1610 ( .A1(ADD_WR[0]), .A2(ADD_WR[1]), .A3(n1825), .ZN(n2602) );
  OAI21_X1 U1611 ( .B1(n2609), .B2(n2603), .A(n51), .ZN(N2695) );
  NAND3_X1 U1612 ( .A1(ADD_WR[2]), .A2(n1826), .A3(n1823), .ZN(n2603) );
  OAI21_X1 U1613 ( .B1(n2609), .B2(n2604), .A(n49), .ZN(N2631) );
  NAND3_X1 U1614 ( .A1(ADD_WR[2]), .A2(ADD_WR[0]), .A3(n1823), .ZN(n2604) );
  OAI21_X1 U1615 ( .B1(n2609), .B2(n2605), .A(n49), .ZN(N2567) );
  NAND3_X1 U1616 ( .A1(ADD_WR[2]), .A2(ADD_WR[1]), .A3(n1826), .ZN(n2605) );
  OAI21_X1 U1617 ( .B1(n2609), .B2(n2606), .A(n51), .ZN(N2503) );
  NAND3_X1 U1618 ( .A1(ADD_WR[0]), .A2(ADD_WR[2]), .A3(ADD_WR[1]), .ZN(n2606)
         );
  NAND3_X1 U1619 ( .A1(ADD_WR[4]), .A2(ADD_WR[3]), .A3(WR), .ZN(n2609) );
endmodule



    module dlx_cu_MICROCODE_MEM_SIZE64_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE13 ( 
        Clk, Rst, IR_IN, stall_exe_i, mispredict_i, D1_i, D2_i, S1_LATCH_EN, 
        S2_LATCH_EN, S3_LATCH_EN, S_MUX_PC_BUS, S_EXT, S_EXT_SIGN, S_EQ_NEQ, 
        S_MUX_DEST, S_MUX_LINK, S_MUX_MEM, S_MEM_W_R, S_MEM_EN, S_RF_W_wb, 
        S_RF_W_mem, S_RF_W_exe, S_MUX_ALUIN, stall_exe_o, stall_dec_o, 
        stall_fetch_o, stall_btb_o, was_branch_o, was_jmp_o, ALU_WORD_o, 
    .ALU_OPCODE({\ALU_OPCODE[4] , \ALU_OPCODE[3] , \ALU_OPCODE[2] , 
        \ALU_OPCODE[1] , \ALU_OPCODE[0] }) );
  input [31:0] IR_IN;
  input [4:0] D1_i;
  input [4:0] D2_i;
  output [1:0] S_MUX_PC_BUS;
  output [1:0] S_MUX_DEST;
  output [12:0] ALU_WORD_o;
  input Clk, Rst, stall_exe_i, mispredict_i;
  output S1_LATCH_EN, S2_LATCH_EN, S3_LATCH_EN, S_EXT, S_EXT_SIGN, S_EQ_NEQ,
         S_MUX_LINK, S_MUX_MEM, S_MEM_W_R, S_MEM_EN, S_RF_W_wb, S_RF_W_mem,
         S_RF_W_exe, S_MUX_ALUIN, stall_exe_o, stall_dec_o, stall_fetch_o,
         stall_btb_o, was_branch_o, was_jmp_o, \ALU_OPCODE[4] ,
         \ALU_OPCODE[3] , \ALU_OPCODE[2] , \ALU_OPCODE[1] , \ALU_OPCODE[0] ;
  wire   IR_IN_10, IR_IN_9, IR_IN_8, IR_IN_7, IR_IN_6, IR_IN_5, IR_IN_4,
         IR_IN_3, IR_IN_2, IR_IN_1, IR_IN_0, stall_exe_i, n122, S_MEM_LOAD,
         S_EXE_LOAD, next_bubble_dec, stall_dec_o_TEMP, stall_btb_o_TEMP,
         stall_fetch_o_TEMP, N20, N21, N22, N23, N24, N25, N26, N27, N29, N30,
         N31, N32, net338222, n2, n3, n4, n5, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n65, n70, n71, n72, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n101, n103, n113, n114, n115, n1,
         n6, n7, n62, n63, n64, n66, n67, n69, n73;
  wire   [12:0] cw_from_mem;
  wire   [4:0] aluOpcode_d;
  assign IR_IN_10 = IR_IN[10];
  assign IR_IN_9 = IR_IN[9];
  assign IR_IN_8 = IR_IN[8];
  assign IR_IN_7 = IR_IN[7];
  assign IR_IN_6 = IR_IN[6];
  assign IR_IN_5 = IR_IN[5];
  assign IR_IN_4 = IR_IN[4];
  assign IR_IN_3 = IR_IN[3];
  assign IR_IN_2 = IR_IN[2];
  assign IR_IN_1 = IR_IN[1];
  assign IR_IN_0 = IR_IN[0];
  assign stall_exe_o = stall_exe_i;

  DFF_X1 bubble_dec_reg ( .D(n113), .CK(Clk), .Q(n69), .QN(n114) );
  DFFR_X1 \cw_e_reg[0]  ( .D(N21), .CK(net338222), .RN(n73), .Q(n122), .QN(n2)
         );
  DFFR_X1 \cw_e_reg[6]  ( .D(N27), .CK(net338222), .RN(n73), .Q(S_MUX_ALUIN)
         );
  DFFR_X1 \cw_e_reg[5]  ( .D(N26), .CK(net338222), .RN(n73), .Q(S_MUX_DEST[1])
         );
  DFFR_X1 \cw_e_reg[4]  ( .D(N25), .CK(net338222), .RN(n73), .Q(S_MUX_DEST[0])
         );
  DFFR_X1 \cw_e_reg[3]  ( .D(N24), .CK(net338222), .RN(n73), .Q(n3) );
  DFFR_X1 \cw_e_reg[2]  ( .D(N23), .CK(net338222), .RN(n73), .QN(n4) );
  DFFR_X1 \cw_e_reg[1]  ( .D(N22), .CK(net338222), .RN(n73), .QN(n5) );
  DFFR_X1 \cw_m_reg[2]  ( .D(N31), .CK(Clk), .RN(n73), .Q(S_MEM_W_R) );
  DFFR_X1 \cw_m_reg[3]  ( .D(N32), .CK(Clk), .RN(n73), .Q(S_MEM_EN), .QN(n115)
         );
  DFFR_X1 \cw_m_reg[0]  ( .D(N29), .CK(Clk), .RN(n73), .Q(S_RF_W_mem), .QN(
        n103) );
  DFFS_X1 \cw_w_reg[0]  ( .D(n103), .CK(Clk), .SN(n73), .QN(S_RF_W_wb) );
  XOR2_X1 U3 ( .A(S_MUX_PC_BUS[1]), .B(S_MUX_PC_BUS[0]), .Z(was_jmp_o) );
  MUX2_X1 U8 ( .A(n69), .B(next_bubble_dec), .S(n73), .Z(n113) );
  NAND3_X1 U13 ( .A1(n19), .A2(IR_IN[28]), .A3(n20), .ZN(n18) );
  NAND3_X1 U24 ( .A1(n34), .A2(n43), .A3(n21), .ZN(n42) );
  NAND3_X1 U60 ( .A1(IR_IN[30]), .A2(IR_IN[29]), .A3(n72), .ZN(n58) );
  NAND3_X1 U78 ( .A1(IR_IN_5), .A2(IR_IN_4), .A3(n61), .ZN(n54) );
  NAND3_X1 U92 ( .A1(n97), .A2(n93), .A3(n21), .ZN(n41) );
  stall_logic_FUNC_SIZE11_OP_CODE_SIZE6 STALL_L ( .OPCODE_i(IR_IN[31:26]), 
        .FUNC_i({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .rA_i(IR_IN[25:21]), .rB_i(IR_IN[20:16]), .D1_i(D1_i), .D2_i(
        D2_i), .S_mem_LOAD_i(S_MEM_LOAD), .S_exe_LOAD_i(S_EXE_LOAD), 
        .S_exe_WRITE_i(n122), .S_MUX_PC_BUS_i({1'b0, 1'b0}), .mispredict_i(
        mispredict_i), .bubble_dec_o(next_bubble_dec), .stall_dec_o(
        stall_dec_o_TEMP), .stall_btb_o(stall_btb_o_TEMP), .stall_fetch_o(
        stall_fetch_o_TEMP) );
  cw_mem_MICROCODE_MEM_SIZE64_OP_CODE_SIZE6_CW_SIZE13 CWM ( .OPCODE_IN(
        IR_IN[31:26]), .CW_OUT(cw_from_mem) );
  alu_ctrl ALU_C ( .OP(aluOpcode_d), .ALU_WORD(ALU_WORD_o) );
  SNPS_CLOCK_GATE_HIGH_dlx_cu_MICROCODE_MEM_SIZE64_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE13_0 clk_gate_cw_e_reg ( 
        .CLK(Clk), .EN(N20), .ENCLK(net338222) );
  AND2_X1 U111 ( .A1(n114), .A2(cw_from_mem[9]), .ZN(S_EXT_SIGN) );
  AND2_X1 U114 ( .A1(n114), .A2(cw_from_mem[8]), .ZN(S_EQ_NEQ) );
  NOR2_X1 U109 ( .A1(n115), .A2(S_MEM_W_R), .ZN(S_MEM_LOAD) );
  NAND2_X1 U47 ( .A1(IR_IN_4), .A2(IR_IN_5), .ZN(n8) );
  NOR3_X1 U98 ( .A1(IR_IN[31]), .A2(IR_IN[28]), .A3(IR_IN[30]), .ZN(n89) );
  NOR4_X1 U97 ( .A1(IR_IN_7), .A2(IR_IN_6), .A3(IR_IN[27]), .A4(IR_IN_10), 
        .ZN(n99) );
  NAND2_X1 U96 ( .A1(n89), .A2(n99), .ZN(n98) );
  NOR4_X1 U95 ( .A1(IR_IN_9), .A2(IR_IN_8), .A3(IR_IN[29]), .A4(n98), .ZN(n92)
         );
  NAND2_X1 U94 ( .A1(n44), .A2(n92), .ZN(n49) );
  NOR3_X1 U74 ( .A1(IR_IN_5), .A2(n39), .A3(n75), .ZN(n82) );
  NAND4_X1 U73 ( .A1(n92), .A2(IR_IN[26]), .A3(n82), .A4(n61), .ZN(n47) );
  AOI221_X1 U26 ( .B1(IR_IN_4), .B2(IR_IN_3), .C1(n45), .C2(n46), .A(n47), 
        .ZN(n29) );
  NOR2_X1 U70 ( .A1(n39), .A2(IR_IN_1), .ZN(n60) );
  NOR2_X1 U68 ( .A1(n46), .A2(n25), .ZN(n34) );
  NAND2_X1 U20 ( .A1(n21), .A2(n34), .ZN(n15) );
  NOR3_X1 U100 ( .A1(IR_IN_2), .A2(n46), .A3(n75), .ZN(n93) );
  NAND2_X1 U77 ( .A1(n21), .A2(n93), .ZN(n31) );
  INV_X1 U61 ( .A(IR_IN[28]), .ZN(n57) );
  NAND2_X1 U85 ( .A1(IR_IN[30]), .A2(IR_IN[29]), .ZN(n96) );
  NOR3_X1 U84 ( .A1(IR_IN[28]), .A2(n72), .A3(n96), .ZN(n33) );
  OAI21_X1 U19 ( .B1(n12), .B2(n33), .A(IR_IN[31]), .ZN(n32) );
  OAI221_X1 U18 ( .B1(n8), .B2(n15), .C1(n8), .C2(n31), .A(n32), .ZN(n30) );
  NOR2_X1 U17 ( .A1(n29), .A2(n30), .ZN(n10) );
  NOR2_X1 U56 ( .A1(n61), .A2(n26), .ZN(n14) );
  AOI22_X1 U10 ( .A1(IR_IN[26]), .A2(n12), .B1(n13), .B2(n14), .ZN(n11) );
  OAI211_X1 U9 ( .C1(n8), .C2(n9), .A(n10), .B(n11), .ZN(aluOpcode_d[4]) );
  INV_X1 U91 ( .A(IR_IN[31]), .ZN(n55) );
  NAND2_X1 U90 ( .A1(IR_IN[29]), .A2(n55), .ZN(n56) );
  NOR2_X1 U35 ( .A1(IR_IN[28]), .A2(n56), .ZN(n27) );
  NOR2_X1 U48 ( .A1(IR_IN_0), .A2(n26), .ZN(n43) );
  NOR2_X1 U46 ( .A1(n8), .A2(n61), .ZN(n50) );
  OAI221_X1 U28 ( .B1(n43), .B2(IR_IN_1), .C1(n43), .C2(n50), .A(n46), .ZN(n48) );
  NOR2_X1 U27 ( .A1(n48), .A2(n49), .ZN(n28) );
  AOI22_X1 U16 ( .A1(IR_IN[30]), .A2(n27), .B1(IR_IN_2), .B2(n28), .ZN(n16) );
  NOR4_X1 U71 ( .A1(IR_IN_1), .A2(IR_IN_2), .A3(n46), .A4(n26), .ZN(n22) );
  NOR3_X1 U15 ( .A1(n25), .A2(n26), .A3(n9), .ZN(n23) );
  AOI21_X1 U25 ( .B1(n12), .B2(n44), .A(n33), .ZN(n40) );
  OAI211_X1 U23 ( .C1(n40), .C2(IR_IN[31]), .A(n41), .B(n42), .ZN(n24) );
  AOI211_X1 U14 ( .C1(n21), .C2(n22), .A(n23), .B(n24), .ZN(n17) );
  NOR2_X1 U89 ( .A1(IR_IN[30]), .A2(n56), .ZN(n19) );
  NAND2_X1 U63 ( .A1(IR_IN[26]), .A2(IR_IN[27]), .ZN(n20) );
  NAND4_X1 U12 ( .A1(n10), .A2(n16), .A3(n17), .A4(n18), .ZN(aluOpcode_d[3])
         );
  NOR3_X1 U65 ( .A1(IR_IN_2), .A2(n61), .A3(n26), .ZN(n59) );
  OAI221_X1 U36 ( .B1(n59), .B2(n60), .C1(n59), .C2(n50), .A(n21), .ZN(n35) );
  OAI221_X1 U33 ( .B1(n27), .B2(IR_IN[31]), .C1(n27), .C2(n12), .A(IR_IN[26]), 
        .ZN(n36) );
  NOR2_X1 U32 ( .A1(IR_IN[28]), .A2(IR_IN[30]), .ZN(n51) );
  OAI21_X1 U31 ( .B1(n55), .B2(n20), .A(n56), .ZN(n52) );
  NOR3_X1 U30 ( .A1(n39), .A2(n54), .A3(n9), .ZN(n53) );
  AOI21_X1 U29 ( .B1(n51), .B2(n52), .A(n53), .ZN(n37) );
  AOI211_X1 U22 ( .C1(n28), .C2(n39), .A(n29), .B(n24), .ZN(n38) );
  NOR2_X1 U87 ( .A1(IR_IN[27]), .A2(n71), .ZN(n94) );
  INV_X1 U83 ( .A(IR_IN[29]), .ZN(n91) );
  NAND4_X1 U82 ( .A1(IR_IN[28]), .A2(IR_IN[30]), .A3(n55), .A4(n91), .ZN(n70)
         );
  AOI221_X1 U81 ( .B1(IR_IN[27]), .B2(n44), .C1(n72), .C2(IR_IN[26]), .A(n70), 
        .ZN(n95) );
  AOI221_X1 U80 ( .B1(n94), .B2(IR_IN[26]), .C1(n33), .C2(n44), .A(n95), .ZN(
        n76) );
  NOR2_X1 U76 ( .A1(n54), .A2(n31), .ZN(n78) );
  NOR3_X1 U72 ( .A1(IR_IN_3), .A2(n45), .A3(n47), .ZN(n79) );
  OAI221_X1 U67 ( .B1(n22), .B2(n34), .C1(n22), .C2(IR_IN_5), .A(n61), .ZN(n85) );
  OAI211_X1 U64 ( .C1(n84), .C2(n59), .A(IR_IN_1), .B(n46), .ZN(n86) );
  NOR2_X1 U62 ( .A1(n91), .A2(n20), .ZN(n88) );
  AOI211_X1 U59 ( .C1(IR_IN[31]), .C2(n57), .A(IR_IN[26]), .B(n58), .ZN(n90)
         );
  AOI21_X1 U58 ( .B1(n88), .B2(n89), .A(n90), .ZN(n87) );
  OAI221_X1 U57 ( .B1(n49), .B2(n85), .C1(n49), .C2(n86), .A(n87), .ZN(n65) );
  NOR4_X1 U55 ( .A1(IR_IN_4), .A2(IR_IN_5), .A3(IR_IN_0), .A4(n25), .ZN(n83)
         );
  AOI211_X1 U54 ( .C1(n14), .C2(n75), .A(n83), .B(n84), .ZN(n81) );
  NAND2_X1 U53 ( .A1(n82), .A2(n45), .ZN(n74) );
  AOI221_X1 U51 ( .B1(n61), .B2(n81), .C1(n74), .C2(n81), .A(n9), .ZN(n80) );
  NOR4_X1 U50 ( .A1(n78), .A2(n79), .A3(n65), .A4(n80), .ZN(n77) );
  OAI211_X1 U49 ( .C1(IR_IN_0), .C2(n41), .A(n76), .B(n77), .ZN(aluOpcode_d[0]) );
  NOR2_X1 U118 ( .A1(n5), .A2(stall_exe_i), .ZN(N30) );
  NOR2_X1 U117 ( .A1(n4), .A2(stall_exe_i), .ZN(N31) );
  NOR2_X1 U119 ( .A1(n2), .A2(stall_exe_i), .ZN(N29) );
  INV_X1 U99 ( .A(IR_IN[26]), .ZN(n44) );
  NAND2_X1 U52 ( .A1(n21), .A2(n46), .ZN(n9) );
  NOR2_X1 U34 ( .A1(n57), .A2(n58), .ZN(n12) );
  NAND2_X1 U104 ( .A1(IR_IN_5), .A2(n45), .ZN(n26) );
  NAND4_X1 U21 ( .A1(n35), .A2(n36), .A3(n37), .A4(n38), .ZN(aluOpcode_d[2])
         );
  NOR2_X1 U127 ( .A1(stall_dec_o_TEMP), .A2(n69), .ZN(n101) );
  AND2_X1 U106 ( .A1(cw_from_mem[12]), .A2(n114), .ZN(S_MUX_PC_BUS[1]) );
  AND2_X1 U112 ( .A1(n114), .A2(cw_from_mem[10]), .ZN(S_EXT) );
  INV_X1 U86 ( .A(IR_IN[27]), .ZN(n72) );
  AND2_X1 U4 ( .A1(S_MUX_PC_BUS[1]), .A2(S_MUX_PC_BUS[0]), .ZN(was_branch_o)
         );
  AND2_X1 U113 ( .A1(n4), .A2(n3), .ZN(S_EXE_LOAD) );
  OR2_X1 U6 ( .A1(stall_exe_i), .A2(stall_dec_o_TEMP), .ZN(stall_dec_o) );
  OR2_X1 U5 ( .A1(stall_exe_i), .A2(stall_fetch_o_TEMP), .ZN(stall_fetch_o) );
  INV_X1 U93 ( .A(n49), .ZN(n21) );
  INV_X1 U102 ( .A(IR_IN_3), .ZN(n46) );
  INV_X1 U105 ( .A(IR_IN_4), .ZN(n45) );
  INV_X1 U75 ( .A(IR_IN_2), .ZN(n39) );
  INV_X1 U101 ( .A(IR_IN_1), .ZN(n75) );
  INV_X1 U79 ( .A(IR_IN_0), .ZN(n61) );
  INV_X1 U69 ( .A(n60), .ZN(n25) );
  INV_X1 U11 ( .A(n15), .ZN(n13) );
  INV_X1 U103 ( .A(n26), .ZN(n97) );
  INV_X1 U88 ( .A(n19), .ZN(n71) );
  INV_X1 U66 ( .A(n54), .ZN(n84) );
  AND2_X1 U122 ( .A1(n101), .A2(cw_from_mem[4]), .ZN(N25) );
  AND2_X1 U125 ( .A1(n101), .A2(cw_from_mem[1]), .ZN(N22) );
  AND2_X1 U120 ( .A1(n101), .A2(cw_from_mem[6]), .ZN(N27) );
  AND2_X1 U121 ( .A1(n101), .A2(cw_from_mem[5]), .ZN(N26) );
  AND2_X1 U123 ( .A1(n101), .A2(cw_from_mem[3]), .ZN(N24) );
  AND2_X1 U124 ( .A1(n101), .A2(cw_from_mem[2]), .ZN(N23) );
  AND2_X1 U126 ( .A1(n101), .A2(cw_from_mem[0]), .ZN(N21) );
  AND2_X1 U116 ( .A1(N20), .A2(n3), .ZN(N32) );
  DFFR_X2 \cw_m_reg[1]  ( .D(N30), .CK(Clk), .RN(n73), .Q(S_MUX_MEM) );
  AND2_X1 U107 ( .A1(n114), .A2(cw_from_mem[11]), .ZN(S_MUX_PC_BUS[0]) );
  OR2_X1 U7 ( .A1(stall_exe_i), .A2(stall_btb_o_TEMP), .ZN(stall_btb_o) );
  OAI21_X1 U37 ( .B1(IR_IN[26]), .B2(n71), .A(n70), .ZN(n1) );
  INV_X1 U38 ( .A(n72), .ZN(n6) );
  INV_X1 U39 ( .A(n31), .ZN(n7) );
  AOI222_X1 U40 ( .A1(n1), .A2(n6), .B1(IR_IN[26]), .B2(n33), .C1(n7), .C2(n50), .ZN(n62) );
  AOI22_X1 U41 ( .A1(IR_IN_1), .A2(n43), .B1(n50), .B2(n75), .ZN(n63) );
  AOI21_X1 U42 ( .B1(n74), .B2(n63), .A(n9), .ZN(n64) );
  NOR3_X1 U43 ( .A1(n46), .A2(n47), .A3(IR_IN_4), .ZN(n66) );
  NOR3_X1 U44 ( .A1(n65), .A2(n64), .A3(n66), .ZN(n67) );
  OAI211_X1 U45 ( .C1(n61), .C2(n41), .A(n62), .B(n67), .ZN(aluOpcode_d[1]) );
  AND2_X2 U108 ( .A1(n114), .A2(cw_from_mem[7]), .ZN(S_MUX_LINK) );
  INV_X1 U110 ( .A(stall_exe_i), .ZN(N20) );
  INV_X1 U115 ( .A(Rst), .ZN(n73) );
endmodule


module jump_logic ( NPCF_i, IR_i, A_i, A_o, rA_o, rB_o, rC_o, branch_target_o, 
        sum_addr_o, extended_imm, taken_o, FW_X_i, FW_W_i, S_FW_Adec_i, 
        S_EXT_i, S_EXT_SIGN_i, S_MUX_LINK_i, S_EQ_NEQ_i );
  input [31:0] NPCF_i;
  input [31:0] IR_i;
  input [31:0] A_i;
  output [31:0] A_o;
  output [4:0] rA_o;
  output [4:0] rB_o;
  output [4:0] rC_o;
  output [31:0] branch_target_o;
  output [31:0] sum_addr_o;
  output [31:0] extended_imm;
  input [31:0] FW_X_i;
  input [31:0] FW_W_i;
  input [1:0] S_FW_Adec_i;
  input S_EXT_i, S_EXT_SIGN_i, S_MUX_LINK_i, S_EQ_NEQ_i;
  output taken_o;
  wire   \IR_i[25] , \IR_i[24] , \IR_i[23] , \IR_i[22] , \IR_i[21] ,
         \IR_i[20] , \IR_i[19] , \IR_i[18] , \IR_i[17] , \IR_i[16] ,
         \IR_i[15] , \IR_i[14] , \IR_i[13] , \IR_i[12] , \IR_i[11] ,
         branch_sel;
  wire   [31:0] ext_imm;
  assign rA_o[4] = \IR_i[25] ;
  assign \IR_i[25]  = IR_i[25];
  assign rA_o[3] = \IR_i[24] ;
  assign \IR_i[24]  = IR_i[24];
  assign rA_o[2] = \IR_i[23] ;
  assign \IR_i[23]  = IR_i[23];
  assign rA_o[1] = \IR_i[22] ;
  assign \IR_i[22]  = IR_i[22];
  assign rA_o[0] = \IR_i[21] ;
  assign \IR_i[21]  = IR_i[21];
  assign rB_o[4] = \IR_i[20] ;
  assign \IR_i[20]  = IR_i[20];
  assign rB_o[3] = \IR_i[19] ;
  assign \IR_i[19]  = IR_i[19];
  assign rB_o[2] = \IR_i[18] ;
  assign \IR_i[18]  = IR_i[18];
  assign rB_o[1] = \IR_i[17] ;
  assign \IR_i[17]  = IR_i[17];
  assign rB_o[0] = \IR_i[16] ;
  assign \IR_i[16]  = IR_i[16];
  assign rC_o[4] = \IR_i[15] ;
  assign \IR_i[15]  = IR_i[15];
  assign rC_o[3] = \IR_i[14] ;
  assign \IR_i[14]  = IR_i[14];
  assign rC_o[2] = \IR_i[13] ;
  assign \IR_i[13]  = IR_i[13];
  assign rC_o[1] = \IR_i[12] ;
  assign \IR_i[12]  = IR_i[12];
  assign rC_o[0] = \IR_i[11] ;
  assign \IR_i[11]  = IR_i[11];

  extender_32 EXTENDER ( .IN1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, \IR_i[25] , 
        \IR_i[24] , \IR_i[23] , \IR_i[22] , \IR_i[21] , \IR_i[20] , \IR_i[19] , 
        \IR_i[18] , \IR_i[17] , \IR_i[16] , \IR_i[15] , \IR_i[14] , \IR_i[13] , 
        \IR_i[12] , \IR_i[11] , IR_i[10:0]}), .CTRL(S_EXT_i), .SIGN(
        S_EXT_SIGN_i), .OUT1(ext_imm) );
  p4add_N32_logN5_0 JUMPADDER ( .A(NPCF_i), .B(ext_imm), .Cin(1'b0), .sign(
        1'b0), .S(sum_addr_o) );
  mux21_0 BRANCHMUX ( .IN0(sum_addr_o), .IN1(NPCF_i), .CTRL(branch_sel), 
        .OUT1(branch_target_o) );
  zerocheck ZC ( .IN0(A_o), .CTRL(S_EQ_NEQ_i), .OUT1(branch_sel) );
  mux21_4 MUXLINK ( .IN0(ext_imm), .IN1(NPCF_i), .CTRL(S_MUX_LINK_i), .OUT1(
        extended_imm) );
  mux41_MUX_SIZE32_0 MUX_FWA ( .IN0(A_i), .IN1(FW_X_i), .IN2(FW_W_i), .IN3({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CTRL(S_FW_Adec_i), 
        .OUT1(A_o) );
  INV_X1 U2 ( .A(branch_sel), .ZN(taken_o) );
endmodule


module fetch_regs ( NPCF_i, IR_i, NPCF_o, IR_o, stall_i, clk, rst );
  input [31:0] NPCF_i;
  input [31:0] IR_i;
  output [31:0] NPCF_o;
  output [31:0] IR_o;
  input stall_i, clk, rst;
  wire   enable;

  ff32_en_1 NPCF ( .D(NPCF_i), .en(enable), .clk(clk), .rst(rst), .Q(NPCF_o)
         );
  ff32_en_IR IR ( .D(IR_i), .en(enable), .clk(clk), .rst(rst), .Q(IR_o) );
  INV_X1 U1 ( .A(stall_i), .ZN(enable) );
endmodule


module btb_N_LINES4_SIZE32 ( clock, reset, stall_i, TAG_i, target_PC_i, 
        was_taken_i, predicted_next_PC_o, taken_o, mispredict_o );
  input [3:0] TAG_i;
  input [31:0] target_PC_i;
  output [31:0] predicted_next_PC_o;
  input clock, reset, stall_i, was_taken_i;
  output taken_o, mispredict_o;
  wire   \predict_PC[0][31] , \predict_PC[0][30] , \predict_PC[0][29] ,
         \predict_PC[0][28] , \predict_PC[0][27] , \predict_PC[0][26] ,
         \predict_PC[0][25] , \predict_PC[0][24] , \predict_PC[0][23] ,
         \predict_PC[0][22] , \predict_PC[0][21] , \predict_PC[0][20] ,
         \predict_PC[0][19] , \predict_PC[0][18] , \predict_PC[0][17] ,
         \predict_PC[0][16] , \predict_PC[0][15] , \predict_PC[0][14] ,
         \predict_PC[0][13] , \predict_PC[0][12] , \predict_PC[0][11] ,
         \predict_PC[0][10] , \predict_PC[0][9] , \predict_PC[0][8] ,
         \predict_PC[0][7] , \predict_PC[0][6] , \predict_PC[0][5] ,
         \predict_PC[0][4] , \predict_PC[0][3] , \predict_PC[0][2] ,
         \predict_PC[0][1] , \predict_PC[0][0] , \predict_PC[1][31] ,
         \predict_PC[1][30] , \predict_PC[1][29] , \predict_PC[1][28] ,
         \predict_PC[1][27] , \predict_PC[1][26] , \predict_PC[1][25] ,
         \predict_PC[1][24] , \predict_PC[1][23] , \predict_PC[1][22] ,
         \predict_PC[1][21] , \predict_PC[1][20] , \predict_PC[1][19] ,
         \predict_PC[1][18] , \predict_PC[1][17] , \predict_PC[1][16] ,
         \predict_PC[1][15] , \predict_PC[1][14] , \predict_PC[1][13] ,
         \predict_PC[1][12] , \predict_PC[1][11] , \predict_PC[1][10] ,
         \predict_PC[1][9] , \predict_PC[1][8] , \predict_PC[1][7] ,
         \predict_PC[1][6] , \predict_PC[1][5] , \predict_PC[1][4] ,
         \predict_PC[1][3] , \predict_PC[1][2] , \predict_PC[1][1] ,
         \predict_PC[1][0] , \predict_PC[2][31] , \predict_PC[2][30] ,
         \predict_PC[2][29] , \predict_PC[2][28] , \predict_PC[2][27] ,
         \predict_PC[2][26] , \predict_PC[2][25] , \predict_PC[2][24] ,
         \predict_PC[2][23] , \predict_PC[2][22] , \predict_PC[2][21] ,
         \predict_PC[2][20] , \predict_PC[2][19] , \predict_PC[2][18] ,
         \predict_PC[2][17] , \predict_PC[2][16] , \predict_PC[2][15] ,
         \predict_PC[2][14] , \predict_PC[2][13] , \predict_PC[2][12] ,
         \predict_PC[2][11] , \predict_PC[2][10] , \predict_PC[2][9] ,
         \predict_PC[2][8] , \predict_PC[2][7] , \predict_PC[2][6] ,
         \predict_PC[2][5] , \predict_PC[2][4] , \predict_PC[2][3] ,
         \predict_PC[2][2] , \predict_PC[2][1] , \predict_PC[2][0] ,
         \predict_PC[3][31] , \predict_PC[3][30] , \predict_PC[3][29] ,
         \predict_PC[3][28] , \predict_PC[3][27] , \predict_PC[3][26] ,
         \predict_PC[3][25] , \predict_PC[3][24] , \predict_PC[3][23] ,
         \predict_PC[3][22] , \predict_PC[3][21] , \predict_PC[3][20] ,
         \predict_PC[3][19] , \predict_PC[3][18] , \predict_PC[3][17] ,
         \predict_PC[3][16] , \predict_PC[3][15] , \predict_PC[3][14] ,
         \predict_PC[3][13] , \predict_PC[3][12] , \predict_PC[3][11] ,
         \predict_PC[3][10] , \predict_PC[3][9] , \predict_PC[3][8] ,
         \predict_PC[3][7] , \predict_PC[3][6] , \predict_PC[3][5] ,
         \predict_PC[3][4] , \predict_PC[3][3] , \predict_PC[3][2] ,
         \predict_PC[3][1] , \predict_PC[3][0] , \predict_PC[4][31] ,
         \predict_PC[4][30] , \predict_PC[4][29] , \predict_PC[4][28] ,
         \predict_PC[4][27] , \predict_PC[4][26] , \predict_PC[4][25] ,
         \predict_PC[4][24] , \predict_PC[4][23] , \predict_PC[4][22] ,
         \predict_PC[4][21] , \predict_PC[4][20] , \predict_PC[4][19] ,
         \predict_PC[4][18] , \predict_PC[4][17] , \predict_PC[4][16] ,
         \predict_PC[4][15] , \predict_PC[4][14] , \predict_PC[4][13] ,
         \predict_PC[4][12] , \predict_PC[4][11] , \predict_PC[4][10] ,
         \predict_PC[4][9] , \predict_PC[4][8] , \predict_PC[4][7] ,
         \predict_PC[4][6] , \predict_PC[4][5] , \predict_PC[4][4] ,
         \predict_PC[4][3] , \predict_PC[4][2] , \predict_PC[4][1] ,
         \predict_PC[4][0] , \predict_PC[5][31] , \predict_PC[5][30] ,
         \predict_PC[5][29] , \predict_PC[5][28] , \predict_PC[5][27] ,
         \predict_PC[5][26] , \predict_PC[5][25] , \predict_PC[5][24] ,
         \predict_PC[5][23] , \predict_PC[5][22] , \predict_PC[5][21] ,
         \predict_PC[5][20] , \predict_PC[5][19] , \predict_PC[5][18] ,
         \predict_PC[5][17] , \predict_PC[5][16] , \predict_PC[5][15] ,
         \predict_PC[5][14] , \predict_PC[5][13] , \predict_PC[5][12] ,
         \predict_PC[5][11] , \predict_PC[5][10] , \predict_PC[5][9] ,
         \predict_PC[5][8] , \predict_PC[5][7] , \predict_PC[5][6] ,
         \predict_PC[5][5] , \predict_PC[5][4] , \predict_PC[5][3] ,
         \predict_PC[5][2] , \predict_PC[5][1] , \predict_PC[5][0] ,
         \predict_PC[6][31] , \predict_PC[6][30] , \predict_PC[6][29] ,
         \predict_PC[6][28] , \predict_PC[6][27] , \predict_PC[6][26] ,
         \predict_PC[6][25] , \predict_PC[6][24] , \predict_PC[6][23] ,
         \predict_PC[6][22] , \predict_PC[6][21] , \predict_PC[6][20] ,
         \predict_PC[6][19] , \predict_PC[6][18] , \predict_PC[6][17] ,
         \predict_PC[6][16] , \predict_PC[6][15] , \predict_PC[6][14] ,
         \predict_PC[6][13] , \predict_PC[6][12] , \predict_PC[6][11] ,
         \predict_PC[6][10] , \predict_PC[6][9] , \predict_PC[6][8] ,
         \predict_PC[6][7] , \predict_PC[6][6] , \predict_PC[6][5] ,
         \predict_PC[6][4] , \predict_PC[6][3] , \predict_PC[6][2] ,
         \predict_PC[6][1] , \predict_PC[6][0] , \predict_PC[7][31] ,
         \predict_PC[7][30] , \predict_PC[7][29] , \predict_PC[7][28] ,
         \predict_PC[7][27] , \predict_PC[7][26] , \predict_PC[7][25] ,
         \predict_PC[7][24] , \predict_PC[7][23] , \predict_PC[7][22] ,
         \predict_PC[7][21] , \predict_PC[7][20] , \predict_PC[7][19] ,
         \predict_PC[7][18] , \predict_PC[7][17] , \predict_PC[7][16] ,
         \predict_PC[7][15] , \predict_PC[7][14] , \predict_PC[7][13] ,
         \predict_PC[7][12] , \predict_PC[7][11] , \predict_PC[7][10] ,
         \predict_PC[7][9] , \predict_PC[7][8] , \predict_PC[7][7] ,
         \predict_PC[7][6] , \predict_PC[7][5] , \predict_PC[7][4] ,
         \predict_PC[7][3] , \predict_PC[7][2] , \predict_PC[7][1] ,
         \predict_PC[7][0] , \predict_PC[8][31] , \predict_PC[8][30] ,
         \predict_PC[8][29] , \predict_PC[8][28] , \predict_PC[8][27] ,
         \predict_PC[8][26] , \predict_PC[8][25] , \predict_PC[8][24] ,
         \predict_PC[8][23] , \predict_PC[8][22] , \predict_PC[8][21] ,
         \predict_PC[8][20] , \predict_PC[8][19] , \predict_PC[8][18] ,
         \predict_PC[8][17] , \predict_PC[8][16] , \predict_PC[8][15] ,
         \predict_PC[8][14] , \predict_PC[8][13] , \predict_PC[8][12] ,
         \predict_PC[8][11] , \predict_PC[8][10] , \predict_PC[8][9] ,
         \predict_PC[8][8] , \predict_PC[8][7] , \predict_PC[8][6] ,
         \predict_PC[8][5] , \predict_PC[8][4] , \predict_PC[8][3] ,
         \predict_PC[8][2] , \predict_PC[8][1] , \predict_PC[8][0] ,
         \predict_PC[9][31] , \predict_PC[9][30] , \predict_PC[9][29] ,
         \predict_PC[9][28] , \predict_PC[9][27] , \predict_PC[9][26] ,
         \predict_PC[9][25] , \predict_PC[9][24] , \predict_PC[9][23] ,
         \predict_PC[9][22] , \predict_PC[9][21] , \predict_PC[9][20] ,
         \predict_PC[9][19] , \predict_PC[9][18] , \predict_PC[9][17] ,
         \predict_PC[9][16] , \predict_PC[9][15] , \predict_PC[9][14] ,
         \predict_PC[9][13] , \predict_PC[9][12] , \predict_PC[9][11] ,
         \predict_PC[9][10] , \predict_PC[9][9] , \predict_PC[9][8] ,
         \predict_PC[9][7] , \predict_PC[9][6] , \predict_PC[9][5] ,
         \predict_PC[9][4] , \predict_PC[9][3] , \predict_PC[9][2] ,
         \predict_PC[9][1] , \predict_PC[9][0] , \predict_PC[10][31] ,
         \predict_PC[10][30] , \predict_PC[10][29] , \predict_PC[10][28] ,
         \predict_PC[10][27] , \predict_PC[10][26] , \predict_PC[10][25] ,
         \predict_PC[10][24] , \predict_PC[10][23] , \predict_PC[10][22] ,
         \predict_PC[10][21] , \predict_PC[10][20] , \predict_PC[10][19] ,
         \predict_PC[10][18] , \predict_PC[10][17] , \predict_PC[10][16] ,
         \predict_PC[10][15] , \predict_PC[10][14] , \predict_PC[10][13] ,
         \predict_PC[10][12] , \predict_PC[10][11] , \predict_PC[10][10] ,
         \predict_PC[10][9] , \predict_PC[10][8] , \predict_PC[10][7] ,
         \predict_PC[10][6] , \predict_PC[10][5] , \predict_PC[10][4] ,
         \predict_PC[10][3] , \predict_PC[10][2] , \predict_PC[10][1] ,
         \predict_PC[10][0] , \predict_PC[11][31] , \predict_PC[11][30] ,
         \predict_PC[11][29] , \predict_PC[11][28] , \predict_PC[11][27] ,
         \predict_PC[11][26] , \predict_PC[11][25] , \predict_PC[11][24] ,
         \predict_PC[11][23] , \predict_PC[11][22] , \predict_PC[11][21] ,
         \predict_PC[11][20] , \predict_PC[11][19] , \predict_PC[11][18] ,
         \predict_PC[11][17] , \predict_PC[11][16] , \predict_PC[11][15] ,
         \predict_PC[11][14] , \predict_PC[11][13] , \predict_PC[11][12] ,
         \predict_PC[11][11] , \predict_PC[11][10] , \predict_PC[11][9] ,
         \predict_PC[11][8] , \predict_PC[11][7] , \predict_PC[11][6] ,
         \predict_PC[11][5] , \predict_PC[11][4] , \predict_PC[11][3] ,
         \predict_PC[11][2] , \predict_PC[11][1] , \predict_PC[11][0] ,
         \predict_PC[12][31] , \predict_PC[12][30] , \predict_PC[12][29] ,
         \predict_PC[12][28] , \predict_PC[12][27] , \predict_PC[12][26] ,
         \predict_PC[12][25] , \predict_PC[12][24] , \predict_PC[12][23] ,
         \predict_PC[12][22] , \predict_PC[12][21] , \predict_PC[12][20] ,
         \predict_PC[12][19] , \predict_PC[12][18] , \predict_PC[12][17] ,
         \predict_PC[12][16] , \predict_PC[12][15] , \predict_PC[12][14] ,
         \predict_PC[12][13] , \predict_PC[12][12] , \predict_PC[12][11] ,
         \predict_PC[12][10] , \predict_PC[12][9] , \predict_PC[12][8] ,
         \predict_PC[12][7] , \predict_PC[12][6] , \predict_PC[12][5] ,
         \predict_PC[12][4] , \predict_PC[12][3] , \predict_PC[12][2] ,
         \predict_PC[12][1] , \predict_PC[12][0] , \predict_PC[13][31] ,
         \predict_PC[13][30] , \predict_PC[13][29] , \predict_PC[13][28] ,
         \predict_PC[13][27] , \predict_PC[13][26] , \predict_PC[13][25] ,
         \predict_PC[13][24] , \predict_PC[13][23] , \predict_PC[13][22] ,
         \predict_PC[13][21] , \predict_PC[13][20] , \predict_PC[13][19] ,
         \predict_PC[13][18] , \predict_PC[13][17] , \predict_PC[13][16] ,
         \predict_PC[13][15] , \predict_PC[13][14] , \predict_PC[13][13] ,
         \predict_PC[13][12] , \predict_PC[13][11] , \predict_PC[13][10] ,
         \predict_PC[13][9] , \predict_PC[13][8] , \predict_PC[13][7] ,
         \predict_PC[13][6] , \predict_PC[13][5] , \predict_PC[13][4] ,
         \predict_PC[13][3] , \predict_PC[13][2] , \predict_PC[13][1] ,
         \predict_PC[13][0] , \predict_PC[14][31] , \predict_PC[14][30] ,
         \predict_PC[14][29] , \predict_PC[14][28] , \predict_PC[14][27] ,
         \predict_PC[14][26] , \predict_PC[14][25] , \predict_PC[14][24] ,
         \predict_PC[14][23] , \predict_PC[14][22] , \predict_PC[14][21] ,
         \predict_PC[14][20] , \predict_PC[14][19] , \predict_PC[14][18] ,
         \predict_PC[14][17] , \predict_PC[14][16] , \predict_PC[14][15] ,
         \predict_PC[14][14] , \predict_PC[14][13] , \predict_PC[14][12] ,
         \predict_PC[14][11] , \predict_PC[14][10] , \predict_PC[14][9] ,
         \predict_PC[14][8] , \predict_PC[14][7] , \predict_PC[14][6] ,
         \predict_PC[14][5] , \predict_PC[14][4] , \predict_PC[14][3] ,
         \predict_PC[14][2] , \predict_PC[14][1] , \predict_PC[14][0] ,
         \predict_PC[15][31] , \predict_PC[15][30] , \predict_PC[15][29] ,
         \predict_PC[15][28] , \predict_PC[15][27] , \predict_PC[15][26] ,
         \predict_PC[15][25] , \predict_PC[15][24] , \predict_PC[15][23] ,
         \predict_PC[15][22] , \predict_PC[15][21] , \predict_PC[15][20] ,
         \predict_PC[15][19] , \predict_PC[15][18] , \predict_PC[15][17] ,
         \predict_PC[15][16] , \predict_PC[15][15] , \predict_PC[15][14] ,
         \predict_PC[15][13] , \predict_PC[15][12] , \predict_PC[15][11] ,
         \predict_PC[15][10] , \predict_PC[15][9] , \predict_PC[15][8] ,
         \predict_PC[15][7] , \predict_PC[15][6] , \predict_PC[15][5] ,
         \predict_PC[15][4] , \predict_PC[15][3] , \predict_PC[15][2] ,
         \predict_PC[15][1] , \predict_PC[15][0] , N38, N39, N40, N41, N42,
         N43, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N86, N118,
         N150, N182, N214, N246, N278, N310, N342, N374, N406, N438, N470,
         N502, N534, N566, N567, net338272, net338277, net338282, net338287,
         net338292, net338297, net338302, net338307, net338312, net338317,
         net338322, net338327, net338332, net338337, net338342, net338347,
         net338352, n483, n485, n487, n489, n491, n493, n495, n497, n499, n501,
         n503, n505, n507, n509, n511, n513, n515, n517, n519, n521, n523,
         n525, n527, n529, n531, n533, n535, n537, n539, n541, n543, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n951, n955, n972, n973,
         n974, n975, n976, n977, n978, n979, n1, n2, n3, n4, n5, n6, n7, n8,
         n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45;
  wire   [15:0] taken;
  wire   [15:0] write_enable;

  DFFS_X1 \last_TAG_reg[3]  ( .D(n972), .CK(net338272), .SN(n31), .Q(n977), 
        .QN(n4) );
  DFFS_X1 \last_TAG_reg[2]  ( .D(n973), .CK(net338272), .SN(n22), .Q(n976), 
        .QN(n2) );
  DFFS_X1 \last_TAG_reg[1]  ( .D(n974), .CK(net338272), .SN(n24), .Q(n979), 
        .QN(n3) );
  DFFR_X1 \last_TAG_reg[0]  ( .D(TAG_i[0]), .CK(net338272), .RN(n32), .Q(n1), 
        .QN(n978) );
  DFFR_X1 \write_enable_reg[15]  ( .D(N53), .CK(net338272), .RN(n26), .Q(
        write_enable[15]) );
  DFFR_X1 \write_enable_reg[14]  ( .D(N52), .CK(net338272), .RN(n24), .Q(
        write_enable[14]) );
  DFFR_X1 \write_enable_reg[13]  ( .D(N51), .CK(net338272), .RN(n27), .Q(
        write_enable[13]) );
  DFFR_X1 \write_enable_reg[12]  ( .D(N50), .CK(net338272), .RN(n28), .Q(
        write_enable[12]) );
  DFFR_X1 \write_enable_reg[11]  ( .D(N49), .CK(net338272), .RN(n30), .Q(
        write_enable[11]) );
  DFFR_X1 \write_enable_reg[10]  ( .D(N48), .CK(net338272), .RN(n31), .Q(
        write_enable[10]) );
  DFFR_X1 \write_enable_reg[9]  ( .D(N47), .CK(net338272), .RN(n30), .Q(
        write_enable[9]) );
  DFFR_X1 \write_enable_reg[8]  ( .D(N46), .CK(net338272), .RN(n29), .Q(
        write_enable[8]) );
  DFFR_X1 \write_enable_reg[7]  ( .D(N45), .CK(net338272), .RN(n32), .Q(
        write_enable[7]) );
  DFFR_X1 \write_enable_reg[6]  ( .D(N44), .CK(net338272), .RN(n29), .Q(
        write_enable[6]) );
  DFFR_X1 \write_enable_reg[5]  ( .D(N43), .CK(net338272), .RN(n31), .Q(
        write_enable[5]) );
  DFFR_X1 \write_enable_reg[4]  ( .D(N42), .CK(net338272), .RN(n30), .Q(
        write_enable[4]) );
  DFFR_X1 \write_enable_reg[3]  ( .D(N41), .CK(net338272), .RN(n29), .Q(
        write_enable[3]) );
  DFFR_X1 \write_enable_reg[2]  ( .D(N40), .CK(net338272), .RN(n32), .Q(
        write_enable[2]) );
  DFFR_X1 \write_enable_reg[1]  ( .D(N39), .CK(net338272), .RN(n32), .Q(
        write_enable[1]) );
  DFFR_X1 \write_enable_reg[0]  ( .D(N38), .CK(net338272), .RN(n31), .Q(
        write_enable[0]) );
  DFF_X1 last_taken_reg ( .D(n955), .CK(clock), .Q(n5), .QN(n975) );
  DFFR_X1 \predict_PC_reg[0][31]  ( .D(target_PC_i[31]), .CK(net338277), .RN(
        n32), .Q(\predict_PC[0][31] ) );
  DFFR_X1 \predict_PC_reg[0][30]  ( .D(target_PC_i[30]), .CK(net338277), .RN(
        n29), .Q(\predict_PC[0][30] ) );
  DFFR_X1 \predict_PC_reg[0][29]  ( .D(target_PC_i[29]), .CK(net338277), .RN(
        n30), .Q(\predict_PC[0][29] ) );
  DFFR_X1 \predict_PC_reg[0][28]  ( .D(target_PC_i[28]), .CK(net338277), .RN(
        n31), .Q(\predict_PC[0][28] ) );
  DFFR_X1 \predict_PC_reg[0][27]  ( .D(target_PC_i[27]), .CK(net338277), .RN(
        n32), .Q(\predict_PC[0][27] ) );
  DFFR_X1 \predict_PC_reg[0][26]  ( .D(target_PC_i[26]), .CK(net338277), .RN(
        n29), .Q(\predict_PC[0][26] ) );
  DFFR_X1 \predict_PC_reg[0][25]  ( .D(target_PC_i[25]), .CK(net338277), .RN(
        n30), .Q(\predict_PC[0][25] ) );
  DFFR_X1 \predict_PC_reg[0][24]  ( .D(target_PC_i[24]), .CK(net338277), .RN(
        n31), .Q(\predict_PC[0][24] ) );
  DFFR_X1 \predict_PC_reg[0][23]  ( .D(target_PC_i[23]), .CK(net338277), .RN(
        n32), .Q(\predict_PC[0][23] ) );
  DFFR_X1 \predict_PC_reg[0][22]  ( .D(target_PC_i[22]), .CK(net338277), .RN(
        n29), .Q(\predict_PC[0][22] ) );
  DFFR_X1 \predict_PC_reg[0][21]  ( .D(target_PC_i[21]), .CK(net338277), .RN(
        n30), .Q(\predict_PC[0][21] ) );
  DFFR_X1 \predict_PC_reg[0][20]  ( .D(target_PC_i[20]), .CK(net338277), .RN(
        n31), .Q(\predict_PC[0][20] ) );
  DFFR_X1 \predict_PC_reg[0][19]  ( .D(target_PC_i[19]), .CK(net338277), .RN(
        n29), .Q(\predict_PC[0][19] ) );
  DFFR_X1 \predict_PC_reg[0][18]  ( .D(target_PC_i[18]), .CK(net338277), .RN(
        n29), .Q(\predict_PC[0][18] ) );
  DFFR_X1 \predict_PC_reg[0][17]  ( .D(target_PC_i[17]), .CK(net338277), .RN(
        n29), .Q(\predict_PC[0][17] ) );
  DFFR_X1 \predict_PC_reg[0][16]  ( .D(target_PC_i[16]), .CK(net338277), .RN(
        n29), .Q(\predict_PC[0][16] ) );
  DFFR_X1 \predict_PC_reg[0][15]  ( .D(target_PC_i[15]), .CK(net338277), .RN(
        n29), .Q(\predict_PC[0][15] ) );
  DFFR_X1 \predict_PC_reg[0][14]  ( .D(target_PC_i[14]), .CK(net338277), .RN(
        n29), .Q(\predict_PC[0][14] ) );
  DFFR_X1 \predict_PC_reg[0][13]  ( .D(target_PC_i[13]), .CK(net338277), .RN(
        n29), .Q(\predict_PC[0][13] ) );
  DFFR_X1 \predict_PC_reg[0][12]  ( .D(target_PC_i[12]), .CK(net338277), .RN(
        n29), .Q(\predict_PC[0][12] ) );
  DFFR_X1 \predict_PC_reg[0][11]  ( .D(target_PC_i[11]), .CK(net338277), .RN(
        n29), .Q(\predict_PC[0][11] ) );
  DFFR_X1 \predict_PC_reg[0][10]  ( .D(target_PC_i[10]), .CK(net338277), .RN(
        n29), .Q(\predict_PC[0][10] ) );
  DFFR_X1 \predict_PC_reg[0][9]  ( .D(target_PC_i[9]), .CK(net338277), .RN(n29), .Q(\predict_PC[0][9] ) );
  DFFR_X1 \predict_PC_reg[0][8]  ( .D(target_PC_i[8]), .CK(net338277), .RN(n29), .Q(\predict_PC[0][8] ) );
  DFFR_X1 \predict_PC_reg[0][7]  ( .D(target_PC_i[7]), .CK(net338277), .RN(n30), .Q(\predict_PC[0][7] ) );
  DFFR_X1 \predict_PC_reg[0][6]  ( .D(target_PC_i[6]), .CK(net338277), .RN(n30), .Q(\predict_PC[0][6] ) );
  DFFR_X1 \predict_PC_reg[0][5]  ( .D(target_PC_i[5]), .CK(net338277), .RN(n30), .Q(\predict_PC[0][5] ) );
  DFFR_X1 \predict_PC_reg[0][4]  ( .D(target_PC_i[4]), .CK(net338277), .RN(n30), .Q(\predict_PC[0][4] ) );
  DFFR_X1 \predict_PC_reg[0][3]  ( .D(target_PC_i[3]), .CK(net338277), .RN(n30), .Q(\predict_PC[0][3] ) );
  DFFR_X1 \predict_PC_reg[0][2]  ( .D(target_PC_i[2]), .CK(net338277), .RN(n30), .Q(\predict_PC[0][2] ) );
  DFFR_X1 \predict_PC_reg[0][1]  ( .D(target_PC_i[1]), .CK(net338277), .RN(n30), .Q(\predict_PC[0][1] ) );
  DFFR_X1 \predict_PC_reg[0][0]  ( .D(target_PC_i[0]), .CK(net338277), .RN(n30), .Q(\predict_PC[0][0] ) );
  DFFR_X1 \predict_PC_reg[1][31]  ( .D(target_PC_i[31]), .CK(net338282), .RN(
        n30), .Q(\predict_PC[1][31] ) );
  DFFR_X1 \predict_PC_reg[1][30]  ( .D(target_PC_i[30]), .CK(net338282), .RN(
        n30), .Q(\predict_PC[1][30] ) );
  DFFR_X1 \predict_PC_reg[1][29]  ( .D(target_PC_i[29]), .CK(net338282), .RN(
        n30), .Q(\predict_PC[1][29] ) );
  DFFR_X1 \predict_PC_reg[1][28]  ( .D(target_PC_i[28]), .CK(net338282), .RN(
        n30), .Q(\predict_PC[1][28] ) );
  DFFR_X1 \predict_PC_reg[1][27]  ( .D(target_PC_i[27]), .CK(net338282), .RN(
        n31), .Q(\predict_PC[1][27] ) );
  DFFR_X1 \predict_PC_reg[1][26]  ( .D(target_PC_i[26]), .CK(net338282), .RN(
        n31), .Q(\predict_PC[1][26] ) );
  DFFR_X1 \predict_PC_reg[1][25]  ( .D(target_PC_i[25]), .CK(net338282), .RN(
        n31), .Q(\predict_PC[1][25] ) );
  DFFR_X1 \predict_PC_reg[1][24]  ( .D(target_PC_i[24]), .CK(net338282), .RN(
        n31), .Q(\predict_PC[1][24] ) );
  DFFR_X1 \predict_PC_reg[1][23]  ( .D(target_PC_i[23]), .CK(net338282), .RN(
        n31), .Q(\predict_PC[1][23] ) );
  DFFR_X1 \predict_PC_reg[1][22]  ( .D(target_PC_i[22]), .CK(net338282), .RN(
        n31), .Q(\predict_PC[1][22] ) );
  DFFR_X1 \predict_PC_reg[1][21]  ( .D(target_PC_i[21]), .CK(net338282), .RN(
        n31), .Q(\predict_PC[1][21] ) );
  DFFR_X1 \predict_PC_reg[1][20]  ( .D(target_PC_i[20]), .CK(net338282), .RN(
        n31), .Q(\predict_PC[1][20] ) );
  DFFR_X1 \predict_PC_reg[1][19]  ( .D(target_PC_i[19]), .CK(net338282), .RN(
        n31), .Q(\predict_PC[1][19] ) );
  DFFR_X1 \predict_PC_reg[1][18]  ( .D(target_PC_i[18]), .CK(net338282), .RN(
        n31), .Q(\predict_PC[1][18] ) );
  DFFR_X1 \predict_PC_reg[1][17]  ( .D(target_PC_i[17]), .CK(net338282), .RN(
        n31), .Q(\predict_PC[1][17] ) );
  DFFR_X1 \predict_PC_reg[1][16]  ( .D(target_PC_i[16]), .CK(net338282), .RN(
        n31), .Q(\predict_PC[1][16] ) );
  DFFR_X1 \predict_PC_reg[1][15]  ( .D(target_PC_i[15]), .CK(net338282), .RN(
        n32), .Q(\predict_PC[1][15] ) );
  DFFR_X1 \predict_PC_reg[1][14]  ( .D(target_PC_i[14]), .CK(net338282), .RN(
        n32), .Q(\predict_PC[1][14] ) );
  DFFR_X1 \predict_PC_reg[1][13]  ( .D(target_PC_i[13]), .CK(net338282), .RN(
        n32), .Q(\predict_PC[1][13] ) );
  DFFR_X1 \predict_PC_reg[1][12]  ( .D(target_PC_i[12]), .CK(net338282), .RN(
        n32), .Q(\predict_PC[1][12] ) );
  DFFR_X1 \predict_PC_reg[1][11]  ( .D(target_PC_i[11]), .CK(net338282), .RN(
        n32), .Q(\predict_PC[1][11] ) );
  DFFR_X1 \predict_PC_reg[1][10]  ( .D(target_PC_i[10]), .CK(net338282), .RN(
        n32), .Q(\predict_PC[1][10] ) );
  DFFR_X1 \predict_PC_reg[1][9]  ( .D(target_PC_i[9]), .CK(net338282), .RN(n32), .Q(\predict_PC[1][9] ) );
  DFFR_X1 \predict_PC_reg[1][8]  ( .D(target_PC_i[8]), .CK(net338282), .RN(n32), .Q(\predict_PC[1][8] ) );
  DFFR_X1 \predict_PC_reg[1][7]  ( .D(target_PC_i[7]), .CK(net338282), .RN(n32), .Q(\predict_PC[1][7] ) );
  DFFR_X1 \predict_PC_reg[1][6]  ( .D(target_PC_i[6]), .CK(net338282), .RN(n32), .Q(\predict_PC[1][6] ) );
  DFFR_X1 \predict_PC_reg[1][5]  ( .D(target_PC_i[5]), .CK(net338282), .RN(n32), .Q(\predict_PC[1][5] ) );
  DFFR_X1 \predict_PC_reg[1][4]  ( .D(target_PC_i[4]), .CK(net338282), .RN(n35), .Q(\predict_PC[1][4] ) );
  DFFR_X1 \predict_PC_reg[1][3]  ( .D(target_PC_i[3]), .CK(net338282), .RN(n39), .Q(\predict_PC[1][3] ) );
  DFFR_X1 \predict_PC_reg[1][2]  ( .D(target_PC_i[2]), .CK(net338282), .RN(n34), .Q(\predict_PC[1][2] ) );
  DFFR_X1 \predict_PC_reg[1][1]  ( .D(target_PC_i[1]), .CK(net338282), .RN(n34), .Q(\predict_PC[1][1] ) );
  DFFR_X1 \predict_PC_reg[1][0]  ( .D(target_PC_i[0]), .CK(net338282), .RN(n35), .Q(\predict_PC[1][0] ) );
  DFFR_X1 \predict_PC_reg[2][31]  ( .D(target_PC_i[31]), .CK(net338287), .RN(
        n45), .Q(\predict_PC[2][31] ) );
  DFFR_X1 \predict_PC_reg[2][30]  ( .D(target_PC_i[30]), .CK(net338287), .RN(
        n33), .Q(\predict_PC[2][30] ) );
  DFFR_X1 \predict_PC_reg[2][29]  ( .D(target_PC_i[29]), .CK(net338287), .RN(
        n38), .Q(\predict_PC[2][29] ) );
  DFFR_X1 \predict_PC_reg[2][28]  ( .D(target_PC_i[28]), .CK(net338287), .RN(
        n45), .Q(\predict_PC[2][28] ) );
  DFFR_X1 \predict_PC_reg[2][27]  ( .D(target_PC_i[27]), .CK(net338287), .RN(
        n44), .Q(\predict_PC[2][27] ) );
  DFFR_X1 \predict_PC_reg[2][26]  ( .D(target_PC_i[26]), .CK(net338287), .RN(
        n30), .Q(\predict_PC[2][26] ) );
  DFFR_X1 \predict_PC_reg[2][25]  ( .D(target_PC_i[25]), .CK(net338287), .RN(
        n30), .Q(\predict_PC[2][25] ) );
  DFFR_X1 \predict_PC_reg[2][24]  ( .D(target_PC_i[24]), .CK(net338287), .RN(
        n34), .Q(\predict_PC[2][24] ) );
  DFFR_X1 \predict_PC_reg[2][23]  ( .D(target_PC_i[23]), .CK(net338287), .RN(
        n32), .Q(\predict_PC[2][23] ) );
  DFFR_X1 \predict_PC_reg[2][22]  ( .D(target_PC_i[22]), .CK(net338287), .RN(
        n32), .Q(\predict_PC[2][22] ) );
  DFFR_X1 \predict_PC_reg[2][21]  ( .D(target_PC_i[21]), .CK(net338287), .RN(
        n29), .Q(\predict_PC[2][21] ) );
  DFFR_X1 \predict_PC_reg[2][20]  ( .D(target_PC_i[20]), .CK(net338287), .RN(
        n41), .Q(\predict_PC[2][20] ) );
  DFFR_X1 \predict_PC_reg[2][19]  ( .D(target_PC_i[19]), .CK(net338287), .RN(
        n43), .Q(\predict_PC[2][19] ) );
  DFFR_X1 \predict_PC_reg[2][18]  ( .D(target_PC_i[18]), .CK(net338287), .RN(
        n42), .Q(\predict_PC[2][18] ) );
  DFFR_X1 \predict_PC_reg[2][17]  ( .D(target_PC_i[17]), .CK(net338287), .RN(
        n41), .Q(\predict_PC[2][17] ) );
  DFFR_X1 \predict_PC_reg[2][16]  ( .D(target_PC_i[16]), .CK(net338287), .RN(
        n40), .Q(\predict_PC[2][16] ) );
  DFFR_X1 \predict_PC_reg[2][15]  ( .D(target_PC_i[15]), .CK(net338287), .RN(
        n39), .Q(\predict_PC[2][15] ) );
  DFFR_X1 \predict_PC_reg[2][14]  ( .D(target_PC_i[14]), .CK(net338287), .RN(
        n37), .Q(\predict_PC[2][14] ) );
  DFFR_X1 \predict_PC_reg[2][13]  ( .D(target_PC_i[13]), .CK(net338287), .RN(
        n36), .Q(\predict_PC[2][13] ) );
  DFFR_X1 \predict_PC_reg[2][12]  ( .D(target_PC_i[12]), .CK(net338287), .RN(
        n26), .Q(\predict_PC[2][12] ) );
  DFFR_X1 \predict_PC_reg[2][11]  ( .D(target_PC_i[11]), .CK(net338287), .RN(
        n29), .Q(\predict_PC[2][11] ) );
  DFFR_X1 \predict_PC_reg[2][10]  ( .D(target_PC_i[10]), .CK(net338287), .RN(
        n27), .Q(\predict_PC[2][10] ) );
  DFFR_X1 \predict_PC_reg[2][9]  ( .D(target_PC_i[9]), .CK(net338287), .RN(n43), .Q(\predict_PC[2][9] ) );
  DFFR_X1 \predict_PC_reg[2][8]  ( .D(target_PC_i[8]), .CK(net338287), .RN(n43), .Q(\predict_PC[2][8] ) );
  DFFR_X1 \predict_PC_reg[2][7]  ( .D(target_PC_i[7]), .CK(net338287), .RN(n44), .Q(\predict_PC[2][7] ) );
  DFFR_X1 \predict_PC_reg[2][6]  ( .D(target_PC_i[6]), .CK(net338287), .RN(n33), .Q(\predict_PC[2][6] ) );
  DFFR_X1 \predict_PC_reg[2][5]  ( .D(target_PC_i[5]), .CK(net338287), .RN(n38), .Q(\predict_PC[2][5] ) );
  DFFR_X1 \predict_PC_reg[2][4]  ( .D(target_PC_i[4]), .CK(net338287), .RN(n45), .Q(\predict_PC[2][4] ) );
  DFFR_X1 \predict_PC_reg[2][3]  ( .D(target_PC_i[3]), .CK(net338287), .RN(n44), .Q(\predict_PC[2][3] ) );
  DFFR_X1 \predict_PC_reg[2][2]  ( .D(target_PC_i[2]), .CK(net338287), .RN(n31), .Q(\predict_PC[2][2] ) );
  DFFR_X1 \predict_PC_reg[2][1]  ( .D(target_PC_i[1]), .CK(net338287), .RN(n31), .Q(\predict_PC[2][1] ) );
  DFFR_X1 \predict_PC_reg[2][0]  ( .D(target_PC_i[0]), .CK(net338287), .RN(n27), .Q(\predict_PC[2][0] ) );
  DFFR_X1 \predict_PC_reg[3][31]  ( .D(target_PC_i[31]), .CK(net338292), .RN(
        n29), .Q(\predict_PC[3][31] ) );
  DFFR_X1 \predict_PC_reg[3][30]  ( .D(target_PC_i[30]), .CK(net338292), .RN(
        n33), .Q(\predict_PC[3][30] ) );
  DFFR_X1 \predict_PC_reg[3][29]  ( .D(target_PC_i[29]), .CK(net338292), .RN(
        n40), .Q(\predict_PC[3][29] ) );
  DFFR_X1 \predict_PC_reg[3][28]  ( .D(target_PC_i[28]), .CK(net338292), .RN(
        n43), .Q(\predict_PC[3][28] ) );
  DFFR_X1 \predict_PC_reg[3][27]  ( .D(target_PC_i[27]), .CK(net338292), .RN(
        n42), .Q(\predict_PC[3][27] ) );
  DFFR_X1 \predict_PC_reg[3][26]  ( .D(target_PC_i[26]), .CK(net338292), .RN(
        n41), .Q(\predict_PC[3][26] ) );
  DFFR_X1 \predict_PC_reg[3][25]  ( .D(target_PC_i[25]), .CK(net338292), .RN(
        n40), .Q(\predict_PC[3][25] ) );
  DFFR_X1 \predict_PC_reg[3][24]  ( .D(target_PC_i[24]), .CK(net338292), .RN(
        n39), .Q(\predict_PC[3][24] ) );
  DFFR_X1 \predict_PC_reg[3][23]  ( .D(target_PC_i[23]), .CK(net338292), .RN(
        n37), .Q(\predict_PC[3][23] ) );
  DFFR_X1 \predict_PC_reg[3][22]  ( .D(target_PC_i[22]), .CK(net338292), .RN(
        n36), .Q(\predict_PC[3][22] ) );
  DFFR_X1 \predict_PC_reg[3][21]  ( .D(target_PC_i[21]), .CK(net338292), .RN(
        n35), .Q(\predict_PC[3][21] ) );
  DFFR_X1 \predict_PC_reg[3][20]  ( .D(target_PC_i[20]), .CK(net338292), .RN(
        n42), .Q(\predict_PC[3][20] ) );
  DFFR_X1 \predict_PC_reg[3][19]  ( .D(target_PC_i[19]), .CK(net338292), .RN(
        n26), .Q(\predict_PC[3][19] ) );
  DFFR_X1 \predict_PC_reg[3][18]  ( .D(target_PC_i[18]), .CK(net338292), .RN(
        n33), .Q(\predict_PC[3][18] ) );
  DFFR_X1 \predict_PC_reg[3][17]  ( .D(target_PC_i[17]), .CK(net338292), .RN(
        n38), .Q(\predict_PC[3][17] ) );
  DFFR_X1 \predict_PC_reg[3][16]  ( .D(target_PC_i[16]), .CK(net338292), .RN(
        n45), .Q(\predict_PC[3][16] ) );
  DFFR_X1 \predict_PC_reg[3][15]  ( .D(target_PC_i[15]), .CK(net338292), .RN(
        n44), .Q(\predict_PC[3][15] ) );
  DFFR_X1 \predict_PC_reg[3][14]  ( .D(target_PC_i[14]), .CK(net338292), .RN(
        n32), .Q(\predict_PC[3][14] ) );
  DFFR_X1 \predict_PC_reg[3][13]  ( .D(target_PC_i[13]), .CK(net338292), .RN(
        n32), .Q(\predict_PC[3][13] ) );
  DFFR_X1 \predict_PC_reg[3][12]  ( .D(target_PC_i[12]), .CK(net338292), .RN(
        n41), .Q(\predict_PC[3][12] ) );
  DFFR_X1 \predict_PC_reg[3][11]  ( .D(target_PC_i[11]), .CK(net338292), .RN(
        n25), .Q(\predict_PC[3][11] ) );
  DFFR_X1 \predict_PC_reg[3][10]  ( .D(target_PC_i[10]), .CK(net338292), .RN(
        n33), .Q(\predict_PC[3][10] ) );
  DFFR_X1 \predict_PC_reg[3][9]  ( .D(target_PC_i[9]), .CK(net338292), .RN(n38), .Q(\predict_PC[3][9] ) );
  DFFR_X1 \predict_PC_reg[3][8]  ( .D(target_PC_i[8]), .CK(net338292), .RN(n26), .Q(\predict_PC[3][8] ) );
  DFFR_X1 \predict_PC_reg[3][7]  ( .D(target_PC_i[7]), .CK(net338292), .RN(n41), .Q(\predict_PC[3][7] ) );
  DFFR_X1 \predict_PC_reg[3][6]  ( .D(target_PC_i[6]), .CK(net338292), .RN(n40), .Q(\predict_PC[3][6] ) );
  DFFR_X1 \predict_PC_reg[3][5]  ( .D(target_PC_i[5]), .CK(net338292), .RN(n36), .Q(\predict_PC[3][5] ) );
  DFFR_X1 \predict_PC_reg[3][4]  ( .D(target_PC_i[4]), .CK(net338292), .RN(n39), .Q(\predict_PC[3][4] ) );
  DFFR_X1 \predict_PC_reg[3][3]  ( .D(target_PC_i[3]), .CK(net338292), .RN(n37), .Q(\predict_PC[3][3] ) );
  DFFR_X1 \predict_PC_reg[3][2]  ( .D(target_PC_i[2]), .CK(net338292), .RN(n25), .Q(\predict_PC[3][2] ) );
  DFFR_X1 \predict_PC_reg[3][1]  ( .D(target_PC_i[1]), .CK(net338292), .RN(n22), .Q(\predict_PC[3][1] ) );
  DFFR_X1 \predict_PC_reg[3][0]  ( .D(target_PC_i[0]), .CK(net338292), .RN(n23), .Q(\predict_PC[3][0] ) );
  DFFR_X1 \predict_PC_reg[4][31]  ( .D(target_PC_i[31]), .CK(net338297), .RN(
        n23), .Q(\predict_PC[4][31] ) );
  DFFR_X1 \predict_PC_reg[4][30]  ( .D(target_PC_i[30]), .CK(net338297), .RN(
        n24), .Q(\predict_PC[4][30] ) );
  DFFR_X1 \predict_PC_reg[4][29]  ( .D(target_PC_i[29]), .CK(net338297), .RN(
        n22), .Q(\predict_PC[4][29] ) );
  DFFR_X1 \predict_PC_reg[4][28]  ( .D(target_PC_i[28]), .CK(net338297), .RN(
        n24), .Q(\predict_PC[4][28] ) );
  DFFR_X1 \predict_PC_reg[4][27]  ( .D(target_PC_i[27]), .CK(net338297), .RN(
        n23), .Q(\predict_PC[4][27] ) );
  DFFR_X1 \predict_PC_reg[4][26]  ( .D(target_PC_i[26]), .CK(net338297), .RN(
        n24), .Q(\predict_PC[4][26] ) );
  DFFR_X1 \predict_PC_reg[4][25]  ( .D(target_PC_i[25]), .CK(net338297), .RN(
        n22), .Q(\predict_PC[4][25] ) );
  DFFR_X1 \predict_PC_reg[4][24]  ( .D(target_PC_i[24]), .CK(net338297), .RN(
        n22), .Q(\predict_PC[4][24] ) );
  DFFR_X1 \predict_PC_reg[4][23]  ( .D(target_PC_i[23]), .CK(net338297), .RN(
        n23), .Q(\predict_PC[4][23] ) );
  DFFR_X1 \predict_PC_reg[4][22]  ( .D(target_PC_i[22]), .CK(net338297), .RN(
        n23), .Q(\predict_PC[4][22] ) );
  DFFR_X1 \predict_PC_reg[4][21]  ( .D(target_PC_i[21]), .CK(net338297), .RN(
        n22), .Q(\predict_PC[4][21] ) );
  DFFR_X1 \predict_PC_reg[4][20]  ( .D(target_PC_i[20]), .CK(net338297), .RN(
        n23), .Q(\predict_PC[4][20] ) );
  DFFR_X1 \predict_PC_reg[4][19]  ( .D(target_PC_i[19]), .CK(net338297), .RN(
        n24), .Q(\predict_PC[4][19] ) );
  DFFR_X1 \predict_PC_reg[4][18]  ( .D(target_PC_i[18]), .CK(net338297), .RN(
        n22), .Q(\predict_PC[4][18] ) );
  DFFR_X1 \predict_PC_reg[4][17]  ( .D(target_PC_i[17]), .CK(net338297), .RN(
        n23), .Q(\predict_PC[4][17] ) );
  DFFR_X1 \predict_PC_reg[4][16]  ( .D(target_PC_i[16]), .CK(net338297), .RN(
        n24), .Q(\predict_PC[4][16] ) );
  DFFR_X1 \predict_PC_reg[4][15]  ( .D(target_PC_i[15]), .CK(net338297), .RN(
        n22), .Q(\predict_PC[4][15] ) );
  DFFR_X1 \predict_PC_reg[4][14]  ( .D(target_PC_i[14]), .CK(net338297), .RN(
        n23), .Q(\predict_PC[4][14] ) );
  DFFR_X1 \predict_PC_reg[4][13]  ( .D(target_PC_i[13]), .CK(net338297), .RN(
        n24), .Q(\predict_PC[4][13] ) );
  DFFR_X1 \predict_PC_reg[4][12]  ( .D(target_PC_i[12]), .CK(net338297), .RN(
        n22), .Q(\predict_PC[4][12] ) );
  DFFR_X1 \predict_PC_reg[4][11]  ( .D(target_PC_i[11]), .CK(net338297), .RN(
        n23), .Q(\predict_PC[4][11] ) );
  DFFR_X1 \predict_PC_reg[4][10]  ( .D(target_PC_i[10]), .CK(net338297), .RN(
        n22), .Q(\predict_PC[4][10] ) );
  DFFR_X1 \predict_PC_reg[4][9]  ( .D(target_PC_i[9]), .CK(net338297), .RN(n22), .Q(\predict_PC[4][9] ) );
  DFFR_X1 \predict_PC_reg[4][8]  ( .D(target_PC_i[8]), .CK(net338297), .RN(n22), .Q(\predict_PC[4][8] ) );
  DFFR_X1 \predict_PC_reg[4][7]  ( .D(target_PC_i[7]), .CK(net338297), .RN(n22), .Q(\predict_PC[4][7] ) );
  DFFR_X1 \predict_PC_reg[4][6]  ( .D(target_PC_i[6]), .CK(net338297), .RN(n22), .Q(\predict_PC[4][6] ) );
  DFFR_X1 \predict_PC_reg[4][5]  ( .D(target_PC_i[5]), .CK(net338297), .RN(n22), .Q(\predict_PC[4][5] ) );
  DFFR_X1 \predict_PC_reg[4][4]  ( .D(target_PC_i[4]), .CK(net338297), .RN(n22), .Q(\predict_PC[4][4] ) );
  DFFR_X1 \predict_PC_reg[4][3]  ( .D(target_PC_i[3]), .CK(net338297), .RN(n22), .Q(\predict_PC[4][3] ) );
  DFFR_X1 \predict_PC_reg[4][2]  ( .D(target_PC_i[2]), .CK(net338297), .RN(n22), .Q(\predict_PC[4][2] ) );
  DFFR_X1 \predict_PC_reg[4][1]  ( .D(target_PC_i[1]), .CK(net338297), .RN(n22), .Q(\predict_PC[4][1] ) );
  DFFR_X1 \predict_PC_reg[4][0]  ( .D(target_PC_i[0]), .CK(net338297), .RN(n22), .Q(\predict_PC[4][0] ) );
  DFFR_X1 \predict_PC_reg[5][31]  ( .D(target_PC_i[31]), .CK(net338302), .RN(
        n22), .Q(\predict_PC[5][31] ) );
  DFFR_X1 \predict_PC_reg[5][30]  ( .D(target_PC_i[30]), .CK(net338302), .RN(
        n23), .Q(\predict_PC[5][30] ) );
  DFFR_X1 \predict_PC_reg[5][29]  ( .D(target_PC_i[29]), .CK(net338302), .RN(
        n23), .Q(\predict_PC[5][29] ) );
  DFFR_X1 \predict_PC_reg[5][28]  ( .D(target_PC_i[28]), .CK(net338302), .RN(
        n23), .Q(\predict_PC[5][28] ) );
  DFFR_X1 \predict_PC_reg[5][27]  ( .D(target_PC_i[27]), .CK(net338302), .RN(
        n23), .Q(\predict_PC[5][27] ) );
  DFFR_X1 \predict_PC_reg[5][26]  ( .D(target_PC_i[26]), .CK(net338302), .RN(
        n23), .Q(\predict_PC[5][26] ) );
  DFFR_X1 \predict_PC_reg[5][25]  ( .D(target_PC_i[25]), .CK(net338302), .RN(
        n23), .Q(\predict_PC[5][25] ) );
  DFFR_X1 \predict_PC_reg[5][24]  ( .D(target_PC_i[24]), .CK(net338302), .RN(
        n23), .Q(\predict_PC[5][24] ) );
  DFFR_X1 \predict_PC_reg[5][23]  ( .D(target_PC_i[23]), .CK(net338302), .RN(
        n23), .Q(\predict_PC[5][23] ) );
  DFFR_X1 \predict_PC_reg[5][22]  ( .D(target_PC_i[22]), .CK(net338302), .RN(
        n23), .Q(\predict_PC[5][22] ) );
  DFFR_X1 \predict_PC_reg[5][21]  ( .D(target_PC_i[21]), .CK(net338302), .RN(
        n23), .Q(\predict_PC[5][21] ) );
  DFFR_X1 \predict_PC_reg[5][20]  ( .D(target_PC_i[20]), .CK(net338302), .RN(
        n23), .Q(\predict_PC[5][20] ) );
  DFFR_X1 \predict_PC_reg[5][19]  ( .D(target_PC_i[19]), .CK(net338302), .RN(
        n23), .Q(\predict_PC[5][19] ) );
  DFFR_X1 \predict_PC_reg[5][18]  ( .D(target_PC_i[18]), .CK(net338302), .RN(
        n24), .Q(\predict_PC[5][18] ) );
  DFFR_X1 \predict_PC_reg[5][17]  ( .D(target_PC_i[17]), .CK(net338302), .RN(
        n24), .Q(\predict_PC[5][17] ) );
  DFFR_X1 \predict_PC_reg[5][16]  ( .D(target_PC_i[16]), .CK(net338302), .RN(
        n24), .Q(\predict_PC[5][16] ) );
  DFFR_X1 \predict_PC_reg[5][15]  ( .D(target_PC_i[15]), .CK(net338302), .RN(
        n24), .Q(\predict_PC[5][15] ) );
  DFFR_X1 \predict_PC_reg[5][14]  ( .D(target_PC_i[14]), .CK(net338302), .RN(
        n24), .Q(\predict_PC[5][14] ) );
  DFFR_X1 \predict_PC_reg[5][13]  ( .D(target_PC_i[13]), .CK(net338302), .RN(
        n24), .Q(\predict_PC[5][13] ) );
  DFFR_X1 \predict_PC_reg[5][12]  ( .D(target_PC_i[12]), .CK(net338302), .RN(
        n24), .Q(\predict_PC[5][12] ) );
  DFFR_X1 \predict_PC_reg[5][11]  ( .D(target_PC_i[11]), .CK(net338302), .RN(
        n24), .Q(\predict_PC[5][11] ) );
  DFFR_X1 \predict_PC_reg[5][10]  ( .D(target_PC_i[10]), .CK(net338302), .RN(
        n24), .Q(\predict_PC[5][10] ) );
  DFFR_X1 \predict_PC_reg[5][9]  ( .D(target_PC_i[9]), .CK(net338302), .RN(n24), .Q(\predict_PC[5][9] ) );
  DFFR_X1 \predict_PC_reg[5][8]  ( .D(target_PC_i[8]), .CK(net338302), .RN(n24), .Q(\predict_PC[5][8] ) );
  DFFR_X1 \predict_PC_reg[5][7]  ( .D(target_PC_i[7]), .CK(net338302), .RN(n24), .Q(\predict_PC[5][7] ) );
  DFFR_X1 \predict_PC_reg[5][6]  ( .D(target_PC_i[6]), .CK(net338302), .RN(n25), .Q(\predict_PC[5][6] ) );
  DFFR_X1 \predict_PC_reg[5][5]  ( .D(target_PC_i[5]), .CK(net338302), .RN(n26), .Q(\predict_PC[5][5] ) );
  DFFR_X1 \predict_PC_reg[5][4]  ( .D(target_PC_i[4]), .CK(net338302), .RN(n27), .Q(\predict_PC[5][4] ) );
  DFFR_X1 \predict_PC_reg[5][3]  ( .D(target_PC_i[3]), .CK(net338302), .RN(n28), .Q(\predict_PC[5][3] ) );
  DFFR_X1 \predict_PC_reg[5][2]  ( .D(target_PC_i[2]), .CK(net338302), .RN(n28), .Q(\predict_PC[5][2] ) );
  DFFR_X1 \predict_PC_reg[5][1]  ( .D(target_PC_i[1]), .CK(net338302), .RN(n25), .Q(\predict_PC[5][1] ) );
  DFFR_X1 \predict_PC_reg[5][0]  ( .D(target_PC_i[0]), .CK(net338302), .RN(n26), .Q(\predict_PC[5][0] ) );
  DFFR_X1 \predict_PC_reg[6][31]  ( .D(target_PC_i[31]), .CK(net338307), .RN(
        n27), .Q(\predict_PC[6][31] ) );
  DFFR_X1 \predict_PC_reg[6][30]  ( .D(target_PC_i[30]), .CK(net338307), .RN(
        n28), .Q(\predict_PC[6][30] ) );
  DFFR_X1 \predict_PC_reg[6][29]  ( .D(target_PC_i[29]), .CK(net338307), .RN(
        n28), .Q(\predict_PC[6][29] ) );
  DFFR_X1 \predict_PC_reg[6][28]  ( .D(target_PC_i[28]), .CK(net338307), .RN(
        n26), .Q(\predict_PC[6][28] ) );
  DFFR_X1 \predict_PC_reg[6][27]  ( .D(target_PC_i[27]), .CK(net338307), .RN(
        n26), .Q(\predict_PC[6][27] ) );
  DFFR_X1 \predict_PC_reg[6][26]  ( .D(target_PC_i[26]), .CK(net338307), .RN(
        n27), .Q(\predict_PC[6][26] ) );
  DFFR_X1 \predict_PC_reg[6][25]  ( .D(target_PC_i[25]), .CK(net338307), .RN(
        n28), .Q(\predict_PC[6][25] ) );
  DFFR_X1 \predict_PC_reg[6][24]  ( .D(target_PC_i[24]), .CK(net338307), .RN(
        n25), .Q(\predict_PC[6][24] ) );
  DFFR_X1 \predict_PC_reg[6][23]  ( .D(target_PC_i[23]), .CK(net338307), .RN(
        n26), .Q(\predict_PC[6][23] ) );
  DFFR_X1 \predict_PC_reg[6][22]  ( .D(target_PC_i[22]), .CK(net338307), .RN(
        n27), .Q(\predict_PC[6][22] ) );
  DFFR_X1 \predict_PC_reg[6][21]  ( .D(target_PC_i[21]), .CK(net338307), .RN(
        n28), .Q(\predict_PC[6][21] ) );
  DFFR_X1 \predict_PC_reg[6][20]  ( .D(target_PC_i[20]), .CK(net338307), .RN(
        n25), .Q(\predict_PC[6][20] ) );
  DFFR_X1 \predict_PC_reg[6][19]  ( .D(target_PC_i[19]), .CK(net338307), .RN(
        n26), .Q(\predict_PC[6][19] ) );
  DFFR_X1 \predict_PC_reg[6][18]  ( .D(target_PC_i[18]), .CK(net338307), .RN(
        n27), .Q(\predict_PC[6][18] ) );
  DFFR_X1 \predict_PC_reg[6][17]  ( .D(target_PC_i[17]), .CK(net338307), .RN(
        n28), .Q(\predict_PC[6][17] ) );
  DFFR_X1 \predict_PC_reg[6][16]  ( .D(target_PC_i[16]), .CK(net338307), .RN(
        n25), .Q(\predict_PC[6][16] ) );
  DFFR_X1 \predict_PC_reg[6][15]  ( .D(target_PC_i[15]), .CK(net338307), .RN(
        n25), .Q(\predict_PC[6][15] ) );
  DFFR_X1 \predict_PC_reg[6][14]  ( .D(target_PC_i[14]), .CK(net338307), .RN(
        n25), .Q(\predict_PC[6][14] ) );
  DFFR_X1 \predict_PC_reg[6][13]  ( .D(target_PC_i[13]), .CK(net338307), .RN(
        n25), .Q(\predict_PC[6][13] ) );
  DFFR_X1 \predict_PC_reg[6][12]  ( .D(target_PC_i[12]), .CK(net338307), .RN(
        n25), .Q(\predict_PC[6][12] ) );
  DFFR_X1 \predict_PC_reg[6][11]  ( .D(target_PC_i[11]), .CK(net338307), .RN(
        n25), .Q(\predict_PC[6][11] ) );
  DFFR_X1 \predict_PC_reg[6][10]  ( .D(target_PC_i[10]), .CK(net338307), .RN(
        n25), .Q(\predict_PC[6][10] ) );
  DFFR_X1 \predict_PC_reg[6][9]  ( .D(target_PC_i[9]), .CK(net338307), .RN(n25), .Q(\predict_PC[6][9] ) );
  DFFR_X1 \predict_PC_reg[6][8]  ( .D(target_PC_i[8]), .CK(net338307), .RN(n25), .Q(\predict_PC[6][8] ) );
  DFFR_X1 \predict_PC_reg[6][7]  ( .D(target_PC_i[7]), .CK(net338307), .RN(n25), .Q(\predict_PC[6][7] ) );
  DFFR_X1 \predict_PC_reg[6][6]  ( .D(target_PC_i[6]), .CK(net338307), .RN(n25), .Q(\predict_PC[6][6] ) );
  DFFR_X1 \predict_PC_reg[6][5]  ( .D(target_PC_i[5]), .CK(net338307), .RN(n25), .Q(\predict_PC[6][5] ) );
  DFFR_X1 \predict_PC_reg[6][4]  ( .D(target_PC_i[4]), .CK(net338307), .RN(n25), .Q(\predict_PC[6][4] ) );
  DFFR_X1 \predict_PC_reg[6][3]  ( .D(target_PC_i[3]), .CK(net338307), .RN(n26), .Q(\predict_PC[6][3] ) );
  DFFR_X1 \predict_PC_reg[6][2]  ( .D(target_PC_i[2]), .CK(net338307), .RN(n26), .Q(\predict_PC[6][2] ) );
  DFFR_X1 \predict_PC_reg[6][1]  ( .D(target_PC_i[1]), .CK(net338307), .RN(n26), .Q(\predict_PC[6][1] ) );
  DFFR_X1 \predict_PC_reg[6][0]  ( .D(target_PC_i[0]), .CK(net338307), .RN(n26), .Q(\predict_PC[6][0] ) );
  DFFR_X1 \predict_PC_reg[7][31]  ( .D(target_PC_i[31]), .CK(net338312), .RN(
        n26), .Q(\predict_PC[7][31] ) );
  DFFR_X1 \predict_PC_reg[7][30]  ( .D(target_PC_i[30]), .CK(net338312), .RN(
        n26), .Q(\predict_PC[7][30] ) );
  DFFR_X1 \predict_PC_reg[7][29]  ( .D(target_PC_i[29]), .CK(net338312), .RN(
        n26), .Q(\predict_PC[7][29] ) );
  DFFR_X1 \predict_PC_reg[7][28]  ( .D(target_PC_i[28]), .CK(net338312), .RN(
        n26), .Q(\predict_PC[7][28] ) );
  DFFR_X1 \predict_PC_reg[7][27]  ( .D(target_PC_i[27]), .CK(net338312), .RN(
        n26), .Q(\predict_PC[7][27] ) );
  DFFR_X1 \predict_PC_reg[7][26]  ( .D(target_PC_i[26]), .CK(net338312), .RN(
        n26), .Q(\predict_PC[7][26] ) );
  DFFR_X1 \predict_PC_reg[7][25]  ( .D(target_PC_i[25]), .CK(net338312), .RN(
        n26), .Q(\predict_PC[7][25] ) );
  DFFR_X1 \predict_PC_reg[7][24]  ( .D(target_PC_i[24]), .CK(net338312), .RN(
        n26), .Q(\predict_PC[7][24] ) );
  DFFR_X1 \predict_PC_reg[7][23]  ( .D(target_PC_i[23]), .CK(net338312), .RN(
        n27), .Q(\predict_PC[7][23] ) );
  DFFR_X1 \predict_PC_reg[7][22]  ( .D(target_PC_i[22]), .CK(net338312), .RN(
        n27), .Q(\predict_PC[7][22] ) );
  DFFR_X1 \predict_PC_reg[7][21]  ( .D(target_PC_i[21]), .CK(net338312), .RN(
        n27), .Q(\predict_PC[7][21] ) );
  DFFR_X1 \predict_PC_reg[7][20]  ( .D(target_PC_i[20]), .CK(net338312), .RN(
        n27), .Q(\predict_PC[7][20] ) );
  DFFR_X1 \predict_PC_reg[7][19]  ( .D(target_PC_i[19]), .CK(net338312), .RN(
        n27), .Q(\predict_PC[7][19] ) );
  DFFR_X1 \predict_PC_reg[7][18]  ( .D(target_PC_i[18]), .CK(net338312), .RN(
        n27), .Q(\predict_PC[7][18] ) );
  DFFR_X1 \predict_PC_reg[7][17]  ( .D(target_PC_i[17]), .CK(net338312), .RN(
        n27), .Q(\predict_PC[7][17] ) );
  DFFR_X1 \predict_PC_reg[7][16]  ( .D(target_PC_i[16]), .CK(net338312), .RN(
        n27), .Q(\predict_PC[7][16] ) );
  DFFR_X1 \predict_PC_reg[7][15]  ( .D(target_PC_i[15]), .CK(net338312), .RN(
        n27), .Q(\predict_PC[7][15] ) );
  DFFR_X1 \predict_PC_reg[7][14]  ( .D(target_PC_i[14]), .CK(net338312), .RN(
        n27), .Q(\predict_PC[7][14] ) );
  DFFR_X1 \predict_PC_reg[7][13]  ( .D(target_PC_i[13]), .CK(net338312), .RN(
        n27), .Q(\predict_PC[7][13] ) );
  DFFR_X1 \predict_PC_reg[7][12]  ( .D(target_PC_i[12]), .CK(net338312), .RN(
        n27), .Q(\predict_PC[7][12] ) );
  DFFR_X1 \predict_PC_reg[7][11]  ( .D(target_PC_i[11]), .CK(net338312), .RN(
        n28), .Q(\predict_PC[7][11] ) );
  DFFR_X1 \predict_PC_reg[7][10]  ( .D(target_PC_i[10]), .CK(net338312), .RN(
        n28), .Q(\predict_PC[7][10] ) );
  DFFR_X1 \predict_PC_reg[7][9]  ( .D(target_PC_i[9]), .CK(net338312), .RN(n28), .Q(\predict_PC[7][9] ) );
  DFFR_X1 \predict_PC_reg[7][8]  ( .D(target_PC_i[8]), .CK(net338312), .RN(n28), .Q(\predict_PC[7][8] ) );
  DFFR_X1 \predict_PC_reg[7][7]  ( .D(target_PC_i[7]), .CK(net338312), .RN(n28), .Q(\predict_PC[7][7] ) );
  DFFR_X1 \predict_PC_reg[7][6]  ( .D(target_PC_i[6]), .CK(net338312), .RN(n28), .Q(\predict_PC[7][6] ) );
  DFFR_X1 \predict_PC_reg[7][5]  ( .D(target_PC_i[5]), .CK(net338312), .RN(n28), .Q(\predict_PC[7][5] ) );
  DFFR_X1 \predict_PC_reg[7][4]  ( .D(target_PC_i[4]), .CK(net338312), .RN(n28), .Q(\predict_PC[7][4] ) );
  DFFR_X1 \predict_PC_reg[7][3]  ( .D(target_PC_i[3]), .CK(net338312), .RN(n28), .Q(\predict_PC[7][3] ) );
  DFFR_X1 \predict_PC_reg[7][2]  ( .D(target_PC_i[2]), .CK(net338312), .RN(n28), .Q(\predict_PC[7][2] ) );
  DFFR_X1 \predict_PC_reg[7][1]  ( .D(target_PC_i[1]), .CK(net338312), .RN(n28), .Q(\predict_PC[7][1] ) );
  DFFR_X1 \predict_PC_reg[7][0]  ( .D(target_PC_i[0]), .CK(net338312), .RN(n28), .Q(\predict_PC[7][0] ) );
  DFFR_X1 \predict_PC_reg[8][31]  ( .D(target_PC_i[31]), .CK(net338317), .RN(
        n27), .Q(\predict_PC[8][31] ) );
  DFFR_X1 \predict_PC_reg[8][30]  ( .D(target_PC_i[30]), .CK(net338317), .RN(
        n26), .Q(\predict_PC[8][30] ) );
  DFFR_X1 \predict_PC_reg[8][29]  ( .D(target_PC_i[29]), .CK(net338317), .RN(
        n25), .Q(\predict_PC[8][29] ) );
  DFFR_X1 \predict_PC_reg[8][28]  ( .D(target_PC_i[28]), .CK(net338317), .RN(
        n26), .Q(\predict_PC[8][28] ) );
  DFFR_X1 \predict_PC_reg[8][27]  ( .D(target_PC_i[27]), .CK(net338317), .RN(
        n27), .Q(\predict_PC[8][27] ) );
  DFFR_X1 \predict_PC_reg[8][26]  ( .D(target_PC_i[26]), .CK(net338317), .RN(
        n28), .Q(\predict_PC[8][26] ) );
  DFFR_X1 \predict_PC_reg[8][25]  ( .D(target_PC_i[25]), .CK(net338317), .RN(
        n25), .Q(\predict_PC[8][25] ) );
  DFFR_X1 \predict_PC_reg[8][24]  ( .D(target_PC_i[24]), .CK(net338317), .RN(
        n27), .Q(\predict_PC[8][24] ) );
  DFFR_X1 \predict_PC_reg[8][23]  ( .D(target_PC_i[23]), .CK(net338317), .RN(
        n25), .Q(\predict_PC[8][23] ) );
  DFFR_X1 \predict_PC_reg[8][22]  ( .D(target_PC_i[22]), .CK(net338317), .RN(
        n33), .Q(\predict_PC[8][22] ) );
  DFFR_X1 \predict_PC_reg[8][21]  ( .D(target_PC_i[21]), .CK(net338317), .RN(
        n38), .Q(\predict_PC[8][21] ) );
  DFFR_X1 \predict_PC_reg[8][20]  ( .D(target_PC_i[20]), .CK(net338317), .RN(
        n45), .Q(\predict_PC[8][20] ) );
  DFFR_X1 \predict_PC_reg[8][19]  ( .D(target_PC_i[19]), .CK(net338317), .RN(
        n44), .Q(\predict_PC[8][19] ) );
  DFFR_X1 \predict_PC_reg[8][18]  ( .D(target_PC_i[18]), .CK(net338317), .RN(
        n25), .Q(\predict_PC[8][18] ) );
  DFFR_X1 \predict_PC_reg[8][17]  ( .D(target_PC_i[17]), .CK(net338317), .RN(
        n25), .Q(\predict_PC[8][17] ) );
  DFFR_X1 \predict_PC_reg[8][16]  ( .D(target_PC_i[16]), .CK(net338317), .RN(
        n27), .Q(\predict_PC[8][16] ) );
  DFFR_X1 \predict_PC_reg[8][15]  ( .D(target_PC_i[15]), .CK(net338317), .RN(
        n45), .Q(\predict_PC[8][15] ) );
  DFFR_X1 \predict_PC_reg[8][14]  ( .D(target_PC_i[14]), .CK(net338317), .RN(
        n44), .Q(\predict_PC[8][14] ) );
  DFFR_X1 \predict_PC_reg[8][13]  ( .D(target_PC_i[13]), .CK(net338317), .RN(
        n43), .Q(\predict_PC[8][13] ) );
  DFFR_X1 \predict_PC_reg[8][12]  ( .D(target_PC_i[12]), .CK(net338317), .RN(
        n42), .Q(\predict_PC[8][12] ) );
  DFFR_X1 \predict_PC_reg[8][11]  ( .D(target_PC_i[11]), .CK(net338317), .RN(
        n40), .Q(\predict_PC[8][11] ) );
  DFFR_X1 \predict_PC_reg[8][10]  ( .D(target_PC_i[10]), .CK(net338317), .RN(
        n35), .Q(\predict_PC[8][10] ) );
  DFFR_X1 \predict_PC_reg[8][9]  ( .D(target_PC_i[9]), .CK(net338317), .RN(n34), .Q(\predict_PC[8][9] ) );
  DFFR_X1 \predict_PC_reg[8][8]  ( .D(target_PC_i[8]), .CK(net338317), .RN(n29), .Q(\predict_PC[8][8] ) );
  DFFR_X1 \predict_PC_reg[8][7]  ( .D(target_PC_i[7]), .CK(net338317), .RN(n33), .Q(\predict_PC[8][7] ) );
  DFFR_X1 \predict_PC_reg[8][6]  ( .D(target_PC_i[6]), .CK(net338317), .RN(n38), .Q(\predict_PC[8][6] ) );
  DFFR_X1 \predict_PC_reg[8][5]  ( .D(target_PC_i[5]), .CK(net338317), .RN(n45), .Q(\predict_PC[8][5] ) );
  DFFR_X1 \predict_PC_reg[8][4]  ( .D(target_PC_i[4]), .CK(net338317), .RN(n44), .Q(\predict_PC[8][4] ) );
  DFFR_X1 \predict_PC_reg[8][3]  ( .D(target_PC_i[3]), .CK(net338317), .RN(n28), .Q(\predict_PC[8][3] ) );
  DFFR_X1 \predict_PC_reg[8][2]  ( .D(target_PC_i[2]), .CK(net338317), .RN(n28), .Q(\predict_PC[8][2] ) );
  DFFR_X1 \predict_PC_reg[8][1]  ( .D(target_PC_i[1]), .CK(net338317), .RN(n29), .Q(\predict_PC[8][1] ) );
  DFFR_X1 \predict_PC_reg[8][0]  ( .D(target_PC_i[0]), .CK(net338317), .RN(n44), .Q(\predict_PC[8][0] ) );
  DFFR_X1 \predict_PC_reg[9][31]  ( .D(target_PC_i[31]), .CK(net338322), .RN(
        n43), .Q(\predict_PC[9][31] ) );
  DFFR_X1 \predict_PC_reg[9][30]  ( .D(target_PC_i[30]), .CK(net338322), .RN(
        n39), .Q(\predict_PC[9][30] ) );
  DFFR_X1 \predict_PC_reg[9][29]  ( .D(target_PC_i[29]), .CK(net338322), .RN(
        n37), .Q(\predict_PC[9][29] ) );
  DFFR_X1 \predict_PC_reg[9][28]  ( .D(target_PC_i[28]), .CK(net338322), .RN(
        n36), .Q(\predict_PC[9][28] ) );
  DFFR_X1 \predict_PC_reg[9][27]  ( .D(target_PC_i[27]), .CK(net338322), .RN(
        n35), .Q(\predict_PC[9][27] ) );
  DFFR_X1 \predict_PC_reg[9][26]  ( .D(target_PC_i[26]), .CK(net338322), .RN(
        n34), .Q(\predict_PC[9][26] ) );
  DFFR_X1 \predict_PC_reg[9][25]  ( .D(target_PC_i[25]), .CK(net338322), .RN(
        n32), .Q(\predict_PC[9][25] ) );
  DFFR_X1 \predict_PC_reg[9][24]  ( .D(target_PC_i[24]), .CK(net338322), .RN(
        n29), .Q(\predict_PC[9][24] ) );
  DFFR_X1 \predict_PC_reg[9][23]  ( .D(target_PC_i[23]), .CK(net338322), .RN(
        n33), .Q(\predict_PC[9][23] ) );
  DFFR_X1 \predict_PC_reg[9][22]  ( .D(target_PC_i[22]), .CK(net338322), .RN(
        n38), .Q(\predict_PC[9][22] ) );
  DFFR_X1 \predict_PC_reg[9][21]  ( .D(target_PC_i[21]), .CK(net338322), .RN(
        n45), .Q(\predict_PC[9][21] ) );
  DFFR_X1 \predict_PC_reg[9][20]  ( .D(target_PC_i[20]), .CK(net338322), .RN(
        n44), .Q(\predict_PC[9][20] ) );
  DFFR_X1 \predict_PC_reg[9][19]  ( .D(target_PC_i[19]), .CK(net338322), .RN(
        n38), .Q(\predict_PC[9][19] ) );
  DFFR_X1 \predict_PC_reg[9][18]  ( .D(target_PC_i[18]), .CK(net338322), .RN(
        n42), .Q(\predict_PC[9][18] ) );
  DFFR_X1 \predict_PC_reg[9][17]  ( .D(target_PC_i[17]), .CK(net338322), .RN(
        n41), .Q(\predict_PC[9][17] ) );
  DFFR_X1 \predict_PC_reg[9][16]  ( .D(target_PC_i[16]), .CK(net338322), .RN(
        n40), .Q(\predict_PC[9][16] ) );
  DFFR_X1 \predict_PC_reg[9][15]  ( .D(target_PC_i[15]), .CK(net338322), .RN(
        n39), .Q(\predict_PC[9][15] ) );
  DFFR_X1 \predict_PC_reg[9][14]  ( .D(target_PC_i[14]), .CK(net338322), .RN(
        n37), .Q(\predict_PC[9][14] ) );
  DFFR_X1 \predict_PC_reg[9][13]  ( .D(target_PC_i[13]), .CK(net338322), .RN(
        n36), .Q(\predict_PC[9][13] ) );
  DFFR_X1 \predict_PC_reg[9][12]  ( .D(target_PC_i[12]), .CK(net338322), .RN(
        n35), .Q(\predict_PC[9][12] ) );
  DFFR_X1 \predict_PC_reg[9][11]  ( .D(target_PC_i[11]), .CK(net338322), .RN(
        n34), .Q(\predict_PC[9][11] ) );
  DFFR_X1 \predict_PC_reg[9][10]  ( .D(target_PC_i[10]), .CK(net338322), .RN(
        n30), .Q(\predict_PC[9][10] ) );
  DFFR_X1 \predict_PC_reg[9][9]  ( .D(target_PC_i[9]), .CK(net338322), .RN(n31), .Q(\predict_PC[9][9] ) );
  DFFR_X1 \predict_PC_reg[9][8]  ( .D(target_PC_i[8]), .CK(net338322), .RN(n32), .Q(\predict_PC[9][8] ) );
  DFFR_X1 \predict_PC_reg[9][7]  ( .D(target_PC_i[7]), .CK(net338322), .RN(n33), .Q(\predict_PC[9][7] ) );
  DFFR_X1 \predict_PC_reg[9][6]  ( .D(target_PC_i[6]), .CK(net338322), .RN(n43), .Q(\predict_PC[9][6] ) );
  DFFR_X1 \predict_PC_reg[9][5]  ( .D(target_PC_i[5]), .CK(net338322), .RN(n42), .Q(\predict_PC[9][5] ) );
  DFFR_X1 \predict_PC_reg[9][4]  ( .D(target_PC_i[4]), .CK(net338322), .RN(n41), .Q(\predict_PC[9][4] ) );
  DFFR_X1 \predict_PC_reg[9][3]  ( .D(target_PC_i[3]), .CK(net338322), .RN(n40), .Q(\predict_PC[9][3] ) );
  DFFR_X1 \predict_PC_reg[9][2]  ( .D(target_PC_i[2]), .CK(net338322), .RN(n39), .Q(\predict_PC[9][2] ) );
  DFFR_X1 \predict_PC_reg[9][1]  ( .D(target_PC_i[1]), .CK(net338322), .RN(n37), .Q(\predict_PC[9][1] ) );
  DFFR_X1 \predict_PC_reg[9][0]  ( .D(target_PC_i[0]), .CK(net338322), .RN(n36), .Q(\predict_PC[9][0] ) );
  DFFR_X1 \predict_PC_reg[10][31]  ( .D(target_PC_i[31]), .CK(net338327), .RN(
        n35), .Q(\predict_PC[10][31] ) );
  DFFR_X1 \predict_PC_reg[10][30]  ( .D(target_PC_i[30]), .CK(net338327), .RN(
        n34), .Q(\predict_PC[10][30] ) );
  DFFR_X1 \predict_PC_reg[10][29]  ( .D(target_PC_i[29]), .CK(net338327), .RN(
        n30), .Q(\predict_PC[10][29] ) );
  DFFR_X1 \predict_PC_reg[10][28]  ( .D(target_PC_i[28]), .CK(net338327), .RN(
        n31), .Q(\predict_PC[10][28] ) );
  DFFR_X1 \predict_PC_reg[10][27]  ( .D(target_PC_i[27]), .CK(net338327), .RN(
        n45), .Q(\predict_PC[10][27] ) );
  DFFR_X1 \predict_PC_reg[10][26]  ( .D(target_PC_i[26]), .CK(net338327), .RN(
        n43), .Q(\predict_PC[10][26] ) );
  DFFR_X1 \predict_PC_reg[10][25]  ( .D(target_PC_i[25]), .CK(net338327), .RN(
        n42), .Q(\predict_PC[10][25] ) );
  DFFR_X1 \predict_PC_reg[10][24]  ( .D(target_PC_i[24]), .CK(net338327), .RN(
        n41), .Q(\predict_PC[10][24] ) );
  DFFR_X1 \predict_PC_reg[10][23]  ( .D(target_PC_i[23]), .CK(net338327), .RN(
        n40), .Q(\predict_PC[10][23] ) );
  DFFR_X1 \predict_PC_reg[10][22]  ( .D(target_PC_i[22]), .CK(net338327), .RN(
        n39), .Q(\predict_PC[10][22] ) );
  DFFR_X1 \predict_PC_reg[10][21]  ( .D(target_PC_i[21]), .CK(net338327), .RN(
        n37), .Q(\predict_PC[10][21] ) );
  DFFR_X1 \predict_PC_reg[10][20]  ( .D(target_PC_i[20]), .CK(net338327), .RN(
        n36), .Q(\predict_PC[10][20] ) );
  DFFR_X1 \predict_PC_reg[10][19]  ( .D(target_PC_i[19]), .CK(net338327), .RN(
        n35), .Q(\predict_PC[10][19] ) );
  DFFR_X1 \predict_PC_reg[10][18]  ( .D(target_PC_i[18]), .CK(net338327), .RN(
        n34), .Q(\predict_PC[10][18] ) );
  DFFR_X1 \predict_PC_reg[10][17]  ( .D(target_PC_i[17]), .CK(net338327), .RN(
        n30), .Q(\predict_PC[10][17] ) );
  DFFR_X1 \predict_PC_reg[10][16]  ( .D(target_PC_i[16]), .CK(net338327), .RN(
        n31), .Q(\predict_PC[10][16] ) );
  DFFR_X1 \predict_PC_reg[10][15]  ( .D(target_PC_i[15]), .CK(net338327), .RN(
        n28), .Q(\predict_PC[10][15] ) );
  DFFR_X1 \predict_PC_reg[10][14]  ( .D(target_PC_i[14]), .CK(net338327), .RN(
        n45), .Q(\predict_PC[10][14] ) );
  DFFR_X1 \predict_PC_reg[10][13]  ( .D(target_PC_i[13]), .CK(net338327), .RN(
        n37), .Q(\predict_PC[10][13] ) );
  DFFR_X1 \predict_PC_reg[10][12]  ( .D(target_PC_i[12]), .CK(net338327), .RN(
        n43), .Q(\predict_PC[10][12] ) );
  DFFR_X1 \predict_PC_reg[10][11]  ( .D(target_PC_i[11]), .CK(net338327), .RN(
        n42), .Q(\predict_PC[10][11] ) );
  DFFR_X1 \predict_PC_reg[10][10]  ( .D(target_PC_i[10]), .CK(net338327), .RN(
        n41), .Q(\predict_PC[10][10] ) );
  DFFR_X1 \predict_PC_reg[10][9]  ( .D(target_PC_i[9]), .CK(net338327), .RN(
        n40), .Q(\predict_PC[10][9] ) );
  DFFR_X1 \predict_PC_reg[10][8]  ( .D(target_PC_i[8]), .CK(net338327), .RN(
        n39), .Q(\predict_PC[10][8] ) );
  DFFR_X1 \predict_PC_reg[10][7]  ( .D(target_PC_i[7]), .CK(net338327), .RN(
        n37), .Q(\predict_PC[10][7] ) );
  DFFR_X1 \predict_PC_reg[10][6]  ( .D(target_PC_i[6]), .CK(net338327), .RN(
        n36), .Q(\predict_PC[10][6] ) );
  DFFR_X1 \predict_PC_reg[10][5]  ( .D(target_PC_i[5]), .CK(net338327), .RN(
        n38), .Q(\predict_PC[10][5] ) );
  DFFR_X1 \predict_PC_reg[10][4]  ( .D(target_PC_i[4]), .CK(net338327), .RN(
        n44), .Q(\predict_PC[10][4] ) );
  DFFR_X1 \predict_PC_reg[10][3]  ( .D(target_PC_i[3]), .CK(net338327), .RN(
        n38), .Q(\predict_PC[10][3] ) );
  DFFR_X1 \predict_PC_reg[10][2]  ( .D(target_PC_i[2]), .CK(net338327), .RN(
        n43), .Q(\predict_PC[10][2] ) );
  DFFR_X1 \predict_PC_reg[10][1]  ( .D(target_PC_i[1]), .CK(net338327), .RN(
        n38), .Q(\predict_PC[10][1] ) );
  DFFR_X1 \predict_PC_reg[10][0]  ( .D(target_PC_i[0]), .CK(net338327), .RN(
        n41), .Q(\predict_PC[10][0] ) );
  DFFR_X1 \predict_PC_reg[11][31]  ( .D(target_PC_i[31]), .CK(net338332), .RN(
        n34), .Q(\predict_PC[11][31] ) );
  DFFR_X1 \predict_PC_reg[11][30]  ( .D(target_PC_i[30]), .CK(net338332), .RN(
        n40), .Q(\predict_PC[11][30] ) );
  DFFR_X1 \predict_PC_reg[11][29]  ( .D(target_PC_i[29]), .CK(net338332), .RN(
        n39), .Q(\predict_PC[11][29] ) );
  DFFR_X1 \predict_PC_reg[11][28]  ( .D(target_PC_i[28]), .CK(net338332), .RN(
        n37), .Q(\predict_PC[11][28] ) );
  DFFR_X1 \predict_PC_reg[11][27]  ( .D(target_PC_i[27]), .CK(net338332), .RN(
        n36), .Q(\predict_PC[11][27] ) );
  DFFR_X1 \predict_PC_reg[11][26]  ( .D(target_PC_i[26]), .CK(net338332), .RN(
        n35), .Q(\predict_PC[11][26] ) );
  DFFR_X1 \predict_PC_reg[11][25]  ( .D(target_PC_i[25]), .CK(net338332), .RN(
        n45), .Q(\predict_PC[11][25] ) );
  DFFR_X1 \predict_PC_reg[11][24]  ( .D(target_PC_i[24]), .CK(net338332), .RN(
        n45), .Q(\predict_PC[11][24] ) );
  DFFR_X1 \predict_PC_reg[11][23]  ( .D(target_PC_i[23]), .CK(net338332), .RN(
        n44), .Q(\predict_PC[11][23] ) );
  DFFR_X1 \predict_PC_reg[11][22]  ( .D(target_PC_i[22]), .CK(net338332), .RN(
        n43), .Q(\predict_PC[11][22] ) );
  DFFR_X1 \predict_PC_reg[11][21]  ( .D(target_PC_i[21]), .CK(net338332), .RN(
        n42), .Q(\predict_PC[11][21] ) );
  DFFR_X1 \predict_PC_reg[11][20]  ( .D(target_PC_i[20]), .CK(net338332), .RN(
        n41), .Q(\predict_PC[11][20] ) );
  DFFR_X1 \predict_PC_reg[11][19]  ( .D(target_PC_i[19]), .CK(net338332), .RN(
        n42), .Q(\predict_PC[11][19] ) );
  DFFR_X1 \predict_PC_reg[11][18]  ( .D(target_PC_i[18]), .CK(net338332), .RN(
        n39), .Q(\predict_PC[11][18] ) );
  DFFR_X1 \predict_PC_reg[11][17]  ( .D(target_PC_i[17]), .CK(net338332), .RN(
        n37), .Q(\predict_PC[11][17] ) );
  DFFR_X1 \predict_PC_reg[11][16]  ( .D(target_PC_i[16]), .CK(net338332), .RN(
        n36), .Q(\predict_PC[11][16] ) );
  DFFR_X1 \predict_PC_reg[11][15]  ( .D(target_PC_i[15]), .CK(net338332), .RN(
        n35), .Q(\predict_PC[11][15] ) );
  DFFR_X1 \predict_PC_reg[11][14]  ( .D(target_PC_i[14]), .CK(net338332), .RN(
        n34), .Q(\predict_PC[11][14] ) );
  DFFR_X1 \predict_PC_reg[11][13]  ( .D(target_PC_i[13]), .CK(net338332), .RN(
        n44), .Q(\predict_PC[11][13] ) );
  DFFR_X1 \predict_PC_reg[11][12]  ( .D(target_PC_i[12]), .CK(net338332), .RN(
        n44), .Q(\predict_PC[11][12] ) );
  DFFR_X1 \predict_PC_reg[11][11]  ( .D(target_PC_i[11]), .CK(net338332), .RN(
        n44), .Q(\predict_PC[11][11] ) );
  DFFR_X1 \predict_PC_reg[11][10]  ( .D(target_PC_i[10]), .CK(net338332), .RN(
        n44), .Q(\predict_PC[11][10] ) );
  DFFR_X1 \predict_PC_reg[11][9]  ( .D(target_PC_i[9]), .CK(net338332), .RN(
        n44), .Q(\predict_PC[11][9] ) );
  DFFR_X1 \predict_PC_reg[11][8]  ( .D(target_PC_i[8]), .CK(net338332), .RN(
        n44), .Q(\predict_PC[11][8] ) );
  DFFR_X1 \predict_PC_reg[11][7]  ( .D(target_PC_i[7]), .CK(net338332), .RN(
        n44), .Q(\predict_PC[11][7] ) );
  DFFR_X1 \predict_PC_reg[11][6]  ( .D(target_PC_i[6]), .CK(net338332), .RN(
        n44), .Q(\predict_PC[11][6] ) );
  DFFR_X1 \predict_PC_reg[11][5]  ( .D(target_PC_i[5]), .CK(net338332), .RN(
        n40), .Q(\predict_PC[11][5] ) );
  DFFR_X1 \predict_PC_reg[11][4]  ( .D(target_PC_i[4]), .CK(net338332), .RN(
        n44), .Q(\predict_PC[11][4] ) );
  DFFR_X1 \predict_PC_reg[11][3]  ( .D(target_PC_i[3]), .CK(net338332), .RN(
        n44), .Q(\predict_PC[11][3] ) );
  DFFR_X1 \predict_PC_reg[11][2]  ( .D(target_PC_i[2]), .CK(net338332), .RN(
        n44), .Q(\predict_PC[11][2] ) );
  DFFR_X1 \predict_PC_reg[11][1]  ( .D(target_PC_i[1]), .CK(net338332), .RN(
        n45), .Q(\predict_PC[11][1] ) );
  DFFR_X1 \predict_PC_reg[11][0]  ( .D(target_PC_i[0]), .CK(net338332), .RN(
        n45), .Q(\predict_PC[11][0] ) );
  DFFR_X1 \predict_PC_reg[12][31]  ( .D(target_PC_i[31]), .CK(net338337), .RN(
        n45), .Q(\predict_PC[12][31] ) );
  DFFR_X1 \predict_PC_reg[12][30]  ( .D(target_PC_i[30]), .CK(net338337), .RN(
        n45), .Q(\predict_PC[12][30] ) );
  DFFR_X1 \predict_PC_reg[12][29]  ( .D(target_PC_i[29]), .CK(net338337), .RN(
        n45), .Q(\predict_PC[12][29] ) );
  DFFR_X1 \predict_PC_reg[12][28]  ( .D(target_PC_i[28]), .CK(net338337), .RN(
        n45), .Q(\predict_PC[12][28] ) );
  DFFR_X1 \predict_PC_reg[12][27]  ( .D(target_PC_i[27]), .CK(net338337), .RN(
        n45), .Q(\predict_PC[12][27] ) );
  DFFR_X1 \predict_PC_reg[12][26]  ( .D(target_PC_i[26]), .CK(net338337), .RN(
        n45), .Q(\predict_PC[12][26] ) );
  DFFR_X1 \predict_PC_reg[12][25]  ( .D(target_PC_i[25]), .CK(net338337), .RN(
        n45), .Q(\predict_PC[12][25] ) );
  DFFR_X1 \predict_PC_reg[12][24]  ( .D(target_PC_i[24]), .CK(net338337), .RN(
        n45), .Q(\predict_PC[12][24] ) );
  DFFR_X1 \predict_PC_reg[12][23]  ( .D(target_PC_i[23]), .CK(net338337), .RN(
        n44), .Q(\predict_PC[12][23] ) );
  DFFR_X1 \predict_PC_reg[12][22]  ( .D(target_PC_i[22]), .CK(net338337), .RN(
        n45), .Q(\predict_PC[12][22] ) );
  DFFR_X1 \predict_PC_reg[12][21]  ( .D(target_PC_i[21]), .CK(net338337), .RN(
        n24), .Q(\predict_PC[12][21] ) );
  DFFR_X1 \predict_PC_reg[12][20]  ( .D(target_PC_i[20]), .CK(net338337), .RN(
        n24), .Q(\predict_PC[12][20] ) );
  DFFR_X1 \predict_PC_reg[12][19]  ( .D(target_PC_i[19]), .CK(net338337), .RN(
        n23), .Q(\predict_PC[12][19] ) );
  DFFR_X1 \predict_PC_reg[12][18]  ( .D(target_PC_i[18]), .CK(net338337), .RN(
        n23), .Q(\predict_PC[12][18] ) );
  DFFR_X1 \predict_PC_reg[12][17]  ( .D(target_PC_i[17]), .CK(net338337), .RN(
        n24), .Q(\predict_PC[12][17] ) );
  DFFR_X1 \predict_PC_reg[12][16]  ( .D(target_PC_i[16]), .CK(net338337), .RN(
        n22), .Q(\predict_PC[12][16] ) );
  DFFR_X1 \predict_PC_reg[12][15]  ( .D(target_PC_i[15]), .CK(net338337), .RN(
        n22), .Q(\predict_PC[12][15] ) );
  DFFR_X1 \predict_PC_reg[12][14]  ( .D(target_PC_i[14]), .CK(net338337), .RN(
        n22), .Q(\predict_PC[12][14] ) );
  DFFR_X1 \predict_PC_reg[12][13]  ( .D(target_PC_i[13]), .CK(net338337), .RN(
        n23), .Q(\predict_PC[12][13] ) );
  DFFR_X1 \predict_PC_reg[12][12]  ( .D(target_PC_i[12]), .CK(net338337), .RN(
        n24), .Q(\predict_PC[12][12] ) );
  DFFR_X1 \predict_PC_reg[12][11]  ( .D(target_PC_i[11]), .CK(net338337), .RN(
        n45), .Q(\predict_PC[12][11] ) );
  DFFR_X1 \predict_PC_reg[12][10]  ( .D(target_PC_i[10]), .CK(net338337), .RN(
        n38), .Q(\predict_PC[12][10] ) );
  DFFR_X1 \predict_PC_reg[12][9]  ( .D(target_PC_i[9]), .CK(net338337), .RN(
        n35), .Q(\predict_PC[12][9] ) );
  DFFR_X1 \predict_PC_reg[12][8]  ( .D(target_PC_i[8]), .CK(net338337), .RN(
        n34), .Q(\predict_PC[12][8] ) );
  DFFR_X1 \predict_PC_reg[12][7]  ( .D(target_PC_i[7]), .CK(net338337), .RN(
        n42), .Q(\predict_PC[12][7] ) );
  DFFR_X1 \predict_PC_reg[12][6]  ( .D(target_PC_i[6]), .CK(net338337), .RN(
        n33), .Q(\predict_PC[12][6] ) );
  DFFR_X1 \predict_PC_reg[12][5]  ( .D(target_PC_i[5]), .CK(net338337), .RN(
        n33), .Q(\predict_PC[12][5] ) );
  DFFR_X1 \predict_PC_reg[12][4]  ( .D(target_PC_i[4]), .CK(net338337), .RN(
        n38), .Q(\predict_PC[12][4] ) );
  DFFR_X1 \predict_PC_reg[12][3]  ( .D(target_PC_i[3]), .CK(net338337), .RN(
        n33), .Q(\predict_PC[12][3] ) );
  DFFR_X1 \predict_PC_reg[12][2]  ( .D(target_PC_i[2]), .CK(net338337), .RN(
        n33), .Q(\predict_PC[12][2] ) );
  DFFR_X1 \predict_PC_reg[12][1]  ( .D(target_PC_i[1]), .CK(net338337), .RN(
        n33), .Q(\predict_PC[12][1] ) );
  DFFR_X1 \predict_PC_reg[12][0]  ( .D(target_PC_i[0]), .CK(net338337), .RN(
        n33), .Q(\predict_PC[12][0] ) );
  DFFR_X1 \predict_PC_reg[13][31]  ( .D(target_PC_i[31]), .CK(net338342), .RN(
        n33), .Q(\predict_PC[13][31] ) );
  DFFR_X1 \predict_PC_reg[13][30]  ( .D(target_PC_i[30]), .CK(net338342), .RN(
        n33), .Q(\predict_PC[13][30] ) );
  DFFR_X1 \predict_PC_reg[13][29]  ( .D(target_PC_i[29]), .CK(net338342), .RN(
        n33), .Q(\predict_PC[13][29] ) );
  DFFR_X1 \predict_PC_reg[13][28]  ( .D(target_PC_i[28]), .CK(net338342), .RN(
        n33), .Q(\predict_PC[13][28] ) );
  DFFR_X1 \predict_PC_reg[13][27]  ( .D(target_PC_i[27]), .CK(net338342), .RN(
        n33), .Q(\predict_PC[13][27] ) );
  DFFR_X1 \predict_PC_reg[13][26]  ( .D(target_PC_i[26]), .CK(net338342), .RN(
        n33), .Q(\predict_PC[13][26] ) );
  DFFR_X1 \predict_PC_reg[13][25]  ( .D(target_PC_i[25]), .CK(net338342), .RN(
        n33), .Q(\predict_PC[13][25] ) );
  DFFR_X1 \predict_PC_reg[13][24]  ( .D(target_PC_i[24]), .CK(net338342), .RN(
        n33), .Q(\predict_PC[13][24] ) );
  DFFR_X1 \predict_PC_reg[13][23]  ( .D(target_PC_i[23]), .CK(net338342), .RN(
        n34), .Q(\predict_PC[13][23] ) );
  DFFR_X1 \predict_PC_reg[13][22]  ( .D(target_PC_i[22]), .CK(net338342), .RN(
        n34), .Q(\predict_PC[13][22] ) );
  DFFR_X1 \predict_PC_reg[13][21]  ( .D(target_PC_i[21]), .CK(net338342), .RN(
        n34), .Q(\predict_PC[13][21] ) );
  DFFR_X1 \predict_PC_reg[13][20]  ( .D(target_PC_i[20]), .CK(net338342), .RN(
        n34), .Q(\predict_PC[13][20] ) );
  DFFR_X1 \predict_PC_reg[13][19]  ( .D(target_PC_i[19]), .CK(net338342), .RN(
        n34), .Q(\predict_PC[13][19] ) );
  DFFR_X1 \predict_PC_reg[13][18]  ( .D(target_PC_i[18]), .CK(net338342), .RN(
        n34), .Q(\predict_PC[13][18] ) );
  DFFR_X1 \predict_PC_reg[13][17]  ( .D(target_PC_i[17]), .CK(net338342), .RN(
        n34), .Q(\predict_PC[13][17] ) );
  DFFR_X1 \predict_PC_reg[13][16]  ( .D(target_PC_i[16]), .CK(net338342), .RN(
        n34), .Q(\predict_PC[13][16] ) );
  DFFR_X1 \predict_PC_reg[13][15]  ( .D(target_PC_i[15]), .CK(net338342), .RN(
        n34), .Q(\predict_PC[13][15] ) );
  DFFR_X1 \predict_PC_reg[13][14]  ( .D(target_PC_i[14]), .CK(net338342), .RN(
        n34), .Q(\predict_PC[13][14] ) );
  DFFR_X1 \predict_PC_reg[13][13]  ( .D(target_PC_i[13]), .CK(net338342), .RN(
        n34), .Q(\predict_PC[13][13] ) );
  DFFR_X1 \predict_PC_reg[13][12]  ( .D(target_PC_i[12]), .CK(net338342), .RN(
        n34), .Q(\predict_PC[13][12] ) );
  DFFR_X1 \predict_PC_reg[13][11]  ( .D(target_PC_i[11]), .CK(net338342), .RN(
        n35), .Q(\predict_PC[13][11] ) );
  DFFR_X1 \predict_PC_reg[13][10]  ( .D(target_PC_i[10]), .CK(net338342), .RN(
        n35), .Q(\predict_PC[13][10] ) );
  DFFR_X1 \predict_PC_reg[13][9]  ( .D(target_PC_i[9]), .CK(net338342), .RN(
        n35), .Q(\predict_PC[13][9] ) );
  DFFR_X1 \predict_PC_reg[13][8]  ( .D(target_PC_i[8]), .CK(net338342), .RN(
        n35), .Q(\predict_PC[13][8] ) );
  DFFR_X1 \predict_PC_reg[13][7]  ( .D(target_PC_i[7]), .CK(net338342), .RN(
        n35), .Q(\predict_PC[13][7] ) );
  DFFR_X1 \predict_PC_reg[13][6]  ( .D(target_PC_i[6]), .CK(net338342), .RN(
        n35), .Q(\predict_PC[13][6] ) );
  DFFR_X1 \predict_PC_reg[13][5]  ( .D(target_PC_i[5]), .CK(net338342), .RN(
        n35), .Q(\predict_PC[13][5] ) );
  DFFR_X1 \predict_PC_reg[13][4]  ( .D(target_PC_i[4]), .CK(net338342), .RN(
        n35), .Q(\predict_PC[13][4] ) );
  DFFR_X1 \predict_PC_reg[13][3]  ( .D(target_PC_i[3]), .CK(net338342), .RN(
        n35), .Q(\predict_PC[13][3] ) );
  DFFR_X1 \predict_PC_reg[13][2]  ( .D(target_PC_i[2]), .CK(net338342), .RN(
        n35), .Q(\predict_PC[13][2] ) );
  DFFR_X1 \predict_PC_reg[13][1]  ( .D(target_PC_i[1]), .CK(net338342), .RN(
        n35), .Q(\predict_PC[13][1] ) );
  DFFR_X1 \predict_PC_reg[13][0]  ( .D(target_PC_i[0]), .CK(net338342), .RN(
        n35), .Q(\predict_PC[13][0] ) );
  DFFR_X1 \predict_PC_reg[14][31]  ( .D(target_PC_i[31]), .CK(net338347), .RN(
        n36), .Q(\predict_PC[14][31] ) );
  DFFR_X1 \predict_PC_reg[14][30]  ( .D(target_PC_i[30]), .CK(net338347), .RN(
        n36), .Q(\predict_PC[14][30] ) );
  DFFR_X1 \predict_PC_reg[14][29]  ( .D(target_PC_i[29]), .CK(net338347), .RN(
        n36), .Q(\predict_PC[14][29] ) );
  DFFR_X1 \predict_PC_reg[14][28]  ( .D(target_PC_i[28]), .CK(net338347), .RN(
        n36), .Q(\predict_PC[14][28] ) );
  DFFR_X1 \predict_PC_reg[14][27]  ( .D(target_PC_i[27]), .CK(net338347), .RN(
        n36), .Q(\predict_PC[14][27] ) );
  DFFR_X1 \predict_PC_reg[14][26]  ( .D(target_PC_i[26]), .CK(net338347), .RN(
        n36), .Q(\predict_PC[14][26] ) );
  DFFR_X1 \predict_PC_reg[14][25]  ( .D(target_PC_i[25]), .CK(net338347), .RN(
        n36), .Q(\predict_PC[14][25] ) );
  DFFR_X1 \predict_PC_reg[14][24]  ( .D(target_PC_i[24]), .CK(net338347), .RN(
        n36), .Q(\predict_PC[14][24] ) );
  DFFR_X1 \predict_PC_reg[14][23]  ( .D(target_PC_i[23]), .CK(net338347), .RN(
        n36), .Q(\predict_PC[14][23] ) );
  DFFR_X1 \predict_PC_reg[14][22]  ( .D(target_PC_i[22]), .CK(net338347), .RN(
        n36), .Q(\predict_PC[14][22] ) );
  DFFR_X1 \predict_PC_reg[14][21]  ( .D(target_PC_i[21]), .CK(net338347), .RN(
        n36), .Q(\predict_PC[14][21] ) );
  DFFR_X1 \predict_PC_reg[14][20]  ( .D(target_PC_i[20]), .CK(net338347), .RN(
        n36), .Q(\predict_PC[14][20] ) );
  DFFR_X1 \predict_PC_reg[14][19]  ( .D(target_PC_i[19]), .CK(net338347), .RN(
        n37), .Q(\predict_PC[14][19] ) );
  DFFR_X1 \predict_PC_reg[14][18]  ( .D(target_PC_i[18]), .CK(net338347), .RN(
        n37), .Q(\predict_PC[14][18] ) );
  DFFR_X1 \predict_PC_reg[14][17]  ( .D(target_PC_i[17]), .CK(net338347), .RN(
        n37), .Q(\predict_PC[14][17] ) );
  DFFR_X1 \predict_PC_reg[14][16]  ( .D(target_PC_i[16]), .CK(net338347), .RN(
        n37), .Q(\predict_PC[14][16] ) );
  DFFR_X1 \predict_PC_reg[14][15]  ( .D(target_PC_i[15]), .CK(net338347), .RN(
        n37), .Q(\predict_PC[14][15] ) );
  DFFR_X1 \predict_PC_reg[14][14]  ( .D(target_PC_i[14]), .CK(net338347), .RN(
        n37), .Q(\predict_PC[14][14] ) );
  DFFR_X1 \predict_PC_reg[14][13]  ( .D(target_PC_i[13]), .CK(net338347), .RN(
        n37), .Q(\predict_PC[14][13] ) );
  DFFR_X1 \predict_PC_reg[14][12]  ( .D(target_PC_i[12]), .CK(net338347), .RN(
        n37), .Q(\predict_PC[14][12] ) );
  DFFR_X1 \predict_PC_reg[14][11]  ( .D(target_PC_i[11]), .CK(net338347), .RN(
        n37), .Q(\predict_PC[14][11] ) );
  DFFR_X1 \predict_PC_reg[14][10]  ( .D(target_PC_i[10]), .CK(net338347), .RN(
        n37), .Q(\predict_PC[14][10] ) );
  DFFR_X1 \predict_PC_reg[14][9]  ( .D(target_PC_i[9]), .CK(net338347), .RN(
        n37), .Q(\predict_PC[14][9] ) );
  DFFR_X1 \predict_PC_reg[14][8]  ( .D(target_PC_i[8]), .CK(net338347), .RN(
        n37), .Q(\predict_PC[14][8] ) );
  DFFR_X1 \predict_PC_reg[14][7]  ( .D(target_PC_i[7]), .CK(net338347), .RN(
        n38), .Q(\predict_PC[14][7] ) );
  DFFR_X1 \predict_PC_reg[14][6]  ( .D(target_PC_i[6]), .CK(net338347), .RN(
        n38), .Q(\predict_PC[14][6] ) );
  DFFR_X1 \predict_PC_reg[14][5]  ( .D(target_PC_i[5]), .CK(net338347), .RN(
        n38), .Q(\predict_PC[14][5] ) );
  DFFR_X1 \predict_PC_reg[14][4]  ( .D(target_PC_i[4]), .CK(net338347), .RN(
        n38), .Q(\predict_PC[14][4] ) );
  DFFR_X1 \predict_PC_reg[14][3]  ( .D(target_PC_i[3]), .CK(net338347), .RN(
        n33), .Q(\predict_PC[14][3] ) );
  DFFR_X1 \predict_PC_reg[14][2]  ( .D(target_PC_i[2]), .CK(net338347), .RN(
        n38), .Q(\predict_PC[14][2] ) );
  DFFR_X1 \predict_PC_reg[14][1]  ( .D(target_PC_i[1]), .CK(net338347), .RN(
        n38), .Q(\predict_PC[14][1] ) );
  DFFR_X1 \predict_PC_reg[14][0]  ( .D(target_PC_i[0]), .CK(net338347), .RN(
        n38), .Q(\predict_PC[14][0] ) );
  DFFR_X1 \predict_PC_reg[15][31]  ( .D(target_PC_i[31]), .CK(net338352), .RN(
        n38), .Q(\predict_PC[15][31] ) );
  DFFR_X1 \last_PC_reg[31]  ( .D(predicted_next_PC_o[31]), .CK(net338272), 
        .RN(n38), .QN(n483) );
  DFFR_X1 \predict_PC_reg[15][30]  ( .D(target_PC_i[30]), .CK(net338352), .RN(
        n38), .Q(\predict_PC[15][30] ) );
  DFFR_X1 \last_PC_reg[30]  ( .D(predicted_next_PC_o[30]), .CK(net338272), 
        .RN(n38), .QN(n485) );
  DFFR_X1 \predict_PC_reg[15][29]  ( .D(target_PC_i[29]), .CK(net338352), .RN(
        n39), .Q(\predict_PC[15][29] ) );
  DFFR_X1 \last_PC_reg[29]  ( .D(predicted_next_PC_o[29]), .CK(net338272), 
        .RN(n39), .QN(n487) );
  DFFR_X1 \predict_PC_reg[15][28]  ( .D(target_PC_i[28]), .CK(net338352), .RN(
        n39), .Q(\predict_PC[15][28] ) );
  DFFR_X1 \last_PC_reg[28]  ( .D(predicted_next_PC_o[28]), .CK(net338272), 
        .RN(n39), .QN(n489) );
  DFFR_X1 \predict_PC_reg[15][27]  ( .D(target_PC_i[27]), .CK(net338352), .RN(
        n39), .Q(\predict_PC[15][27] ) );
  DFFR_X1 \last_PC_reg[27]  ( .D(predicted_next_PC_o[27]), .CK(net338272), 
        .RN(n39), .QN(n491) );
  DFFR_X1 \predict_PC_reg[15][26]  ( .D(target_PC_i[26]), .CK(net338352), .RN(
        n39), .Q(\predict_PC[15][26] ) );
  DFFR_X1 \last_PC_reg[26]  ( .D(predicted_next_PC_o[26]), .CK(net338272), 
        .RN(n39), .QN(n493) );
  DFFR_X1 \predict_PC_reg[15][25]  ( .D(target_PC_i[25]), .CK(net338352), .RN(
        n39), .Q(\predict_PC[15][25] ) );
  DFFR_X1 \last_PC_reg[25]  ( .D(predicted_next_PC_o[25]), .CK(net338272), 
        .RN(n39), .QN(n495) );
  DFFR_X1 \predict_PC_reg[15][24]  ( .D(target_PC_i[24]), .CK(net338352), .RN(
        n39), .Q(\predict_PC[15][24] ) );
  DFFR_X1 \last_PC_reg[24]  ( .D(predicted_next_PC_o[24]), .CK(net338272), 
        .RN(n39), .QN(n497) );
  DFFR_X1 \predict_PC_reg[15][23]  ( .D(target_PC_i[23]), .CK(net338352), .RN(
        n40), .Q(\predict_PC[15][23] ) );
  DFFR_X1 \last_PC_reg[23]  ( .D(predicted_next_PC_o[23]), .CK(net338272), 
        .RN(n40), .QN(n499) );
  DFFR_X1 \predict_PC_reg[15][22]  ( .D(target_PC_i[22]), .CK(net338352), .RN(
        n40), .Q(\predict_PC[15][22] ) );
  DFFR_X1 \last_PC_reg[22]  ( .D(predicted_next_PC_o[22]), .CK(net338272), 
        .RN(n40), .QN(n501) );
  DFFR_X1 \predict_PC_reg[15][21]  ( .D(target_PC_i[21]), .CK(net338352), .RN(
        n40), .Q(\predict_PC[15][21] ) );
  DFFR_X1 \last_PC_reg[21]  ( .D(predicted_next_PC_o[21]), .CK(net338272), 
        .RN(n40), .QN(n503) );
  DFFR_X1 \predict_PC_reg[15][20]  ( .D(target_PC_i[20]), .CK(net338352), .RN(
        n40), .Q(\predict_PC[15][20] ) );
  DFFR_X1 \last_PC_reg[20]  ( .D(predicted_next_PC_o[20]), .CK(net338272), 
        .RN(n40), .QN(n505) );
  DFFR_X1 \predict_PC_reg[15][19]  ( .D(target_PC_i[19]), .CK(net338352), .RN(
        n40), .Q(\predict_PC[15][19] ) );
  DFFR_X1 \last_PC_reg[19]  ( .D(predicted_next_PC_o[19]), .CK(net338272), 
        .RN(n40), .QN(n507) );
  DFFR_X1 \predict_PC_reg[15][18]  ( .D(target_PC_i[18]), .CK(net338352), .RN(
        n40), .Q(\predict_PC[15][18] ) );
  DFFR_X1 \last_PC_reg[18]  ( .D(predicted_next_PC_o[18]), .CK(net338272), 
        .RN(n40), .QN(n509) );
  DFFR_X1 \predict_PC_reg[15][17]  ( .D(target_PC_i[17]), .CK(net338352), .RN(
        n41), .Q(\predict_PC[15][17] ) );
  DFFR_X1 \last_PC_reg[17]  ( .D(predicted_next_PC_o[17]), .CK(net338272), 
        .RN(n41), .QN(n511) );
  DFFR_X1 \predict_PC_reg[15][16]  ( .D(target_PC_i[16]), .CK(net338352), .RN(
        n41), .Q(\predict_PC[15][16] ) );
  DFFR_X1 \last_PC_reg[16]  ( .D(predicted_next_PC_o[16]), .CK(net338272), 
        .RN(n41), .QN(n513) );
  DFFR_X1 \predict_PC_reg[15][15]  ( .D(target_PC_i[15]), .CK(net338352), .RN(
        n41), .Q(\predict_PC[15][15] ) );
  DFFR_X1 \last_PC_reg[15]  ( .D(predicted_next_PC_o[15]), .CK(net338272), 
        .RN(n41), .QN(n515) );
  DFFR_X1 \predict_PC_reg[15][14]  ( .D(target_PC_i[14]), .CK(net338352), .RN(
        n41), .Q(\predict_PC[15][14] ) );
  DFFR_X1 \last_PC_reg[14]  ( .D(predicted_next_PC_o[14]), .CK(net338272), 
        .RN(n41), .QN(n517) );
  DFFR_X1 \predict_PC_reg[15][13]  ( .D(target_PC_i[13]), .CK(net338352), .RN(
        n41), .Q(\predict_PC[15][13] ) );
  DFFR_X1 \last_PC_reg[13]  ( .D(predicted_next_PC_o[13]), .CK(net338272), 
        .RN(n41), .QN(n519) );
  DFFR_X1 \predict_PC_reg[15][12]  ( .D(target_PC_i[12]), .CK(net338352), .RN(
        n41), .Q(\predict_PC[15][12] ) );
  DFFR_X1 \last_PC_reg[12]  ( .D(predicted_next_PC_o[12]), .CK(net338272), 
        .RN(n41), .QN(n521) );
  DFFR_X1 \predict_PC_reg[15][11]  ( .D(target_PC_i[11]), .CK(net338352), .RN(
        n42), .Q(\predict_PC[15][11] ) );
  DFFR_X1 \last_PC_reg[11]  ( .D(predicted_next_PC_o[11]), .CK(net338272), 
        .RN(n42), .QN(n523) );
  DFFR_X1 \predict_PC_reg[15][10]  ( .D(target_PC_i[10]), .CK(net338352), .RN(
        n42), .Q(\predict_PC[15][10] ) );
  DFFR_X1 \last_PC_reg[10]  ( .D(predicted_next_PC_o[10]), .CK(net338272), 
        .RN(n42), .QN(n525) );
  DFFR_X1 \predict_PC_reg[15][9]  ( .D(target_PC_i[9]), .CK(net338352), .RN(
        n42), .Q(\predict_PC[15][9] ) );
  DFFR_X1 \last_PC_reg[9]  ( .D(predicted_next_PC_o[9]), .CK(net338272), .RN(
        n42), .QN(n527) );
  DFFR_X1 \predict_PC_reg[15][8]  ( .D(target_PC_i[8]), .CK(net338352), .RN(
        n42), .Q(\predict_PC[15][8] ) );
  DFFR_X1 \last_PC_reg[8]  ( .D(predicted_next_PC_o[8]), .CK(net338272), .RN(
        n42), .QN(n529) );
  DFFR_X1 \predict_PC_reg[15][7]  ( .D(target_PC_i[7]), .CK(net338352), .RN(
        n42), .Q(\predict_PC[15][7] ) );
  DFFR_X1 \last_PC_reg[7]  ( .D(predicted_next_PC_o[7]), .CK(net338272), .RN(
        n42), .QN(n531) );
  DFFR_X1 \predict_PC_reg[15][6]  ( .D(target_PC_i[6]), .CK(net338352), .RN(
        n42), .Q(\predict_PC[15][6] ) );
  DFFR_X1 \last_PC_reg[6]  ( .D(predicted_next_PC_o[6]), .CK(net338272), .RN(
        n42), .QN(n533) );
  DFFR_X1 \predict_PC_reg[15][5]  ( .D(target_PC_i[5]), .CK(net338352), .RN(
        n43), .Q(\predict_PC[15][5] ) );
  DFFR_X1 \last_PC_reg[5]  ( .D(predicted_next_PC_o[5]), .CK(net338272), .RN(
        n43), .QN(n535) );
  DFFR_X1 \predict_PC_reg[15][4]  ( .D(target_PC_i[4]), .CK(net338352), .RN(
        n43), .Q(\predict_PC[15][4] ) );
  DFFR_X1 \last_PC_reg[4]  ( .D(predicted_next_PC_o[4]), .CK(net338272), .RN(
        n43), .QN(n537) );
  DFFR_X1 \predict_PC_reg[15][3]  ( .D(target_PC_i[3]), .CK(net338352), .RN(
        n43), .Q(\predict_PC[15][3] ) );
  DFFR_X1 \last_PC_reg[3]  ( .D(predicted_next_PC_o[3]), .CK(net338272), .RN(
        n43), .QN(n539) );
  DFFR_X1 \predict_PC_reg[15][2]  ( .D(target_PC_i[2]), .CK(net338352), .RN(
        n43), .Q(\predict_PC[15][2] ) );
  DFFR_X1 \last_PC_reg[2]  ( .D(predicted_next_PC_o[2]), .CK(net338272), .RN(
        n43), .QN(n541) );
  DFFR_X1 \predict_PC_reg[15][1]  ( .D(target_PC_i[1]), .CK(net338352), .RN(
        n43), .Q(\predict_PC[15][1] ) );
  DFFR_X1 \last_PC_reg[1]  ( .D(predicted_next_PC_o[1]), .CK(net338272), .RN(
        n43), .QN(n543) );
  DFFR_X1 \predict_PC_reg[15][0]  ( .D(target_PC_i[0]), .CK(net338352), .RN(
        n43), .Q(\predict_PC[15][0] ) );
  DFFR_X1 \last_PC_reg[0]  ( .D(predicted_next_PC_o[0]), .CK(net338272), .RN(
        n43), .QN(n545) );
  DFFR_X1 last_mispredict_reg ( .D(mispredict_o), .CK(net338272), .RN(n36), 
        .QN(n546) );
  predictor_2_0 pred_x_0 ( .clock(clock), .reset(reset), .enable(
        write_enable[0]), .taken_i(was_taken_i), .prediction_o(taken[0]) );
  predictor_2_15 pred_x_1 ( .clock(clock), .reset(reset), .enable(
        write_enable[1]), .taken_i(was_taken_i), .prediction_o(taken[1]) );
  predictor_2_14 pred_x_2 ( .clock(clock), .reset(reset), .enable(
        write_enable[2]), .taken_i(was_taken_i), .prediction_o(taken[2]) );
  predictor_2_13 pred_x_3 ( .clock(clock), .reset(reset), .enable(
        write_enable[3]), .taken_i(was_taken_i), .prediction_o(taken[3]) );
  predictor_2_12 pred_x_4 ( .clock(clock), .reset(reset), .enable(
        write_enable[4]), .taken_i(was_taken_i), .prediction_o(taken[4]) );
  predictor_2_11 pred_x_5 ( .clock(clock), .reset(reset), .enable(
        write_enable[5]), .taken_i(was_taken_i), .prediction_o(taken[5]) );
  predictor_2_10 pred_x_6 ( .clock(clock), .reset(reset), .enable(
        write_enable[6]), .taken_i(was_taken_i), .prediction_o(taken[6]) );
  predictor_2_9 pred_x_7 ( .clock(clock), .reset(reset), .enable(
        write_enable[7]), .taken_i(was_taken_i), .prediction_o(taken[7]) );
  predictor_2_8 pred_x_8 ( .clock(clock), .reset(reset), .enable(
        write_enable[8]), .taken_i(was_taken_i), .prediction_o(taken[8]) );
  predictor_2_7 pred_x_9 ( .clock(clock), .reset(reset), .enable(
        write_enable[9]), .taken_i(was_taken_i), .prediction_o(taken[9]) );
  predictor_2_6 pred_x_10 ( .clock(clock), .reset(reset), .enable(
        write_enable[10]), .taken_i(was_taken_i), .prediction_o(taken[10]) );
  predictor_2_5 pred_x_11 ( .clock(clock), .reset(reset), .enable(
        write_enable[11]), .taken_i(was_taken_i), .prediction_o(taken[11]) );
  predictor_2_4 pred_x_12 ( .clock(clock), .reset(reset), .enable(
        write_enable[12]), .taken_i(was_taken_i), .prediction_o(taken[12]) );
  predictor_2_3 pred_x_13 ( .clock(clock), .reset(reset), .enable(
        write_enable[13]), .taken_i(was_taken_i), .prediction_o(taken[13]) );
  predictor_2_2 pred_x_14 ( .clock(clock), .reset(reset), .enable(
        write_enable[14]), .taken_i(was_taken_i), .prediction_o(taken[14]) );
  predictor_2_1 pred_x_15 ( .clock(clock), .reset(reset), .enable(
        write_enable[15]), .taken_i(was_taken_i), .prediction_o(taken[15]) );
  SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_0 clk_gate_last_TAG_reg ( .CLK(
        clock), .EN(N567), .ENCLK(net338272) );
  SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_16 \clk_gate_predict_PC_reg[0]  ( 
        .CLK(clock), .EN(N566), .ENCLK(net338277) );
  SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_15 \clk_gate_predict_PC_reg[1]  ( 
        .CLK(clock), .EN(N534), .ENCLK(net338282) );
  SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_14 \clk_gate_predict_PC_reg[2]  ( 
        .CLK(clock), .EN(N502), .ENCLK(net338287) );
  SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_13 \clk_gate_predict_PC_reg[3]  ( 
        .CLK(clock), .EN(N470), .ENCLK(net338292) );
  SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_12 \clk_gate_predict_PC_reg[4]  ( 
        .CLK(clock), .EN(N438), .ENCLK(net338297) );
  SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_11 \clk_gate_predict_PC_reg[5]  ( 
        .CLK(clock), .EN(N406), .ENCLK(net338302) );
  SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_10 \clk_gate_predict_PC_reg[6]  ( 
        .CLK(clock), .EN(N374), .ENCLK(net338307) );
  SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_9 \clk_gate_predict_PC_reg[7]  ( 
        .CLK(clock), .EN(N342), .ENCLK(net338312) );
  SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_8 \clk_gate_predict_PC_reg[8]  ( 
        .CLK(clock), .EN(N310), .ENCLK(net338317) );
  SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_7 \clk_gate_predict_PC_reg[9]  ( 
        .CLK(clock), .EN(N278), .ENCLK(net338322) );
  SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_6 \clk_gate_predict_PC_reg[10]  ( 
        .CLK(clock), .EN(N246), .ENCLK(net338327) );
  SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_5 \clk_gate_predict_PC_reg[11]  ( 
        .CLK(clock), .EN(N214), .ENCLK(net338332) );
  SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_4 \clk_gate_predict_PC_reg[12]  ( 
        .CLK(clock), .EN(N182), .ENCLK(net338337) );
  SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_3 \clk_gate_predict_PC_reg[13]  ( 
        .CLK(clock), .EN(N150), .ENCLK(net338342) );
  SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_2 \clk_gate_predict_PC_reg[14]  ( 
        .CLK(clock), .EN(N118), .ENCLK(net338347) );
  SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_1 \clk_gate_predict_PC_reg[15]  ( 
        .CLK(clock), .EN(N86), .ENCLK(net338352) );
  OAI22_X1 U434 ( .A1(target_PC_i[29]), .A2(n487), .B1(target_PC_i[28]), .B2(
        n489), .ZN(n942) );
  AOI221_X1 U433 ( .B1(target_PC_i[29]), .B2(n487), .C1(n489), .C2(
        target_PC_i[28]), .A(n942), .ZN(n935) );
  OAI22_X1 U432 ( .A1(target_PC_i[19]), .A2(n507), .B1(target_PC_i[18]), .B2(
        n509), .ZN(n941) );
  AOI221_X1 U431 ( .B1(target_PC_i[19]), .B2(n507), .C1(n509), .C2(
        target_PC_i[18]), .A(n941), .ZN(n936) );
  OAI22_X1 U430 ( .A1(target_PC_i[17]), .A2(n511), .B1(target_PC_i[16]), .B2(
        n513), .ZN(n940) );
  AOI221_X1 U429 ( .B1(target_PC_i[17]), .B2(n511), .C1(n513), .C2(
        target_PC_i[16]), .A(n940), .ZN(n937) );
  OAI22_X1 U428 ( .A1(target_PC_i[11]), .A2(n523), .B1(target_PC_i[10]), .B2(
        n525), .ZN(n939) );
  AOI221_X1 U427 ( .B1(target_PC_i[11]), .B2(n523), .C1(n525), .C2(
        target_PC_i[10]), .A(n939), .ZN(n938) );
  NAND4_X1 U426 ( .A1(n935), .A2(n936), .A3(n937), .A4(n938), .ZN(n907) );
  OAI22_X1 U425 ( .A1(target_PC_i[9]), .A2(n527), .B1(target_PC_i[8]), .B2(
        n529), .ZN(n934) );
  AOI221_X1 U424 ( .B1(target_PC_i[9]), .B2(n527), .C1(n529), .C2(
        target_PC_i[8]), .A(n934), .ZN(n927) );
  OAI22_X1 U423 ( .A1(target_PC_i[15]), .A2(n515), .B1(target_PC_i[14]), .B2(
        n517), .ZN(n933) );
  AOI221_X1 U422 ( .B1(target_PC_i[15]), .B2(n515), .C1(n517), .C2(
        target_PC_i[14]), .A(n933), .ZN(n928) );
  OAI22_X1 U421 ( .A1(target_PC_i[13]), .A2(n519), .B1(target_PC_i[12]), .B2(
        n521), .ZN(n932) );
  AOI221_X1 U420 ( .B1(target_PC_i[13]), .B2(n519), .C1(n521), .C2(
        target_PC_i[12]), .A(n932), .ZN(n929) );
  OAI22_X1 U419 ( .A1(target_PC_i[3]), .A2(n539), .B1(target_PC_i[2]), .B2(
        n541), .ZN(n931) );
  AOI221_X1 U418 ( .B1(target_PC_i[3]), .B2(n539), .C1(n541), .C2(
        target_PC_i[2]), .A(n931), .ZN(n930) );
  NAND4_X1 U417 ( .A1(n927), .A2(n928), .A3(n929), .A4(n930), .ZN(n908) );
  OAI22_X1 U416 ( .A1(target_PC_i[1]), .A2(n543), .B1(target_PC_i[0]), .B2(
        n545), .ZN(n926) );
  AOI221_X1 U415 ( .B1(target_PC_i[1]), .B2(n543), .C1(n545), .C2(
        target_PC_i[0]), .A(n926), .ZN(n919) );
  OAI22_X1 U414 ( .A1(target_PC_i[7]), .A2(n531), .B1(target_PC_i[6]), .B2(
        n533), .ZN(n925) );
  AOI221_X1 U413 ( .B1(target_PC_i[7]), .B2(n531), .C1(n533), .C2(
        target_PC_i[6]), .A(n925), .ZN(n920) );
  OAI22_X1 U412 ( .A1(target_PC_i[5]), .A2(n535), .B1(target_PC_i[4]), .B2(
        n537), .ZN(n924) );
  AOI221_X1 U411 ( .B1(target_PC_i[5]), .B2(n535), .C1(n537), .C2(
        target_PC_i[4]), .A(n924), .ZN(n921) );
  OAI22_X1 U410 ( .A1(target_PC_i[23]), .A2(n499), .B1(target_PC_i[22]), .B2(
        n501), .ZN(n923) );
  AOI221_X1 U409 ( .B1(target_PC_i[23]), .B2(n499), .C1(n501), .C2(
        target_PC_i[22]), .A(n923), .ZN(n922) );
  NAND4_X1 U408 ( .A1(n919), .A2(n920), .A3(n921), .A4(n922), .ZN(n909) );
  OAI22_X1 U407 ( .A1(target_PC_i[31]), .A2(n483), .B1(target_PC_i[30]), .B2(
        n485), .ZN(n918) );
  AOI221_X1 U406 ( .B1(target_PC_i[31]), .B2(n483), .C1(n485), .C2(
        target_PC_i[30]), .A(n918), .ZN(n911) );
  OAI22_X1 U405 ( .A1(target_PC_i[27]), .A2(n491), .B1(target_PC_i[26]), .B2(
        n493), .ZN(n917) );
  AOI221_X1 U404 ( .B1(target_PC_i[27]), .B2(n491), .C1(n493), .C2(
        target_PC_i[26]), .A(n917), .ZN(n912) );
  OAI22_X1 U403 ( .A1(target_PC_i[25]), .A2(n495), .B1(target_PC_i[24]), .B2(
        n497), .ZN(n916) );
  AOI221_X1 U402 ( .B1(target_PC_i[25]), .B2(n495), .C1(n497), .C2(
        target_PC_i[24]), .A(n916), .ZN(n913) );
  OAI22_X1 U401 ( .A1(target_PC_i[21]), .A2(n503), .B1(target_PC_i[20]), .B2(
        n505), .ZN(n915) );
  AOI221_X1 U400 ( .B1(target_PC_i[21]), .B2(n503), .C1(n505), .C2(
        target_PC_i[20]), .A(n915), .ZN(n914) );
  NAND4_X1 U399 ( .A1(n911), .A2(n912), .A3(n913), .A4(n914), .ZN(n910) );
  OAI21_X1 U397 ( .B1(was_taken_i), .B2(n5), .A(n546), .ZN(n906) );
  NAND2_X1 U391 ( .A1(TAG_i[1]), .A2(n903), .ZN(n895) );
  NAND2_X1 U390 ( .A1(TAG_i[3]), .A2(n973), .ZN(n902) );
  NAND2_X1 U388 ( .A1(TAG_i[0]), .A2(TAG_i[1]), .ZN(n894) );
  AOI22_X1 U386 ( .A1(n17), .A2(taken[10]), .B1(n16), .B2(taken[11]), .ZN(n897) );
  NAND2_X1 U383 ( .A1(TAG_i[0]), .A2(n974), .ZN(n891) );
  AOI22_X1 U381 ( .A1(n15), .A2(taken[8]), .B1(n14), .B2(taken[9]), .ZN(n898)
         );
  NAND2_X1 U380 ( .A1(TAG_i[2]), .A2(TAG_i[3]), .ZN(n901) );
  AOI22_X1 U377 ( .A1(n21), .A2(taken[14]), .B1(n20), .B2(taken[15]), .ZN(n899) );
  AOI22_X1 U374 ( .A1(n19), .A2(taken[12]), .B1(n18), .B2(taken[13]), .ZN(n900) );
  AOI22_X1 U369 ( .A1(n9), .A2(taken[2]), .B1(n8), .B2(taken[3]), .ZN(n887) );
  AOI22_X1 U366 ( .A1(n7), .A2(taken[0]), .B1(n6), .B2(taken[1]), .ZN(n888) );
  NAND2_X1 U365 ( .A1(TAG_i[2]), .A2(n972), .ZN(n892) );
  AOI22_X1 U362 ( .A1(n13), .A2(taken[6]), .B1(n12), .B2(taken[7]), .ZN(n889)
         );
  AOI22_X1 U359 ( .A1(n11), .A2(taken[4]), .B1(n10), .B2(taken[5]), .ZN(n890)
         );
  AOI22_X1 U166 ( .A1(n7), .A2(\predict_PC[0][25] ), .B1(n572), .B2(
        \predict_PC[1][25] ), .ZN(n709) );
  AOI22_X1 U165 ( .A1(n9), .A2(\predict_PC[2][25] ), .B1(n570), .B2(
        \predict_PC[3][25] ), .ZN(n710) );
  AOI22_X1 U164 ( .A1(n11), .A2(\predict_PC[4][25] ), .B1(n568), .B2(
        \predict_PC[5][25] ), .ZN(n711) );
  AOI22_X1 U163 ( .A1(n13), .A2(\predict_PC[6][25] ), .B1(n566), .B2(
        \predict_PC[7][25] ), .ZN(n712) );
  NAND4_X1 U162 ( .A1(n709), .A2(n710), .A3(n711), .A4(n712), .ZN(n703) );
  AOI22_X1 U161 ( .A1(n15), .A2(\predict_PC[8][25] ), .B1(n560), .B2(
        \predict_PC[9][25] ), .ZN(n705) );
  AOI22_X1 U160 ( .A1(n17), .A2(\predict_PC[10][25] ), .B1(n558), .B2(
        \predict_PC[11][25] ), .ZN(n706) );
  AOI22_X1 U159 ( .A1(n19), .A2(\predict_PC[12][25] ), .B1(n556), .B2(
        \predict_PC[13][25] ), .ZN(n707) );
  AOI22_X1 U158 ( .A1(n21), .A2(\predict_PC[14][25] ), .B1(n554), .B2(
        \predict_PC[15][25] ), .ZN(n708) );
  NAND4_X1 U157 ( .A1(n705), .A2(n706), .A3(n707), .A4(n708), .ZN(n704) );
  AOI22_X1 U320 ( .A1(n7), .A2(\predict_PC[0][12] ), .B1(n6), .B2(
        \predict_PC[1][12] ), .ZN(n849) );
  AOI22_X1 U319 ( .A1(n9), .A2(\predict_PC[2][12] ), .B1(n8), .B2(
        \predict_PC[3][12] ), .ZN(n850) );
  AOI22_X1 U318 ( .A1(n11), .A2(\predict_PC[4][12] ), .B1(n10), .B2(
        \predict_PC[5][12] ), .ZN(n851) );
  AOI22_X1 U317 ( .A1(n13), .A2(\predict_PC[6][12] ), .B1(n12), .B2(
        \predict_PC[7][12] ), .ZN(n852) );
  NAND4_X1 U316 ( .A1(n849), .A2(n850), .A3(n851), .A4(n852), .ZN(n843) );
  AOI22_X1 U315 ( .A1(n15), .A2(\predict_PC[8][12] ), .B1(n14), .B2(
        \predict_PC[9][12] ), .ZN(n845) );
  AOI22_X1 U314 ( .A1(n17), .A2(\predict_PC[10][12] ), .B1(n16), .B2(
        \predict_PC[11][12] ), .ZN(n846) );
  AOI22_X1 U313 ( .A1(n19), .A2(\predict_PC[12][12] ), .B1(n18), .B2(
        \predict_PC[13][12] ), .ZN(n847) );
  AOI22_X1 U312 ( .A1(n21), .A2(\predict_PC[14][12] ), .B1(n20), .B2(
        \predict_PC[15][12] ), .ZN(n848) );
  NAND4_X1 U311 ( .A1(n845), .A2(n846), .A3(n847), .A4(n848), .ZN(n844) );
  AOI22_X1 U144 ( .A1(n7), .A2(\predict_PC[0][27] ), .B1(n572), .B2(
        \predict_PC[1][27] ), .ZN(n689) );
  AOI22_X1 U143 ( .A1(n9), .A2(\predict_PC[2][27] ), .B1(n570), .B2(
        \predict_PC[3][27] ), .ZN(n690) );
  AOI22_X1 U142 ( .A1(n11), .A2(\predict_PC[4][27] ), .B1(n10), .B2(
        \predict_PC[5][27] ), .ZN(n691) );
  AOI22_X1 U141 ( .A1(n13), .A2(\predict_PC[6][27] ), .B1(n12), .B2(
        \predict_PC[7][27] ), .ZN(n692) );
  NAND4_X1 U140 ( .A1(n689), .A2(n690), .A3(n691), .A4(n692), .ZN(n683) );
  AOI22_X1 U139 ( .A1(n15), .A2(\predict_PC[8][27] ), .B1(n560), .B2(
        \predict_PC[9][27] ), .ZN(n685) );
  AOI22_X1 U138 ( .A1(n17), .A2(\predict_PC[10][27] ), .B1(n558), .B2(
        \predict_PC[11][27] ), .ZN(n686) );
  AOI22_X1 U137 ( .A1(n19), .A2(\predict_PC[12][27] ), .B1(n556), .B2(
        \predict_PC[13][27] ), .ZN(n687) );
  AOI22_X1 U136 ( .A1(n21), .A2(\predict_PC[14][27] ), .B1(n20), .B2(
        \predict_PC[15][27] ), .ZN(n688) );
  NAND4_X1 U135 ( .A1(n685), .A2(n686), .A3(n687), .A4(n688), .ZN(n684) );
  AOI22_X1 U342 ( .A1(n7), .A2(\predict_PC[0][10] ), .B1(n6), .B2(
        \predict_PC[1][10] ), .ZN(n869) );
  AOI22_X1 U341 ( .A1(n9), .A2(\predict_PC[2][10] ), .B1(n8), .B2(
        \predict_PC[3][10] ), .ZN(n870) );
  AOI22_X1 U340 ( .A1(n11), .A2(\predict_PC[4][10] ), .B1(n10), .B2(
        \predict_PC[5][10] ), .ZN(n871) );
  AOI22_X1 U339 ( .A1(n13), .A2(\predict_PC[6][10] ), .B1(n12), .B2(
        \predict_PC[7][10] ), .ZN(n872) );
  NAND4_X1 U338 ( .A1(n869), .A2(n870), .A3(n871), .A4(n872), .ZN(n863) );
  AOI22_X1 U337 ( .A1(n15), .A2(\predict_PC[8][10] ), .B1(n14), .B2(
        \predict_PC[9][10] ), .ZN(n865) );
  AOI22_X1 U336 ( .A1(n17), .A2(\predict_PC[10][10] ), .B1(n16), .B2(
        \predict_PC[11][10] ), .ZN(n866) );
  AOI22_X1 U335 ( .A1(n19), .A2(\predict_PC[12][10] ), .B1(n18), .B2(
        \predict_PC[13][10] ), .ZN(n867) );
  AOI22_X1 U334 ( .A1(n21), .A2(\predict_PC[14][10] ), .B1(n20), .B2(
        \predict_PC[15][10] ), .ZN(n868) );
  NAND4_X1 U333 ( .A1(n865), .A2(n866), .A3(n867), .A4(n868), .ZN(n864) );
  AOI22_X1 U111 ( .A1(n7), .A2(\predict_PC[0][2] ), .B1(n6), .B2(
        \predict_PC[1][2] ), .ZN(n659) );
  AOI22_X1 U110 ( .A1(n9), .A2(\predict_PC[2][2] ), .B1(n8), .B2(
        \predict_PC[3][2] ), .ZN(n660) );
  AOI22_X1 U109 ( .A1(n11), .A2(\predict_PC[4][2] ), .B1(n10), .B2(
        \predict_PC[5][2] ), .ZN(n661) );
  AOI22_X1 U108 ( .A1(n13), .A2(\predict_PC[6][2] ), .B1(n12), .B2(
        \predict_PC[7][2] ), .ZN(n662) );
  NAND4_X1 U107 ( .A1(n659), .A2(n660), .A3(n661), .A4(n662), .ZN(n653) );
  AOI22_X1 U106 ( .A1(n15), .A2(\predict_PC[8][2] ), .B1(n14), .B2(
        \predict_PC[9][2] ), .ZN(n655) );
  AOI22_X1 U105 ( .A1(n17), .A2(\predict_PC[10][2] ), .B1(n16), .B2(
        \predict_PC[11][2] ), .ZN(n656) );
  AOI22_X1 U104 ( .A1(n19), .A2(\predict_PC[12][2] ), .B1(n18), .B2(
        \predict_PC[13][2] ), .ZN(n657) );
  AOI22_X1 U103 ( .A1(n21), .A2(\predict_PC[14][2] ), .B1(n20), .B2(
        \predict_PC[15][2] ), .ZN(n658) );
  NAND4_X1 U102 ( .A1(n655), .A2(n656), .A3(n657), .A4(n658), .ZN(n654) );
  AOI22_X1 U287 ( .A1(n7), .A2(\predict_PC[0][15] ), .B1(n6), .B2(
        \predict_PC[1][15] ), .ZN(n819) );
  AOI22_X1 U286 ( .A1(n9), .A2(\predict_PC[2][15] ), .B1(n8), .B2(
        \predict_PC[3][15] ), .ZN(n820) );
  AOI22_X1 U285 ( .A1(n11), .A2(\predict_PC[4][15] ), .B1(n10), .B2(
        \predict_PC[5][15] ), .ZN(n821) );
  AOI22_X1 U284 ( .A1(n13), .A2(\predict_PC[6][15] ), .B1(n12), .B2(
        \predict_PC[7][15] ), .ZN(n822) );
  NAND4_X1 U283 ( .A1(n819), .A2(n820), .A3(n821), .A4(n822), .ZN(n813) );
  AOI22_X1 U282 ( .A1(n15), .A2(\predict_PC[8][15] ), .B1(n14), .B2(
        \predict_PC[9][15] ), .ZN(n815) );
  AOI22_X1 U281 ( .A1(n17), .A2(\predict_PC[10][15] ), .B1(n16), .B2(
        \predict_PC[11][15] ), .ZN(n816) );
  AOI22_X1 U280 ( .A1(n19), .A2(\predict_PC[12][15] ), .B1(n18), .B2(
        \predict_PC[13][15] ), .ZN(n817) );
  AOI22_X1 U279 ( .A1(n21), .A2(\predict_PC[14][15] ), .B1(n20), .B2(
        \predict_PC[15][15] ), .ZN(n818) );
  NAND4_X1 U278 ( .A1(n815), .A2(n816), .A3(n817), .A4(n818), .ZN(n814) );
  AOI22_X1 U78 ( .A1(n571), .A2(\predict_PC[0][3] ), .B1(n6), .B2(
        \predict_PC[1][3] ), .ZN(n629) );
  AOI22_X1 U77 ( .A1(n569), .A2(\predict_PC[2][3] ), .B1(n8), .B2(
        \predict_PC[3][3] ), .ZN(n630) );
  AOI22_X1 U76 ( .A1(n11), .A2(\predict_PC[4][3] ), .B1(n10), .B2(
        \predict_PC[5][3] ), .ZN(n631) );
  AOI22_X1 U75 ( .A1(n565), .A2(\predict_PC[6][3] ), .B1(n12), .B2(
        \predict_PC[7][3] ), .ZN(n632) );
  NAND4_X1 U74 ( .A1(n629), .A2(n630), .A3(n631), .A4(n632), .ZN(n623) );
  AOI22_X1 U73 ( .A1(n559), .A2(\predict_PC[8][3] ), .B1(n14), .B2(
        \predict_PC[9][3] ), .ZN(n625) );
  AOI22_X1 U72 ( .A1(n557), .A2(\predict_PC[10][3] ), .B1(n16), .B2(
        \predict_PC[11][3] ), .ZN(n626) );
  AOI22_X1 U71 ( .A1(n555), .A2(\predict_PC[12][3] ), .B1(n18), .B2(
        \predict_PC[13][3] ), .ZN(n627) );
  AOI22_X1 U70 ( .A1(n553), .A2(\predict_PC[14][3] ), .B1(n20), .B2(
        \predict_PC[15][3] ), .ZN(n628) );
  NAND4_X1 U69 ( .A1(n625), .A2(n626), .A3(n627), .A4(n628), .ZN(n624) );
  AOI22_X1 U188 ( .A1(n7), .A2(\predict_PC[0][23] ), .B1(n6), .B2(
        \predict_PC[1][23] ), .ZN(n729) );
  AOI22_X1 U187 ( .A1(n9), .A2(\predict_PC[2][23] ), .B1(n8), .B2(
        \predict_PC[3][23] ), .ZN(n730) );
  AOI22_X1 U186 ( .A1(n567), .A2(\predict_PC[4][23] ), .B1(n10), .B2(
        \predict_PC[5][23] ), .ZN(n731) );
  AOI22_X1 U185 ( .A1(n565), .A2(\predict_PC[6][23] ), .B1(n12), .B2(
        \predict_PC[7][23] ), .ZN(n732) );
  NAND4_X1 U184 ( .A1(n729), .A2(n730), .A3(n731), .A4(n732), .ZN(n723) );
  AOI22_X1 U183 ( .A1(n15), .A2(\predict_PC[8][23] ), .B1(n14), .B2(
        \predict_PC[9][23] ), .ZN(n725) );
  AOI22_X1 U182 ( .A1(n17), .A2(\predict_PC[10][23] ), .B1(n16), .B2(
        \predict_PC[11][23] ), .ZN(n726) );
  AOI22_X1 U181 ( .A1(n19), .A2(\predict_PC[12][23] ), .B1(n18), .B2(
        \predict_PC[13][23] ), .ZN(n727) );
  AOI22_X1 U180 ( .A1(n553), .A2(\predict_PC[14][23] ), .B1(n20), .B2(
        \predict_PC[15][23] ), .ZN(n728) );
  NAND4_X1 U179 ( .A1(n725), .A2(n726), .A3(n727), .A4(n728), .ZN(n724) );
  AOI22_X1 U56 ( .A1(n571), .A2(\predict_PC[0][5] ), .B1(n6), .B2(
        \predict_PC[1][5] ), .ZN(n609) );
  AOI22_X1 U55 ( .A1(n569), .A2(\predict_PC[2][5] ), .B1(n8), .B2(
        \predict_PC[3][5] ), .ZN(n610) );
  AOI22_X1 U54 ( .A1(n11), .A2(\predict_PC[4][5] ), .B1(n10), .B2(
        \predict_PC[5][5] ), .ZN(n611) );
  AOI22_X1 U53 ( .A1(n13), .A2(\predict_PC[6][5] ), .B1(n12), .B2(
        \predict_PC[7][5] ), .ZN(n612) );
  NAND4_X1 U52 ( .A1(n609), .A2(n610), .A3(n611), .A4(n612), .ZN(n603) );
  AOI22_X1 U51 ( .A1(n559), .A2(\predict_PC[8][5] ), .B1(n14), .B2(
        \predict_PC[9][5] ), .ZN(n605) );
  AOI22_X1 U50 ( .A1(n557), .A2(\predict_PC[10][5] ), .B1(n16), .B2(
        \predict_PC[11][5] ), .ZN(n606) );
  AOI22_X1 U49 ( .A1(n555), .A2(\predict_PC[12][5] ), .B1(n18), .B2(
        \predict_PC[13][5] ), .ZN(n607) );
  AOI22_X1 U48 ( .A1(n21), .A2(\predict_PC[14][5] ), .B1(n20), .B2(
        \predict_PC[15][5] ), .ZN(n608) );
  NAND4_X1 U47 ( .A1(n605), .A2(n606), .A3(n607), .A4(n608), .ZN(n604) );
  AOI22_X1 U210 ( .A1(n571), .A2(\predict_PC[0][21] ), .B1(n6), .B2(
        \predict_PC[1][21] ), .ZN(n749) );
  AOI22_X1 U209 ( .A1(n569), .A2(\predict_PC[2][21] ), .B1(n8), .B2(
        \predict_PC[3][21] ), .ZN(n750) );
  AOI22_X1 U208 ( .A1(n567), .A2(\predict_PC[4][21] ), .B1(n10), .B2(
        \predict_PC[5][21] ), .ZN(n751) );
  AOI22_X1 U207 ( .A1(n565), .A2(\predict_PC[6][21] ), .B1(n12), .B2(
        \predict_PC[7][21] ), .ZN(n752) );
  NAND4_X1 U206 ( .A1(n749), .A2(n750), .A3(n751), .A4(n752), .ZN(n743) );
  AOI22_X1 U205 ( .A1(n559), .A2(\predict_PC[8][21] ), .B1(n14), .B2(
        \predict_PC[9][21] ), .ZN(n745) );
  AOI22_X1 U204 ( .A1(n557), .A2(\predict_PC[10][21] ), .B1(n16), .B2(
        \predict_PC[11][21] ), .ZN(n746) );
  AOI22_X1 U203 ( .A1(n555), .A2(\predict_PC[12][21] ), .B1(n18), .B2(
        \predict_PC[13][21] ), .ZN(n747) );
  AOI22_X1 U202 ( .A1(n553), .A2(\predict_PC[14][21] ), .B1(n20), .B2(
        \predict_PC[15][21] ), .ZN(n748) );
  NAND4_X1 U201 ( .A1(n745), .A2(n746), .A3(n747), .A4(n748), .ZN(n744) );
  AOI22_X1 U276 ( .A1(n7), .A2(\predict_PC[0][16] ), .B1(n6), .B2(
        \predict_PC[1][16] ), .ZN(n809) );
  AOI22_X1 U275 ( .A1(n9), .A2(\predict_PC[2][16] ), .B1(n8), .B2(
        \predict_PC[3][16] ), .ZN(n810) );
  AOI22_X1 U274 ( .A1(n11), .A2(\predict_PC[4][16] ), .B1(n10), .B2(
        \predict_PC[5][16] ), .ZN(n811) );
  AOI22_X1 U273 ( .A1(n13), .A2(\predict_PC[6][16] ), .B1(n12), .B2(
        \predict_PC[7][16] ), .ZN(n812) );
  NAND4_X1 U272 ( .A1(n809), .A2(n810), .A3(n811), .A4(n812), .ZN(n803) );
  AOI22_X1 U271 ( .A1(n15), .A2(\predict_PC[8][16] ), .B1(n14), .B2(
        \predict_PC[9][16] ), .ZN(n805) );
  AOI22_X1 U270 ( .A1(n17), .A2(\predict_PC[10][16] ), .B1(n16), .B2(
        \predict_PC[11][16] ), .ZN(n806) );
  AOI22_X1 U269 ( .A1(n19), .A2(\predict_PC[12][16] ), .B1(n18), .B2(
        \predict_PC[13][16] ), .ZN(n807) );
  AOI22_X1 U268 ( .A1(n21), .A2(\predict_PC[14][16] ), .B1(n20), .B2(
        \predict_PC[15][16] ), .ZN(n808) );
  NAND4_X1 U267 ( .A1(n805), .A2(n806), .A3(n807), .A4(n808), .ZN(n804) );
  AOI22_X1 U243 ( .A1(n7), .A2(\predict_PC[0][19] ), .B1(n572), .B2(
        \predict_PC[1][19] ), .ZN(n779) );
  AOI22_X1 U242 ( .A1(n9), .A2(\predict_PC[2][19] ), .B1(n570), .B2(
        \predict_PC[3][19] ), .ZN(n780) );
  AOI22_X1 U241 ( .A1(n11), .A2(\predict_PC[4][19] ), .B1(n568), .B2(
        \predict_PC[5][19] ), .ZN(n781) );
  AOI22_X1 U240 ( .A1(n13), .A2(\predict_PC[6][19] ), .B1(n566), .B2(
        \predict_PC[7][19] ), .ZN(n782) );
  NAND4_X1 U239 ( .A1(n779), .A2(n780), .A3(n781), .A4(n782), .ZN(n773) );
  AOI22_X1 U238 ( .A1(n15), .A2(\predict_PC[8][19] ), .B1(n560), .B2(
        \predict_PC[9][19] ), .ZN(n775) );
  AOI22_X1 U237 ( .A1(n17), .A2(\predict_PC[10][19] ), .B1(n558), .B2(
        \predict_PC[11][19] ), .ZN(n776) );
  AOI22_X1 U236 ( .A1(n19), .A2(\predict_PC[12][19] ), .B1(n556), .B2(
        \predict_PC[13][19] ), .ZN(n777) );
  AOI22_X1 U235 ( .A1(n21), .A2(\predict_PC[14][19] ), .B1(n554), .B2(
        \predict_PC[15][19] ), .ZN(n778) );
  NAND4_X1 U234 ( .A1(n775), .A2(n776), .A3(n777), .A4(n778), .ZN(n774) );
  AOI22_X1 U199 ( .A1(n571), .A2(\predict_PC[0][22] ), .B1(n6), .B2(
        \predict_PC[1][22] ), .ZN(n739) );
  AOI22_X1 U198 ( .A1(n569), .A2(\predict_PC[2][22] ), .B1(n8), .B2(
        \predict_PC[3][22] ), .ZN(n740) );
  AOI22_X1 U197 ( .A1(n567), .A2(\predict_PC[4][22] ), .B1(n10), .B2(
        \predict_PC[5][22] ), .ZN(n741) );
  AOI22_X1 U196 ( .A1(n565), .A2(\predict_PC[6][22] ), .B1(n12), .B2(
        \predict_PC[7][22] ), .ZN(n742) );
  NAND4_X1 U195 ( .A1(n739), .A2(n740), .A3(n741), .A4(n742), .ZN(n733) );
  AOI22_X1 U194 ( .A1(n559), .A2(\predict_PC[8][22] ), .B1(n14), .B2(
        \predict_PC[9][22] ), .ZN(n735) );
  AOI22_X1 U193 ( .A1(n557), .A2(\predict_PC[10][22] ), .B1(n16), .B2(
        \predict_PC[11][22] ), .ZN(n736) );
  AOI22_X1 U192 ( .A1(n555), .A2(\predict_PC[12][22] ), .B1(n18), .B2(
        \predict_PC[13][22] ), .ZN(n737) );
  AOI22_X1 U191 ( .A1(n553), .A2(\predict_PC[14][22] ), .B1(n20), .B2(
        \predict_PC[15][22] ), .ZN(n738) );
  NAND4_X1 U190 ( .A1(n735), .A2(n736), .A3(n737), .A4(n738), .ZN(n734) );
  AOI22_X1 U265 ( .A1(n571), .A2(\predict_PC[0][17] ), .B1(n6), .B2(
        \predict_PC[1][17] ), .ZN(n799) );
  AOI22_X1 U264 ( .A1(n569), .A2(\predict_PC[2][17] ), .B1(n8), .B2(
        \predict_PC[3][17] ), .ZN(n800) );
  AOI22_X1 U263 ( .A1(n567), .A2(\predict_PC[4][17] ), .B1(n10), .B2(
        \predict_PC[5][17] ), .ZN(n801) );
  AOI22_X1 U262 ( .A1(n565), .A2(\predict_PC[6][17] ), .B1(n12), .B2(
        \predict_PC[7][17] ), .ZN(n802) );
  NAND4_X1 U261 ( .A1(n799), .A2(n800), .A3(n801), .A4(n802), .ZN(n793) );
  AOI22_X1 U260 ( .A1(n559), .A2(\predict_PC[8][17] ), .B1(n14), .B2(
        \predict_PC[9][17] ), .ZN(n795) );
  AOI22_X1 U259 ( .A1(n557), .A2(\predict_PC[10][17] ), .B1(n16), .B2(
        \predict_PC[11][17] ), .ZN(n796) );
  AOI22_X1 U258 ( .A1(n555), .A2(\predict_PC[12][17] ), .B1(n18), .B2(
        \predict_PC[13][17] ), .ZN(n797) );
  AOI22_X1 U257 ( .A1(n553), .A2(\predict_PC[14][17] ), .B1(n20), .B2(
        \predict_PC[15][17] ), .ZN(n798) );
  NAND4_X1 U256 ( .A1(n795), .A2(n796), .A3(n797), .A4(n798), .ZN(n794) );
  AOI22_X1 U254 ( .A1(n7), .A2(\predict_PC[0][18] ), .B1(n572), .B2(
        \predict_PC[1][18] ), .ZN(n789) );
  AOI22_X1 U253 ( .A1(n9), .A2(\predict_PC[2][18] ), .B1(n570), .B2(
        \predict_PC[3][18] ), .ZN(n790) );
  AOI22_X1 U252 ( .A1(n11), .A2(\predict_PC[4][18] ), .B1(n568), .B2(
        \predict_PC[5][18] ), .ZN(n791) );
  AOI22_X1 U251 ( .A1(n13), .A2(\predict_PC[6][18] ), .B1(n566), .B2(
        \predict_PC[7][18] ), .ZN(n792) );
  NAND4_X1 U250 ( .A1(n789), .A2(n790), .A3(n791), .A4(n792), .ZN(n783) );
  AOI22_X1 U249 ( .A1(n15), .A2(\predict_PC[8][18] ), .B1(n560), .B2(
        \predict_PC[9][18] ), .ZN(n785) );
  AOI22_X1 U248 ( .A1(n17), .A2(\predict_PC[10][18] ), .B1(n558), .B2(
        \predict_PC[11][18] ), .ZN(n786) );
  AOI22_X1 U247 ( .A1(n19), .A2(\predict_PC[12][18] ), .B1(n556), .B2(
        \predict_PC[13][18] ), .ZN(n787) );
  AOI22_X1 U246 ( .A1(n21), .A2(\predict_PC[14][18] ), .B1(n554), .B2(
        \predict_PC[15][18] ), .ZN(n788) );
  NAND4_X1 U245 ( .A1(n785), .A2(n786), .A3(n787), .A4(n788), .ZN(n784) );
  AOI22_X1 U331 ( .A1(n7), .A2(\predict_PC[0][11] ), .B1(n6), .B2(
        \predict_PC[1][11] ), .ZN(n859) );
  AOI22_X1 U330 ( .A1(n9), .A2(\predict_PC[2][11] ), .B1(n8), .B2(
        \predict_PC[3][11] ), .ZN(n860) );
  AOI22_X1 U329 ( .A1(n11), .A2(\predict_PC[4][11] ), .B1(n10), .B2(
        \predict_PC[5][11] ), .ZN(n861) );
  AOI22_X1 U328 ( .A1(n13), .A2(\predict_PC[6][11] ), .B1(n12), .B2(
        \predict_PC[7][11] ), .ZN(n862) );
  NAND4_X1 U327 ( .A1(n859), .A2(n860), .A3(n861), .A4(n862), .ZN(n853) );
  AOI22_X1 U326 ( .A1(n15), .A2(\predict_PC[8][11] ), .B1(n14), .B2(
        \predict_PC[9][11] ), .ZN(n855) );
  AOI22_X1 U325 ( .A1(n17), .A2(\predict_PC[10][11] ), .B1(n16), .B2(
        \predict_PC[11][11] ), .ZN(n856) );
  AOI22_X1 U324 ( .A1(n19), .A2(\predict_PC[12][11] ), .B1(n18), .B2(
        \predict_PC[13][11] ), .ZN(n857) );
  AOI22_X1 U323 ( .A1(n21), .A2(\predict_PC[14][11] ), .B1(n20), .B2(
        \predict_PC[15][11] ), .ZN(n858) );
  NAND4_X1 U322 ( .A1(n855), .A2(n856), .A3(n857), .A4(n858), .ZN(n854) );
  AOI22_X1 U122 ( .A1(n7), .A2(\predict_PC[0][29] ), .B1(n6), .B2(
        \predict_PC[1][29] ), .ZN(n669) );
  AOI22_X1 U121 ( .A1(n9), .A2(\predict_PC[2][29] ), .B1(n8), .B2(
        \predict_PC[3][29] ), .ZN(n670) );
  AOI22_X1 U120 ( .A1(n11), .A2(\predict_PC[4][29] ), .B1(n10), .B2(
        \predict_PC[5][29] ), .ZN(n671) );
  AOI22_X1 U119 ( .A1(n13), .A2(\predict_PC[6][29] ), .B1(n12), .B2(
        \predict_PC[7][29] ), .ZN(n672) );
  NAND4_X1 U118 ( .A1(n669), .A2(n670), .A3(n671), .A4(n672), .ZN(n663) );
  AOI22_X1 U117 ( .A1(n15), .A2(\predict_PC[8][29] ), .B1(n14), .B2(
        \predict_PC[9][29] ), .ZN(n665) );
  AOI22_X1 U116 ( .A1(n17), .A2(\predict_PC[10][29] ), .B1(n16), .B2(
        \predict_PC[11][29] ), .ZN(n666) );
  AOI22_X1 U115 ( .A1(n19), .A2(\predict_PC[12][29] ), .B1(n18), .B2(
        \predict_PC[13][29] ), .ZN(n667) );
  AOI22_X1 U114 ( .A1(n21), .A2(\predict_PC[14][29] ), .B1(n20), .B2(
        \predict_PC[15][29] ), .ZN(n668) );
  NAND4_X1 U113 ( .A1(n665), .A2(n666), .A3(n667), .A4(n668), .ZN(n664) );
  AOI22_X1 U309 ( .A1(n7), .A2(\predict_PC[0][13] ), .B1(n6), .B2(
        \predict_PC[1][13] ), .ZN(n839) );
  AOI22_X1 U308 ( .A1(n9), .A2(\predict_PC[2][13] ), .B1(n8), .B2(
        \predict_PC[3][13] ), .ZN(n840) );
  AOI22_X1 U307 ( .A1(n11), .A2(\predict_PC[4][13] ), .B1(n10), .B2(
        \predict_PC[5][13] ), .ZN(n841) );
  AOI22_X1 U306 ( .A1(n13), .A2(\predict_PC[6][13] ), .B1(n12), .B2(
        \predict_PC[7][13] ), .ZN(n842) );
  NAND4_X1 U305 ( .A1(n839), .A2(n840), .A3(n841), .A4(n842), .ZN(n833) );
  AOI22_X1 U304 ( .A1(n15), .A2(\predict_PC[8][13] ), .B1(n14), .B2(
        \predict_PC[9][13] ), .ZN(n835) );
  AOI22_X1 U303 ( .A1(n17), .A2(\predict_PC[10][13] ), .B1(n16), .B2(
        \predict_PC[11][13] ), .ZN(n836) );
  AOI22_X1 U302 ( .A1(n19), .A2(\predict_PC[12][13] ), .B1(n18), .B2(
        \predict_PC[13][13] ), .ZN(n837) );
  AOI22_X1 U301 ( .A1(n21), .A2(\predict_PC[14][13] ), .B1(n20), .B2(
        \predict_PC[15][13] ), .ZN(n838) );
  NAND4_X1 U300 ( .A1(n835), .A2(n836), .A3(n837), .A4(n838), .ZN(n834) );
  AOI22_X1 U298 ( .A1(n7), .A2(\predict_PC[0][14] ), .B1(n6), .B2(
        \predict_PC[1][14] ), .ZN(n829) );
  AOI22_X1 U297 ( .A1(n9), .A2(\predict_PC[2][14] ), .B1(n8), .B2(
        \predict_PC[3][14] ), .ZN(n830) );
  AOI22_X1 U296 ( .A1(n11), .A2(\predict_PC[4][14] ), .B1(n10), .B2(
        \predict_PC[5][14] ), .ZN(n831) );
  AOI22_X1 U295 ( .A1(n13), .A2(\predict_PC[6][14] ), .B1(n12), .B2(
        \predict_PC[7][14] ), .ZN(n832) );
  NAND4_X1 U294 ( .A1(n829), .A2(n830), .A3(n831), .A4(n832), .ZN(n823) );
  AOI22_X1 U293 ( .A1(n15), .A2(\predict_PC[8][14] ), .B1(n14), .B2(
        \predict_PC[9][14] ), .ZN(n825) );
  AOI22_X1 U292 ( .A1(n17), .A2(\predict_PC[10][14] ), .B1(n16), .B2(
        \predict_PC[11][14] ), .ZN(n826) );
  AOI22_X1 U291 ( .A1(n19), .A2(\predict_PC[12][14] ), .B1(n18), .B2(
        \predict_PC[13][14] ), .ZN(n827) );
  AOI22_X1 U290 ( .A1(n21), .A2(\predict_PC[14][14] ), .B1(n20), .B2(
        \predict_PC[15][14] ), .ZN(n828) );
  NAND4_X1 U289 ( .A1(n825), .A2(n826), .A3(n827), .A4(n828), .ZN(n824) );
  AOI22_X1 U221 ( .A1(n7), .A2(\predict_PC[0][20] ), .B1(n572), .B2(
        \predict_PC[1][20] ), .ZN(n759) );
  AOI22_X1 U220 ( .A1(n9), .A2(\predict_PC[2][20] ), .B1(n570), .B2(
        \predict_PC[3][20] ), .ZN(n760) );
  AOI22_X1 U219 ( .A1(n11), .A2(\predict_PC[4][20] ), .B1(n568), .B2(
        \predict_PC[5][20] ), .ZN(n761) );
  AOI22_X1 U218 ( .A1(n13), .A2(\predict_PC[6][20] ), .B1(n566), .B2(
        \predict_PC[7][20] ), .ZN(n762) );
  NAND4_X1 U217 ( .A1(n759), .A2(n760), .A3(n761), .A4(n762), .ZN(n753) );
  AOI22_X1 U216 ( .A1(n15), .A2(\predict_PC[8][20] ), .B1(n560), .B2(
        \predict_PC[9][20] ), .ZN(n755) );
  AOI22_X1 U215 ( .A1(n17), .A2(\predict_PC[10][20] ), .B1(n558), .B2(
        \predict_PC[11][20] ), .ZN(n756) );
  AOI22_X1 U214 ( .A1(n19), .A2(\predict_PC[12][20] ), .B1(n556), .B2(
        \predict_PC[13][20] ), .ZN(n757) );
  AOI22_X1 U213 ( .A1(n21), .A2(\predict_PC[14][20] ), .B1(n554), .B2(
        \predict_PC[15][20] ), .ZN(n758) );
  NAND4_X1 U212 ( .A1(n755), .A2(n756), .A3(n757), .A4(n758), .ZN(n754) );
  AOI22_X1 U177 ( .A1(n7), .A2(\predict_PC[0][24] ), .B1(n572), .B2(
        \predict_PC[1][24] ), .ZN(n719) );
  AOI22_X1 U176 ( .A1(n9), .A2(\predict_PC[2][24] ), .B1(n570), .B2(
        \predict_PC[3][24] ), .ZN(n720) );
  AOI22_X1 U175 ( .A1(n11), .A2(\predict_PC[4][24] ), .B1(n568), .B2(
        \predict_PC[5][24] ), .ZN(n721) );
  AOI22_X1 U174 ( .A1(n13), .A2(\predict_PC[6][24] ), .B1(n566), .B2(
        \predict_PC[7][24] ), .ZN(n722) );
  NAND4_X1 U173 ( .A1(n719), .A2(n720), .A3(n721), .A4(n722), .ZN(n713) );
  AOI22_X1 U172 ( .A1(n15), .A2(\predict_PC[8][24] ), .B1(n560), .B2(
        \predict_PC[9][24] ), .ZN(n715) );
  AOI22_X1 U171 ( .A1(n17), .A2(\predict_PC[10][24] ), .B1(n558), .B2(
        \predict_PC[11][24] ), .ZN(n716) );
  AOI22_X1 U170 ( .A1(n19), .A2(\predict_PC[12][24] ), .B1(n556), .B2(
        \predict_PC[13][24] ), .ZN(n717) );
  AOI22_X1 U169 ( .A1(n21), .A2(\predict_PC[14][24] ), .B1(n554), .B2(
        \predict_PC[15][24] ), .ZN(n718) );
  NAND4_X1 U168 ( .A1(n715), .A2(n716), .A3(n717), .A4(n718), .ZN(n714) );
  AOI22_X1 U133 ( .A1(n7), .A2(\predict_PC[0][28] ), .B1(n6), .B2(
        \predict_PC[1][28] ), .ZN(n679) );
  AOI22_X1 U132 ( .A1(n9), .A2(\predict_PC[2][28] ), .B1(n8), .B2(
        \predict_PC[3][28] ), .ZN(n680) );
  AOI22_X1 U131 ( .A1(n11), .A2(\predict_PC[4][28] ), .B1(n568), .B2(
        \predict_PC[5][28] ), .ZN(n681) );
  AOI22_X1 U130 ( .A1(n13), .A2(\predict_PC[6][28] ), .B1(n566), .B2(
        \predict_PC[7][28] ), .ZN(n682) );
  NAND4_X1 U129 ( .A1(n679), .A2(n680), .A3(n681), .A4(n682), .ZN(n673) );
  AOI22_X1 U128 ( .A1(n15), .A2(\predict_PC[8][28] ), .B1(n14), .B2(
        \predict_PC[9][28] ), .ZN(n675) );
  AOI22_X1 U127 ( .A1(n17), .A2(\predict_PC[10][28] ), .B1(n16), .B2(
        \predict_PC[11][28] ), .ZN(n676) );
  AOI22_X1 U126 ( .A1(n19), .A2(\predict_PC[12][28] ), .B1(n18), .B2(
        \predict_PC[13][28] ), .ZN(n677) );
  AOI22_X1 U125 ( .A1(n21), .A2(\predict_PC[14][28] ), .B1(n554), .B2(
        \predict_PC[15][28] ), .ZN(n678) );
  NAND4_X1 U124 ( .A1(n675), .A2(n676), .A3(n677), .A4(n678), .ZN(n674) );
  AOI22_X1 U155 ( .A1(n7), .A2(\predict_PC[0][26] ), .B1(n572), .B2(
        \predict_PC[1][26] ), .ZN(n699) );
  AOI22_X1 U154 ( .A1(n9), .A2(\predict_PC[2][26] ), .B1(n570), .B2(
        \predict_PC[3][26] ), .ZN(n700) );
  AOI22_X1 U153 ( .A1(n11), .A2(\predict_PC[4][26] ), .B1(n568), .B2(
        \predict_PC[5][26] ), .ZN(n701) );
  AOI22_X1 U152 ( .A1(n13), .A2(\predict_PC[6][26] ), .B1(n566), .B2(
        \predict_PC[7][26] ), .ZN(n702) );
  NAND4_X1 U151 ( .A1(n699), .A2(n700), .A3(n701), .A4(n702), .ZN(n693) );
  AOI22_X1 U150 ( .A1(n15), .A2(\predict_PC[8][26] ), .B1(n560), .B2(
        \predict_PC[9][26] ), .ZN(n695) );
  AOI22_X1 U149 ( .A1(n17), .A2(\predict_PC[10][26] ), .B1(n558), .B2(
        \predict_PC[11][26] ), .ZN(n696) );
  AOI22_X1 U148 ( .A1(n19), .A2(\predict_PC[12][26] ), .B1(n556), .B2(
        \predict_PC[13][26] ), .ZN(n697) );
  AOI22_X1 U147 ( .A1(n21), .A2(\predict_PC[14][26] ), .B1(n554), .B2(
        \predict_PC[15][26] ), .ZN(n698) );
  NAND4_X1 U146 ( .A1(n695), .A2(n696), .A3(n697), .A4(n698), .ZN(n694) );
  AOI22_X1 U353 ( .A1(n7), .A2(\predict_PC[0][0] ), .B1(n6), .B2(
        \predict_PC[1][0] ), .ZN(n879) );
  AOI22_X1 U352 ( .A1(n9), .A2(\predict_PC[2][0] ), .B1(n8), .B2(
        \predict_PC[3][0] ), .ZN(n880) );
  AOI22_X1 U351 ( .A1(n11), .A2(\predict_PC[4][0] ), .B1(n10), .B2(
        \predict_PC[5][0] ), .ZN(n881) );
  AOI22_X1 U350 ( .A1(n13), .A2(\predict_PC[6][0] ), .B1(n12), .B2(
        \predict_PC[7][0] ), .ZN(n882) );
  NAND4_X1 U349 ( .A1(n879), .A2(n880), .A3(n881), .A4(n882), .ZN(n873) );
  AOI22_X1 U348 ( .A1(n15), .A2(\predict_PC[8][0] ), .B1(n14), .B2(
        \predict_PC[9][0] ), .ZN(n875) );
  AOI22_X1 U347 ( .A1(n17), .A2(\predict_PC[10][0] ), .B1(n16), .B2(
        \predict_PC[11][0] ), .ZN(n876) );
  AOI22_X1 U346 ( .A1(n19), .A2(\predict_PC[12][0] ), .B1(n18), .B2(
        \predict_PC[13][0] ), .ZN(n877) );
  AOI22_X1 U345 ( .A1(n21), .A2(\predict_PC[14][0] ), .B1(n20), .B2(
        \predict_PC[15][0] ), .ZN(n878) );
  NAND4_X1 U344 ( .A1(n875), .A2(n876), .A3(n877), .A4(n878), .ZN(n874) );
  AOI22_X1 U232 ( .A1(n571), .A2(\predict_PC[0][1] ), .B1(n6), .B2(
        \predict_PC[1][1] ), .ZN(n769) );
  AOI22_X1 U231 ( .A1(n569), .A2(\predict_PC[2][1] ), .B1(n8), .B2(
        \predict_PC[3][1] ), .ZN(n770) );
  AOI22_X1 U230 ( .A1(n11), .A2(\predict_PC[4][1] ), .B1(n10), .B2(
        \predict_PC[5][1] ), .ZN(n771) );
  AOI22_X1 U229 ( .A1(n13), .A2(\predict_PC[6][1] ), .B1(n12), .B2(
        \predict_PC[7][1] ), .ZN(n772) );
  NAND4_X1 U228 ( .A1(n769), .A2(n770), .A3(n771), .A4(n772), .ZN(n763) );
  AOI22_X1 U227 ( .A1(n559), .A2(\predict_PC[8][1] ), .B1(n14), .B2(
        \predict_PC[9][1] ), .ZN(n765) );
  AOI22_X1 U226 ( .A1(n17), .A2(\predict_PC[10][1] ), .B1(n16), .B2(
        \predict_PC[11][1] ), .ZN(n766) );
  AOI22_X1 U225 ( .A1(n555), .A2(\predict_PC[12][1] ), .B1(n18), .B2(
        \predict_PC[13][1] ), .ZN(n767) );
  AOI22_X1 U224 ( .A1(n21), .A2(\predict_PC[14][1] ), .B1(n20), .B2(
        \predict_PC[15][1] ), .ZN(n768) );
  NAND4_X1 U223 ( .A1(n765), .A2(n766), .A3(n767), .A4(n768), .ZN(n764) );
  AOI22_X1 U100 ( .A1(n7), .A2(\predict_PC[0][30] ), .B1(n6), .B2(
        \predict_PC[1][30] ), .ZN(n649) );
  AOI22_X1 U99 ( .A1(n9), .A2(\predict_PC[2][30] ), .B1(n8), .B2(
        \predict_PC[3][30] ), .ZN(n650) );
  AOI22_X1 U98 ( .A1(n567), .A2(\predict_PC[4][30] ), .B1(n10), .B2(
        \predict_PC[5][30] ), .ZN(n651) );
  AOI22_X1 U97 ( .A1(n565), .A2(\predict_PC[6][30] ), .B1(n12), .B2(
        \predict_PC[7][30] ), .ZN(n652) );
  NAND4_X1 U96 ( .A1(n649), .A2(n650), .A3(n651), .A4(n652), .ZN(n643) );
  AOI22_X1 U95 ( .A1(n15), .A2(\predict_PC[8][30] ), .B1(n14), .B2(
        \predict_PC[9][30] ), .ZN(n645) );
  AOI22_X1 U94 ( .A1(n557), .A2(\predict_PC[10][30] ), .B1(n16), .B2(
        \predict_PC[11][30] ), .ZN(n646) );
  AOI22_X1 U93 ( .A1(n19), .A2(\predict_PC[12][30] ), .B1(n18), .B2(
        \predict_PC[13][30] ), .ZN(n647) );
  AOI22_X1 U92 ( .A1(n553), .A2(\predict_PC[14][30] ), .B1(n20), .B2(
        \predict_PC[15][30] ), .ZN(n648) );
  NAND4_X1 U91 ( .A1(n645), .A2(n646), .A3(n647), .A4(n648), .ZN(n644) );
  AOI22_X1 U23 ( .A1(n7), .A2(\predict_PC[0][8] ), .B1(n6), .B2(
        \predict_PC[1][8] ), .ZN(n579) );
  AOI22_X1 U22 ( .A1(n9), .A2(\predict_PC[2][8] ), .B1(n8), .B2(
        \predict_PC[3][8] ), .ZN(n580) );
  AOI22_X1 U21 ( .A1(n11), .A2(\predict_PC[4][8] ), .B1(n10), .B2(
        \predict_PC[5][8] ), .ZN(n581) );
  AOI22_X1 U20 ( .A1(n13), .A2(\predict_PC[6][8] ), .B1(n12), .B2(
        \predict_PC[7][8] ), .ZN(n582) );
  NAND4_X1 U19 ( .A1(n579), .A2(n580), .A3(n581), .A4(n582), .ZN(n573) );
  AOI22_X1 U18 ( .A1(n15), .A2(\predict_PC[8][8] ), .B1(n14), .B2(
        \predict_PC[9][8] ), .ZN(n575) );
  AOI22_X1 U17 ( .A1(n17), .A2(\predict_PC[10][8] ), .B1(n16), .B2(
        \predict_PC[11][8] ), .ZN(n576) );
  AOI22_X1 U16 ( .A1(n19), .A2(\predict_PC[12][8] ), .B1(n18), .B2(
        \predict_PC[13][8] ), .ZN(n577) );
  AOI22_X1 U15 ( .A1(n21), .A2(\predict_PC[14][8] ), .B1(n20), .B2(
        \predict_PC[15][8] ), .ZN(n578) );
  NAND4_X1 U14 ( .A1(n575), .A2(n576), .A3(n577), .A4(n578), .ZN(n574) );
  AOI22_X1 U89 ( .A1(n7), .A2(\predict_PC[0][31] ), .B1(n6), .B2(
        \predict_PC[1][31] ), .ZN(n639) );
  AOI22_X1 U88 ( .A1(n9), .A2(\predict_PC[2][31] ), .B1(n8), .B2(
        \predict_PC[3][31] ), .ZN(n640) );
  AOI22_X1 U87 ( .A1(n11), .A2(\predict_PC[4][31] ), .B1(n10), .B2(
        \predict_PC[5][31] ), .ZN(n641) );
  AOI22_X1 U86 ( .A1(n13), .A2(\predict_PC[6][31] ), .B1(n12), .B2(
        \predict_PC[7][31] ), .ZN(n642) );
  NAND4_X1 U85 ( .A1(n639), .A2(n640), .A3(n641), .A4(n642), .ZN(n633) );
  AOI22_X1 U84 ( .A1(n15), .A2(\predict_PC[8][31] ), .B1(n14), .B2(
        \predict_PC[9][31] ), .ZN(n635) );
  AOI22_X1 U83 ( .A1(n17), .A2(\predict_PC[10][31] ), .B1(n16), .B2(
        \predict_PC[11][31] ), .ZN(n636) );
  AOI22_X1 U82 ( .A1(n19), .A2(\predict_PC[12][31] ), .B1(n18), .B2(
        \predict_PC[13][31] ), .ZN(n637) );
  AOI22_X1 U81 ( .A1(n21), .A2(\predict_PC[14][31] ), .B1(n20), .B2(
        \predict_PC[15][31] ), .ZN(n638) );
  NAND4_X1 U80 ( .A1(n635), .A2(n636), .A3(n637), .A4(n638), .ZN(n634) );
  AOI22_X1 U34 ( .A1(n7), .A2(\predict_PC[0][7] ), .B1(n6), .B2(
        \predict_PC[1][7] ), .ZN(n589) );
  AOI22_X1 U33 ( .A1(n9), .A2(\predict_PC[2][7] ), .B1(n8), .B2(
        \predict_PC[3][7] ), .ZN(n590) );
  AOI22_X1 U32 ( .A1(n11), .A2(\predict_PC[4][7] ), .B1(n10), .B2(
        \predict_PC[5][7] ), .ZN(n591) );
  AOI22_X1 U31 ( .A1(n13), .A2(\predict_PC[6][7] ), .B1(n12), .B2(
        \predict_PC[7][7] ), .ZN(n592) );
  NAND4_X1 U30 ( .A1(n589), .A2(n590), .A3(n591), .A4(n592), .ZN(n583) );
  AOI22_X1 U29 ( .A1(n15), .A2(\predict_PC[8][7] ), .B1(n14), .B2(
        \predict_PC[9][7] ), .ZN(n585) );
  AOI22_X1 U28 ( .A1(n17), .A2(\predict_PC[10][7] ), .B1(n16), .B2(
        \predict_PC[11][7] ), .ZN(n586) );
  AOI22_X1 U27 ( .A1(n19), .A2(\predict_PC[12][7] ), .B1(n18), .B2(
        \predict_PC[13][7] ), .ZN(n587) );
  AOI22_X1 U26 ( .A1(n21), .A2(\predict_PC[14][7] ), .B1(n20), .B2(
        \predict_PC[15][7] ), .ZN(n588) );
  NAND4_X1 U25 ( .A1(n585), .A2(n586), .A3(n587), .A4(n588), .ZN(n584) );
  AOI22_X1 U45 ( .A1(n7), .A2(\predict_PC[0][6] ), .B1(n6), .B2(
        \predict_PC[1][6] ), .ZN(n599) );
  AOI22_X1 U44 ( .A1(n9), .A2(\predict_PC[2][6] ), .B1(n8), .B2(
        \predict_PC[3][6] ), .ZN(n600) );
  AOI22_X1 U43 ( .A1(n11), .A2(\predict_PC[4][6] ), .B1(n10), .B2(
        \predict_PC[5][6] ), .ZN(n601) );
  AOI22_X1 U42 ( .A1(n13), .A2(\predict_PC[6][6] ), .B1(n12), .B2(
        \predict_PC[7][6] ), .ZN(n602) );
  NAND4_X1 U41 ( .A1(n599), .A2(n600), .A3(n601), .A4(n602), .ZN(n593) );
  AOI22_X1 U40 ( .A1(n15), .A2(\predict_PC[8][6] ), .B1(n14), .B2(
        \predict_PC[9][6] ), .ZN(n595) );
  AOI22_X1 U39 ( .A1(n17), .A2(\predict_PC[10][6] ), .B1(n16), .B2(
        \predict_PC[11][6] ), .ZN(n596) );
  AOI22_X1 U38 ( .A1(n19), .A2(\predict_PC[12][6] ), .B1(n18), .B2(
        \predict_PC[13][6] ), .ZN(n597) );
  AOI22_X1 U37 ( .A1(n21), .A2(\predict_PC[14][6] ), .B1(n20), .B2(
        \predict_PC[15][6] ), .ZN(n598) );
  NAND4_X1 U36 ( .A1(n595), .A2(n596), .A3(n597), .A4(n598), .ZN(n594) );
  AOI22_X1 U12 ( .A1(n7), .A2(\predict_PC[0][9] ), .B1(n6), .B2(
        \predict_PC[1][9] ), .ZN(n561) );
  AOI22_X1 U11 ( .A1(n9), .A2(\predict_PC[2][9] ), .B1(n8), .B2(
        \predict_PC[3][9] ), .ZN(n562) );
  AOI22_X1 U10 ( .A1(n11), .A2(\predict_PC[4][9] ), .B1(n10), .B2(
        \predict_PC[5][9] ), .ZN(n563) );
  AOI22_X1 U9 ( .A1(n13), .A2(\predict_PC[6][9] ), .B1(n12), .B2(
        \predict_PC[7][9] ), .ZN(n564) );
  NAND4_X1 U8 ( .A1(n561), .A2(n562), .A3(n563), .A4(n564), .ZN(n547) );
  AOI22_X1 U7 ( .A1(n15), .A2(\predict_PC[8][9] ), .B1(n14), .B2(
        \predict_PC[9][9] ), .ZN(n549) );
  AOI22_X1 U6 ( .A1(n17), .A2(\predict_PC[10][9] ), .B1(n16), .B2(
        \predict_PC[11][9] ), .ZN(n550) );
  AOI22_X1 U5 ( .A1(n19), .A2(\predict_PC[12][9] ), .B1(n18), .B2(
        \predict_PC[13][9] ), .ZN(n551) );
  AOI22_X1 U4 ( .A1(n21), .A2(\predict_PC[14][9] ), .B1(n20), .B2(
        \predict_PC[15][9] ), .ZN(n552) );
  NAND4_X1 U3 ( .A1(n549), .A2(n550), .A3(n551), .A4(n552), .ZN(n548) );
  AOI22_X1 U67 ( .A1(n7), .A2(\predict_PC[0][4] ), .B1(n6), .B2(
        \predict_PC[1][4] ), .ZN(n619) );
  AOI22_X1 U66 ( .A1(n9), .A2(\predict_PC[2][4] ), .B1(n8), .B2(
        \predict_PC[3][4] ), .ZN(n620) );
  AOI22_X1 U65 ( .A1(n567), .A2(\predict_PC[4][4] ), .B1(n10), .B2(
        \predict_PC[5][4] ), .ZN(n621) );
  AOI22_X1 U64 ( .A1(n13), .A2(\predict_PC[6][4] ), .B1(n12), .B2(
        \predict_PC[7][4] ), .ZN(n622) );
  NAND4_X1 U63 ( .A1(n619), .A2(n620), .A3(n621), .A4(n622), .ZN(n613) );
  AOI22_X1 U62 ( .A1(n15), .A2(\predict_PC[8][4] ), .B1(n14), .B2(
        \predict_PC[9][4] ), .ZN(n615) );
  AOI22_X1 U61 ( .A1(n17), .A2(\predict_PC[10][4] ), .B1(n16), .B2(
        \predict_PC[11][4] ), .ZN(n616) );
  AOI22_X1 U60 ( .A1(n19), .A2(\predict_PC[12][4] ), .B1(n18), .B2(
        \predict_PC[13][4] ), .ZN(n617) );
  AOI22_X1 U59 ( .A1(n21), .A2(\predict_PC[14][4] ), .B1(n20), .B2(
        \predict_PC[15][4] ), .ZN(n618) );
  NAND4_X1 U58 ( .A1(n615), .A2(n616), .A3(n617), .A4(n618), .ZN(n614) );
  NAND2_X1 U469 ( .A1(n979), .A2(n978), .ZN(n945) );
  NOR2_X1 U450 ( .A1(n945), .A2(n947), .ZN(N38) );
  NAND2_X1 U456 ( .A1(n977), .A2(n2), .ZN(n946) );
  NOR2_X1 U447 ( .A1(n948), .A2(n946), .ZN(N43) );
  NOR2_X1 U449 ( .A1(n948), .A2(n947), .ZN(N39) );
  NAND2_X1 U477 ( .A1(n978), .A2(n3), .ZN(n949) );
  NOR2_X1 U448 ( .A1(n949), .A2(n947), .ZN(N40) );
  NAND2_X1 U466 ( .A1(n3), .A2(n1), .ZN(n944) );
  NOR2_X1 U445 ( .A1(n944), .A2(n947), .ZN(N41) );
  NOR2_X1 U444 ( .A1(n945), .A2(n946), .ZN(N42) );
  NAND2_X1 U465 ( .A1(n976), .A2(n4), .ZN(n951) );
  NOR2_X1 U464 ( .A1(n944), .A2(n951), .ZN(N49) );
  NOR2_X1 U453 ( .A1(n949), .A2(n946), .ZN(N44) );
  NOR2_X1 U455 ( .A1(n944), .A2(n946), .ZN(N45) );
  NOR2_X1 U458 ( .A1(n945), .A2(n951), .ZN(N46) );
  NOR2_X1 U460 ( .A1(n948), .A2(n951), .ZN(N47) );
  NOR2_X1 U462 ( .A1(n949), .A2(n951), .ZN(N48) );
  NAND2_X1 U479 ( .A1(n4), .A2(n2), .ZN(n943) );
  NOR2_X1 U471 ( .A1(n943), .A2(n948), .ZN(N51) );
  NOR2_X1 U468 ( .A1(n943), .A2(n945), .ZN(N50) );
  NOR2_X1 U440 ( .A1(n943), .A2(n944), .ZN(N53) );
  NOR2_X1 U476 ( .A1(n943), .A2(n949), .ZN(N52) );
  NOR2_X1 U355 ( .A1(stall_i), .A2(reset), .ZN(n884) );
  OAI22_X1 U354 ( .A1(stall_i), .A2(n883), .B1(n884), .B2(n975), .ZN(n955) );
  INV_X1 U392 ( .A(TAG_i[0]), .ZN(n903) );
  NAND2_X1 U451 ( .A1(n977), .A2(n976), .ZN(n947) );
  NAND2_X1 U472 ( .A1(n979), .A2(n1), .ZN(n948) );
  INV_X1 U394 ( .A(TAG_i[2]), .ZN(n973) );
  INV_X1 U393 ( .A(TAG_i[1]), .ZN(n974) );
  NAND2_X1 U385 ( .A1(n903), .A2(n974), .ZN(n893) );
  INV_X1 U395 ( .A(TAG_i[3]), .ZN(n972) );
  NAND2_X1 U372 ( .A1(n973), .A2(n972), .ZN(n896) );
  AOI21_X1 U357 ( .B1(n885), .B2(n886), .A(reset), .ZN(taken_o) );
  NOR4_X1 U398 ( .A1(n907), .A2(n908), .A3(n909), .A4(n910), .ZN(n905) );
  AOI21_X1 U396 ( .B1(n5), .B2(n905), .A(n906), .ZN(mispredict_o) );
  AND4_X1 U373 ( .A1(n897), .A2(n898), .A3(n899), .A4(n900), .ZN(n885) );
  AND4_X1 U358 ( .A1(n887), .A2(n888), .A3(n889), .A4(n890), .ZN(n886) );
  OR2_X1 U156 ( .A1(n703), .A2(n704), .ZN(predicted_next_PC_o[25]) );
  OR2_X1 U310 ( .A1(n843), .A2(n844), .ZN(predicted_next_PC_o[12]) );
  OR2_X1 U134 ( .A1(n683), .A2(n684), .ZN(predicted_next_PC_o[27]) );
  OR2_X1 U332 ( .A1(n863), .A2(n864), .ZN(predicted_next_PC_o[10]) );
  OR2_X1 U101 ( .A1(n653), .A2(n654), .ZN(predicted_next_PC_o[2]) );
  OR2_X1 U277 ( .A1(n813), .A2(n814), .ZN(predicted_next_PC_o[15]) );
  OR2_X1 U68 ( .A1(n623), .A2(n624), .ZN(predicted_next_PC_o[3]) );
  OR2_X1 U178 ( .A1(n723), .A2(n724), .ZN(predicted_next_PC_o[23]) );
  OR2_X1 U46 ( .A1(n603), .A2(n604), .ZN(predicted_next_PC_o[5]) );
  OR2_X1 U200 ( .A1(n743), .A2(n744), .ZN(predicted_next_PC_o[21]) );
  OR2_X1 U266 ( .A1(n803), .A2(n804), .ZN(predicted_next_PC_o[16]) );
  OR2_X1 U233 ( .A1(n773), .A2(n774), .ZN(predicted_next_PC_o[19]) );
  OR2_X1 U189 ( .A1(n733), .A2(n734), .ZN(predicted_next_PC_o[22]) );
  OR2_X1 U255 ( .A1(n793), .A2(n794), .ZN(predicted_next_PC_o[17]) );
  OR2_X1 U244 ( .A1(n783), .A2(n784), .ZN(predicted_next_PC_o[18]) );
  OR2_X1 U321 ( .A1(n853), .A2(n854), .ZN(predicted_next_PC_o[11]) );
  OR2_X1 U112 ( .A1(n663), .A2(n664), .ZN(predicted_next_PC_o[29]) );
  OR2_X1 U299 ( .A1(n833), .A2(n834), .ZN(predicted_next_PC_o[13]) );
  OR2_X1 U288 ( .A1(n823), .A2(n824), .ZN(predicted_next_PC_o[14]) );
  OR2_X1 U211 ( .A1(n753), .A2(n754), .ZN(predicted_next_PC_o[20]) );
  OR2_X1 U167 ( .A1(n713), .A2(n714), .ZN(predicted_next_PC_o[24]) );
  OR2_X1 U123 ( .A1(n673), .A2(n674), .ZN(predicted_next_PC_o[28]) );
  OR2_X1 U145 ( .A1(n693), .A2(n694), .ZN(predicted_next_PC_o[26]) );
  OR2_X1 U343 ( .A1(n873), .A2(n874), .ZN(predicted_next_PC_o[0]) );
  OR2_X1 U222 ( .A1(n763), .A2(n764), .ZN(predicted_next_PC_o[1]) );
  OR2_X1 U90 ( .A1(n643), .A2(n644), .ZN(predicted_next_PC_o[30]) );
  OR2_X1 U13 ( .A1(n573), .A2(n574), .ZN(predicted_next_PC_o[8]) );
  OR2_X1 U79 ( .A1(n633), .A2(n634), .ZN(predicted_next_PC_o[31]) );
  OR2_X1 U24 ( .A1(n583), .A2(n584), .ZN(predicted_next_PC_o[7]) );
  OR2_X1 U35 ( .A1(n593), .A2(n594), .ZN(predicted_next_PC_o[6]) );
  OR2_X1 U2 ( .A1(n547), .A2(n548), .ZN(predicted_next_PC_o[9]) );
  OR2_X1 U57 ( .A1(n613), .A2(n614), .ZN(predicted_next_PC_o[4]) );
  INV_X1 U475 ( .A(stall_i), .ZN(N567) );
  AND2_X1 U438 ( .A1(N38), .A2(N567), .ZN(N566) );
  AND2_X1 U446 ( .A1(N43), .A2(N567), .ZN(N406) );
  AND2_X1 U439 ( .A1(N39), .A2(N567), .ZN(N534) );
  AND2_X1 U441 ( .A1(N40), .A2(N567), .ZN(N502) );
  AND2_X1 U442 ( .A1(N41), .A2(N567), .ZN(N470) );
  AND2_X1 U443 ( .A1(N42), .A2(N567), .ZN(N438) );
  AND2_X1 U463 ( .A1(N49), .A2(N567), .ZN(N214) );
  AND2_X1 U452 ( .A1(N44), .A2(N567), .ZN(N374) );
  AND2_X1 U454 ( .A1(N45), .A2(N567), .ZN(N342) );
  AND2_X1 U457 ( .A1(N46), .A2(N567), .ZN(N310) );
  AND2_X1 U459 ( .A1(N47), .A2(N567), .ZN(N278) );
  AND2_X1 U461 ( .A1(N48), .A2(N567), .ZN(N246) );
  AND2_X1 U470 ( .A1(N51), .A2(N567), .ZN(N150) );
  AND2_X1 U467 ( .A1(N50), .A2(N567), .ZN(N182) );
  AND2_X1 U436 ( .A1(N53), .A2(N567), .ZN(N86) );
  AND2_X1 U474 ( .A1(N52), .A2(N567), .ZN(N118) );
  INV_X1 U356 ( .A(taken_o), .ZN(n883) );
  BUF_X1 U360 ( .A(n572), .Z(n6) );
  BUF_X2 U361 ( .A(n571), .Z(n7) );
  BUF_X1 U363 ( .A(n570), .Z(n8) );
  BUF_X2 U364 ( .A(n569), .Z(n9) );
  BUF_X1 U367 ( .A(n556), .Z(n18) );
  BUF_X2 U368 ( .A(n555), .Z(n19) );
  BUF_X2 U370 ( .A(n553), .Z(n21) );
  BUF_X1 U371 ( .A(n560), .Z(n14) );
  BUF_X2 U375 ( .A(n559), .Z(n15) );
  BUF_X1 U376 ( .A(n558), .Z(n16) );
  BUF_X2 U378 ( .A(n557), .Z(n17) );
  BUF_X1 U379 ( .A(n568), .Z(n10) );
  BUF_X2 U382 ( .A(n567), .Z(n11) );
  BUF_X1 U384 ( .A(n566), .Z(n12) );
  BUF_X2 U387 ( .A(n565), .Z(n13) );
  BUF_X1 U389 ( .A(n554), .Z(n20) );
  INV_X1 U435 ( .A(reset), .ZN(n34) );
  INV_X1 U437 ( .A(reset), .ZN(n35) );
  INV_X1 U473 ( .A(reset), .ZN(n36) );
  INV_X1 U478 ( .A(reset), .ZN(n37) );
  INV_X1 U480 ( .A(reset), .ZN(n39) );
  INV_X1 U481 ( .A(reset), .ZN(n40) );
  INV_X1 U482 ( .A(reset), .ZN(n41) );
  INV_X1 U483 ( .A(reset), .ZN(n42) );
  INV_X1 U484 ( .A(reset), .ZN(n43) );
  INV_X1 U485 ( .A(reset), .ZN(n44) );
  INV_X1 U486 ( .A(reset), .ZN(n45) );
  INV_X1 U487 ( .A(reset), .ZN(n38) );
  INV_X1 U488 ( .A(reset), .ZN(n33) );
  INV_X1 U489 ( .A(reset), .ZN(n29) );
  INV_X1 U490 ( .A(reset), .ZN(n27) );
  INV_X1 U491 ( .A(reset), .ZN(n28) );
  INV_X1 U492 ( .A(reset), .ZN(n25) );
  INV_X1 U493 ( .A(reset), .ZN(n26) );
  INV_X1 U494 ( .A(reset), .ZN(n22) );
  INV_X1 U495 ( .A(reset), .ZN(n23) );
  INV_X1 U496 ( .A(reset), .ZN(n24) );
  INV_X1 U497 ( .A(reset), .ZN(n32) );
  INV_X1 U498 ( .A(reset), .ZN(n31) );
  INV_X1 U499 ( .A(reset), .ZN(n30) );
  NOR2_X1 U500 ( .A1(n891), .A2(n892), .ZN(n568) );
  NOR2_X1 U501 ( .A1(n894), .A2(n892), .ZN(n566) );
  NOR2_X1 U502 ( .A1(n891), .A2(n896), .ZN(n572) );
  NOR2_X1 U503 ( .A1(n894), .A2(n896), .ZN(n570) );
  NOR2_X1 U504 ( .A1(n891), .A2(n901), .ZN(n556) );
  NOR2_X1 U505 ( .A1(n894), .A2(n901), .ZN(n554) );
  NOR2_X1 U506 ( .A1(n895), .A2(n901), .ZN(n553) );
  NOR2_X1 U507 ( .A1(n902), .A2(n891), .ZN(n560) );
  NOR2_X1 U508 ( .A1(n902), .A2(n894), .ZN(n558) );
  NOR2_X1 U509 ( .A1(n893), .A2(n892), .ZN(n567) );
  NOR2_X1 U510 ( .A1(n895), .A2(n892), .ZN(n565) );
  NOR2_X1 U511 ( .A1(n893), .A2(n896), .ZN(n571) );
  NOR2_X1 U512 ( .A1(n895), .A2(n896), .ZN(n569) );
  NOR2_X1 U513 ( .A1(n893), .A2(n901), .ZN(n555) );
  NOR2_X1 U514 ( .A1(n902), .A2(n893), .ZN(n559) );
  NOR2_X1 U515 ( .A1(n895), .A2(n902), .ZN(n557) );
endmodule


module fetch_block ( branch_target_i, sum_addr_i, A_i, NPC4_i, S_MUX_PC_BUS_i, 
        PC_o, PC4_o, PC_BUS_pre_BTB, stall_i, take_prediction_i, mispredict_i, 
        predicted_PC, clk, rst );
  input [31:0] branch_target_i;
  input [31:0] sum_addr_i;
  input [31:0] A_i;
  input [31:0] NPC4_i;
  input [1:0] S_MUX_PC_BUS_i;
  output [31:0] PC_o;
  output [31:0] PC4_o;
  output [31:0] PC_BUS_pre_BTB;
  input [31:0] predicted_PC;
  input stall_i, take_prediction_i, mispredict_i, clk, rst;
  wire   en_IR;
  wire   [31:0] PC_BUS;

  ff32_en_0 PC ( .D(PC_BUS), .en(en_IR), .clk(clk), .rst(rst), .Q(PC_o) );
  add4 PCADD ( .IN1(PC_o), .OUT1(PC4_o) );
  mux41_0 MUXTARGET ( .IN0(NPC4_i), .IN1(A_i), .IN2(sum_addr_i), .IN3(
        branch_target_i), .CTRL(S_MUX_PC_BUS_i), .OUT1(PC_BUS_pre_BTB) );
  mux41_1 MUXPREDICTION ( .IN0(PC4_o), .IN1(predicted_PC), .IN2(PC_BUS_pre_BTB), .IN3(PC_BUS_pre_BTB), .CTRL({mispredict_i, take_prediction_i}), .OUT1(PC_BUS) );
  INV_X1 U1 ( .A(stall_i), .ZN(en_IR) );
endmodule


module top_level ( clock, rst, IRAM_Addr_o, IRAM_Dout_i, DRAM_Enable_o, 
        DRAM_WR_o, DRAM_Din_o, DRAM_Addr_o, DRAM_Dout_i );
  output [31:0] IRAM_Addr_o;
  input [31:0] IRAM_Dout_i;
  output [31:0] DRAM_Din_o;
  output [31:0] DRAM_Addr_o;
  input [31:0] DRAM_Dout_i;
  input clock, rst;
  output DRAM_Enable_o, DRAM_WR_o;
  wire   was_taken_from_jl, was_branch, was_jmp, was_taken, stall_fetch,
         mispredict, take_prediction, stall_btb, stall_decode, dummy_S_EXT,
         dummy_S_EXT_SIGN, dummy_S_EQ_NEQ, exe_stall_cu, dummy_S_MUX_MEM,
         dummy_S_RF_W_wb, dummy_S_RF_W_mem, dummy_S_MUX_ALUIN, stall_exe,
         enable_regfile, n3, n4;
  wire   [31:0] dummy_branch_target;
  wire   [31:0] dummy_sum_addr;
  wire   [31:0] dummy_A;
  wire   [31:0] NPCF;
  wire   [1:0] dummy_S_MUX_PC_BUS;
  wire   [31:0] PC4;
  wire   [31:0] TARGET_PC;
  wire   [31:0] predicted_PC;
  wire   [31:0] IR;
  wire   [31:0] AtoComp;
  wire   [4:0] rA2reg;
  wire   [4:0] rB2reg;
  wire   [4:0] rC2reg;
  wire   [31:0] help_IMM;
  wire   [31:0] wb2reg;
  wire   [1:0] dummy_S_FWAdec;
  wire   [4:0] muxed_dest2exe;
  wire   [4:0] D22D3;
  wire   [1:0] dummy_S_MUX_DEST;
  wire   [12:0] ALUW_dec;
  wire   [31:0] W2wb;
  wire   [31:0] dummy_B;
  wire   [31:0] A2exe;
  wire   [31:0] B2exe;
  wire   [4:0] rA2fw;
  wire   [4:0] rB2mux;
  wire   [4:0] rC2mux;
  wire   [31:0] IMM2exe;
  wire   [12:0] ALUW;
  wire   [31:0] X2mem;
  wire   [31:0] S2mem;
  wire   [1:0] dummy_S_FWA2exe;
  wire   [1:0] dummy_S_FWB2exe;
  wire   [4:0] D32reg;

  fetch_block UFETCH_BLOCK ( .branch_target_i(dummy_branch_target), 
        .sum_addr_i(dummy_sum_addr), .A_i(dummy_A), .NPC4_i(NPCF), 
        .S_MUX_PC_BUS_i(dummy_S_MUX_PC_BUS), .PC_o(IRAM_Addr_o), .PC4_o(PC4), 
        .PC_BUS_pre_BTB(TARGET_PC), .stall_i(stall_fetch), .take_prediction_i(
        take_prediction), .mispredict_i(mispredict), .predicted_PC(
        predicted_PC), .clk(clock), .rst(rst) );
  btb_N_LINES4_SIZE32 UBTB ( .clock(clock), .reset(rst), .stall_i(stall_btb), 
        .TAG_i(IRAM_Addr_o[5:2]), .target_PC_i(TARGET_PC), .was_taken_i(
        was_taken), .predicted_next_PC_o(predicted_PC), .taken_o(
        take_prediction), .mispredict_o(mispredict) );
  fetch_regs UFEETCH_REGS ( .NPCF_i(PC4), .IR_i(IRAM_Dout_i), .NPCF_o(NPCF), 
        .IR_o(IR), .stall_i(stall_decode), .clk(clock), .rst(rst) );
  jump_logic UJUMP_LOGIC ( .NPCF_i(NPCF), .IR_i({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, IR[25:0]}), .A_i(AtoComp), .A_o(dummy_A), .rA_o(rA2reg), .rB_o(
        rB2reg), .rC_o(rC2reg), .branch_target_o(dummy_branch_target), 
        .sum_addr_o(dummy_sum_addr), .extended_imm(help_IMM), .taken_o(
        was_taken_from_jl), .FW_X_i(DRAM_Addr_o), .FW_W_i(wb2reg), 
        .S_FW_Adec_i(dummy_S_FWAdec), .S_EXT_i(dummy_S_EXT), .S_EXT_SIGN_i(
        dummy_S_EXT_SIGN), .S_MUX_LINK_i(n4), .S_EQ_NEQ_i(dummy_S_EQ_NEQ) );
  dlx_cu_MICROCODE_MEM_SIZE64_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE13 UCU ( 
        .Clk(clock), .Rst(rst), .IR_IN({IR[31:16], 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, IR[10:0]}), .stall_exe_i(exe_stall_cu), .mispredict_i(mispredict), .D1_i(muxed_dest2exe), .D2_i(D22D3), .S_MUX_PC_BUS(dummy_S_MUX_PC_BUS), 
        .S_EXT(dummy_S_EXT), .S_EXT_SIGN(dummy_S_EXT_SIGN), .S_EQ_NEQ(
        dummy_S_EQ_NEQ), .S_MUX_DEST(dummy_S_MUX_DEST), .S_MUX_LINK(n4), 
        .S_MUX_MEM(dummy_S_MUX_MEM), .S_MEM_W_R(DRAM_WR_o), .S_MEM_EN(
        DRAM_Enable_o), .S_RF_W_wb(dummy_S_RF_W_wb), .S_RF_W_mem(
        dummy_S_RF_W_mem), .S_MUX_ALUIN(dummy_S_MUX_ALUIN), .stall_exe_o(
        stall_exe), .stall_dec_o(stall_decode), .stall_fetch_o(stall_fetch), 
        .stall_btb_o(stall_btb), .was_branch_o(was_branch), .was_jmp_o(was_jmp), .ALU_WORD_o(ALUW_dec) );
  dlx_regfile RF ( .Clk(clock), .Rst(rst), .ENABLE(enable_regfile), .RD1(1'b1), 
        .RD2(1'b1), .WR(dummy_S_RF_W_mem), .ADD_WR(D22D3), .ADD_RD1(
        IRAM_Dout_i[25:21]), .ADD_RD2(IRAM_Dout_i[20:16]), .DATAIN(W2wb), 
        .OUT1(AtoComp), .OUT2(dummy_B) );
  decode_regs UDECODE_REGS ( .A_i(AtoComp), .B_i(dummy_B), .rA_i(rA2reg), 
        .rB_i(rB2reg), .rC_i(rC2reg), .IMM_i(help_IMM), .ALUW_i(ALUW_dec), 
        .A_o(A2exe), .B_o(B2exe), .rA_o(rA2fw), .rB_o(rB2mux), .rC_o(rC2mux), 
        .IMM_o(IMM2exe), .ALUW_o(ALUW), .stall_i(stall_exe), .clk(clock), 
        .rst(rst) );
  execute_regs UEXECUTE_REGS ( .X_i(X2mem), .S_i(S2mem), .D2_i(muxed_dest2exe), 
        .X_o(DRAM_Addr_o), .S_o(DRAM_Din_o), .D2_o(D22D3), .stall_i(1'b0), 
        .clk(clock), .rst(rst) );
  execute_block UEXECUTE_BLOCK ( .IMM_i(IMM2exe), .A_i(A2exe), .rB_i(rB2mux), 
        .rC_i(rC2mux), .MUXED_B_i(B2exe), .S_MUX_ALUIN_i(dummy_S_MUX_ALUIN), 
        .FW_X_i(DRAM_Addr_o), .FW_W_i(wb2reg), .S_FW_A_i(dummy_S_FWA2exe), 
        .S_FW_B_i(dummy_S_FWB2exe), .muxed_dest(muxed_dest2exe), .muxed_B(
        S2mem), .S_MUX_DEST_i(dummy_S_MUX_DEST), .OP({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .ALUW_i(ALUW), .DOUT(X2mem), .stall_o(exe_stall_cu), .Clock(
        clock), .Reset(rst) );
  mem_regs UMEM_REGS ( .W_i(W2wb), .D3_i(D22D3), .W_o(wb2reg), .D3_o(D32reg), 
        .clk(clock), .rst(rst) );
  mem_block UMEM_BLOCK ( .X_i(DRAM_Addr_o), .LOAD_i(DRAM_Dout_i), 
        .S_MUX_MEM_i(dummy_S_MUX_MEM), .W_o(W2wb) );
  fw_logic UFW_LOGIC ( .D1_i({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .rAdec_i(
        IR[25:21]), .D2_i(D22D3), .D3_i(D32reg), .rA_i(rA2fw), .rB_i(rB2mux), 
        .S_mem_W(dummy_S_RF_W_mem), .S_mem_LOAD(dummy_S_MUX_MEM), .S_wb_W(
        dummy_S_RF_W_wb), .S_exe_W(1'b0), .S_FWAdec(dummy_S_FWAdec), .S_FWA(
        dummy_S_FWA2exe), .S_FWB(dummy_S_FWB2exe) );
  AOI21_X1 U4 ( .B1(was_taken_from_jl), .B2(was_branch), .A(was_jmp), .ZN(n3)
         );
  INV_X1 U5 ( .A(stall_decode), .ZN(enable_regfile) );
  INV_X2 U6 ( .A(n3), .ZN(was_taken) );
endmodule

