
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_top_level is

-- define attributes
attribute ENUM_ENCODING : STRING;

-- define any necessary types
type aluOp is (NOP, SLLS, SRLS, SRAS, ADDS, ADDUS, SUBS, SUBUS, ANDS, ORS, 
   XORS, SEQS, SNES, SLTS, SGTS, SLES, SGES, MOVI2SS, MOVS2IS, MOVFS, MOVDS, 
   MOVFP2IS, MOVI2FP, MOVI2TS, MOVT2IS, SLTUS, SGTUS, SLEUS, SGEUS, MULTU, 
   MULTS);
attribute ENUM_ENCODING of aluOp : type is 
   "00000 00001 00010 00011 00100 00101 00110 00111 01000 01001 01010 01011 01100 01101 01110 01111 10000 10001 10010 10011 10100 10101 10110 10111 11000 11001 11010 11011 11100 11101 11110";
type UNSIGNED is array (INTEGER range <>) of std_logic;
   
   -- Declarations for conversion functions.
   function std_logic_vector_to_aluOp(arg : in std_logic_vector( 1 to 5 )) 
               return aluOp;
   function aluOp_to_std_logic_vector(arg : in aluOp) return std_logic_vector;

end CONV_PACK_top_level;

package body CONV_PACK_top_level is
   
   -- std_logic_vector to enum type function
   function std_logic_vector_to_aluOp(arg : in std_logic_vector( 1 to 5 )) 
   return aluOp is
   -- synopsys built_in SYN_FEED_THRU;
   begin
      case arg is
         when "00000" => return NOP;
         when "00001" => return SLLS;
         when "00010" => return SRLS;
         when "00011" => return SRAS;
         when "00100" => return ADDS;
         when "00101" => return ADDUS;
         when "00110" => return SUBS;
         when "00111" => return SUBUS;
         when "01000" => return ANDS;
         when "01001" => return ORS;
         when "01010" => return XORS;
         when "01011" => return SEQS;
         when "01100" => return SNES;
         when "01101" => return SLTS;
         when "01110" => return SGTS;
         when "01111" => return SLES;
         when "10000" => return SGES;
         when "10001" => return MOVI2SS;
         when "10010" => return MOVS2IS;
         when "10011" => return MOVFS;
         when "10100" => return MOVDS;
         when "10101" => return MOVFP2IS;
         when "10110" => return MOVI2FP;
         when "10111" => return MOVI2TS;
         when "11000" => return MOVT2IS;
         when "11001" => return SLTUS;
         when "11010" => return SGTUS;
         when "11011" => return SLEUS;
         when "11100" => return SGEUS;
         when "11101" => return MULTU;
         when "11110" => return MULTS;
         when others => assert FALSE -- this should not happen.
               report "un-convertible value"
               severity warning;
               return NOP;
      end case;
   end;
   
   -- enum type to std_logic_vector function
   function aluOp_to_std_logic_vector(arg : in aluOp) return std_logic_vector 
   is
   -- synopsys built_in SYN_FEED_THRU;
   begin
      case arg is
         when NOP => return "00000";
         when SLLS => return "00001";
         when SRLS => return "00010";
         when SRAS => return "00011";
         when ADDS => return "00100";
         when ADDUS => return "00101";
         when SUBS => return "00110";
         when SUBUS => return "00111";
         when ANDS => return "01000";
         when ORS => return "01001";
         when XORS => return "01010";
         when SEQS => return "01011";
         when SNES => return "01100";
         when SLTS => return "01101";
         when SGTS => return "01110";
         when SLES => return "01111";
         when SGES => return "10000";
         when MOVI2SS => return "10001";
         when MOVS2IS => return "10010";
         when MOVFS => return "10011";
         when MOVDS => return "10100";
         when MOVFP2IS => return "10101";
         when MOVI2FP => return "10110";
         when MOVI2TS => return "10111";
         when MOVT2IS => return "11000";
         when SLTUS => return "11001";
         when SGTUS => return "11010";
         when SLEUS => return "11011";
         when SGEUS => return "11100";
         when MULTU => return "11101";
         when MULTS => return "11110";
         when others => assert FALSE -- this should not happen.
               report "un-convertible value"
               severity warning;
               return "00000";
      end case;
   end;

end CONV_PACK_top_level;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity mux21_4 is

   port( IN0, IN1 : in std_logic_vector (31 downto 0);  CTRL : in std_logic;  
         OUT1 : out std_logic_vector (31 downto 0));

end mux21_4;

architecture SYN_Bhe of mux21_4 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => IN0(9), B => IN1(9), S => CTRL, Z => OUT1(9));
   U2 : MUX2_X1 port map( A => IN0(8), B => IN1(8), S => CTRL, Z => OUT1(8));
   U3 : MUX2_X1 port map( A => IN0(7), B => IN1(7), S => CTRL, Z => OUT1(7));
   U4 : MUX2_X1 port map( A => IN0(6), B => IN1(6), S => CTRL, Z => OUT1(6));
   U5 : MUX2_X1 port map( A => IN0(5), B => IN1(5), S => CTRL, Z => OUT1(5));
   U6 : MUX2_X1 port map( A => IN0(4), B => IN1(4), S => CTRL, Z => OUT1(4));
   U7 : MUX2_X1 port map( A => IN0(3), B => IN1(3), S => CTRL, Z => OUT1(3));
   U8 : MUX2_X1 port map( A => IN0(31), B => IN1(31), S => CTRL, Z => OUT1(31))
                           ;
   U9 : MUX2_X1 port map( A => IN0(30), B => IN1(30), S => CTRL, Z => OUT1(30))
                           ;
   U10 : MUX2_X1 port map( A => IN0(2), B => IN1(2), S => CTRL, Z => OUT1(2));
   U11 : MUX2_X1 port map( A => IN0(29), B => IN1(29), S => CTRL, Z => OUT1(29)
                           );
   U12 : MUX2_X1 port map( A => IN0(28), B => IN1(28), S => CTRL, Z => OUT1(28)
                           );
   U13 : MUX2_X1 port map( A => IN0(27), B => IN1(27), S => CTRL, Z => OUT1(27)
                           );
   U14 : MUX2_X1 port map( A => IN0(26), B => IN1(26), S => CTRL, Z => OUT1(26)
                           );
   U15 : MUX2_X1 port map( A => IN0(25), B => IN1(25), S => CTRL, Z => OUT1(25)
                           );
   U16 : MUX2_X1 port map( A => IN0(24), B => IN1(24), S => CTRL, Z => OUT1(24)
                           );
   U17 : MUX2_X1 port map( A => IN0(23), B => IN1(23), S => CTRL, Z => OUT1(23)
                           );
   U18 : MUX2_X1 port map( A => IN0(22), B => IN1(22), S => CTRL, Z => OUT1(22)
                           );
   U19 : MUX2_X1 port map( A => IN0(21), B => IN1(21), S => CTRL, Z => OUT1(21)
                           );
   U20 : MUX2_X1 port map( A => IN0(20), B => IN1(20), S => CTRL, Z => OUT1(20)
                           );
   U21 : MUX2_X1 port map( A => IN0(1), B => IN1(1), S => CTRL, Z => OUT1(1));
   U22 : MUX2_X1 port map( A => IN0(19), B => IN1(19), S => CTRL, Z => OUT1(19)
                           );
   U23 : MUX2_X1 port map( A => IN0(18), B => IN1(18), S => CTRL, Z => OUT1(18)
                           );
   U24 : MUX2_X1 port map( A => IN0(17), B => IN1(17), S => CTRL, Z => OUT1(17)
                           );
   U25 : MUX2_X1 port map( A => IN0(16), B => IN1(16), S => CTRL, Z => OUT1(16)
                           );
   U26 : MUX2_X1 port map( A => IN0(15), B => IN1(15), S => CTRL, Z => OUT1(15)
                           );
   U27 : MUX2_X1 port map( A => IN0(14), B => IN1(14), S => CTRL, Z => OUT1(14)
                           );
   U28 : MUX2_X1 port map( A => IN0(13), B => IN1(13), S => CTRL, Z => OUT1(13)
                           );
   U29 : MUX2_X1 port map( A => IN0(12), B => IN1(12), S => CTRL, Z => OUT1(12)
                           );
   U30 : MUX2_X1 port map( A => IN0(11), B => IN1(11), S => CTRL, Z => OUT1(11)
                           );
   U31 : MUX2_X1 port map( A => IN0(10), B => IN1(10), S => CTRL, Z => OUT1(10)
                           );
   U32 : MUX2_X1 port map( A => IN0(0), B => IN1(0), S => CTRL, Z => OUT1(0));

end SYN_Bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity mux21_3 is

   port( IN0, IN1 : in std_logic_vector (31 downto 0);  OUT1 : out 
         std_logic_vector (31 downto 0);  CTRL_BAR : in std_logic);

end mux21_3;

architecture SYN_Bhe of mux21_3 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U32 : MUX2_X1 port map( A => IN0(0), B => IN1(0), S => n1, Z => OUT1(0));
   U9 : MUX2_X1 port map( A => IN0(30), B => IN1(30), S => n2, Z => OUT1(30));
   U11 : MUX2_X1 port map( A => IN0(29), B => IN1(29), S => n2, Z => OUT1(29));
   U12 : MUX2_X1 port map( A => IN0(28), B => IN1(28), S => n2, Z => OUT1(28));
   U8 : MUX2_X1 port map( A => IN0(31), B => IN1(31), S => n2, Z => OUT1(31));
   U15 : MUX2_X1 port map( A => IN0(25), B => IN1(25), S => n3, Z => OUT1(25));
   U26 : MUX2_X1 port map( A => IN0(15), B => IN1(15), S => n1, Z => OUT1(15));
   U27 : MUX2_X1 port map( A => IN0(14), B => IN1(14), S => n1, Z => OUT1(14));
   U1 : MUX2_X1 port map( A => IN0(9), B => IN1(9), S => n2, Z => OUT1(9));
   U28 : MUX2_X1 port map( A => IN0(13), B => IN1(13), S => n1, Z => OUT1(13));
   U24 : MUX2_X1 port map( A => IN0(17), B => IN1(17), S => n3, Z => OUT1(17));
   U10 : MUX2_X1 port map( A => IN0(2), B => IN1(2), S => n2, Z => OUT1(2));
   U29 : MUX2_X1 port map( A => IN0(12), B => IN1(12), S => n1, Z => OUT1(12));
   U31 : MUX2_X1 port map( A => IN0(10), B => IN1(10), S => n1, Z => OUT1(10));
   U30 : MUX2_X1 port map( A => IN0(11), B => IN1(11), S => n1, Z => OUT1(11));
   U7 : MUX2_X1 port map( A => IN0(3), B => IN1(3), S => n2, Z => OUT1(3));
   U22 : MUX2_X1 port map( A => IN0(19), B => IN1(19), S => n3, Z => OUT1(19));
   U20 : MUX2_X1 port map( A => IN0(20), B => IN1(20), S => n3, Z => OUT1(20));
   U23 : MUX2_X1 port map( A => IN0(18), B => IN1(18), S => n3, Z => OUT1(18));
   U16 : MUX2_X1 port map( A => IN0(24), B => IN1(24), S => n3, Z => OUT1(24));
   U19 : MUX2_X1 port map( A => IN0(21), B => IN1(21), S => n3, Z => OUT1(21));
   U25 : MUX2_X1 port map( A => IN0(16), B => IN1(16), S => n1, Z => OUT1(16));
   U2 : MUX2_X1 port map( A => IN0(8), B => IN1(8), S => n2, Z => OUT1(8));
   U4 : MUX2_X1 port map( A => IN0(6), B => IN1(6), S => n2, Z => OUT1(6));
   U18 : MUX2_X1 port map( A => IN0(22), B => IN1(22), S => n3, Z => OUT1(22));
   U13 : MUX2_X1 port map( A => IN0(27), B => IN1(27), S => n3, Z => OUT1(27));
   U17 : MUX2_X1 port map( A => IN0(23), B => IN1(23), S => n3, Z => OUT1(23));
   U5 : MUX2_X1 port map( A => IN0(5), B => IN1(5), S => n2, Z => OUT1(5));
   U21 : MUX2_X1 port map( A => IN0(1), B => IN1(1), S => n3, Z => OUT1(1));
   U6 : MUX2_X1 port map( A => IN0(4), B => IN1(4), S => n2, Z => OUT1(4));
   U3 : MUX2_X1 port map( A => IN0(7), B => IN1(7), S => n2, Z => OUT1(7));
   U14 : MUX2_X1 port map( A => IN0(26), B => IN1(26), S => n3, Z => OUT1(26));
   U33 : INV_X1 port map( A => CTRL_BAR, ZN => n1);
   U34 : INV_X1 port map( A => CTRL_BAR, ZN => n3);
   U35 : INV_X1 port map( A => CTRL_BAR, ZN => n2);

end SYN_Bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_47 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_47;

architecture SYN_BEHAVIORAL of FA_47 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n10, n11, n12 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n12, ZN => S);
   U3 : NAND2_X1 port map( A1 => n11, A2 => n10, ZN => Co);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n12);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n10);
   U5 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n11);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_96 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_96;

architecture SYN_BEHAVIORAL of FA_96 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n6 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U1 : XNOR2_X1 port map( A => n6, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_37 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_37;

architecture SYN_BEHAVIORAL of FA_37 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n6 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U1 : XNOR2_X1 port map( A => n6, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_33 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_33;

architecture SYN_BEHAVIORAL of FA_33 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n6 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U1 : XNOR2_X1 port map( A => n6, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_111 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_111;

architecture SYN_BEHAVIORAL of FA_111 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_103 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_103;

architecture SYN_BEHAVIORAL of FA_103 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_95 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_95;

architecture SYN_BEHAVIORAL of FA_95 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_87 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_87;

architecture SYN_BEHAVIORAL of FA_87 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_79 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_79;

architecture SYN_BEHAVIORAL of FA_79 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_71 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_71;

architecture SYN_BEHAVIORAL of FA_71 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_56 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_56;

architecture SYN_BEHAVIORAL of FA_56 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_48 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_48;

architecture SYN_BEHAVIORAL of FA_48 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_40 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_40;

architecture SYN_BEHAVIORAL of FA_40 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_32 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_32;

architecture SYN_BEHAVIORAL of FA_32 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_24 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_24;

architecture SYN_BEHAVIORAL of FA_24 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_16 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_16;

architecture SYN_BEHAVIORAL of FA_16 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_8 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_8;

architecture SYN_BEHAVIORAL of FA_8 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_115 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_115;

architecture SYN_BEHAVIORAL of FA_115 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => S);
   U2 : OR2_X1 port map( A1 => A, A2 => B, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_107 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_107;

architecture SYN_BEHAVIORAL of FA_107 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => S);
   U2 : OR2_X1 port map( A1 => A, A2 => B, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_99 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_99;

architecture SYN_BEHAVIORAL of FA_99 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => S);
   U2 : OR2_X1 port map( A1 => A, A2 => B, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_91 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_91;

architecture SYN_BEHAVIORAL of FA_91 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => S);
   U2 : OR2_X1 port map( A1 => A, A2 => B, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_83 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_83;

architecture SYN_BEHAVIORAL of FA_83 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => S);
   U2 : OR2_X1 port map( A1 => A, A2 => B, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_75 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_75;

architecture SYN_BEHAVIORAL of FA_75 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => S);
   U2 : OR2_X1 port map( A1 => A, A2 => B, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_67 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_67;

architecture SYN_BEHAVIORAL of FA_67 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => A, A2 => B, ZN => Co);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_60 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_60;

architecture SYN_BEHAVIORAL of FA_60 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => A, A2 => B, ZN => Co);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_52 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_52;

architecture SYN_BEHAVIORAL of FA_52 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => S);
   U2 : OR2_X1 port map( A1 => A, A2 => B, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_44 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_44;

architecture SYN_BEHAVIORAL of FA_44 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => A, A2 => B, ZN => Co);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_36 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_36;

architecture SYN_BEHAVIORAL of FA_36 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => A, A2 => B, ZN => Co);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_28 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_28;

architecture SYN_BEHAVIORAL of FA_28 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => S);
   U2 : OR2_X1 port map( A1 => A, A2 => B, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_20 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_20;

architecture SYN_BEHAVIORAL of FA_20 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => S);
   U2 : OR2_X1 port map( A1 => A, A2 => B, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_12 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_12;

architecture SYN_BEHAVIORAL of FA_12 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => S);
   U2 : OR2_X1 port map( A1 => A, A2 => B, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_4 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_4;

architecture SYN_BEHAVIORAL of FA_4 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => S);
   U2 : OR2_X1 port map( A1 => A, A2 => B, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_125 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_125;

architecture SYN_BEHAVIORAL of FA_125 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n9, n10, n11 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n11);
   U1 : XNOR2_X1 port map( A => Ci, B => n11, ZN => S);
   U5 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n10);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n9);
   U3 : NAND2_X1 port map( A1 => n10, A2 => n9, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_118 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_118;

architecture SYN_BEHAVIORAL of FA_118 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n9, n10, n11 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n11);
   U1 : XNOR2_X1 port map( A => Ci, B => n11, ZN => S);
   U5 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n10);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n9);
   U3 : NAND2_X1 port map( A1 => n10, A2 => n9, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_117 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_117;

architecture SYN_BEHAVIORAL of FA_117 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n9, n10, n11 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n11);
   U1 : XNOR2_X1 port map( A => Ci, B => n11, ZN => S);
   U5 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n10);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n9);
   U3 : NAND2_X1 port map( A1 => n10, A2 => n9, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_114 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_114;

architecture SYN_BEHAVIORAL of FA_114 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n9, n10, n11 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n11);
   U1 : XNOR2_X1 port map( A => Ci, B => n11, ZN => S);
   U5 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n10);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n9);
   U3 : NAND2_X1 port map( A1 => n10, A2 => n9, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_113 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_113;

architecture SYN_BEHAVIORAL of FA_113 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n9, n10, n11 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n11);
   U1 : XNOR2_X1 port map( A => Ci, B => n11, ZN => S);
   U5 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n10);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n9);
   U3 : NAND2_X1 port map( A1 => n10, A2 => n9, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_109 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_109;

architecture SYN_BEHAVIORAL of FA_109 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n9, n10, n11 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n11);
   U1 : XNOR2_X1 port map( A => Ci, B => n11, ZN => S);
   U5 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n10);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n9);
   U3 : NAND2_X1 port map( A1 => n10, A2 => n9, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_106 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_106;

architecture SYN_BEHAVIORAL of FA_106 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n9, n10, n11 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n11);
   U1 : XNOR2_X1 port map( A => Ci, B => n11, ZN => S);
   U5 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n10);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n9);
   U3 : NAND2_X1 port map( A1 => n10, A2 => n9, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_105 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_105;

architecture SYN_BEHAVIORAL of FA_105 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n9, n10, n11 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n11);
   U1 : XNOR2_X1 port map( A => Ci, B => n11, ZN => S);
   U5 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n10);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n9);
   U3 : NAND2_X1 port map( A1 => n10, A2 => n9, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_102 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_102;

architecture SYN_BEHAVIORAL of FA_102 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n9, n10, n11 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n11);
   U1 : XNOR2_X1 port map( A => Ci, B => n11, ZN => S);
   U5 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n10);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n9);
   U3 : NAND2_X1 port map( A1 => n10, A2 => n9, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_101 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_101;

architecture SYN_BEHAVIORAL of FA_101 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n9, n10, n11 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n11);
   U1 : XNOR2_X1 port map( A => Ci, B => n11, ZN => S);
   U5 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n10);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n9);
   U3 : NAND2_X1 port map( A1 => n10, A2 => n9, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_98 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_98;

architecture SYN_BEHAVIORAL of FA_98 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n9, n10, n11 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n11);
   U1 : XNOR2_X1 port map( A => Ci, B => n11, ZN => S);
   U5 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n10);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n9);
   U3 : NAND2_X1 port map( A1 => n10, A2 => n9, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_97 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_97;

architecture SYN_BEHAVIORAL of FA_97 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n9, n10, n11 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n11);
   U1 : XNOR2_X1 port map( A => Ci, B => n11, ZN => S);
   U5 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n10);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n9);
   U3 : NAND2_X1 port map( A1 => n10, A2 => n9, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_94 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_94;

architecture SYN_BEHAVIORAL of FA_94 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n9, n10, n11 : std_logic;

begin
   
   U3 : NAND2_X1 port map( A1 => n10, A2 => n9, ZN => Co);
   U1 : XNOR2_X1 port map( A => Ci, B => n11, ZN => S);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n11);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n9);
   U5 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_93 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_93;

architecture SYN_BEHAVIORAL of FA_93 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n9, n10, n11 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n11, ZN => S);
   U3 : NAND2_X1 port map( A1 => n10, A2 => n9, ZN => Co);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n11);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n9);
   U5 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_90 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_90;

architecture SYN_BEHAVIORAL of FA_90 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n9, n10, n11 : std_logic;

begin
   
   U3 : NAND2_X1 port map( A1 => n10, A2 => n9, ZN => Co);
   U1 : XNOR2_X1 port map( A => Ci, B => n11, ZN => S);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n11);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n9);
   U5 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_89 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_89;

architecture SYN_BEHAVIORAL of FA_89 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n9, n10, n11 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n11, ZN => S);
   U3 : NAND2_X1 port map( A1 => n10, A2 => n9, ZN => Co);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n11);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n9);
   U5 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_86 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_86;

architecture SYN_BEHAVIORAL of FA_86 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n9, n10, n11 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n11, ZN => S);
   U3 : NAND2_X1 port map( A1 => n10, A2 => n9, ZN => Co);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n11);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n9);
   U5 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_85 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_85;

architecture SYN_BEHAVIORAL of FA_85 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n9, n10, n11 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n11, ZN => S);
   U3 : NAND2_X1 port map( A1 => n10, A2 => n9, ZN => Co);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n11);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n9);
   U5 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_82 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_82;

architecture SYN_BEHAVIORAL of FA_82 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n9, n10, n11 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n11, ZN => S);
   U3 : NAND2_X1 port map( A1 => n10, A2 => n9, ZN => Co);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n11);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n9);
   U5 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_81 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_81;

architecture SYN_BEHAVIORAL of FA_81 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n9, n10, n11 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n11, ZN => S);
   U3 : NAND2_X1 port map( A1 => n10, A2 => n9, ZN => Co);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n11);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n9);
   U5 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_78 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_78;

architecture SYN_BEHAVIORAL of FA_78 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n9, n10, n11 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n11, ZN => S);
   U3 : NAND2_X1 port map( A1 => n10, A2 => n9, ZN => Co);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n11);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n9);
   U5 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_77 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_77;

architecture SYN_BEHAVIORAL of FA_77 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n9, n10, n11 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n11, ZN => S);
   U3 : NAND2_X1 port map( A1 => n10, A2 => n9, ZN => Co);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n11);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n9);
   U5 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_74 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_74;

architecture SYN_BEHAVIORAL of FA_74 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n9, n10, n11 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n11, ZN => S);
   U3 : NAND2_X1 port map( A1 => n10, A2 => n9, ZN => Co);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n11);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n9);
   U5 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_73 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_73;

architecture SYN_BEHAVIORAL of FA_73 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n9, n10, n11 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n11, ZN => S);
   U3 : NAND2_X1 port map( A1 => n10, A2 => n9, ZN => Co);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n11);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n9);
   U5 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_70 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_70;

architecture SYN_BEHAVIORAL of FA_70 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n9, n10, n11 : std_logic;

begin
   
   U3 : NAND2_X1 port map( A1 => n10, A2 => n9, ZN => Co);
   U1 : XNOR2_X1 port map( A => Ci, B => n11, ZN => S);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n11);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n9);
   U5 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_69 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_69;

architecture SYN_BEHAVIORAL of FA_69 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n9, n10, n11 : std_logic;

begin
   
   U3 : NAND2_X1 port map( A1 => n10, A2 => n9, ZN => Co);
   U1 : XNOR2_X1 port map( A => Ci, B => n11, ZN => S);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n11);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n9);
   U5 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_66 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_66;

architecture SYN_BEHAVIORAL of FA_66 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n9, n10, n11 : std_logic;

begin
   
   U3 : NAND2_X1 port map( A1 => n10, A2 => n9, ZN => Co);
   U1 : XNOR2_X1 port map( A => Ci, B => n11, ZN => S);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n11);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n9);
   U5 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_65 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_65;

architecture SYN_BEHAVIORAL of FA_65 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n9, n10, n11 : std_logic;

begin
   
   U3 : NAND2_X1 port map( A1 => n10, A2 => n9, ZN => Co);
   U1 : XNOR2_X1 port map( A => Ci, B => n11, ZN => S);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n11);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n9);
   U5 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_63 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_63;

architecture SYN_BEHAVIORAL of FA_63 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n9, n10, n11 : std_logic;

begin
   
   U3 : NAND2_X1 port map( A1 => n10, A2 => n9, ZN => Co);
   U1 : XNOR2_X1 port map( A => Ci, B => n11, ZN => S);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n11);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n9);
   U5 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_62 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_62;

architecture SYN_BEHAVIORAL of FA_62 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n9, n10, n11 : std_logic;

begin
   
   U3 : NAND2_X1 port map( A1 => n10, A2 => n9, ZN => Co);
   U1 : XNOR2_X1 port map( A => Ci, B => n11, ZN => S);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n11);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n9);
   U5 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_59 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_59;

architecture SYN_BEHAVIORAL of FA_59 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n9, n10, n11 : std_logic;

begin
   
   U3 : NAND2_X1 port map( A1 => n10, A2 => n9, ZN => Co);
   U1 : XNOR2_X1 port map( A => Ci, B => n11, ZN => S);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n11);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n9);
   U5 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_58 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_58;

architecture SYN_BEHAVIORAL of FA_58 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n9, n10, n11 : std_logic;

begin
   
   U3 : NAND2_X1 port map( A1 => n10, A2 => n9, ZN => Co);
   U1 : XNOR2_X1 port map( A => Ci, B => n11, ZN => S);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n11);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n9);
   U5 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_55 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_55;

architecture SYN_BEHAVIORAL of FA_55 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n9, n10, n11 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n11, ZN => S);
   U3 : NAND2_X1 port map( A1 => n10, A2 => n9, ZN => Co);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n11);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n9);
   U5 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_54 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_54;

architecture SYN_BEHAVIORAL of FA_54 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n9, n10, n11 : std_logic;

begin
   
   U3 : NAND2_X1 port map( A1 => n10, A2 => n9, ZN => Co);
   U1 : XNOR2_X1 port map( A => Ci, B => n11, ZN => S);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n11);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n9);
   U5 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_51 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_51;

architecture SYN_BEHAVIORAL of FA_51 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n9, n10, n11 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n11, ZN => S);
   U3 : NAND2_X1 port map( A1 => n10, A2 => n9, ZN => Co);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n11);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n9);
   U5 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_50 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_50;

architecture SYN_BEHAVIORAL of FA_50 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n9, n10, n11 : std_logic;

begin
   
   U3 : NAND2_X1 port map( A1 => n10, A2 => n9, ZN => Co);
   U1 : XNOR2_X1 port map( A => Ci, B => n11, ZN => S);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n11);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n9);
   U5 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_46 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_46;

architecture SYN_BEHAVIORAL of FA_46 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n9, n10, n11 : std_logic;

begin
   
   U3 : NAND2_X1 port map( A1 => n10, A2 => n9, ZN => Co);
   U1 : XNOR2_X1 port map( A => Ci, B => n11, ZN => S);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n11);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n9);
   U5 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_43 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_43;

architecture SYN_BEHAVIORAL of FA_43 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n9, n10, n11 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n11, ZN => S);
   U3 : NAND2_X1 port map( A1 => n10, A2 => n9, ZN => Co);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n11);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n9);
   U5 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_42 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_42;

architecture SYN_BEHAVIORAL of FA_42 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n9, n10, n11 : std_logic;

begin
   
   U3 : NAND2_X1 port map( A1 => n10, A2 => n9, ZN => Co);
   U1 : XNOR2_X1 port map( A => Ci, B => n11, ZN => S);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n11);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n9);
   U5 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_39 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_39;

architecture SYN_BEHAVIORAL of FA_39 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n9, n10, n11 : std_logic;

begin
   
   U3 : NAND2_X1 port map( A1 => n10, A2 => n9, ZN => Co);
   U1 : XNOR2_X1 port map( A => Ci, B => n11, ZN => S);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n9);
   U4 : XNOR2_X1 port map( A => B, B => A, ZN => n11);
   U5 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_38 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_38;

architecture SYN_BEHAVIORAL of FA_38 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n9, n10, n11 : std_logic;

begin
   
   U3 : NAND2_X1 port map( A1 => n10, A2 => n9, ZN => Co);
   U1 : XNOR2_X1 port map( A => Ci, B => n11, ZN => S);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n11);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n9);
   U5 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_35 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_35;

architecture SYN_BEHAVIORAL of FA_35 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n9, n10, n11 : std_logic;

begin
   
   U3 : NAND2_X1 port map( A1 => n10, A2 => n9, ZN => Co);
   U1 : XNOR2_X1 port map( A => Ci, B => n11, ZN => S);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n9);
   U4 : XNOR2_X1 port map( A => B, B => A, ZN => n11);
   U5 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_34 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_34;

architecture SYN_BEHAVIORAL of FA_34 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n9, n10, n11 : std_logic;

begin
   
   U3 : NAND2_X1 port map( A1 => n10, A2 => n9, ZN => Co);
   U1 : XNOR2_X1 port map( A => Ci, B => n11, ZN => S);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n11);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n9);
   U5 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_31 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_31;

architecture SYN_BEHAVIORAL of FA_31 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n9, n10, n11 : std_logic;

begin
   
   U3 : NAND2_X1 port map( A1 => n10, A2 => n9, ZN => Co);
   U1 : XNOR2_X1 port map( A => Ci, B => n11, ZN => S);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n11);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n9);
   U5 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_30 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_30;

architecture SYN_BEHAVIORAL of FA_30 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n9, n10, n11 : std_logic;

begin
   
   U5 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n10);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n9);
   U3 : NAND2_X1 port map( A1 => n10, A2 => n9, ZN => Co);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n11);
   U1 : XNOR2_X1 port map( A => Ci, B => n11, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_27 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_27;

architecture SYN_BEHAVIORAL of FA_27 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n9, n10, n11 : std_logic;

begin
   
   U3 : NAND2_X1 port map( A1 => n10, A2 => n9, ZN => Co);
   U1 : XNOR2_X1 port map( A => Ci, B => n11, ZN => S);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n11);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n9);
   U5 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_26 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_26;

architecture SYN_BEHAVIORAL of FA_26 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n9, n10, n11 : std_logic;

begin
   
   U5 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n10);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n9);
   U3 : NAND2_X1 port map( A1 => n10, A2 => n9, ZN => Co);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n11);
   U1 : XNOR2_X1 port map( A => Ci, B => n11, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_23 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_23;

architecture SYN_BEHAVIORAL of FA_23 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n9, n10, n11 : std_logic;

begin
   
   U5 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n10);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n9);
   U3 : NAND2_X1 port map( A1 => n10, A2 => n9, ZN => Co);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n11);
   U1 : XNOR2_X1 port map( A => Ci, B => n11, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_22 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_22;

architecture SYN_BEHAVIORAL of FA_22 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n9, n10, n11 : std_logic;

begin
   
   U3 : NAND2_X1 port map( A1 => n10, A2 => n9, ZN => Co);
   U1 : XNOR2_X1 port map( A => Ci, B => n11, ZN => S);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n11);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n9);
   U5 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_19 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_19;

architecture SYN_BEHAVIORAL of FA_19 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n9, n10, n11 : std_logic;

begin
   
   U5 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n10);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n9);
   U3 : NAND2_X1 port map( A1 => n10, A2 => n9, ZN => Co);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n11);
   U1 : XNOR2_X1 port map( A => Ci, B => n11, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_18 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_18;

architecture SYN_BEHAVIORAL of FA_18 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n9, n10, n11 : std_logic;

begin
   
   U3 : NAND2_X1 port map( A1 => n10, A2 => n9, ZN => Co);
   U1 : XNOR2_X1 port map( A => Ci, B => n11, ZN => S);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n11);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n9);
   U5 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_15 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_15;

architecture SYN_BEHAVIORAL of FA_15 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n9, n10, n11 : std_logic;

begin
   
   U5 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n10);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n9);
   U3 : NAND2_X1 port map( A1 => n10, A2 => n9, ZN => Co);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n11);
   U1 : XNOR2_X1 port map( A => Ci, B => n11, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_14 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_14;

architecture SYN_BEHAVIORAL of FA_14 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n9, n10, n11 : std_logic;

begin
   
   U3 : NAND2_X1 port map( A1 => n10, A2 => n9, ZN => Co);
   U1 : XNOR2_X1 port map( A => Ci, B => n11, ZN => S);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n11);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n9);
   U5 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_11 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_11;

architecture SYN_BEHAVIORAL of FA_11 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n9, n10, n11 : std_logic;

begin
   
   U5 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n10);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n9);
   U3 : NAND2_X1 port map( A1 => n10, A2 => n9, ZN => Co);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n11);
   U1 : XNOR2_X1 port map( A => Ci, B => n11, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_10 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_10;

architecture SYN_BEHAVIORAL of FA_10 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n9, n10, n11 : std_logic;

begin
   
   U3 : NAND2_X1 port map( A1 => n10, A2 => n9, ZN => Co);
   U1 : XNOR2_X1 port map( A => Ci, B => n11, ZN => S);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n11);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n9);
   U5 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_7 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_7;

architecture SYN_BEHAVIORAL of FA_7 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n9, n10, n11 : std_logic;

begin
   
   U5 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n10);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n9);
   U3 : NAND2_X1 port map( A1 => n10, A2 => n9, ZN => Co);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n11);
   U1 : XNOR2_X1 port map( A => Ci, B => n11, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_6 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_6;

architecture SYN_BEHAVIORAL of FA_6 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n9, n10, n11 : std_logic;

begin
   
   U5 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n10);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n9);
   U3 : NAND2_X1 port map( A1 => n10, A2 => n9, ZN => Co);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n11);
   U1 : XNOR2_X1 port map( A => Ci, B => n11, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_3 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_3;

architecture SYN_BEHAVIORAL of FA_3 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n9, n10, n11 : std_logic;

begin
   
   U5 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n10);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n9);
   U3 : NAND2_X1 port map( A1 => n10, A2 => n9, ZN => Co);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n11);
   U1 : XNOR2_X1 port map( A => Ci, B => n11, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_2 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_2;

architecture SYN_BEHAVIORAL of FA_2 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n9, n10, n11 : std_logic;

begin
   
   U5 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n10);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n9);
   U3 : NAND2_X1 port map( A1 => n10, A2 => n9, ZN => Co);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n11);
   U1 : XNOR2_X1 port map( A => Ci, B => n11, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_116 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_116;

architecture SYN_BEHAVIORAL of FA_116 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n5);
   U1 : XNOR2_X1 port map( A => n5, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_112 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_112;

architecture SYN_BEHAVIORAL of FA_112 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n5);
   U1 : XNOR2_X1 port map( A => n5, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_108 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_108;

architecture SYN_BEHAVIORAL of FA_108 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n5);
   U1 : XNOR2_X1 port map( A => n5, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_104 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_104;

architecture SYN_BEHAVIORAL of FA_104 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n5);
   U1 : XNOR2_X1 port map( A => n5, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_92 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_92;

architecture SYN_BEHAVIORAL of FA_92 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n6 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U1 : XNOR2_X1 port map( A => n6, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_88 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_88;

architecture SYN_BEHAVIORAL of FA_88 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n6 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U1 : XNOR2_X1 port map( A => n6, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_84 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_84;

architecture SYN_BEHAVIORAL of FA_84 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n5);
   U1 : XNOR2_X1 port map( A => n5, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_80 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_80;

architecture SYN_BEHAVIORAL of FA_80 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n5);
   U1 : XNOR2_X1 port map( A => n5, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_76 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_76;

architecture SYN_BEHAVIORAL of FA_76 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n5);
   U1 : XNOR2_X1 port map( A => n5, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_72 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_72;

architecture SYN_BEHAVIORAL of FA_72 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n5);
   U1 : XNOR2_X1 port map( A => n5, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_68 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_68;

architecture SYN_BEHAVIORAL of FA_68 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n5);
   U1 : XNOR2_X1 port map( A => n5, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_64 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_64;

architecture SYN_BEHAVIORAL of FA_64 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n5);
   U1 : XNOR2_X1 port map( A => n5, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_61 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_61;

architecture SYN_BEHAVIORAL of FA_61 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n5);
   U1 : XNOR2_X1 port map( A => n5, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_57 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_57;

architecture SYN_BEHAVIORAL of FA_57 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n5);
   U1 : XNOR2_X1 port map( A => n5, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_53 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_53;

architecture SYN_BEHAVIORAL of FA_53 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n5);
   U1 : XNOR2_X1 port map( A => n5, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_49 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_49;

architecture SYN_BEHAVIORAL of FA_49 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n5);
   U1 : XNOR2_X1 port map( A => n5, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_45 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_45;

architecture SYN_BEHAVIORAL of FA_45 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n5);
   U1 : XNOR2_X1 port map( A => n5, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_41 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_41;

architecture SYN_BEHAVIORAL of FA_41 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n5);
   U1 : XNOR2_X1 port map( A => n5, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_29 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_29;

architecture SYN_BEHAVIORAL of FA_29 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n5);
   U1 : XNOR2_X1 port map( A => n5, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_25 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_25;

architecture SYN_BEHAVIORAL of FA_25 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n5);
   U1 : XNOR2_X1 port map( A => n5, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_21 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_21;

architecture SYN_BEHAVIORAL of FA_21 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n5);
   U1 : XNOR2_X1 port map( A => n5, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_17 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_17;

architecture SYN_BEHAVIORAL of FA_17 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n5);
   U1 : XNOR2_X1 port map( A => n5, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_13 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_13;

architecture SYN_BEHAVIORAL of FA_13 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n5);
   U1 : XNOR2_X1 port map( A => n5, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_9 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_9;

architecture SYN_BEHAVIORAL of FA_9 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n5);
   U1 : XNOR2_X1 port map( A => n5, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_5 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_5;

architecture SYN_BEHAVIORAL of FA_5 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n5);
   U2 : XNOR2_X1 port map( A => Ci, B => n5, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_1 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1;

architecture SYN_BEHAVIORAL of FA_1 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n5);
   U2 : XNOR2_X1 port map( A => Ci, B => n5, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity mux21_SIZE4_13 is

   port( IN0, IN1 : in std_logic_vector (3 downto 0);  CTRL : in std_logic;  
         OUT1 : out std_logic_vector (3 downto 0));

end mux21_SIZE4_13;

architecture SYN_Bhe of mux21_SIZE4_13 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => IN0(3), B => IN1(3), S => CTRL, Z => OUT1(3));
   U2 : MUX2_X1 port map( A => IN0(2), B => IN1(2), S => CTRL, Z => OUT1(2));
   U3 : MUX2_X1 port map( A => IN0(1), B => IN1(1), S => CTRL, Z => OUT1(1));
   U4 : MUX2_X1 port map( A => IN0(0), B => IN1(0), S => CTRL, Z => OUT1(0));

end SYN_Bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity mux21_SIZE4_12 is

   port( IN0, IN1 : in std_logic_vector (3 downto 0);  CTRL : in std_logic;  
         OUT1 : out std_logic_vector (3 downto 0));

end mux21_SIZE4_12;

architecture SYN_Bhe of mux21_SIZE4_12 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => IN0(3), B => IN1(3), S => CTRL, Z => OUT1(3));
   U2 : MUX2_X1 port map( A => IN0(2), B => IN1(2), S => CTRL, Z => OUT1(2));
   U3 : MUX2_X1 port map( A => IN0(1), B => IN1(1), S => CTRL, Z => OUT1(1));
   U4 : MUX2_X1 port map( A => IN0(0), B => IN1(0), S => CTRL, Z => OUT1(0));

end SYN_Bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity mux21_SIZE4_11 is

   port( IN0, IN1 : in std_logic_vector (3 downto 0);  CTRL : in std_logic;  
         OUT1 : out std_logic_vector (3 downto 0));

end mux21_SIZE4_11;

architecture SYN_Bhe of mux21_SIZE4_11 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => IN0(3), B => IN1(3), S => CTRL, Z => OUT1(3));
   U2 : MUX2_X1 port map( A => IN0(2), B => IN1(2), S => CTRL, Z => OUT1(2));
   U3 : MUX2_X1 port map( A => IN0(1), B => IN1(1), S => CTRL, Z => OUT1(1));
   U4 : MUX2_X1 port map( A => IN0(0), B => IN1(0), S => CTRL, Z => OUT1(0));

end SYN_Bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity mux21_SIZE4_10 is

   port( IN0, IN1 : in std_logic_vector (3 downto 0);  CTRL : in std_logic;  
         OUT1 : out std_logic_vector (3 downto 0));

end mux21_SIZE4_10;

architecture SYN_Bhe of mux21_SIZE4_10 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => IN0(3), B => IN1(3), S => CTRL, Z => OUT1(3));
   U2 : MUX2_X1 port map( A => IN0(2), B => IN1(2), S => CTRL, Z => OUT1(2));
   U3 : MUX2_X1 port map( A => IN0(1), B => IN1(1), S => CTRL, Z => OUT1(1));
   U4 : MUX2_X1 port map( A => IN0(0), B => IN1(0), S => CTRL, Z => OUT1(0));

end SYN_Bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity mux21_SIZE4_9 is

   port( IN0, IN1 : in std_logic_vector (3 downto 0);  CTRL : in std_logic;  
         OUT1 : out std_logic_vector (3 downto 0));

end mux21_SIZE4_9;

architecture SYN_Bhe of mux21_SIZE4_9 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => IN0(3), B => IN1(3), S => CTRL, Z => OUT1(3));
   U3 : MUX2_X1 port map( A => IN0(1), B => IN1(1), S => CTRL, Z => OUT1(1));
   U4 : MUX2_X1 port map( A => IN0(0), B => IN1(0), S => CTRL, Z => OUT1(0));
   U2 : MUX2_X1 port map( A => IN0(2), B => IN1(2), S => CTRL, Z => OUT1(2));

end SYN_Bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity mux21_SIZE4_8 is

   port( IN0, IN1 : in std_logic_vector (3 downto 0);  CTRL : in std_logic;  
         OUT1 : out std_logic_vector (3 downto 0));

end mux21_SIZE4_8;

architecture SYN_Bhe of mux21_SIZE4_8 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => IN0(3), B => IN1(3), S => CTRL, Z => OUT1(3));
   U2 : MUX2_X1 port map( A => IN0(2), B => IN1(2), S => CTRL, Z => OUT1(2));
   U3 : MUX2_X1 port map( A => IN0(1), B => IN1(1), S => CTRL, Z => OUT1(1));
   U4 : MUX2_X1 port map( A => IN0(0), B => IN1(0), S => CTRL, Z => OUT1(0));

end SYN_Bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity mux21_SIZE4_7 is

   port( IN0, IN1 : in std_logic_vector (3 downto 0);  CTRL : in std_logic;  
         OUT1 : out std_logic_vector (3 downto 0));

end mux21_SIZE4_7;

architecture SYN_Bhe of mux21_SIZE4_7 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => IN0(3), B => IN1(3), S => CTRL, Z => OUT1(3));
   U2 : MUX2_X1 port map( A => IN0(2), B => IN1(2), S => CTRL, Z => OUT1(2));
   U3 : MUX2_X1 port map( A => IN0(1), B => IN1(1), S => CTRL, Z => OUT1(1));
   U4 : MUX2_X1 port map( A => IN0(0), B => IN1(0), S => CTRL, Z => OUT1(0));

end SYN_Bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity mux21_SIZE4_6 is

   port( IN0, IN1 : in std_logic_vector (3 downto 0);  CTRL : in std_logic;  
         OUT1 : out std_logic_vector (3 downto 0));

end mux21_SIZE4_6;

architecture SYN_Bhe of mux21_SIZE4_6 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => IN0(3), B => IN1(3), S => CTRL, Z => OUT1(3));
   U2 : MUX2_X1 port map( A => IN0(2), B => IN1(2), S => CTRL, Z => OUT1(2));
   U3 : MUX2_X1 port map( A => IN0(1), B => IN1(1), S => CTRL, Z => OUT1(1));
   U4 : MUX2_X1 port map( A => IN0(0), B => IN1(0), S => CTRL, Z => OUT1(0));

end SYN_Bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity mux21_SIZE4_5 is

   port( IN0, IN1 : in std_logic_vector (3 downto 0);  CTRL : in std_logic;  
         OUT1 : out std_logic_vector (3 downto 0));

end mux21_SIZE4_5;

architecture SYN_Bhe of mux21_SIZE4_5 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => IN0(3), B => IN1(3), S => CTRL, Z => OUT1(3));
   U2 : MUX2_X1 port map( A => IN0(2), B => IN1(2), S => CTRL, Z => OUT1(2));
   U3 : MUX2_X1 port map( A => IN0(1), B => IN1(1), S => CTRL, Z => OUT1(1));
   U4 : MUX2_X1 port map( A => IN0(0), B => IN1(0), S => CTRL, Z => OUT1(0));

end SYN_Bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity mux21_SIZE4_4 is

   port( IN0, IN1 : in std_logic_vector (3 downto 0);  CTRL : in std_logic;  
         OUT1 : out std_logic_vector (3 downto 0));

end mux21_SIZE4_4;

architecture SYN_Bhe of mux21_SIZE4_4 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => IN0(3), B => IN1(3), S => CTRL, Z => OUT1(3));
   U2 : MUX2_X1 port map( A => IN0(2), B => IN1(2), S => CTRL, Z => OUT1(2));
   U3 : MUX2_X1 port map( A => IN0(1), B => IN1(1), S => CTRL, Z => OUT1(1));
   U4 : MUX2_X1 port map( A => IN0(0), B => IN1(0), S => CTRL, Z => OUT1(0));

end SYN_Bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity mux21_SIZE4_3 is

   port( IN0, IN1 : in std_logic_vector (3 downto 0);  CTRL : in std_logic;  
         OUT1 : out std_logic_vector (3 downto 0));

end mux21_SIZE4_3;

architecture SYN_Bhe of mux21_SIZE4_3 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => IN0(3), B => IN1(3), S => CTRL, Z => OUT1(3));
   U2 : MUX2_X1 port map( A => IN0(2), B => IN1(2), S => CTRL, Z => OUT1(2));
   U3 : MUX2_X1 port map( A => IN0(1), B => IN1(1), S => CTRL, Z => OUT1(1));
   U4 : MUX2_X1 port map( A => IN0(0), B => IN1(0), S => CTRL, Z => OUT1(0));

end SYN_Bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity mux21_SIZE4_2 is

   port( IN0, IN1 : in std_logic_vector (3 downto 0);  CTRL : in std_logic;  
         OUT1 : out std_logic_vector (3 downto 0));

end mux21_SIZE4_2;

architecture SYN_Bhe of mux21_SIZE4_2 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => IN0(3), B => IN1(3), S => CTRL, Z => OUT1(3));
   U2 : MUX2_X1 port map( A => IN0(2), B => IN1(2), S => CTRL, Z => OUT1(2));
   U3 : MUX2_X1 port map( A => IN0(0), B => IN1(0), S => CTRL, Z => OUT1(0));
   U4 : MUX2_X1 port map( A => IN0(1), B => IN1(1), S => CTRL, Z => OUT1(1));

end SYN_Bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity mux21_SIZE4_1 is

   port( IN0, IN1 : in std_logic_vector (3 downto 0);  CTRL : in std_logic;  
         OUT1 : out std_logic_vector (3 downto 0));

end mux21_SIZE4_1;

architecture SYN_Bhe of mux21_SIZE4_1 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : MUX2_X1 port map( A => IN0(2), B => IN1(2), S => CTRL, Z => OUT1(2));
   U1 : MUX2_X1 port map( A => IN0(0), B => IN1(0), S => CTRL, Z => OUT1(0));
   U3 : MUX2_X1 port map( A => IN0(3), B => IN1(3), S => CTRL, Z => OUT1(3));
   U4 : MUX2_X1 port map( A => IN0(1), B => IN1(1), S => CTRL, Z => OUT1(1));

end SYN_Bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity RCA_N4_12 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_12;

architecture SYN_STRUCTURAL of RCA_N4_12 is

   component FA_45
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_46
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_47
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_48
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal n2, CTMP_3_port, CTMP_2_port, n1, net684402 : std_logic;

begin
   
   n2 <= '0';
   FAI_1 : FA_48 port map( A => A(0), B => B(0), Ci => n2, S => S(0), Co => n1)
                           ;
   FAI_2 : FA_47 port map( A => A(1), B => B(1), Ci => n1, S => S(1), Co => 
                           CTMP_2_port);
   FAI_3 : FA_46 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_45 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => net684402);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity RCA_N4_10 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_10;

architecture SYN_STRUCTURAL of RCA_N4_10 is

   component FA_37
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_38
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_39
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_40
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal n2, CTMP_3_port, CTMP_2_port, CTMP_1_port, net684401 : std_logic;

begin
   
   n2 <= '0';
   FAI_1 : FA_40 port map( A => A(0), B => B(0), Ci => n2, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_39 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_38 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_37 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => net684401);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity RCA_N4_9 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_9;

architecture SYN_STRUCTURAL of RCA_N4_9 is

   component FA_33
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_34
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_35
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_36
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal n2, CTMP_3_port, CTMP_2_port, CTMP_1_port, net684400 : std_logic;

begin
   
   n2 <= '1';
   FAI_1 : FA_36 port map( A => A(0), B => B(0), Ci => n2, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_35 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_34 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_33 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => net684400);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity RCA_N4_23 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_23;

architecture SYN_STRUCTURAL of RCA_N4_23 is

   component FA_92
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_93
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_94
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_95
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal n1, CTMP_3_port, CTMP_2_port, CTMP_1_port, net684399 : std_logic;

begin
   
   n1 <= '0';
   FAI_1 : FA_95 port map( A => A(0), B => B(0), Ci => n1, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_94 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_93 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_92 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => net684399);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity RCA_N4_21 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_21;

architecture SYN_STRUCTURAL of RCA_N4_21 is

   component FA_84
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_85
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_86
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_87
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal n1, CTMP_3_port, CTMP_2_port, CTMP_1_port, net684398 : std_logic;

begin
   
   n1 <= '0';
   FAI_1 : FA_87 port map( A => A(0), B => B(0), Ci => n1, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_86 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_85 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_84 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => net684398);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity RCA_N4_19 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_19;

architecture SYN_STRUCTURAL of RCA_N4_19 is

   component FA_76
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_77
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_78
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_79
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal n1, CTMP_3_port, CTMP_2_port, CTMP_1_port, net684397 : std_logic;

begin
   
   n1 <= '0';
   FAI_1 : FA_79 port map( A => A(0), B => B(0), Ci => n1, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_78 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_77 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_76 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => net684397);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity RCA_N4_17 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_17;

architecture SYN_STRUCTURAL of RCA_N4_17 is

   component FA_68
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_69
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_70
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_71
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal n1, CTMP_3_port, CTMP_2_port, CTMP_1_port, net684396 : std_logic;

begin
   
   n1 <= '0';
   FAI_1 : FA_71 port map( A => A(0), B => B(0), Ci => n1, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_70 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_69 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_68 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => net684396);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity RCA_N4_14 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_14;

architecture SYN_STRUCTURAL of RCA_N4_14 is

   component FA_53
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_54
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_55
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_56
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal n1, CTMP_3_port, CTMP_2_port, CTMP_1_port, net684395 : std_logic;

begin
   
   n1 <= '0';
   FAI_1 : FA_56 port map( A => A(0), B => B(0), Ci => n1, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_55 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_54 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_53 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => net684395);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity RCA_N4_8 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_8;

architecture SYN_STRUCTURAL of RCA_N4_8 is

   component FA_29
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_30
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_31
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_32
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal n1, CTMP_3_port, CTMP_2_port, CTMP_1_port, net684394 : std_logic;

begin
   
   n1 <= '0';
   FAI_1 : FA_32 port map( A => A(0), B => B(0), Ci => n1, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_31 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_30 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_29 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => net684394);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity RCA_N4_6 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_6;

architecture SYN_STRUCTURAL of RCA_N4_6 is

   component FA_21
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_22
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_23
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_24
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal n1, CTMP_3_port, CTMP_2_port, CTMP_1_port, net684393 : std_logic;

begin
   
   n1 <= '0';
   FAI_1 : FA_24 port map( A => A(0), B => B(0), Ci => n1, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_23 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_22 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_21 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => net684393);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity RCA_N4_4 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_4;

architecture SYN_STRUCTURAL of RCA_N4_4 is

   component FA_13
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_14
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_15
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_16
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal n1, CTMP_3_port, CTMP_2_port, CTMP_1_port, net684392 : std_logic;

begin
   
   n1 <= '0';
   FAI_1 : FA_16 port map( A => A(0), B => B(0), Ci => n1, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_15 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_14 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_13 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => net684392);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity RCA_N4_2 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_2;

architecture SYN_STRUCTURAL of RCA_N4_2 is

   component FA_5
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_6
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_7
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_8
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal n1, CTMP_3_port, CTMP_2_port, CTMP_1_port, net684391 : std_logic;

begin
   
   n1 <= '0';
   FAI_1 : FA_8 port map( A => A(0), B => B(0), Ci => n1, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_7 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_6 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_5 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => net684391);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity RCA_N4_28 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_28;

architecture SYN_STRUCTURAL of RCA_N4_28 is

   component FA_112
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_113
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_114
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_115
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal n1, CTMP_3_port, CTMP_2_port, CTMP_1_port, net684390 : std_logic;

begin
   
   n1 <= '1';
   FAI_1 : FA_115 port map( A => A(0), B => B(0), Ci => n1, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_114 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_113 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_112 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => net684390);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity RCA_N4_26 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_26;

architecture SYN_STRUCTURAL of RCA_N4_26 is

   component FA_104
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_105
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_106
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_107
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal n1, CTMP_3_port, CTMP_2_port, CTMP_1_port, net684389 : std_logic;

begin
   
   n1 <= '1';
   FAI_1 : FA_107 port map( A => A(0), B => B(0), Ci => n1, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_106 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_105 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_104 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => net684389);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity RCA_N4_22 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_22;

architecture SYN_STRUCTURAL of RCA_N4_22 is

   component FA_88
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_89
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_90
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_91
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal n1, CTMP_3_port, CTMP_2_port, CTMP_1_port, net684388 : std_logic;

begin
   
   n1 <= '1';
   FAI_1 : FA_91 port map( A => A(0), B => B(0), Ci => n1, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_90 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_89 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_88 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => net684388);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity RCA_N4_20 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_20;

architecture SYN_STRUCTURAL of RCA_N4_20 is

   component FA_80
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_81
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_82
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_83
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal n1, CTMP_3_port, CTMP_2_port, CTMP_1_port, net684387 : std_logic;

begin
   
   n1 <= '1';
   FAI_1 : FA_83 port map( A => A(0), B => B(0), Ci => n1, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_82 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_81 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_80 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => net684387);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity RCA_N4_18 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_18;

architecture SYN_STRUCTURAL of RCA_N4_18 is

   component FA_72
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_73
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_74
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_75
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal n1, CTMP_3_port, CTMP_2_port, CTMP_1_port, net684386 : std_logic;

begin
   
   n1 <= '1';
   FAI_1 : FA_75 port map( A => A(0), B => B(0), Ci => n1, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_74 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_73 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_72 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => net684386);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity RCA_N4_16 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_16;

architecture SYN_STRUCTURAL of RCA_N4_16 is

   component FA_64
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_65
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_66
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_67
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal n1, CTMP_3_port, CTMP_2_port, CTMP_1_port, net684385 : std_logic;

begin
   
   n1 <= '1';
   FAI_1 : FA_67 port map( A => A(0), B => B(0), Ci => n1, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_66 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_65 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_64 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => net684385);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity RCA_N4_15 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_15;

architecture SYN_STRUCTURAL of RCA_N4_15 is

   component FA_57
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_58
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_59
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_60
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal n1, CTMP_3_port, CTMP_2_port, CTMP_1_port, net684384 : std_logic;

begin
   
   n1 <= '1';
   FAI_1 : FA_60 port map( A => A(0), B => B(0), Ci => n1, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_59 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_58 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_57 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => net684384);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity RCA_N4_13 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_13;

architecture SYN_STRUCTURAL of RCA_N4_13 is

   component FA_49
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_50
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_51
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_52
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal n1, CTMP_3_port, CTMP_2_port, CTMP_1_port, net684383 : std_logic;

begin
   
   n1 <= '1';
   FAI_1 : FA_52 port map( A => A(0), B => B(0), Ci => n1, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_51 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_50 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_49 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => net684383);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity RCA_N4_11 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_11;

architecture SYN_STRUCTURAL of RCA_N4_11 is

   component FA_41
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_42
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_43
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_44
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal n1, CTMP_3_port, CTMP_2_port, CTMP_1_port, net684382 : std_logic;

begin
   
   n1 <= '1';
   FAI_1 : FA_44 port map( A => A(0), B => B(0), Ci => n1, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_43 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_42 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_41 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => net684382);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity RCA_N4_7 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_7;

architecture SYN_STRUCTURAL of RCA_N4_7 is

   component FA_25
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_26
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_27
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_28
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal n1, CTMP_3_port, CTMP_2_port, CTMP_1_port, net684381 : std_logic;

begin
   
   n1 <= '1';
   FAI_1 : FA_28 port map( A => A(0), B => B(0), Ci => n1, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_27 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_26 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_25 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => net684381);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity RCA_N4_5 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_5;

architecture SYN_STRUCTURAL of RCA_N4_5 is

   component FA_17
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_18
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_19
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_20
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal n1, CTMP_3_port, CTMP_2_port, CTMP_1_port, net684380 : std_logic;

begin
   
   n1 <= '1';
   FAI_1 : FA_20 port map( A => A(0), B => B(0), Ci => n1, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_19 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_18 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_17 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => net684380);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity RCA_N4_3 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_3;

architecture SYN_STRUCTURAL of RCA_N4_3 is

   component FA_9
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_10
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_11
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_12
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal n1, CTMP_3_port, CTMP_2_port, CTMP_1_port, net684379 : std_logic;

begin
   
   n1 <= '1';
   FAI_1 : FA_12 port map( A => A(0), B => B(0), Ci => n1, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_11 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_10 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_9 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => net684379);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity RCA_N4_1 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_1;

architecture SYN_STRUCTURAL of RCA_N4_1 is

   component FA_1
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_2
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_3
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_4
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal n1, CTMP_3_port, CTMP_2_port, CTMP_1_port, net684378 : std_logic;

begin
   
   n1 <= '1';
   FAI_1 : FA_4 port map( A => A(0), B => B(0), Ci => n1, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_3 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_2 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_1 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => net684378);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity carry_sel_gen_N4_6 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end carry_sel_gen_N4_6;

architecture SYN_STRUCTURAL of carry_sel_gen_N4_6 is

   component mux21_SIZE4_6
      port( IN0, IN1 : in std_logic_vector (3 downto 0);  CTRL : in std_logic; 
            OUT1 : out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_N4_11
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_12
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, nocarry_sum_to_mux_3_port, 
      nocarry_sum_to_mux_2_port, nocarry_sum_to_mux_1_port, 
      nocarry_sum_to_mux_0_port, carry_sum_to_mux_3_port, 
      carry_sum_to_mux_2_port, carry_sum_to_mux_1_port, carry_sum_to_mux_0_port
      , net684376, net684377 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   rca_nocarry : RCA_N4_12 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           nocarry_sum_to_mux_3_port, S(2) => 
                           nocarry_sum_to_mux_2_port, S(1) => 
                           nocarry_sum_to_mux_1_port, S(0) => 
                           nocarry_sum_to_mux_0_port, Co => net684377);
   rca_carry : RCA_N4_11 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           carry_sum_to_mux_3_port, S(2) => 
                           carry_sum_to_mux_2_port, S(1) => 
                           carry_sum_to_mux_1_port, S(0) => 
                           carry_sum_to_mux_0_port, Co => net684376);
   outmux : mux21_SIZE4_6 port map( IN0(3) => nocarry_sum_to_mux_3_port, IN0(2)
                           => nocarry_sum_to_mux_2_port, IN0(1) => 
                           nocarry_sum_to_mux_1_port, IN0(0) => 
                           nocarry_sum_to_mux_0_port, IN1(3) => 
                           carry_sum_to_mux_3_port, IN1(2) => 
                           carry_sum_to_mux_2_port, IN1(1) => 
                           carry_sum_to_mux_1_port, IN1(0) => 
                           carry_sum_to_mux_0_port, CTRL => Ci, OUT1(3) => S(3)
                           , OUT1(2) => S(2), OUT1(1) => S(1), OUT1(0) => S(0))
                           ;

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity carry_sel_gen_N4_5 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end carry_sel_gen_N4_5;

architecture SYN_STRUCTURAL of carry_sel_gen_N4_5 is

   component mux21_SIZE4_5
      port( IN0, IN1 : in std_logic_vector (3 downto 0);  CTRL : in std_logic; 
            OUT1 : out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_N4_9
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_10
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, nocarry_sum_to_mux_3_port, 
      nocarry_sum_to_mux_2_port, nocarry_sum_to_mux_1_port, 
      nocarry_sum_to_mux_0_port, carry_sum_to_mux_3_port, 
      carry_sum_to_mux_2_port, carry_sum_to_mux_1_port, carry_sum_to_mux_0_port
      , net684374, net684375 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   rca_nocarry : RCA_N4_10 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           nocarry_sum_to_mux_3_port, S(2) => 
                           nocarry_sum_to_mux_2_port, S(1) => 
                           nocarry_sum_to_mux_1_port, S(0) => 
                           nocarry_sum_to_mux_0_port, Co => net684375);
   rca_carry : RCA_N4_9 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           carry_sum_to_mux_3_port, S(2) => 
                           carry_sum_to_mux_2_port, S(1) => 
                           carry_sum_to_mux_1_port, S(0) => 
                           carry_sum_to_mux_0_port, Co => net684374);
   outmux : mux21_SIZE4_5 port map( IN0(3) => nocarry_sum_to_mux_3_port, IN0(2)
                           => nocarry_sum_to_mux_2_port, IN0(1) => 
                           nocarry_sum_to_mux_1_port, IN0(0) => 
                           nocarry_sum_to_mux_0_port, IN1(3) => 
                           carry_sum_to_mux_3_port, IN1(2) => 
                           carry_sum_to_mux_2_port, IN1(1) => 
                           carry_sum_to_mux_1_port, IN1(0) => 
                           carry_sum_to_mux_0_port, CTRL => Ci, OUT1(3) => S(3)
                           , OUT1(2) => S(2), OUT1(1) => S(1), OUT1(0) => S(0))
                           ;

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity carry_sel_gen_N4_4 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end carry_sel_gen_N4_4;

architecture SYN_STRUCTURAL of carry_sel_gen_N4_4 is

   component mux21_SIZE4_4
      port( IN0, IN1 : in std_logic_vector (3 downto 0);  CTRL : in std_logic; 
            OUT1 : out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_N4_7
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_8
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, nocarry_sum_to_mux_3_port, 
      nocarry_sum_to_mux_2_port, nocarry_sum_to_mux_1_port, 
      nocarry_sum_to_mux_0_port, carry_sum_to_mux_3_port, 
      carry_sum_to_mux_2_port, carry_sum_to_mux_1_port, carry_sum_to_mux_0_port
      , net684372, net684373 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   rca_nocarry : RCA_N4_8 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           nocarry_sum_to_mux_3_port, S(2) => 
                           nocarry_sum_to_mux_2_port, S(1) => 
                           nocarry_sum_to_mux_1_port, S(0) => 
                           nocarry_sum_to_mux_0_port, Co => net684373);
   rca_carry : RCA_N4_7 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           carry_sum_to_mux_3_port, S(2) => 
                           carry_sum_to_mux_2_port, S(1) => 
                           carry_sum_to_mux_1_port, S(0) => 
                           carry_sum_to_mux_0_port, Co => net684372);
   outmux : mux21_SIZE4_4 port map( IN0(3) => nocarry_sum_to_mux_3_port, IN0(2)
                           => nocarry_sum_to_mux_2_port, IN0(1) => 
                           nocarry_sum_to_mux_1_port, IN0(0) => 
                           nocarry_sum_to_mux_0_port, IN1(3) => 
                           carry_sum_to_mux_3_port, IN1(2) => 
                           carry_sum_to_mux_2_port, IN1(1) => 
                           carry_sum_to_mux_1_port, IN1(0) => 
                           carry_sum_to_mux_0_port, CTRL => Ci, OUT1(3) => S(3)
                           , OUT1(2) => S(2), OUT1(1) => S(1), OUT1(0) => S(0))
                           ;

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity carry_sel_gen_N4_10 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end carry_sel_gen_N4_10;

architecture SYN_STRUCTURAL of carry_sel_gen_N4_10 is

   component mux21_SIZE4_10
      port( IN0, IN1 : in std_logic_vector (3 downto 0);  CTRL : in std_logic; 
            OUT1 : out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_N4_20
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_21
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, nocarry_sum_to_mux_3_port, 
      nocarry_sum_to_mux_2_port, nocarry_sum_to_mux_1_port, 
      nocarry_sum_to_mux_0_port, carry_sum_to_mux_3_port, 
      carry_sum_to_mux_2_port, carry_sum_to_mux_1_port, carry_sum_to_mux_0_port
      , net684370, net684371 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   rca_nocarry : RCA_N4_21 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           nocarry_sum_to_mux_3_port, S(2) => 
                           nocarry_sum_to_mux_2_port, S(1) => 
                           nocarry_sum_to_mux_1_port, S(0) => 
                           nocarry_sum_to_mux_0_port, Co => net684371);
   rca_carry : RCA_N4_20 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           carry_sum_to_mux_3_port, S(2) => 
                           carry_sum_to_mux_2_port, S(1) => 
                           carry_sum_to_mux_1_port, S(0) => 
                           carry_sum_to_mux_0_port, Co => net684370);
   outmux : mux21_SIZE4_10 port map( IN0(3) => nocarry_sum_to_mux_3_port, 
                           IN0(2) => nocarry_sum_to_mux_2_port, IN0(1) => 
                           nocarry_sum_to_mux_1_port, IN0(0) => 
                           nocarry_sum_to_mux_0_port, IN1(3) => 
                           carry_sum_to_mux_3_port, IN1(2) => 
                           carry_sum_to_mux_2_port, IN1(1) => 
                           carry_sum_to_mux_1_port, IN1(0) => 
                           carry_sum_to_mux_0_port, CTRL => Ci, OUT1(3) => S(3)
                           , OUT1(2) => S(2), OUT1(1) => S(1), OUT1(0) => S(0))
                           ;

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity carry_sel_gen_N4_9 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end carry_sel_gen_N4_9;

architecture SYN_STRUCTURAL of carry_sel_gen_N4_9 is

   component mux21_SIZE4_9
      port( IN0, IN1 : in std_logic_vector (3 downto 0);  CTRL : in std_logic; 
            OUT1 : out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_N4_18
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_19
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, nocarry_sum_to_mux_3_port, 
      nocarry_sum_to_mux_2_port, nocarry_sum_to_mux_1_port, 
      nocarry_sum_to_mux_0_port, carry_sum_to_mux_3_port, 
      carry_sum_to_mux_2_port, carry_sum_to_mux_1_port, carry_sum_to_mux_0_port
      , net684368, net684369 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   rca_nocarry : RCA_N4_19 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           nocarry_sum_to_mux_3_port, S(2) => 
                           nocarry_sum_to_mux_2_port, S(1) => 
                           nocarry_sum_to_mux_1_port, S(0) => 
                           nocarry_sum_to_mux_0_port, Co => net684369);
   rca_carry : RCA_N4_18 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           carry_sum_to_mux_3_port, S(2) => 
                           carry_sum_to_mux_2_port, S(1) => 
                           carry_sum_to_mux_1_port, S(0) => 
                           carry_sum_to_mux_0_port, Co => net684368);
   outmux : mux21_SIZE4_9 port map( IN0(3) => nocarry_sum_to_mux_3_port, IN0(2)
                           => nocarry_sum_to_mux_2_port, IN0(1) => 
                           nocarry_sum_to_mux_1_port, IN0(0) => 
                           nocarry_sum_to_mux_0_port, IN1(3) => 
                           carry_sum_to_mux_3_port, IN1(2) => 
                           carry_sum_to_mux_2_port, IN1(1) => 
                           carry_sum_to_mux_1_port, IN1(0) => 
                           carry_sum_to_mux_0_port, CTRL => Ci, OUT1(3) => S(3)
                           , OUT1(2) => S(2), OUT1(1) => S(1), OUT1(0) => S(0))
                           ;

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity carry_sel_gen_N4_8 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end carry_sel_gen_N4_8;

architecture SYN_STRUCTURAL of carry_sel_gen_N4_8 is

   component mux21_SIZE4_8
      port( IN0, IN1 : in std_logic_vector (3 downto 0);  CTRL : in std_logic; 
            OUT1 : out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_N4_16
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_17
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, nocarry_sum_to_mux_3_port, 
      nocarry_sum_to_mux_2_port, nocarry_sum_to_mux_1_port, 
      nocarry_sum_to_mux_0_port, carry_sum_to_mux_3_port, 
      carry_sum_to_mux_2_port, carry_sum_to_mux_1_port, carry_sum_to_mux_0_port
      , net684366, net684367 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   rca_nocarry : RCA_N4_17 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           nocarry_sum_to_mux_3_port, S(2) => 
                           nocarry_sum_to_mux_2_port, S(1) => 
                           nocarry_sum_to_mux_1_port, S(0) => 
                           nocarry_sum_to_mux_0_port, Co => net684367);
   rca_carry : RCA_N4_16 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           carry_sum_to_mux_3_port, S(2) => 
                           carry_sum_to_mux_2_port, S(1) => 
                           carry_sum_to_mux_1_port, S(0) => 
                           carry_sum_to_mux_0_port, Co => net684366);
   outmux : mux21_SIZE4_8 port map( IN0(3) => nocarry_sum_to_mux_3_port, IN0(2)
                           => nocarry_sum_to_mux_2_port, IN0(1) => 
                           nocarry_sum_to_mux_1_port, IN0(0) => 
                           nocarry_sum_to_mux_0_port, IN1(3) => 
                           carry_sum_to_mux_3_port, IN1(2) => 
                           carry_sum_to_mux_2_port, IN1(1) => 
                           carry_sum_to_mux_1_port, IN1(0) => 
                           carry_sum_to_mux_0_port, CTRL => Ci, OUT1(3) => S(3)
                           , OUT1(2) => S(2), OUT1(1) => S(1), OUT1(0) => S(0))
                           ;

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity carry_sel_gen_N4_7 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end carry_sel_gen_N4_7;

architecture SYN_STRUCTURAL of carry_sel_gen_N4_7 is

   component mux21_SIZE4_7
      port( IN0, IN1 : in std_logic_vector (3 downto 0);  CTRL : in std_logic; 
            OUT1 : out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_N4_13
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_14
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, nocarry_sum_to_mux_3_port, 
      nocarry_sum_to_mux_2_port, nocarry_sum_to_mux_1_port, 
      nocarry_sum_to_mux_0_port, carry_sum_to_mux_3_port, 
      carry_sum_to_mux_2_port, carry_sum_to_mux_1_port, carry_sum_to_mux_0_port
      , net684364, net684365 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   rca_nocarry : RCA_N4_14 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           nocarry_sum_to_mux_3_port, S(2) => 
                           nocarry_sum_to_mux_2_port, S(1) => 
                           nocarry_sum_to_mux_1_port, S(0) => 
                           nocarry_sum_to_mux_0_port, Co => net684365);
   rca_carry : RCA_N4_13 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           carry_sum_to_mux_3_port, S(2) => 
                           carry_sum_to_mux_2_port, S(1) => 
                           carry_sum_to_mux_1_port, S(0) => 
                           carry_sum_to_mux_0_port, Co => net684364);
   outmux : mux21_SIZE4_7 port map( IN0(3) => nocarry_sum_to_mux_3_port, IN0(2)
                           => nocarry_sum_to_mux_2_port, IN0(1) => 
                           nocarry_sum_to_mux_1_port, IN0(0) => 
                           nocarry_sum_to_mux_0_port, IN1(3) => 
                           carry_sum_to_mux_3_port, IN1(2) => 
                           carry_sum_to_mux_2_port, IN1(1) => 
                           carry_sum_to_mux_1_port, IN1(0) => 
                           carry_sum_to_mux_0_port, CTRL => Ci, OUT1(3) => S(3)
                           , OUT1(2) => S(2), OUT1(1) => S(1), OUT1(0) => S(0))
                           ;

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity carry_sel_gen_N4_3 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end carry_sel_gen_N4_3;

architecture SYN_STRUCTURAL of carry_sel_gen_N4_3 is

   component mux21_SIZE4_3
      port( IN0, IN1 : in std_logic_vector (3 downto 0);  CTRL : in std_logic; 
            OUT1 : out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_N4_5
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_6
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, nocarry_sum_to_mux_3_port, 
      nocarry_sum_to_mux_2_port, nocarry_sum_to_mux_1_port, 
      nocarry_sum_to_mux_0_port, carry_sum_to_mux_3_port, 
      carry_sum_to_mux_2_port, carry_sum_to_mux_1_port, carry_sum_to_mux_0_port
      , net684362, net684363 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   rca_nocarry : RCA_N4_6 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           nocarry_sum_to_mux_3_port, S(2) => 
                           nocarry_sum_to_mux_2_port, S(1) => 
                           nocarry_sum_to_mux_1_port, S(0) => 
                           nocarry_sum_to_mux_0_port, Co => net684363);
   rca_carry : RCA_N4_5 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           carry_sum_to_mux_3_port, S(2) => 
                           carry_sum_to_mux_2_port, S(1) => 
                           carry_sum_to_mux_1_port, S(0) => 
                           carry_sum_to_mux_0_port, Co => net684362);
   outmux : mux21_SIZE4_3 port map( IN0(3) => nocarry_sum_to_mux_3_port, IN0(2)
                           => nocarry_sum_to_mux_2_port, IN0(1) => 
                           nocarry_sum_to_mux_1_port, IN0(0) => 
                           nocarry_sum_to_mux_0_port, IN1(3) => 
                           carry_sum_to_mux_3_port, IN1(2) => 
                           carry_sum_to_mux_2_port, IN1(1) => 
                           carry_sum_to_mux_1_port, IN1(0) => 
                           carry_sum_to_mux_0_port, CTRL => Ci, OUT1(3) => S(3)
                           , OUT1(2) => S(2), OUT1(1) => S(1), OUT1(0) => S(0))
                           ;

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity carry_sel_gen_N4_2 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end carry_sel_gen_N4_2;

architecture SYN_STRUCTURAL of carry_sel_gen_N4_2 is

   component mux21_SIZE4_2
      port( IN0, IN1 : in std_logic_vector (3 downto 0);  CTRL : in std_logic; 
            OUT1 : out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_N4_3
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_4
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, nocarry_sum_to_mux_3_port, 
      nocarry_sum_to_mux_2_port, nocarry_sum_to_mux_1_port, 
      nocarry_sum_to_mux_0_port, carry_sum_to_mux_3_port, 
      carry_sum_to_mux_2_port, carry_sum_to_mux_1_port, carry_sum_to_mux_0_port
      , net684360, net684361 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   rca_nocarry : RCA_N4_4 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           nocarry_sum_to_mux_3_port, S(2) => 
                           nocarry_sum_to_mux_2_port, S(1) => 
                           nocarry_sum_to_mux_1_port, S(0) => 
                           nocarry_sum_to_mux_0_port, Co => net684361);
   rca_carry : RCA_N4_3 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           carry_sum_to_mux_3_port, S(2) => 
                           carry_sum_to_mux_2_port, S(1) => 
                           carry_sum_to_mux_1_port, S(0) => 
                           carry_sum_to_mux_0_port, Co => net684360);
   outmux : mux21_SIZE4_2 port map( IN0(3) => nocarry_sum_to_mux_3_port, IN0(2)
                           => nocarry_sum_to_mux_2_port, IN0(1) => 
                           nocarry_sum_to_mux_1_port, IN0(0) => 
                           nocarry_sum_to_mux_0_port, IN1(3) => 
                           carry_sum_to_mux_3_port, IN1(2) => 
                           carry_sum_to_mux_2_port, IN1(1) => 
                           carry_sum_to_mux_1_port, IN1(0) => 
                           carry_sum_to_mux_0_port, CTRL => Ci, OUT1(3) => S(3)
                           , OUT1(2) => S(2), OUT1(1) => S(1), OUT1(0) => S(0))
                           ;

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity carry_sel_gen_N4_1 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end carry_sel_gen_N4_1;

architecture SYN_STRUCTURAL of carry_sel_gen_N4_1 is

   component mux21_SIZE4_1
      port( IN0, IN1 : in std_logic_vector (3 downto 0);  CTRL : in std_logic; 
            OUT1 : out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_N4_1
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_2
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, nocarry_sum_to_mux_3_port, 
      nocarry_sum_to_mux_2_port, nocarry_sum_to_mux_1_port, 
      nocarry_sum_to_mux_0_port, carry_sum_to_mux_3_port, 
      carry_sum_to_mux_2_port, carry_sum_to_mux_1_port, carry_sum_to_mux_0_port
      , net684358, net684359 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   rca_nocarry : RCA_N4_2 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           nocarry_sum_to_mux_3_port, S(2) => 
                           nocarry_sum_to_mux_2_port, S(1) => 
                           nocarry_sum_to_mux_1_port, S(0) => 
                           nocarry_sum_to_mux_0_port, Co => net684359);
   rca_carry : RCA_N4_1 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           carry_sum_to_mux_3_port, S(2) => 
                           carry_sum_to_mux_2_port, S(1) => 
                           carry_sum_to_mux_1_port, S(0) => 
                           carry_sum_to_mux_0_port, Co => net684358);
   outmux : mux21_SIZE4_1 port map( IN0(3) => nocarry_sum_to_mux_3_port, IN0(2)
                           => nocarry_sum_to_mux_2_port, IN0(1) => 
                           nocarry_sum_to_mux_1_port, IN0(0) => 
                           nocarry_sum_to_mux_0_port, IN1(3) => 
                           carry_sum_to_mux_3_port, IN1(2) => 
                           carry_sum_to_mux_2_port, IN1(1) => 
                           carry_sum_to_mux_1_port, IN1(0) => 
                           carry_sum_to_mux_0_port, CTRL => Ci, OUT1(3) => S(3)
                           , OUT1(2) => S(2), OUT1(1) => S(1), OUT1(0) => S(0))
                           ;

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_20 is

   port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic);

end pg_20;

architecture SYN_beh of pg_20 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n6, n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => g, ZN => n7);
   U2 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);
   U3 : NAND2_X1 port map( A1 => p, A2 => g_prec, ZN => n6);
   U4 : NAND2_X1 port map( A1 => n6, A2 => n7, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_12 is

   port( p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic;  
         g_BAR : in std_logic);

end pg_12;

architecture SYN_beh of pg_12 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);
   U2 : NAND2_X1 port map( A1 => p, A2 => g_prec, ZN => n5);
   U3 : NAND2_X1 port map( A1 => n5, A2 => g_BAR, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_49 is

   port( g, p, g_prec, p_prec : in std_logic;  p_out, g_out_BAR : out std_logic
         );

end pg_49;

architecture SYN_beh of pg_49 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U2 : AOI21_X1 port map( B1 => g_prec, B2 => p, A => g, ZN => g_out_BAR);
   U1 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_47 is

   port( g, p, g_prec, p_prec : in std_logic;  p_out, g_out_BAR : out std_logic
         );

end pg_47;

architecture SYN_beh of pg_47 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U2 : AOI21_X1 port map( B1 => g_prec, B2 => p, A => g, ZN => g_out_BAR);
   U1 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_45 is

   port( g, p, g_prec, p_prec : in std_logic;  p_out, g_out_BAR : out std_logic
         );

end pg_45;

architecture SYN_beh of pg_45 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U2 : AOI21_X1 port map( B1 => g_prec, B2 => p, A => g, ZN => g_out_BAR);
   U1 : AND2_X1 port map( A1 => p_prec, A2 => p, ZN => p_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_34 is

   port( g, p, g_prec, p_prec : in std_logic;  p_out, g_out_BAR : out std_logic
         );

end pg_34;

architecture SYN_beh of pg_34 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U2 : AOI21_X1 port map( B1 => g_prec, B2 => p, A => g, ZN => g_out_BAR);
   U1 : AND2_X1 port map( A1 => p_prec, A2 => p, ZN => p_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_25 is

   port( g, p, g_prec, p_prec : in std_logic;  p_out, g_out_BAR : out std_logic
         );

end pg_25;

architecture SYN_beh of pg_25 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U2 : AOI21_X1 port map( B1 => p, B2 => g_prec, A => g, ZN => g_out_BAR);
   U1 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_23 is

   port( g, p, g_prec, p_prec : in std_logic;  p_out, g_out_BAR : out std_logic
         );

end pg_23;

architecture SYN_beh of pg_23 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U2 : AOI21_X1 port map( B1 => p, B2 => g_prec, A => g, ZN => g_out_BAR);
   U1 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_21 is

   port( g, p, g_prec, p_prec : in std_logic;  p_out, g_out_BAR : out std_logic
         );

end pg_21;

architecture SYN_beh of pg_21 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);
   U2 : AOI21_X1 port map( B1 => p, B2 => g_prec, A => g, ZN => g_out_BAR);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_19 is

   port( g, p, g_prec, p_prec : in std_logic;  p_out, g_out_BAR : out std_logic
         );

end pg_19;

architecture SYN_beh of pg_19 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p_prec, A2 => p, ZN => p_out);
   U2 : AOI21_X1 port map( B1 => g_prec, B2 => p, A => g, ZN => g_out_BAR);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_8 is

   port( g, p, g_prec, p_prec : in std_logic;  p_out, g_out_BAR : out std_logic
         );

end pg_8;

architecture SYN_beh of pg_8 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p_prec, A2 => p, ZN => p_out);
   U2 : AOI21_X1 port map( B1 => g_prec, B2 => p, A => g, ZN => g_out_BAR);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_36 is

   port( p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic;  
         g_BAR : in std_logic);

end pg_36;

architecture SYN_beh of pg_36 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U3 : NAND2_X1 port map( A1 => p, A2 => g_prec, ZN => n4);
   U2 : NAND2_X1 port map( A1 => g_BAR, A2 => n4, ZN => g_out);
   U1 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_35 is

   port( p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic;  
         g_BAR : in std_logic);

end pg_35;

architecture SYN_beh of pg_35 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);
   U2 : NAND2_X1 port map( A1 => g_prec, A2 => p, ZN => n4);
   U3 : NAND2_X1 port map( A1 => n4, A2 => g_BAR, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_30 is

   port( p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic;  
         g_BAR : in std_logic);

end pg_30;

architecture SYN_beh of pg_30 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);
   U2 : NAND2_X1 port map( A1 => g_prec, A2 => p, ZN => n4);
   U3 : NAND2_X1 port map( A1 => n4, A2 => g_BAR, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_11 is

   port( p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic;  
         g_BAR : in std_logic);

end pg_11;

architecture SYN_beh of pg_11 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);
   U2 : NAND2_X1 port map( A1 => g_prec, A2 => p, ZN => n4);
   U3 : NAND2_X1 port map( A1 => n4, A2 => g_BAR, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_10 is

   port( p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic;  
         g_BAR : in std_logic);

end pg_10;

architecture SYN_beh of pg_10 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);
   U2 : NAND2_X1 port map( A1 => p, A2 => g_prec, ZN => n4);
   U3 : NAND2_X1 port map( A1 => n4, A2 => g_BAR, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_9 is

   port( p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic;  
         g_BAR : in std_logic);

end pg_9;

architecture SYN_beh of pg_9 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);
   U2 : NAND2_X1 port map( A1 => g_prec, A2 => p, ZN => n4);
   U3 : NAND2_X1 port map( A1 => n4, A2 => g_BAR, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_4 is

   port( p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic;  
         g_BAR : in std_logic);

end pg_4;

architecture SYN_beh of pg_4 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);
   U2 : NAND2_X1 port map( A1 => p, A2 => g_prec, ZN => n4);
   U3 : NAND2_X1 port map( A1 => n4, A2 => g_BAR, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_50 is

   port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic);

end pg_50;

architecture SYN_beh of pg_50 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U3 : AOI21_X1 port map( B1 => g_prec, B2 => p, A => g, ZN => n5);
   U1 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);
   U2 : INV_X1 port map( A => n5, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_48 is

   port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic);

end pg_48;

architecture SYN_beh of pg_48 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U3 : AOI21_X1 port map( B1 => g_prec, B2 => p, A => g, ZN => n5);
   U1 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);
   U2 : INV_X1 port map( A => n5, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_44 is

   port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic);

end pg_44;

architecture SYN_beh of pg_44 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U3 : AOI21_X1 port map( B1 => g_prec, B2 => p, A => g, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => g_out);
   U1 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_43 is

   port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic);

end pg_43;

architecture SYN_beh of pg_43 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U3 : AOI21_X1 port map( B1 => g_prec, B2 => p, A => g, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => g_out);
   U1 : AND2_X1 port map( A1 => p_prec, A2 => p, ZN => p_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_42 is

   port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic);

end pg_42;

architecture SYN_beh of pg_42 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);
   U2 : INV_X1 port map( A => n5, ZN => g_out);
   U3 : AOI21_X1 port map( B1 => g_prec, B2 => p, A => g, ZN => n5);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_41 is

   port( g, p, g_prec, p_prec : in std_logic;  p_out, g_out_BAR : out std_logic
         );

end pg_41;

architecture SYN_beh of pg_41 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p_prec, A2 => p, ZN => p_out);
   U2 : AOI21_X1 port map( B1 => p, B2 => g_prec, A => g, ZN => g_out_BAR);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_33 is

   port( p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic;  
         g_BAR : in std_logic);

end pg_33;

architecture SYN_beh of pg_33 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);
   U2 : NAND2_X1 port map( A1 => g_prec, A2 => p, ZN => n5);
   U3 : NAND2_X1 port map( A1 => n5, A2 => g_BAR, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_31 is

   port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic);

end pg_31;

architecture SYN_beh of pg_31 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U3 : AOI21_X1 port map( B1 => g_prec, B2 => p, A => g, ZN => n5);
   U1 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);
   U2 : INV_X1 port map( A => n5, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_28 is

   port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic);

end pg_28;

architecture SYN_beh of pg_28 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p_prec, A2 => p, ZN => p_out);
   U2 : INV_X1 port map( A => g, ZN => n6);
   U3 : NAND2_X1 port map( A1 => g_prec, A2 => p, ZN => n5);
   U4 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_26 is

   port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic);

end pg_26;

architecture SYN_beh of pg_26 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => g_prec, B2 => p, A => g, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => g_out);
   U3 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_24 is

   port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic);

end pg_24;

architecture SYN_beh of pg_24 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => p, B2 => g_prec, A => g, ZN => n5);
   U2 : INV_X1 port map( A => n5, ZN => g_out);
   U3 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_22 is

   port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic);

end pg_22;

architecture SYN_beh of pg_22 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U1 : INV_X1 port map( A => g, ZN => n6);
   U2 : AND2_X1 port map( A1 => p_prec, A2 => p, ZN => p_out);
   U3 : NAND2_X1 port map( A1 => p, A2 => g_prec, ZN => n5);
   U4 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_18 is

   port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic);

end pg_18;

architecture SYN_beh of pg_18 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U3 : AOI21_X1 port map( B1 => p, B2 => g_prec, A => g, ZN => n5);
   U1 : INV_X1 port map( A => n5, ZN => g_out);
   U2 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_17 is

   port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic);

end pg_17;

architecture SYN_beh of pg_17 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U3 : AOI21_X1 port map( B1 => p, B2 => g_prec, A => g, ZN => n5);
   U1 : INV_X1 port map( A => n5, ZN => g_out);
   U2 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_16 is

   port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic);

end pg_16;

architecture SYN_beh of pg_16 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n6 : std_logic;

begin
   
   U3 : AOI21_X1 port map( B1 => p, B2 => g_prec, A => g, ZN => n6);
   U1 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);
   U2 : INV_X1 port map( A => n6, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_15 is

   port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic);

end pg_15;

architecture SYN_beh of pg_15 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U3 : AOI21_X1 port map( B1 => g_prec, B2 => p, A => g, ZN => n5);
   U1 : INV_X1 port map( A => n5, ZN => g_out);
   U2 : AND2_X1 port map( A1 => p_prec, A2 => p, ZN => p_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_14 is

   port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic);

end pg_14;

architecture SYN_beh of pg_14 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U3 : AOI21_X1 port map( B1 => g_prec, B2 => p, A => g, ZN => n5);
   U1 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);
   U2 : INV_X1 port map( A => n5, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_13 is

   port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic);

end pg_13;

architecture SYN_beh of pg_13 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U3 : AOI21_X1 port map( B1 => g_prec, B2 => p, A => g, ZN => n5);
   U1 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);
   U2 : INV_X1 port map( A => n5, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_7 is

   port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic);

end pg_7;

architecture SYN_beh of pg_7 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);
   U2 : INV_X1 port map( A => n5, ZN => g_out);
   U3 : AOI21_X1 port map( B1 => g_prec, B2 => p, A => g, ZN => n5);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_6 is

   port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic);

end pg_6;

architecture SYN_beh of pg_6 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U3 : AOI21_X1 port map( B1 => g_prec, B2 => p, A => g, ZN => n5);
   U1 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);
   U2 : INV_X1 port map( A => n5, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_5 is

   port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic);

end pg_5;

architecture SYN_beh of pg_5 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);
   U2 : INV_X1 port map( A => g, ZN => n6);
   U3 : NAND2_X1 port map( A1 => g_prec, A2 => p, ZN => n5);
   U4 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_3 is

   port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic);

end pg_3;

architecture SYN_beh of pg_3 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U3 : AOI21_X1 port map( B1 => g_prec, B2 => p, A => g, ZN => n5);
   U1 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);
   U2 : INV_X1 port map( A => n5, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_2 is

   port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic);

end pg_2;

architecture SYN_beh of pg_2 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);
   U2 : INV_X1 port map( A => g, ZN => n6);
   U3 : NAND2_X1 port map( A1 => g_prec, A2 => p, ZN => n5);
   U4 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_1 is

   port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic);

end pg_1;

architecture SYN_beh of pg_1 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);
   U2 : INV_X1 port map( A => n5, ZN => g_out);
   U3 : AOI21_X1 port map( B1 => g_prec, B2 => p, A => g, ZN => n5);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity g_9 is

   port( g, p, g_prec : in std_logic;  g_out : out std_logic);

end g_9;

architecture SYN_beh of g_9 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => p, B2 => g_prec, A => g, ZN => n4);
   U2 : INV_X1 port map( A => n4, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity g_16 is

   port( g, p, g_prec : in std_logic;  g_out : out std_logic);

end g_16;

architecture SYN_beh of g_16 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U2 : AOI21_X1 port map( B1 => p, B2 => g_prec, A => g, ZN => n5);
   U1 : INV_X1 port map( A => n5, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity g_15 is

   port( g, p, g_prec : in std_logic;  g_out : out std_logic);

end g_15;

architecture SYN_beh of g_15 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U2 : AOI21_X1 port map( B1 => p, B2 => g_prec, A => g, ZN => n5);
   U1 : INV_X1 port map( A => n5, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity g_14 is

   port( g, p, g_prec : in std_logic;  g_out : out std_logic);

end g_14;

architecture SYN_beh of g_14 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U2 : AOI21_X1 port map( B1 => p, B2 => g_prec, A => g, ZN => n5);
   U1 : INV_X1 port map( A => n5, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity g_13 is

   port( g, p, g_prec : in std_logic;  g_out : out std_logic);

end g_13;

architecture SYN_beh of g_13 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => g_out);
   U2 : AOI21_X1 port map( B1 => p, B2 => g_prec, A => g, ZN => n5);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity g_12 is

   port( g, p, g_prec : in std_logic;  g_out : out std_logic);

end g_12;

architecture SYN_beh of g_12 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p, A2 => g_prec, ZN => n5);
   U2 : OR2_X1 port map( A1 => g, A2 => n5, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity g_11 is

   port( g, p, g_prec : in std_logic;  g_out : out std_logic);

end g_11;

architecture SYN_beh of g_11 is

   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p, A2 => g_prec, ZN => n5);
   U2 : OR2_X2 port map( A1 => g, A2 => n5, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity g_8 is

   port( g, p, g_prec : in std_logic;  g_out : out std_logic);

end g_8;

architecture SYN_beh of g_8 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U1 : INV_X1 port map( A => g, ZN => n5);
   U2 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => g_out);
   U3 : NAND2_X1 port map( A1 => g_prec, A2 => p, ZN => n6);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity g_7 is

   port( g, p, g_prec : in std_logic;  g_out : out std_logic);

end g_7;

architecture SYN_beh of g_7 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => g_out);
   U2 : INV_X1 port map( A => g, ZN => n5);
   U3 : NAND2_X1 port map( A1 => g_prec, A2 => p, ZN => n6);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity g_6 is

   port( g, p, g_prec : in std_logic;  g_out : out std_logic);

end g_6;

architecture SYN_beh of g_6 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => g_out);
   U2 : AOI21_X1 port map( B1 => p, B2 => g_prec, A => g, ZN => n5);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity g_5 is

   port( g, p, g_prec : in std_logic;  g_out : out std_logic);

end g_5;

architecture SYN_beh of g_5 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => g_out);
   U2 : AOI21_X1 port map( B1 => g_prec, B2 => p, A => g, ZN => n5);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity g_4 is

   port( g, p, g_prec : in std_logic;  g_out : out std_logic);

end g_4;

architecture SYN_beh of g_4 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => g_out);
   U2 : INV_X1 port map( A => g, ZN => n6);
   U3 : NAND2_X1 port map( A1 => g_prec, A2 => p, ZN => n5);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity g_3 is

   port( g, p, g_prec : in std_logic;  g_out : out std_logic);

end g_3;

architecture SYN_beh of g_3 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U1 : INV_X1 port map( A => g, ZN => n6);
   U2 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => g_out);
   U3 : NAND2_X1 port map( A1 => g_prec, A2 => p, ZN => n5);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity g_2 is

   port( g, p, g_prec : in std_logic;  g_out : out std_logic);

end g_2;

architecture SYN_beh of g_2 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => g_out);
   U2 : AOI21_X1 port map( B1 => g_prec, B2 => p, A => g, ZN => n5);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity g_1 is

   port( g, p, g_prec : in std_logic;  g_out : out std_logic);

end g_1;

architecture SYN_beh of g_1 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => g_out);
   U2 : AOI21_X1 port map( B1 => p, B2 => g_prec, A => g, ZN => n5);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_18 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_18;

architecture SYN_beh of pg_net_18 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_61 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_61;

architecture SYN_beh of pg_net_61 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_60 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_60;

architecture SYN_beh of pg_net_60 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_59 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_59;

architecture SYN_beh of pg_net_59 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_58 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_58;

architecture SYN_beh of pg_net_58 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_57 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_57;

architecture SYN_beh of pg_net_57 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_56 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_56;

architecture SYN_beh of pg_net_56 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_55 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_55;

architecture SYN_beh of pg_net_55 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_54 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_54;

architecture SYN_beh of pg_net_54 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_53 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_53;

architecture SYN_beh of pg_net_53 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_52 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_52;

architecture SYN_beh of pg_net_52 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_51 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_51;

architecture SYN_beh of pg_net_51 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_50 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_50;

architecture SYN_beh of pg_net_50 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_48 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_48;

architecture SYN_beh of pg_net_48 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_47 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_47;

architecture SYN_beh of pg_net_47 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => a, ZN => n2);
   U2 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);
   U3 : XNOR2_X1 port map( A => b, B => n2, ZN => p_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_46 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_46;

architecture SYN_beh of pg_net_46 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_45 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_45;

architecture SYN_beh of pg_net_45 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_44 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_44;

architecture SYN_beh of pg_net_44 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_43 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_43;

architecture SYN_beh of pg_net_43 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);
   U2 : INV_X1 port map( A => a, ZN => n2);
   U3 : XNOR2_X1 port map( A => b, B => n2, ZN => p_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_42 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_42;

architecture SYN_beh of pg_net_42 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_41 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_41;

architecture SYN_beh of pg_net_41 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);
   U2 : INV_X1 port map( A => a, ZN => n2);
   U3 : XNOR2_X1 port map( A => b, B => n2, ZN => p_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_40 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_40;

architecture SYN_beh of pg_net_40 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_39 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_39;

architecture SYN_beh of pg_net_39 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_38 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_38;

architecture SYN_beh of pg_net_38 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => a, B => b, Z => p_out);
   U2 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_37 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_37;

architecture SYN_beh of pg_net_37 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_32 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_32;

architecture SYN_beh of pg_net_32 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_31 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_31;

architecture SYN_beh of pg_net_31 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => a, ZN => n2);
   U2 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);
   U3 : XNOR2_X1 port map( A => b, B => n2, ZN => p_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_30 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_30;

architecture SYN_beh of pg_net_30 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => a, B => b, Z => p_out);
   U2 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_29 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_29;

architecture SYN_beh of pg_net_29 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => a, A2 => b, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_28 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_28;

architecture SYN_beh of pg_net_28 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => a, ZN => n2);
   U2 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);
   U3 : XNOR2_X1 port map( A => b, B => n2, ZN => p_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_27 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_27;

architecture SYN_beh of pg_net_27 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => a, ZN => n3);
   U2 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);
   U3 : XNOR2_X1 port map( A => b, B => n3, ZN => p_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_26 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_26;

architecture SYN_beh of pg_net_26 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_25 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_25;

architecture SYN_beh of pg_net_25 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_24 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_24;

architecture SYN_beh of pg_net_24 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_23 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_23;

architecture SYN_beh of pg_net_23 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => a, ZN => n2);
   U2 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);
   U3 : XNOR2_X1 port map( A => b, B => n2, ZN => p_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_22 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_22;

architecture SYN_beh of pg_net_22 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_21 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_21;

architecture SYN_beh of pg_net_21 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_20 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_20;

architecture SYN_beh of pg_net_20 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => a, ZN => n2);
   U2 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);
   U3 : XNOR2_X1 port map( A => b, B => n2, ZN => p_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_19 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_19;

architecture SYN_beh of pg_net_19 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_17 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_17;

architecture SYN_beh of pg_net_17 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_16 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_16;

architecture SYN_beh of pg_net_16 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_15 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_15;

architecture SYN_beh of pg_net_15 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => a, B => b, Z => p_out);
   U2 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_14 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_14;

architecture SYN_beh of pg_net_14 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_13 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_13;

architecture SYN_beh of pg_net_13 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_12 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_12;

architecture SYN_beh of pg_net_12 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => a, ZN => n2);
   U2 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);
   U3 : XNOR2_X1 port map( A => b, B => n2, ZN => p_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_11 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_11;

architecture SYN_beh of pg_net_11 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_10 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_10;

architecture SYN_beh of pg_net_10 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_9 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_9;

architecture SYN_beh of pg_net_9 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_8 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_8;

architecture SYN_beh of pg_net_8 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_7 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_7;

architecture SYN_beh of pg_net_7 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_6 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_6;

architecture SYN_beh of pg_net_6 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_5 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_5;

architecture SYN_beh of pg_net_5 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_4 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_4;

architecture SYN_beh of pg_net_4 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_3 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_3;

architecture SYN_beh of pg_net_3 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_2 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_2;

architecture SYN_beh of pg_net_2 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_1 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_1;

architecture SYN_beh of pg_net_1 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => a, ZN => n2);
   U2 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);
   U3 : XNOR2_X1 port map( A => b, B => n2, ZN => p_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_0_1 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_0_1;

architecture SYN_BEHAVIORAL of FA_0_1 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity mux21_SIZE4_0_1 is

   port( IN0, IN1 : in std_logic_vector (3 downto 0);  CTRL : in std_logic;  
         OUT1 : out std_logic_vector (3 downto 0));

end mux21_SIZE4_0_1;

architecture SYN_Bhe of mux21_SIZE4_0_1 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => IN0(3), B => IN1(3), S => CTRL, Z => OUT1(3));
   U2 : MUX2_X1 port map( A => IN0(2), B => IN1(2), S => CTRL, Z => OUT1(2));
   U3 : MUX2_X1 port map( A => IN0(1), B => IN1(1), S => CTRL, Z => OUT1(1));
   U4 : MUX2_X1 port map( A => IN0(0), B => IN1(0), S => CTRL, Z => OUT1(0));

end SYN_Bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity RCA_N4_0_1 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_0_1;

architecture SYN_STRUCTURAL of RCA_N4_0_1 is

   component FA_61
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_62
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_63
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_0_1
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal n1, CTMP_3_port, CTMP_2_port, CTMP_1_port, net684357 : std_logic;

begin
   
   n1 <= '0';
   FAI_1 : FA_0_1 port map( A => A(0), B => B(0), Ci => n1, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_63 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_62 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_61 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => net684357);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity carry_sel_gen_N4_0_1 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end carry_sel_gen_N4_0_1;

architecture SYN_STRUCTURAL of carry_sel_gen_N4_0_1 is

   component mux21_SIZE4_0_1
      port( IN0, IN1 : in std_logic_vector (3 downto 0);  CTRL : in std_logic; 
            OUT1 : out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_N4_15
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_0_1
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, nocarry_sum_to_mux_3_port, 
      nocarry_sum_to_mux_2_port, nocarry_sum_to_mux_1_port, 
      nocarry_sum_to_mux_0_port, carry_sum_to_mux_3_port, 
      carry_sum_to_mux_2_port, carry_sum_to_mux_1_port, carry_sum_to_mux_0_port
      , net684355, net684356 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   rca_nocarry : RCA_N4_0_1 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1),
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           nocarry_sum_to_mux_3_port, S(2) => 
                           nocarry_sum_to_mux_2_port, S(1) => 
                           nocarry_sum_to_mux_1_port, S(0) => 
                           nocarry_sum_to_mux_0_port, Co => net684356);
   rca_carry : RCA_N4_15 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           carry_sum_to_mux_3_port, S(2) => 
                           carry_sum_to_mux_2_port, S(1) => 
                           carry_sum_to_mux_1_port, S(0) => 
                           carry_sum_to_mux_0_port, Co => net684355);
   outmux : mux21_SIZE4_0_1 port map( IN0(3) => nocarry_sum_to_mux_3_port, 
                           IN0(2) => nocarry_sum_to_mux_2_port, IN0(1) => 
                           nocarry_sum_to_mux_1_port, IN0(0) => 
                           nocarry_sum_to_mux_0_port, IN1(3) => 
                           carry_sum_to_mux_3_port, IN1(2) => 
                           carry_sum_to_mux_2_port, IN1(1) => 
                           carry_sum_to_mux_1_port, IN1(0) => 
                           carry_sum_to_mux_0_port, CTRL => Ci, OUT1(3) => S(3)
                           , OUT1(2) => S(2), OUT1(1) => S(1), OUT1(0) => S(0))
                           ;

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_0_1 is

   port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic);

end pg_0_1;

architecture SYN_beh of pg_0_1 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U1 : INV_X1 port map( A => g, ZN => n6);
   U2 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);
   U3 : NAND2_X1 port map( A1 => p, A2 => g_prec, ZN => n5);
   U4 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity g_0_1 is

   port( g, p, g_prec : in std_logic;  g_out : out std_logic);

end g_0_1;

architecture SYN_beh of g_0_1 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => p, B2 => g_prec, A => g, ZN => n4);
   U2 : INV_X1 port map( A => n4, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_0_1 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_0_1;

architecture SYN_beh of pg_net_0_1 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => a, ZN => n3);
   U2 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);
   U3 : XNOR2_X1 port map( A => n3, B => b, ZN => p_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity sum_gen_N32_1 is

   port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic_vector 
         (8 downto 0);  S : out std_logic_vector (31 downto 0));

end sum_gen_N32_1;

architecture SYN_STRUCTURAL of sum_gen_N32_1 is

   component carry_sel_gen_N4_1
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component carry_sel_gen_N4_2
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component carry_sel_gen_N4_3
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component carry_sel_gen_N4_4
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component carry_sel_gen_N4_5
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component carry_sel_gen_N4_6
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component carry_sel_gen_N4_7
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component carry_sel_gen_N4_0_1
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal net684347, net684348, net684349, net684350, net684351, net684352, 
      net684353, net684354 : std_logic;

begin
   
   csel_N_0 : carry_sel_gen_N4_0_1 port map( A(3) => A(3), A(2) => A(2), A(1) 
                           => A(1), A(0) => A(0), B(3) => B(3), B(2) => B(2), 
                           B(1) => B(1), B(0) => B(0), Ci => Cin(0), S(3) => 
                           S(3), S(2) => S(2), S(1) => S(1), S(0) => S(0), Co 
                           => net684354);
   csel_N_1 : carry_sel_gen_N4_7 port map( A(3) => A(7), A(2) => A(6), A(1) => 
                           A(5), A(0) => A(4), B(3) => B(7), B(2) => B(6), B(1)
                           => B(5), B(0) => B(4), Ci => Cin(1), S(3) => S(7), 
                           S(2) => S(6), S(1) => S(5), S(0) => S(4), Co => 
                           net684353);
   csel_N_2 : carry_sel_gen_N4_6 port map( A(3) => A(11), A(2) => A(10), A(1) 
                           => A(9), A(0) => A(8), B(3) => B(11), B(2) => B(10),
                           B(1) => B(9), B(0) => B(8), Ci => Cin(2), S(3) => 
                           S(11), S(2) => S(10), S(1) => S(9), S(0) => S(8), Co
                           => net684352);
   csel_N_3 : carry_sel_gen_N4_5 port map( A(3) => A(15), A(2) => A(14), A(1) 
                           => A(13), A(0) => A(12), B(3) => B(15), B(2) => 
                           B(14), B(1) => B(13), B(0) => B(12), Ci => Cin(3), 
                           S(3) => S(15), S(2) => S(14), S(1) => S(13), S(0) =>
                           S(12), Co => net684351);
   csel_N_4 : carry_sel_gen_N4_4 port map( A(3) => A(19), A(2) => A(18), A(1) 
                           => A(17), A(0) => A(16), B(3) => B(19), B(2) => 
                           B(18), B(1) => B(17), B(0) => B(16), Ci => Cin(4), 
                           S(3) => S(19), S(2) => S(18), S(1) => S(17), S(0) =>
                           S(16), Co => net684350);
   csel_N_5 : carry_sel_gen_N4_3 port map( A(3) => A(23), A(2) => A(22), A(1) 
                           => A(21), A(0) => A(20), B(3) => B(23), B(2) => 
                           B(22), B(1) => B(21), B(0) => B(20), Ci => Cin(5), 
                           S(3) => S(23), S(2) => S(22), S(1) => S(21), S(0) =>
                           S(20), Co => net684349);
   csel_N_6 : carry_sel_gen_N4_2 port map( A(3) => A(27), A(2) => A(26), A(1) 
                           => A(25), A(0) => A(24), B(3) => B(27), B(2) => 
                           B(26), B(1) => B(25), B(0) => B(24), Ci => Cin(6), 
                           S(3) => S(27), S(2) => S(26), S(1) => S(25), S(0) =>
                           S(24), Co => net684348);
   csel_N_7 : carry_sel_gen_N4_1 port map( A(3) => A(31), A(2) => A(30), A(1) 
                           => A(29), A(0) => A(28), B(3) => B(31), B(2) => 
                           B(30), B(1) => B(29), B(0) => B(28), Ci => Cin(7), 
                           S(3) => S(31), S(2) => S(30), S(1) => S(29), S(0) =>
                           S(28), Co => net684347);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity carry_tree_N32_logN5_1 is

   port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  Cout :
         out std_logic_vector (7 downto 0));

end carry_tree_N32_logN5_1;

architecture SYN_arch of carry_tree_N32_logN5_1 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component pg_1
      port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic
            );
   end component;
   
   component pg_2
      port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic
            );
   end component;
   
   component pg_3
      port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic
            );
   end component;
   
   component pg_4
      port( p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic;  
            g_BAR : in std_logic);
   end component;
   
   component pg_5
      port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic
            );
   end component;
   
   component g_1
      port( g, p, g_prec : in std_logic;  g_out : out std_logic);
   end component;
   
   component g_2
      port( g, p, g_prec : in std_logic;  g_out : out std_logic);
   end component;
   
   component g_3
      port( g, p, g_prec : in std_logic;  g_out : out std_logic);
   end component;
   
   component g_4
      port( g, p, g_prec : in std_logic;  g_out : out std_logic);
   end component;
   
   component g_5
      port( g, p, g_prec : in std_logic;  g_out : out std_logic);
   end component;
   
   component g_6
      port( g, p, g_prec : in std_logic;  g_out : out std_logic);
   end component;
   
   component g_7
      port( g, p, g_prec : in std_logic;  g_out : out std_logic);
   end component;
   
   component pg_6
      port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic
            );
   end component;
   
   component pg_7
      port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic
            );
   end component;
   
   component pg_8
      port( g, p, g_prec, p_prec : in std_logic;  p_out, g_out_BAR : out 
            std_logic);
   end component;
   
   component pg_9
      port( p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic;  
            g_BAR : in std_logic);
   end component;
   
   component pg_10
      port( p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic;  
            g_BAR : in std_logic);
   end component;
   
   component pg_11
      port( p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic;  
            g_BAR : in std_logic);
   end component;
   
   component pg_12
      port( p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic;  
            g_BAR : in std_logic);
   end component;
   
   component g_8
      port( g, p, g_prec : in std_logic;  g_out : out std_logic);
   end component;
   
   component pg_13
      port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic
            );
   end component;
   
   component pg_14
      port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic
            );
   end component;
   
   component pg_15
      port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic
            );
   end component;
   
   component pg_16
      port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic
            );
   end component;
   
   component pg_17
      port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic
            );
   end component;
   
   component pg_18
      port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic
            );
   end component;
   
   component pg_19
      port( g, p, g_prec, p_prec : in std_logic;  p_out, g_out_BAR : out 
            std_logic);
   end component;
   
   component pg_20
      port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic
            );
   end component;
   
   component pg_21
      port( g, p, g_prec, p_prec : in std_logic;  p_out, g_out_BAR : out 
            std_logic);
   end component;
   
   component pg_22
      port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic
            );
   end component;
   
   component pg_23
      port( g, p, g_prec, p_prec : in std_logic;  p_out, g_out_BAR : out 
            std_logic);
   end component;
   
   component pg_24
      port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic
            );
   end component;
   
   component pg_25
      port( g, p, g_prec, p_prec : in std_logic;  p_out, g_out_BAR : out 
            std_logic);
   end component;
   
   component pg_26
      port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic
            );
   end component;
   
   component pg_0_1
      port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic
            );
   end component;
   
   component g_9
      port( g, p, g_prec : in std_logic;  g_out : out std_logic);
   end component;
   
   component g_0_1
      port( g, p, g_prec : in std_logic;  g_out : out std_logic);
   end component;
   
   component pg_net_1
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_2
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_3
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_4
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_5
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_6
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_7
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_8
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_9
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_10
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_11
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_12
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_13
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_14
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_15
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_16
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_17
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_18
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_19
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_20
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_21
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_22
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_23
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_24
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_25
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_26
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_27
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_28
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_29
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_30
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_31
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_0_1
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   signal Cout_7_port, Cout_6_port, Cout_5_port, Cout_4_port, Cout_2_port, 
      p_net_31_port, p_net_30_port, p_net_29_port, p_net_28_port, p_net_27_port
      , p_net_26_port, p_net_24_port, p_net_23_port, p_net_22_port, 
      p_net_21_port, p_net_20_port, p_net_19_port, p_net_18_port, p_net_17_port
      , p_net_16_port, p_net_15_port, p_net_14_port, p_net_13_port, 
      p_net_12_port, p_net_11_port, p_net_10_port, p_net_9_port, p_net_8_port, 
      p_net_7_port, p_net_6_port, p_net_5_port, p_net_4_port, p_net_3_port, 
      p_net_2_port, p_net_1_port, g_net_31_port, g_net_30_port, g_net_29_port, 
      g_net_28_port, g_net_27_port, g_net_26_port, g_net_25_port, g_net_24_port
      , g_net_23_port, g_net_22_port, g_net_21_port, g_net_20_port, 
      g_net_19_port, g_net_18_port, g_net_17_port, g_net_16_port, g_net_15_port
      , g_net_14_port, g_net_13_port, g_net_12_port, g_net_11_port, 
      g_net_10_port, g_net_9_port, g_net_8_port, g_net_7_port, g_net_6_port, 
      g_net_5_port, g_net_4_port, g_net_3_port, g_net_2_port, g_net_1_port, 
      g_net_0_port, magic_pro_1_port, magic_pro_0_port, pg_1_15_1_port, 
      pg_1_15_0_port, pg_1_14_1_port, pg_1_14_0_port, pg_1_13_1_port, 
      pg_1_13_0_port, pg_1_12_1_port, pg_1_12_0_port, pg_1_11_1_port, 
      pg_1_11_0_port, pg_1_10_1_port, pg_1_10_0_port, pg_1_9_1_port, 
      pg_1_9_0_port, pg_1_8_1_port, pg_1_8_0_port, pg_1_7_1_port, pg_1_7_0_port
      , pg_1_6_1_port, pg_1_6_0_port, pg_1_5_1_port, pg_1_5_0_port, 
      pg_1_4_1_port, pg_1_4_0_port, pg_1_3_1_port, pg_1_3_0_port, pg_1_2_1_port
      , pg_1_2_0_port, pg_1_1_1_port, pg_1_1_0_port, pg_1_0_0_port, 
      pg_n_4_7_1_port, pg_n_4_7_0_port, pg_n_4_6_1_port, pg_n_4_6_0_port, 
      pg_n_3_7_1_port, pg_n_3_7_0_port, pg_n_3_5_1_port, pg_n_3_3_1_port, 
      pg_n_3_3_0_port, pg_n_2_7_1_port, pg_n_2_7_0_port, pg_n_2_6_1_port, 
      pg_n_2_6_0_port, pg_n_2_5_1_port, pg_n_2_5_0_port, pg_n_2_4_1_port, 
      pg_n_2_3_1_port, pg_n_2_3_0_port, pg_n_2_2_1_port, pg_n_2_2_0_port, 
      pg_n_2_1_1_port, pg_n_2_1_0_port, n1, n5, n26, n7, n8, n12, n18, n20, 
      Cout_3_port, n22, n23, Cout_0_port, Cout_1_port : std_logic;

begin
   Cout <= ( Cout_7_port, Cout_6_port, Cout_5_port, Cout_4_port, Cout_3_port, 
      Cout_2_port, Cout_1_port, Cout_0_port );
   
   pg_net_x_1 : pg_net_0_1 port map( a => A(1), b => B(1), g_out => 
                           g_net_1_port, p_out => p_net_1_port);
   pg_net_x_2 : pg_net_31 port map( a => A(2), b => B(2), g_out => g_net_2_port
                           , p_out => p_net_2_port);
   pg_net_x_3 : pg_net_30 port map( a => A(3), b => B(3), g_out => g_net_3_port
                           , p_out => p_net_3_port);
   pg_net_x_4 : pg_net_29 port map( a => A(4), b => B(4), g_out => g_net_4_port
                           , p_out => p_net_4_port);
   pg_net_x_5 : pg_net_28 port map( a => A(5), b => B(5), g_out => g_net_5_port
                           , p_out => p_net_5_port);
   pg_net_x_6 : pg_net_27 port map( a => A(6), b => B(6), g_out => g_net_6_port
                           , p_out => p_net_6_port);
   pg_net_x_7 : pg_net_26 port map( a => A(7), b => B(7), g_out => g_net_7_port
                           , p_out => p_net_7_port);
   pg_net_x_8 : pg_net_25 port map( a => A(8), b => B(8), g_out => g_net_8_port
                           , p_out => p_net_8_port);
   pg_net_x_9 : pg_net_24 port map( a => A(9), b => B(9), g_out => g_net_9_port
                           , p_out => p_net_9_port);
   pg_net_x_10 : pg_net_23 port map( a => A(10), b => B(10), g_out => 
                           g_net_10_port, p_out => p_net_10_port);
   pg_net_x_11 : pg_net_22 port map( a => A(11), b => B(11), g_out => 
                           g_net_11_port, p_out => p_net_11_port);
   pg_net_x_12 : pg_net_21 port map( a => A(12), b => B(12), g_out => 
                           g_net_12_port, p_out => p_net_12_port);
   pg_net_x_13 : pg_net_20 port map( a => A(13), b => B(13), g_out => 
                           g_net_13_port, p_out => p_net_13_port);
   pg_net_x_14 : pg_net_19 port map( a => A(14), b => B(14), g_out => 
                           g_net_14_port, p_out => p_net_14_port);
   pg_net_x_15 : pg_net_18 port map( a => A(15), b => B(15), g_out => 
                           g_net_15_port, p_out => p_net_15_port);
   pg_net_x_16 : pg_net_17 port map( a => A(16), b => B(16), g_out => 
                           g_net_16_port, p_out => p_net_16_port);
   pg_net_x_17 : pg_net_16 port map( a => A(17), b => B(17), g_out => 
                           g_net_17_port, p_out => p_net_17_port);
   pg_net_x_18 : pg_net_15 port map( a => A(18), b => B(18), g_out => 
                           g_net_18_port, p_out => p_net_18_port);
   pg_net_x_19 : pg_net_14 port map( a => A(19), b => B(19), g_out => 
                           g_net_19_port, p_out => p_net_19_port);
   pg_net_x_20 : pg_net_13 port map( a => A(20), b => B(20), g_out => 
                           g_net_20_port, p_out => p_net_20_port);
   pg_net_x_21 : pg_net_12 port map( a => A(21), b => B(21), g_out => 
                           g_net_21_port, p_out => p_net_21_port);
   pg_net_x_22 : pg_net_11 port map( a => A(22), b => B(22), g_out => 
                           g_net_22_port, p_out => p_net_22_port);
   pg_net_x_23 : pg_net_10 port map( a => A(23), b => B(23), g_out => 
                           g_net_23_port, p_out => p_net_23_port);
   pg_net_x_24 : pg_net_9 port map( a => A(24), b => B(24), g_out => 
                           g_net_24_port, p_out => p_net_24_port);
   pg_net_x_25 : pg_net_8 port map( a => A(25), b => B(25), g_out => 
                           g_net_25_port, p_out => n18);
   pg_net_x_26 : pg_net_7 port map( a => A(26), b => B(26), g_out => 
                           g_net_26_port, p_out => p_net_26_port);
   pg_net_x_27 : pg_net_6 port map( a => A(27), b => B(27), g_out => 
                           g_net_27_port, p_out => p_net_27_port);
   pg_net_x_28 : pg_net_5 port map( a => A(28), b => B(28), g_out => 
                           g_net_28_port, p_out => p_net_28_port);
   pg_net_x_29 : pg_net_4 port map( a => A(29), b => B(29), g_out => 
                           g_net_29_port, p_out => p_net_29_port);
   pg_net_x_30 : pg_net_3 port map( a => A(30), b => B(30), g_out => 
                           g_net_30_port, p_out => p_net_30_port);
   pg_net_x_31 : pg_net_2 port map( a => A(31), b => B(31), g_out => 
                           g_net_31_port, p_out => p_net_31_port);
   pg_net_0_MAGIC : pg_net_1 port map( a => A(0), b => B(0), g_out => 
                           magic_pro_0_port, p_out => magic_pro_1_port);
   xG_0_0_MAGIC : g_0_1 port map( g => magic_pro_0_port, p => magic_pro_1_port,
                           g_prec => Cin, g_out => g_net_0_port);
   xG_1_0 : g_9 port map( g => g_net_1_port, p => p_net_1_port, g_prec => 
                           g_net_0_port, g_out => pg_1_0_0_port);
   xPG_1_1 : pg_0_1 port map( g => g_net_3_port, p => p_net_3_port, g_prec => 
                           g_net_2_port, p_prec => p_net_2_port, g_out => 
                           pg_1_1_0_port, p_out => pg_1_1_1_port);
   xPG_1_2 : pg_26 port map( g => g_net_5_port, p => p_net_5_port, g_prec => 
                           g_net_4_port, p_prec => p_net_4_port, g_out => 
                           pg_1_2_0_port, p_out => pg_1_2_1_port);
   xPG_1_3 : pg_25 port map( g => g_net_7_port, p => p_net_7_port, g_prec => 
                           g_net_6_port, p_prec => p_net_6_port, p_out => 
                           pg_1_3_1_port, g_out_BAR => pg_1_3_0_port);
   xPG_1_4 : pg_24 port map( g => g_net_9_port, p => p_net_9_port, g_prec => 
                           g_net_8_port, p_prec => p_net_8_port, g_out => 
                           pg_1_4_0_port, p_out => pg_1_4_1_port);
   xPG_1_5 : pg_23 port map( g => g_net_11_port, p => p_net_11_port, g_prec => 
                           g_net_10_port, p_prec => p_net_10_port, p_out => 
                           pg_1_5_1_port, g_out_BAR => pg_1_5_0_port);
   xPG_1_6 : pg_22 port map( g => g_net_13_port, p => p_net_13_port, g_prec => 
                           g_net_12_port, p_prec => p_net_12_port, g_out => 
                           pg_1_6_0_port, p_out => pg_1_6_1_port);
   xPG_1_7 : pg_21 port map( g => g_net_15_port, p => p_net_15_port, g_prec => 
                           g_net_14_port, p_prec => p_net_14_port, p_out => 
                           pg_1_7_1_port, g_out_BAR => pg_1_7_0_port);
   xPG_1_8 : pg_20 port map( g => g_net_17_port, p => p_net_17_port, g_prec => 
                           g_net_16_port, p_prec => p_net_16_port, g_out => 
                           pg_1_8_0_port, p_out => pg_1_8_1_port);
   xPG_1_9 : pg_19 port map( g => g_net_19_port, p => p_net_19_port, g_prec => 
                           g_net_18_port, p_prec => p_net_18_port, p_out => 
                           pg_1_9_1_port, g_out_BAR => pg_1_9_0_port);
   xPG_1_10 : pg_18 port map( g => g_net_21_port, p => p_net_21_port, g_prec =>
                           g_net_20_port, p_prec => p_net_20_port, g_out => 
                           pg_1_10_0_port, p_out => pg_1_10_1_port);
   xPG_1_11 : pg_17 port map( g => g_net_23_port, p => p_net_23_port, g_prec =>
                           g_net_22_port, p_prec => p_net_22_port, g_out => 
                           pg_1_11_0_port, p_out => pg_1_11_1_port);
   xPG_1_12 : pg_16 port map( g => g_net_25_port, p => n18, g_prec => 
                           g_net_24_port, p_prec => p_net_24_port, g_out => 
                           pg_1_12_0_port, p_out => pg_1_12_1_port);
   xPG_1_13 : pg_15 port map( g => g_net_27_port, p => p_net_27_port, g_prec =>
                           g_net_26_port, p_prec => p_net_26_port, g_out => 
                           pg_1_13_0_port, p_out => pg_1_13_1_port);
   xPG_1_14 : pg_14 port map( g => g_net_29_port, p => p_net_29_port, g_prec =>
                           g_net_28_port, p_prec => p_net_28_port, g_out => 
                           pg_1_14_0_port, p_out => pg_1_14_1_port);
   xPG_1_15 : pg_13 port map( g => g_net_31_port, p => p_net_31_port, g_prec =>
                           g_net_30_port, p_prec => p_net_30_port, g_out => 
                           pg_1_15_0_port, p_out => pg_1_15_1_port);
   xG_2_0 : g_8 port map( g => pg_1_1_0_port, p => pg_1_1_1_port, g_prec => 
                           pg_1_0_0_port, g_out => n26);
   xPG_2_1 : pg_12 port map( p => pg_1_3_1_port, g_prec => pg_1_2_0_port, 
                           p_prec => pg_1_2_1_port, g_out => pg_n_2_1_0_port, 
                           p_out => pg_n_2_1_1_port, g_BAR => pg_1_3_0_port);
   xPG_2_2 : pg_11 port map( p => pg_1_5_1_port, g_prec => pg_1_4_0_port, 
                           p_prec => pg_1_4_1_port, g_out => pg_n_2_2_0_port, 
                           p_out => pg_n_2_2_1_port, g_BAR => pg_1_5_0_port);
   xPG_2_3 : pg_10 port map( p => pg_1_7_1_port, g_prec => pg_1_6_0_port, 
                           p_prec => pg_1_6_1_port, g_out => pg_n_2_3_0_port, 
                           p_out => pg_n_2_3_1_port, g_BAR => pg_1_7_0_port);
   xPG_2_4 : pg_9 port map( p => pg_1_9_1_port, g_prec => pg_1_8_0_port, p_prec
                           => pg_1_8_1_port, g_out => n5, p_out => 
                           pg_n_2_4_1_port, g_BAR => pg_1_9_0_port);
   xPG_2_5 : pg_8 port map( g => pg_1_11_0_port, p => pg_1_11_1_port, g_prec =>
                           pg_1_10_0_port, p_prec => pg_1_10_1_port, p_out => 
                           pg_n_2_5_1_port, g_out_BAR => pg_n_2_5_0_port);
   xPG_2_6 : pg_7 port map( g => pg_1_13_0_port, p => pg_1_13_1_port, g_prec =>
                           pg_1_12_0_port, p_prec => pg_1_12_1_port, g_out => 
                           pg_n_2_6_0_port, p_out => pg_n_2_6_1_port);
   xPG_2_7 : pg_6 port map( g => pg_1_15_0_port, p => pg_1_15_1_port, g_prec =>
                           pg_1_14_0_port, p_prec => pg_1_14_1_port, g_out => 
                           pg_n_2_7_0_port, p_out => pg_n_2_7_1_port);
   xG_3_1 : g_7 port map( g => pg_n_2_1_0_port, p => pg_n_2_1_1_port, g_prec =>
                           n26, g_out => n8);
   xG_4_2 : g_6 port map( g => n20, p => pg_n_2_2_1_port, g_prec => n23, g_out 
                           => Cout_2_port);
   xG_4_3 : g_5 port map( g => pg_n_3_3_0_port, p => pg_n_3_3_1_port, g_prec =>
                           n8, g_out => n1);
   xG_5_4 : g_4 port map( g => n12, p => pg_n_2_4_1_port, g_prec => n1, g_out 
                           => Cout_4_port);
   xG_5_5 : g_3 port map( g => n22, p => pg_n_3_5_1_port, g_prec => n1, g_out 
                           => Cout_5_port);
   xG_5_6 : g_2 port map( g => pg_n_4_6_0_port, p => pg_n_4_6_1_port, g_prec =>
                           n1, g_out => Cout_6_port);
   xG_5_7 : g_1 port map( g => pg_n_4_7_0_port, p => pg_n_4_7_1_port, g_prec =>
                           Cout_3_port, g_out => Cout_7_port);
   xPG_3_3 : pg_5 port map( g => pg_n_2_3_0_port, p => pg_n_2_3_1_port, g_prec 
                           => pg_n_2_2_0_port, p_prec => pg_n_2_2_1_port, g_out
                           => pg_n_3_3_0_port, p_out => pg_n_3_3_1_port);
   xPG_3_5 : pg_4 port map( p => pg_n_2_5_1_port, g_prec => n5, p_prec => 
                           pg_n_2_4_1_port, g_out => n7, p_out => 
                           pg_n_3_5_1_port, g_BAR => pg_n_2_5_0_port);
   xPG_3_7 : pg_3 port map( g => pg_n_2_7_0_port, p => pg_n_2_7_1_port, g_prec 
                           => pg_n_2_6_0_port, p_prec => pg_n_2_6_1_port, g_out
                           => pg_n_3_7_0_port, p_out => pg_n_3_7_1_port);
   xPG_4_6 : pg_2 port map( g => pg_n_2_6_0_port, p => pg_n_2_6_1_port, g_prec 
                           => n7, p_prec => pg_n_3_5_1_port, g_out => 
                           pg_n_4_6_0_port, p_out => pg_n_4_6_1_port);
   xPG_4_7 : pg_1 port map( g => pg_n_3_7_0_port, p => pg_n_3_7_1_port, g_prec 
                           => n22, p_prec => pg_n_3_5_1_port, g_out => 
                           pg_n_4_7_0_port, p_out => pg_n_4_7_1_port);
   U1 : CLKBUF_X1 port map( A => n5, Z => n12);
   U2 : CLKBUF_X1 port map( A => n7, Z => n22);
   U3 : CLKBUF_X1 port map( A => pg_n_2_2_0_port, Z => n20);
   U4 : BUF_X1 port map( A => n8, Z => n23);
   U5 : BUF_X1 port map( A => n1, Z => Cout_3_port);
   U6 : CLKBUF_X1 port map( A => n26, Z => Cout_0_port);
   U7 : BUF_X1 port map( A => n23, Z => Cout_1_port);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity xor_gen_N32_1 is

   port( A : in std_logic_vector (31 downto 0);  B : in std_logic;  S : out 
         std_logic_vector (31 downto 0));

end xor_gen_N32_1;

architecture SYN_bhe of xor_gen_N32_1 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21_X2
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X2
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   signal n15, n16, n17, n19, n20, n21, n22, n23 : std_logic;

begin
   
   U8 : XOR2_X1 port map( A => B, B => A(31), Z => S(31));
   U9 : XOR2_X1 port map( A => B, B => A(30), Z => S(30));
   U12 : XOR2_X1 port map( A => B, B => A(28), Z => S(28));
   U13 : XOR2_X1 port map( A => B, B => A(27), Z => S(27));
   U14 : XOR2_X1 port map( A => B, B => A(26), Z => S(26));
   U16 : XOR2_X1 port map( A => B, B => A(24), Z => S(24));
   U17 : XOR2_X1 port map( A => B, B => A(23), Z => S(23));
   U20 : XOR2_X1 port map( A => B, B => A(20), Z => S(20));
   U29 : XOR2_X1 port map( A => B, B => A(12), Z => S(12));
   U1 : XNOR2_X1 port map( A => A(0), B => n19, ZN => S(0));
   U2 : XNOR2_X1 port map( A => A(3), B => n19, ZN => S(3));
   U3 : MUX2_X1 port map( A => B, B => n19, S => A(9), Z => S(9));
   U4 : XOR2_X1 port map( A => B, B => A(14), Z => S(14));
   U5 : XOR2_X1 port map( A => B, B => A(21), Z => S(21));
   U6 : XOR2_X1 port map( A => B, B => A(29), Z => S(29));
   U7 : MUX2_X1 port map( A => B, B => n19, S => A(5), Z => S(5));
   U10 : XOR2_X2 port map( A => A(18), B => B, Z => S(18));
   U11 : XOR2_X1 port map( A => A(8), B => B, Z => S(8));
   U15 : XOR2_X1 port map( A => B, B => A(16), Z => S(16));
   U18 : INV_X1 port map( A => B, ZN => n19);
   U19 : INV_X1 port map( A => A(13), ZN => n21);
   U21 : XNOR2_X1 port map( A => A(19), B => n19, ZN => S(19));
   U22 : NAND2_X1 port map( A1 => n16, A2 => n17, ZN => S(10));
   U23 : XOR2_X1 port map( A => B, B => A(25), Z => S(25));
   U24 : XOR2_X1 port map( A => B, B => A(22), Z => S(22));
   U25 : NAND2_X1 port map( A1 => n22, A2 => n23, ZN => S(13));
   U26 : XOR2_X1 port map( A => B, B => A(6), Z => S(6));
   U27 : XOR2_X1 port map( A => B, B => A(17), Z => S(17));
   U28 : XOR2_X1 port map( A => A(2), B => B, Z => S(2));
   U30 : NAND2_X1 port map( A1 => A(10), A2 => n19, ZN => n16);
   U31 : NAND2_X1 port map( A1 => n15, A2 => B, ZN => n17);
   U32 : INV_X1 port map( A => A(10), ZN => n15);
   U33 : OAI21_X2 port map( B1 => A(1), B2 => n19, A => n20, ZN => S(1));
   U34 : XOR2_X1 port map( A => A(11), B => B, Z => S(11));
   U35 : XOR2_X1 port map( A => A(15), B => B, Z => S(15));
   U36 : XOR2_X1 port map( A => A(4), B => B, Z => S(4));
   U37 : XOR2_X1 port map( A => A(7), B => B, Z => S(7));
   U38 : NAND2_X1 port map( A1 => A(1), A2 => n19, ZN => n20);
   U39 : NAND2_X1 port map( A1 => n21, A2 => B, ZN => n22);
   U40 : NAND2_X1 port map( A1 => A(13), A2 => n19, ZN => n23);

end SYN_bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity ff32_en_SIZE5_2 is

   port( D : in std_logic_vector (4 downto 0);  en, clk, rst : in std_logic;  Q
         : out std_logic_vector (4 downto 0));

end ff32_en_SIZE5_2;

architecture SYN_behavioral of ff32_en_SIZE5_2 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n3, n4, n5, n6, net645267, net645268, net645269, net645270, 
      net645271, n13, n14, n15, n16, n17, n18, n19 : std_logic;

begin
   
   Q_reg_4_inst : DFFR_X1 port map( D => n1, CK => clk, RN => n14, Q => Q(4), 
                           QN => net645271);
   Q_reg_3_inst : DFFR_X1 port map( D => n3, CK => clk, RN => n14, Q => Q(3), 
                           QN => net645270);
   Q_reg_2_inst : DFFR_X1 port map( D => n4, CK => clk, RN => n14, Q => Q(2), 
                           QN => net645269);
   Q_reg_1_inst : DFFR_X1 port map( D => n5, CK => clk, RN => n14, Q => Q(1), 
                           QN => net645268);
   Q_reg_0_inst : DFFR_X1 port map( D => n6, CK => clk, RN => n14, Q => Q(0), 
                           QN => net645267);
   U7 : NAND2_X1 port map( A1 => n13, A2 => D(2), ZN => n17);
   U6 : OAI21_X1 port map( B1 => n13, B2 => net645269, A => n17, ZN => n4);
   U9 : NAND2_X1 port map( A1 => n13, A2 => D(3), ZN => n16);
   U8 : OAI21_X1 port map( B1 => n13, B2 => net645270, A => n16, ZN => n3);
   U12 : NAND2_X1 port map( A1 => n13, A2 => D(4), ZN => n15);
   U11 : OAI21_X1 port map( B1 => n13, B2 => net645271, A => n15, ZN => n1);
   U3 : NAND2_X1 port map( A1 => n13, A2 => D(0), ZN => n19);
   U2 : OAI21_X1 port map( B1 => n13, B2 => net645267, A => n19, ZN => n6);
   U5 : NAND2_X1 port map( A1 => n13, A2 => D(1), ZN => n18);
   U4 : OAI21_X1 port map( B1 => n13, B2 => net645268, A => n18, ZN => n5);
   U10 : INV_X1 port map( A => rst, ZN => n14);
   U13 : BUF_X1 port map( A => en, Z => n13);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity ff32_en_SIZE5_1 is

   port( D : in std_logic_vector (4 downto 0);  en, clk, rst : in std_logic;  Q
         : out std_logic_vector (4 downto 0));

end ff32_en_SIZE5_1;

architecture SYN_behavioral of ff32_en_SIZE5_1 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFS_X2
      port( D, CK, SN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFS_X1
      port( D, CK, SN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n7, n9, n13, n14, n19, n20, n21, n22, n23, net684346 : std_logic;

begin
   
   Q_reg_1_inst : DFFR_X1 port map( D => D(1), CK => clk, RN => n19, Q => Q(1),
                           QN => net684346);
   Q_reg_0_inst : DFFS_X1 port map( D => n23, CK => clk, SN => n19, Q => n14, 
                           QN => Q(0));
   Q_reg_3_inst : DFFS_X1 port map( D => n21, CK => clk, SN => n19, Q => n13, 
                           QN => Q(3));
   Q_reg_2_inst : DFFS_X1 port map( D => n22, CK => clk, SN => n19, Q => n9, QN
                           => Q(2));
   Q_reg_4_inst : DFFS_X2 port map( D => n20, CK => clk, SN => n19, Q => n7, QN
                           => Q(4));
   U2 : INV_X1 port map( A => D(0), ZN => n23);
   U3 : INV_X1 port map( A => rst, ZN => n19);
   U4 : INV_X1 port map( A => D(4), ZN => n20);
   U5 : INV_X1 port map( A => D(3), ZN => n21);
   U6 : INV_X1 port map( A => D(2), ZN => n22);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity ff32_en_SIZE32_5 is

   port( D : in std_logic_vector (31 downto 0);  en, clk, rst : in std_logic;  
         Q : out std_logic_vector (31 downto 0));

end ff32_en_SIZE32_5;

architecture SYN_behavioral of ff32_en_SIZE32_5 is

   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
      n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93
      , n94, n95, n97, net645107, net645108, net645109, net645110, net645111, 
      net645112, net645113, net645114, net645115, net645116, net645117, 
      net645118, net645119, net645120, net645121, net645122, net645123, 
      net645124, net645125, net645126, net645127, net645128, net645129, 
      net645130, net645131, net645132, net645133, net645134, net645135, 
      net645136, net645137, net645138, n36, n37, n38, n39, n40, n41, n42, n43, 
      n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58
      , n59, n60, n61, n62, n63, n64, n96, n98, n99, n100 : std_logic;

begin
   
   Q_reg_31_inst : DFFR_X1 port map( D => n97, CK => clk, RN => n36, Q => Q(31)
                           , QN => net645138);
   Q_reg_30_inst : DFFR_X1 port map( D => n95, CK => clk, RN => n36, Q => Q(30)
                           , QN => net645137);
   Q_reg_29_inst : DFFR_X1 port map( D => n94, CK => clk, RN => n36, Q => Q(29)
                           , QN => net645136);
   Q_reg_28_inst : DFFR_X1 port map( D => n93, CK => clk, RN => n36, Q => Q(28)
                           , QN => net645135);
   Q_reg_27_inst : DFFR_X1 port map( D => n92, CK => clk, RN => n36, Q => Q(27)
                           , QN => net645134);
   Q_reg_26_inst : DFFR_X1 port map( D => n91, CK => clk, RN => n36, Q => Q(26)
                           , QN => net645133);
   Q_reg_25_inst : DFFR_X1 port map( D => n90, CK => clk, RN => n36, Q => Q(25)
                           , QN => net645132);
   Q_reg_24_inst : DFFR_X1 port map( D => n89, CK => clk, RN => n36, Q => Q(24)
                           , QN => net645131);
   Q_reg_23_inst : DFFR_X1 port map( D => n88, CK => clk, RN => n36, Q => Q(23)
                           , QN => net645130);
   Q_reg_22_inst : DFFR_X1 port map( D => n87, CK => clk, RN => n36, Q => Q(22)
                           , QN => net645129);
   Q_reg_21_inst : DFFR_X1 port map( D => n86, CK => clk, RN => n36, Q => Q(21)
                           , QN => net645128);
   Q_reg_19_inst : DFFR_X1 port map( D => n84, CK => clk, RN => n36, Q => Q(19)
                           , QN => net645127);
   Q_reg_18_inst : DFFR_X1 port map( D => n83, CK => clk, RN => n36, Q => Q(18)
                           , QN => net645126);
   Q_reg_17_inst : DFFR_X1 port map( D => n82, CK => clk, RN => n36, Q => Q(17)
                           , QN => net645125);
   Q_reg_16_inst : DFFR_X1 port map( D => n81, CK => clk, RN => n36, Q => Q(16)
                           , QN => net645124);
   Q_reg_15_inst : DFFR_X1 port map( D => n80, CK => clk, RN => n36, Q => Q(15)
                           , QN => net645123);
   Q_reg_14_inst : DFFR_X1 port map( D => n79, CK => clk, RN => n36, Q => Q(14)
                           , QN => net645122);
   Q_reg_13_inst : DFFR_X1 port map( D => n78, CK => clk, RN => n36, Q => Q(13)
                           , QN => net645121);
   Q_reg_12_inst : DFFR_X1 port map( D => n77, CK => clk, RN => n36, Q => Q(12)
                           , QN => net645120);
   Q_reg_11_inst : DFFR_X1 port map( D => n76, CK => clk, RN => n36, Q => Q(11)
                           , QN => net645119);
   Q_reg_10_inst : DFFR_X1 port map( D => n75, CK => clk, RN => n36, Q => Q(10)
                           , QN => net645118);
   Q_reg_9_inst : DFFR_X1 port map( D => n74, CK => clk, RN => n36, Q => Q(9), 
                           QN => net645117);
   Q_reg_8_inst : DFFR_X1 port map( D => n73, CK => clk, RN => n36, Q => Q(8), 
                           QN => net645116);
   Q_reg_7_inst : DFFR_X1 port map( D => n72, CK => clk, RN => n36, Q => Q(7), 
                           QN => net645115);
   Q_reg_6_inst : DFFR_X1 port map( D => n71, CK => clk, RN => n36, Q => Q(6), 
                           QN => net645114);
   Q_reg_5_inst : DFFR_X1 port map( D => n70, CK => clk, RN => n36, Q => Q(5), 
                           QN => net645113);
   Q_reg_4_inst : DFFR_X1 port map( D => n69, CK => clk, RN => n36, Q => Q(4), 
                           QN => net645112);
   Q_reg_3_inst : DFFR_X1 port map( D => n68, CK => clk, RN => n36, Q => Q(3), 
                           QN => net645111);
   Q_reg_2_inst : DFFR_X1 port map( D => n67, CK => clk, RN => n36, Q => Q(2), 
                           QN => net645110);
   Q_reg_1_inst : DFFR_X1 port map( D => n66, CK => clk, RN => n36, Q => Q(1), 
                           QN => net645109);
   Q_reg_0_inst : DFFR_X1 port map( D => n65, CK => clk, RN => n36, Q => Q(0), 
                           QN => net645108);
   Q_reg_20_inst : DFFR_X1 port map( D => n85, CK => clk, RN => n36, Q => Q(20)
                           , QN => net645107);
   U43 : NAND2_X1 port map( A1 => en, A2 => D(11), ZN => n48);
   U42 : OAI21_X1 port map( B1 => en, B2 => net645119, A => n48, ZN => n76);
   U45 : NAND2_X1 port map( A1 => en, A2 => D(10), ZN => n47);
   U44 : OAI21_X1 port map( B1 => en, B2 => net645118, A => n47, ZN => n75);
   U37 : NAND2_X1 port map( A1 => en, A2 => D(14), ZN => n51);
   U36 : OAI21_X1 port map( B1 => en, B2 => net645122, A => n51, ZN => n79);
   U39 : NAND2_X1 port map( A1 => en, A2 => D(13), ZN => n50);
   U38 : OAI21_X1 port map( B1 => en, B2 => net645121, A => n50, ZN => n78);
   U55 : NAND2_X1 port map( A1 => en, A2 => D(5), ZN => n42);
   U54 : OAI21_X1 port map( B1 => en, B2 => net645113, A => n42, ZN => n70);
   U57 : NAND2_X1 port map( A1 => en, A2 => D(4), ZN => n41);
   U56 : OAI21_X1 port map( B1 => en, B2 => net645112, A => n41, ZN => n69);
   U13 : NAND2_X1 port map( A1 => en, A2 => D(26), ZN => n63);
   U12 : OAI21_X1 port map( B1 => en, B2 => net645133, A => n63, ZN => n91);
   U49 : NAND2_X1 port map( A1 => en, A2 => D(8), ZN => n45);
   U48 : OAI21_X1 port map( B1 => en, B2 => net645116, A => n45, ZN => n73);
   U23 : NAND2_X1 port map( A1 => en, A2 => D(21), ZN => n58);
   U22 : OAI21_X1 port map( B1 => en, B2 => net645128, A => n58, ZN => n86);
   U61 : NAND2_X1 port map( A1 => en, A2 => D(2), ZN => n39);
   U60 : OAI21_X1 port map( B1 => en, B2 => net645110, A => n39, ZN => n67);
   U59 : NAND2_X1 port map( A1 => en, A2 => D(3), ZN => n40);
   U58 : OAI21_X1 port map( B1 => en, B2 => net645111, A => n40, ZN => n68);
   U53 : NAND2_X1 port map( A1 => en, A2 => D(6), ZN => n43);
   U52 : OAI21_X1 port map( B1 => en, B2 => net645114, A => n43, ZN => n71);
   U21 : NAND2_X1 port map( A1 => en, A2 => D(22), ZN => n59);
   U20 : OAI21_X1 port map( B1 => en, B2 => net645129, A => n59, ZN => n87);
   U17 : NAND2_X1 port map( A1 => en, A2 => D(24), ZN => n61);
   U16 : OAI21_X1 port map( B1 => en, B2 => net645131, A => n61, ZN => n89);
   U25 : NAND2_X1 port map( A1 => en, A2 => D(20), ZN => n57);
   U24 : OAI21_X1 port map( B1 => en, B2 => net645107, A => n57, ZN => n85);
   U27 : NAND2_X1 port map( A1 => en, A2 => D(19), ZN => n56);
   U26 : OAI21_X1 port map( B1 => en, B2 => net645127, A => n56, ZN => n84);
   U51 : NAND2_X1 port map( A1 => en, A2 => D(7), ZN => n44);
   U50 : OAI21_X1 port map( B1 => en, B2 => net645115, A => n44, ZN => n72);
   U7 : NAND2_X1 port map( A1 => en, A2 => D(29), ZN => n98);
   U6 : OAI21_X1 port map( B1 => en, B2 => net645136, A => n98, ZN => n94);
   U9 : NAND2_X1 port map( A1 => en, A2 => D(28), ZN => n96);
   U8 : OAI21_X1 port map( B1 => en, B2 => net645135, A => n96, ZN => n93);
   U11 : NAND2_X1 port map( A1 => en, A2 => D(27), ZN => n64);
   U10 : OAI21_X1 port map( B1 => en, B2 => net645134, A => n64, ZN => n92);
   U19 : NAND2_X1 port map( A1 => en, A2 => D(23), ZN => n60);
   U18 : OAI21_X1 port map( B1 => en, B2 => net645130, A => n60, ZN => n88);
   U15 : NAND2_X1 port map( A1 => en, A2 => D(25), ZN => n62);
   U14 : OAI21_X1 port map( B1 => en, B2 => net645132, A => n62, ZN => n90);
   U35 : NAND2_X1 port map( A1 => en, A2 => D(15), ZN => n52);
   U34 : OAI21_X1 port map( B1 => en, B2 => net645123, A => n52, ZN => n80);
   U33 : NAND2_X1 port map( A1 => en, A2 => D(16), ZN => n53);
   U32 : OAI21_X1 port map( B1 => en, B2 => net645124, A => n53, ZN => n81);
   U31 : NAND2_X1 port map( A1 => en, A2 => D(17), ZN => n54);
   U30 : OAI21_X1 port map( B1 => en, B2 => net645125, A => n54, ZN => n82);
   U29 : NAND2_X1 port map( A1 => en, A2 => D(18), ZN => n55);
   U28 : OAI21_X1 port map( B1 => en, B2 => net645126, A => n55, ZN => n83);
   U47 : NAND2_X1 port map( A1 => en, A2 => D(9), ZN => n46);
   U46 : OAI21_X1 port map( B1 => en, B2 => net645117, A => n46, ZN => n74);
   U41 : NAND2_X1 port map( A1 => en, A2 => D(12), ZN => n49);
   U40 : OAI21_X1 port map( B1 => en, B2 => net645120, A => n49, ZN => n77);
   U63 : NAND2_X1 port map( A1 => en, A2 => D(1), ZN => n38);
   U62 : OAI21_X1 port map( B1 => en, B2 => net645109, A => n38, ZN => n66);
   U65 : NAND2_X1 port map( A1 => en, A2 => D(0), ZN => n37);
   U64 : OAI21_X1 port map( B1 => en, B2 => net645108, A => n37, ZN => n65);
   U3 : NAND2_X1 port map( A1 => en, A2 => D(31), ZN => n100);
   U2 : OAI21_X1 port map( B1 => en, B2 => net645138, A => n100, ZN => n97);
   U5 : NAND2_X1 port map( A1 => en, A2 => D(30), ZN => n99);
   U4 : OAI21_X1 port map( B1 => en, B2 => net645137, A => n99, ZN => n95);
   U66 : INV_X2 port map( A => rst, ZN => n36);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity ff32_en_SIZE32_4 is

   port( D : in std_logic_vector (31 downto 0);  en, clk, rst : in std_logic;  
         Q : out std_logic_vector (31 downto 0));

end ff32_en_SIZE32_4;

architecture SYN_behavioral of ff32_en_SIZE32_4 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
      n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93
      , n94, n95, n97, net645107, net645108, net645109, net645110, net645111, 
      net645112, net645113, net645114, net645115, net645116, net645117, 
      net645118, net645119, net645120, net645121, net645122, net645123, 
      net645124, net645125, net645126, net645127, net645128, net645129, 
      net645130, net645131, net645132, net645133, net645134, net645135, 
      net645136, net645137, net645138, n36, n37, n38, n39, n40, n41, n42, n43, 
      n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58
      , n59, n60, n61, n62, n63, n64, n96, n98, n99, n100, n101, n102, n103, 
      n104 : std_logic;

begin
   
   Q_reg_31_inst : DFFR_X1 port map( D => n97, CK => clk, RN => n40, Q => Q(31)
                           , QN => net645138);
   Q_reg_30_inst : DFFR_X1 port map( D => n95, CK => clk, RN => n40, Q => Q(30)
                           , QN => net645137);
   Q_reg_29_inst : DFFR_X1 port map( D => n94, CK => clk, RN => n40, Q => Q(29)
                           , QN => net645136);
   Q_reg_28_inst : DFFR_X1 port map( D => n93, CK => clk, RN => n40, Q => Q(28)
                           , QN => net645135);
   Q_reg_27_inst : DFFR_X1 port map( D => n92, CK => clk, RN => n40, Q => Q(27)
                           , QN => net645134);
   Q_reg_26_inst : DFFR_X1 port map( D => n91, CK => clk, RN => n40, Q => Q(26)
                           , QN => net645133);
   Q_reg_25_inst : DFFR_X1 port map( D => n90, CK => clk, RN => n40, Q => Q(25)
                           , QN => net645132);
   Q_reg_24_inst : DFFR_X1 port map( D => n89, CK => clk, RN => n40, Q => Q(24)
                           , QN => net645131);
   Q_reg_23_inst : DFFR_X1 port map( D => n88, CK => clk, RN => n40, Q => Q(23)
                           , QN => net645130);
   Q_reg_22_inst : DFFR_X1 port map( D => n87, CK => clk, RN => n40, Q => Q(22)
                           , QN => net645129);
   Q_reg_21_inst : DFFR_X1 port map( D => n86, CK => clk, RN => n40, Q => Q(21)
                           , QN => net645128);
   Q_reg_19_inst : DFFR_X1 port map( D => n84, CK => clk, RN => n40, Q => Q(19)
                           , QN => net645127);
   Q_reg_18_inst : DFFR_X1 port map( D => n83, CK => clk, RN => n40, Q => Q(18)
                           , QN => net645126);
   Q_reg_17_inst : DFFR_X1 port map( D => n82, CK => clk, RN => n40, Q => Q(17)
                           , QN => net645125);
   Q_reg_16_inst : DFFR_X1 port map( D => n81, CK => clk, RN => n40, Q => Q(16)
                           , QN => net645124);
   Q_reg_15_inst : DFFR_X1 port map( D => n80, CK => clk, RN => n40, Q => Q(15)
                           , QN => net645123);
   Q_reg_14_inst : DFFR_X1 port map( D => n79, CK => clk, RN => n40, Q => Q(14)
                           , QN => net645122);
   Q_reg_13_inst : DFFR_X1 port map( D => n78, CK => clk, RN => n40, Q => Q(13)
                           , QN => net645121);
   Q_reg_12_inst : DFFR_X1 port map( D => n77, CK => clk, RN => n40, Q => Q(12)
                           , QN => net645120);
   Q_reg_11_inst : DFFR_X1 port map( D => n76, CK => clk, RN => n40, Q => Q(11)
                           , QN => net645119);
   Q_reg_10_inst : DFFR_X1 port map( D => n75, CK => clk, RN => n40, Q => Q(10)
                           , QN => net645118);
   Q_reg_9_inst : DFFR_X1 port map( D => n74, CK => clk, RN => n40, Q => Q(9), 
                           QN => net645117);
   Q_reg_8_inst : DFFR_X1 port map( D => n73, CK => clk, RN => n40, Q => Q(8), 
                           QN => net645116);
   Q_reg_7_inst : DFFR_X1 port map( D => n72, CK => clk, RN => n40, Q => Q(7), 
                           QN => net645115);
   Q_reg_6_inst : DFFR_X1 port map( D => n71, CK => clk, RN => n40, Q => Q(6), 
                           QN => net645114);
   Q_reg_5_inst : DFFR_X1 port map( D => n70, CK => clk, RN => n40, Q => Q(5), 
                           QN => net645113);
   Q_reg_4_inst : DFFR_X1 port map( D => n69, CK => clk, RN => n40, Q => Q(4), 
                           QN => net645112);
   Q_reg_3_inst : DFFR_X1 port map( D => n68, CK => clk, RN => n40, Q => Q(3), 
                           QN => net645111);
   Q_reg_2_inst : DFFR_X1 port map( D => n67, CK => clk, RN => n40, Q => Q(2), 
                           QN => net645110);
   Q_reg_1_inst : DFFR_X1 port map( D => n66, CK => clk, RN => n40, Q => Q(1), 
                           QN => net645109);
   Q_reg_0_inst : DFFR_X1 port map( D => n65, CK => clk, RN => n40, Q => Q(0), 
                           QN => net645108);
   Q_reg_20_inst : DFFR_X1 port map( D => n85, CK => clk, RN => n40, Q => Q(20)
                           , QN => net645107);
   U39 : NAND2_X1 port map( A1 => n39, A2 => D(13), ZN => n54);
   U38 : OAI21_X1 port map( B1 => n37, B2 => net645121, A => n54, ZN => n78);
   U3 : NAND2_X1 port map( A1 => n39, A2 => D(31), ZN => n104);
   U2 : OAI21_X1 port map( B1 => n37, B2 => net645138, A => n104, ZN => n97);
   U43 : NAND2_X1 port map( A1 => n39, A2 => D(11), ZN => n52);
   U42 : OAI21_X1 port map( B1 => n37, B2 => net645119, A => n52, ZN => n76);
   U63 : NAND2_X1 port map( A1 => n39, A2 => D(1), ZN => n42);
   U62 : OAI21_X1 port map( B1 => n36, B2 => net645109, A => n42, ZN => n66);
   U5 : NAND2_X1 port map( A1 => n39, A2 => D(30), ZN => n103);
   U4 : OAI21_X1 port map( B1 => n36, B2 => net645137, A => n103, ZN => n95);
   U45 : NAND2_X1 port map( A1 => n39, A2 => D(10), ZN => n51);
   U44 : OAI21_X1 port map( B1 => n37, B2 => net645118, A => n51, ZN => n75);
   U37 : NAND2_X1 port map( A1 => n39, A2 => D(14), ZN => n55);
   U36 : OAI21_X1 port map( B1 => n37, B2 => net645122, A => n55, ZN => n79);
   U33 : NAND2_X1 port map( A1 => en, A2 => D(16), ZN => n57);
   U32 : OAI21_X1 port map( B1 => n37, B2 => net645124, A => n57, ZN => n81);
   U27 : NAND2_X1 port map( A1 => en, A2 => D(19), ZN => n60);
   U26 : OAI21_X1 port map( B1 => n36, B2 => net645127, A => n60, ZN => n84);
   U41 : NAND2_X1 port map( A1 => en, A2 => D(12), ZN => n53);
   U40 : OAI21_X1 port map( B1 => n37, B2 => net645120, A => n53, ZN => n77);
   U19 : NAND2_X1 port map( A1 => n38, A2 => D(23), ZN => n64);
   U18 : OAI21_X1 port map( B1 => n36, B2 => net645130, A => n64, ZN => n88);
   U9 : NAND2_X1 port map( A1 => n38, A2 => D(28), ZN => n101);
   U8 : OAI21_X1 port map( B1 => n36, B2 => net645135, A => n101, ZN => n93);
   U23 : NAND2_X1 port map( A1 => n38, A2 => D(21), ZN => n62);
   U22 : OAI21_X1 port map( B1 => n36, B2 => net645128, A => n62, ZN => n86);
   U31 : NAND2_X1 port map( A1 => en, A2 => D(17), ZN => n58);
   U30 : OAI21_X1 port map( B1 => n37, B2 => net645125, A => n58, ZN => n82);
   U17 : NAND2_X1 port map( A1 => n38, A2 => D(24), ZN => n96);
   U16 : OAI21_X1 port map( B1 => n36, B2 => net645131, A => n96, ZN => n89);
   U29 : NAND2_X1 port map( A1 => en, A2 => D(18), ZN => n59);
   U28 : OAI21_X1 port map( B1 => n37, B2 => net645126, A => n59, ZN => n83);
   U21 : NAND2_X1 port map( A1 => en, A2 => D(22), ZN => n63);
   U20 : OAI21_X1 port map( B1 => n36, B2 => net645129, A => n63, ZN => n87);
   U61 : NAND2_X1 port map( A1 => n38, A2 => D(2), ZN => n43);
   U60 : OAI21_X1 port map( B1 => n37, B2 => net645110, A => n43, ZN => n67);
   U51 : NAND2_X1 port map( A1 => en, A2 => D(7), ZN => n48);
   U50 : OAI21_X1 port map( B1 => n37, B2 => net645115, A => n48, ZN => n72);
   U7 : NAND2_X1 port map( A1 => n38, A2 => D(29), ZN => n102);
   U6 : OAI21_X1 port map( B1 => n36, B2 => net645136, A => n102, ZN => n94);
   U49 : NAND2_X1 port map( A1 => en, A2 => D(8), ZN => n49);
   U48 : OAI21_X1 port map( B1 => n36, B2 => net645116, A => n49, ZN => n73);
   U25 : NAND2_X1 port map( A1 => en, A2 => D(20), ZN => n61);
   U24 : OAI21_X1 port map( B1 => n36, B2 => net645107, A => n61, ZN => n85);
   U13 : NAND2_X1 port map( A1 => n38, A2 => D(26), ZN => n99);
   U12 : OAI21_X1 port map( B1 => n36, B2 => net645133, A => n99, ZN => n91);
   U15 : NAND2_X1 port map( A1 => n38, A2 => D(25), ZN => n98);
   U14 : OAI21_X1 port map( B1 => n36, B2 => net645132, A => n98, ZN => n90);
   U11 : NAND2_X1 port map( A1 => n38, A2 => D(27), ZN => n100);
   U10 : OAI21_X1 port map( B1 => n36, B2 => net645134, A => n100, ZN => n92);
   U35 : NAND2_X1 port map( A1 => en, A2 => D(15), ZN => n56);
   U34 : OAI21_X1 port map( B1 => n37, B2 => net645123, A => n56, ZN => n80);
   U53 : NAND2_X1 port map( A1 => n38, A2 => D(6), ZN => n47);
   U52 : OAI21_X1 port map( B1 => n37, B2 => net645114, A => n47, ZN => n71);
   U47 : NAND2_X1 port map( A1 => en, A2 => D(9), ZN => n50);
   U46 : OAI21_X1 port map( B1 => n37, B2 => net645117, A => n50, ZN => n74);
   U65 : NAND2_X1 port map( A1 => n39, A2 => D(0), ZN => n41);
   U64 : OAI21_X1 port map( B1 => n39, B2 => net645108, A => n41, ZN => n65);
   U57 : NAND2_X1 port map( A1 => n38, A2 => D(4), ZN => n45);
   U56 : OAI21_X1 port map( B1 => n39, B2 => net645112, A => n45, ZN => n69);
   U59 : NAND2_X1 port map( A1 => n38, A2 => D(3), ZN => n44);
   U58 : OAI21_X1 port map( B1 => n39, B2 => net645111, A => n44, ZN => n68);
   U55 : NAND2_X1 port map( A1 => en, A2 => D(5), ZN => n46);
   U54 : OAI21_X1 port map( B1 => n39, B2 => net645113, A => n46, ZN => n70);
   U66 : INV_X2 port map( A => rst, ZN => n40);
   U67 : BUF_X1 port map( A => en, Z => n36);
   U68 : BUF_X1 port map( A => en, Z => n37);
   U69 : BUF_X1 port map( A => en, Z => n38);
   U70 : BUF_X1 port map( A => en, Z => n39);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity ff32_en_SIZE32_3 is

   port( D : in std_logic_vector (31 downto 0);  en, clk, rst : in std_logic;  
         Q : out std_logic_vector (31 downto 0));

end ff32_en_SIZE32_3;

architecture SYN_behavioral of ff32_en_SIZE32_3 is

   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal net645107, net645108, net645109, net645110, net645111, net645112, 
      net645113, net645114, net645115, net645116, net645117, net645118, 
      net645119, net645120, net645121, net645122, net645123, net645124, 
      net645125, net645126, net645127, net645128, net645129, net645130, 
      net645131, net645132, net645133, net645134, net645135, net645136, 
      net645137, net645138, n35 : std_logic;

begin
   
   Q_reg_31_inst : DFFR_X1 port map( D => D(31), CK => clk, RN => n35, Q => 
                           Q(31), QN => net645138);
   Q_reg_30_inst : DFFR_X1 port map( D => D(30), CK => clk, RN => n35, Q => 
                           Q(30), QN => net645137);
   Q_reg_29_inst : DFFR_X1 port map( D => D(29), CK => clk, RN => n35, Q => 
                           Q(29), QN => net645136);
   Q_reg_28_inst : DFFR_X1 port map( D => D(28), CK => clk, RN => n35, Q => 
                           Q(28), QN => net645135);
   Q_reg_27_inst : DFFR_X1 port map( D => D(27), CK => clk, RN => n35, Q => 
                           Q(27), QN => net645134);
   Q_reg_26_inst : DFFR_X1 port map( D => D(26), CK => clk, RN => n35, Q => 
                           Q(26), QN => net645133);
   Q_reg_25_inst : DFFR_X1 port map( D => D(25), CK => clk, RN => n35, Q => 
                           Q(25), QN => net645132);
   Q_reg_24_inst : DFFR_X1 port map( D => D(24), CK => clk, RN => n35, Q => 
                           Q(24), QN => net645131);
   Q_reg_23_inst : DFFR_X1 port map( D => D(23), CK => clk, RN => n35, Q => 
                           Q(23), QN => net645130);
   Q_reg_22_inst : DFFR_X1 port map( D => D(22), CK => clk, RN => n35, Q => 
                           Q(22), QN => net645129);
   Q_reg_21_inst : DFFR_X1 port map( D => D(21), CK => clk, RN => n35, Q => 
                           Q(21), QN => net645128);
   Q_reg_19_inst : DFFR_X1 port map( D => D(19), CK => clk, RN => n35, Q => 
                           Q(19), QN => net645127);
   Q_reg_18_inst : DFFR_X1 port map( D => D(18), CK => clk, RN => n35, Q => 
                           Q(18), QN => net645126);
   Q_reg_17_inst : DFFR_X1 port map( D => D(17), CK => clk, RN => n35, Q => 
                           Q(17), QN => net645125);
   Q_reg_16_inst : DFFR_X1 port map( D => D(16), CK => clk, RN => n35, Q => 
                           Q(16), QN => net645124);
   Q_reg_15_inst : DFFR_X1 port map( D => D(15), CK => clk, RN => n35, Q => 
                           Q(15), QN => net645123);
   Q_reg_14_inst : DFFR_X1 port map( D => D(14), CK => clk, RN => n35, Q => 
                           Q(14), QN => net645122);
   Q_reg_13_inst : DFFR_X1 port map( D => D(13), CK => clk, RN => n35, Q => 
                           Q(13), QN => net645121);
   Q_reg_12_inst : DFFR_X1 port map( D => D(12), CK => clk, RN => n35, Q => 
                           Q(12), QN => net645120);
   Q_reg_11_inst : DFFR_X1 port map( D => D(11), CK => clk, RN => n35, Q => 
                           Q(11), QN => net645119);
   Q_reg_10_inst : DFFR_X1 port map( D => D(10), CK => clk, RN => n35, Q => 
                           Q(10), QN => net645118);
   Q_reg_9_inst : DFFR_X1 port map( D => D(9), CK => clk, RN => n35, Q => Q(9),
                           QN => net645117);
   Q_reg_8_inst : DFFR_X1 port map( D => D(8), CK => clk, RN => n35, Q => Q(8),
                           QN => net645116);
   Q_reg_7_inst : DFFR_X1 port map( D => D(7), CK => clk, RN => n35, Q => Q(7),
                           QN => net645115);
   Q_reg_6_inst : DFFR_X1 port map( D => D(6), CK => clk, RN => n35, Q => Q(6),
                           QN => net645114);
   Q_reg_5_inst : DFFR_X1 port map( D => D(5), CK => clk, RN => n35, Q => Q(5),
                           QN => net645113);
   Q_reg_4_inst : DFFR_X1 port map( D => D(4), CK => clk, RN => n35, Q => Q(4),
                           QN => net645112);
   Q_reg_3_inst : DFFR_X1 port map( D => D(3), CK => clk, RN => n35, Q => Q(3),
                           QN => net645111);
   Q_reg_2_inst : DFFR_X1 port map( D => D(2), CK => clk, RN => n35, Q => Q(2),
                           QN => net645110);
   Q_reg_1_inst : DFFR_X1 port map( D => D(1), CK => clk, RN => n35, Q => Q(1),
                           QN => net645109);
   Q_reg_0_inst : DFFR_X1 port map( D => D(0), CK => clk, RN => n35, Q => Q(0),
                           QN => net645108);
   Q_reg_20_inst : DFFR_X1 port map( D => D(20), CK => clk, RN => n35, Q => 
                           Q(20), QN => net645107);
   U2 : INV_X2 port map( A => rst, ZN => n35);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity ff32_en_SIZE32_2 is

   port( D : in std_logic_vector (31 downto 0);  en, clk, rst : in std_logic;  
         Q : out std_logic_vector (31 downto 0));

end ff32_en_SIZE32_2;

architecture SYN_behavioral of ff32_en_SIZE32_2 is

   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal net645107, net645108, net645109, net645110, net645111, net645112, 
      net645113, net645114, net645115, net645116, net645117, net645118, 
      net645119, net645120, net645121, net645122, net645123, net645124, 
      net645125, net645126, net645127, net645128, net645129, net645130, 
      net645131, net645132, net645133, net645134, net645135, net645136, 
      net645137, net645138, n37 : std_logic;

begin
   
   Q_reg_31_inst : DFFR_X1 port map( D => D(31), CK => clk, RN => n37, Q => 
                           Q(31), QN => net645138);
   Q_reg_30_inst : DFFR_X1 port map( D => D(30), CK => clk, RN => n37, Q => 
                           Q(30), QN => net645137);
   Q_reg_29_inst : DFFR_X1 port map( D => D(29), CK => clk, RN => n37, Q => 
                           Q(29), QN => net645136);
   Q_reg_28_inst : DFFR_X1 port map( D => D(28), CK => clk, RN => n37, Q => 
                           Q(28), QN => net645135);
   Q_reg_27_inst : DFFR_X1 port map( D => D(27), CK => clk, RN => n37, Q => 
                           Q(27), QN => net645134);
   Q_reg_26_inst : DFFR_X1 port map( D => D(26), CK => clk, RN => n37, Q => 
                           Q(26), QN => net645133);
   Q_reg_25_inst : DFFR_X1 port map( D => D(25), CK => clk, RN => n37, Q => 
                           Q(25), QN => net645132);
   Q_reg_24_inst : DFFR_X1 port map( D => D(24), CK => clk, RN => n37, Q => 
                           Q(24), QN => net645131);
   Q_reg_23_inst : DFFR_X1 port map( D => D(23), CK => clk, RN => n37, Q => 
                           Q(23), QN => net645130);
   Q_reg_22_inst : DFFR_X1 port map( D => D(22), CK => clk, RN => n37, Q => 
                           Q(22), QN => net645129);
   Q_reg_21_inst : DFFR_X1 port map( D => D(21), CK => clk, RN => n37, Q => 
                           Q(21), QN => net645128);
   Q_reg_19_inst : DFFR_X1 port map( D => D(19), CK => clk, RN => n37, Q => 
                           Q(19), QN => net645127);
   Q_reg_18_inst : DFFR_X1 port map( D => D(18), CK => clk, RN => n37, Q => 
                           Q(18), QN => net645126);
   Q_reg_17_inst : DFFR_X1 port map( D => D(17), CK => clk, RN => n37, Q => 
                           Q(17), QN => net645125);
   Q_reg_16_inst : DFFR_X1 port map( D => D(16), CK => clk, RN => n37, Q => 
                           Q(16), QN => net645124);
   Q_reg_15_inst : DFFR_X1 port map( D => D(15), CK => clk, RN => n37, Q => 
                           Q(15), QN => net645123);
   Q_reg_14_inst : DFFR_X1 port map( D => D(14), CK => clk, RN => n37, Q => 
                           Q(14), QN => net645122);
   Q_reg_13_inst : DFFR_X1 port map( D => D(13), CK => clk, RN => n37, Q => 
                           Q(13), QN => net645121);
   Q_reg_12_inst : DFFR_X1 port map( D => D(12), CK => clk, RN => n37, Q => 
                           Q(12), QN => net645120);
   Q_reg_11_inst : DFFR_X1 port map( D => D(11), CK => clk, RN => n37, Q => 
                           Q(11), QN => net645119);
   Q_reg_10_inst : DFFR_X1 port map( D => D(10), CK => clk, RN => n37, Q => 
                           Q(10), QN => net645118);
   Q_reg_9_inst : DFFR_X1 port map( D => D(9), CK => clk, RN => n37, Q => Q(9),
                           QN => net645117);
   Q_reg_8_inst : DFFR_X1 port map( D => D(8), CK => clk, RN => n37, Q => Q(8),
                           QN => net645116);
   Q_reg_7_inst : DFFR_X1 port map( D => D(7), CK => clk, RN => n37, Q => Q(7),
                           QN => net645115);
   Q_reg_6_inst : DFFR_X1 port map( D => D(6), CK => clk, RN => n37, Q => Q(6),
                           QN => net645114);
   Q_reg_5_inst : DFFR_X1 port map( D => D(5), CK => clk, RN => n37, Q => Q(5),
                           QN => net645113);
   Q_reg_4_inst : DFFR_X1 port map( D => D(4), CK => clk, RN => n37, Q => Q(4),
                           QN => net645112);
   Q_reg_3_inst : DFFR_X1 port map( D => D(3), CK => clk, RN => n37, Q => Q(3),
                           QN => net645111);
   Q_reg_2_inst : DFFR_X1 port map( D => D(2), CK => clk, RN => n37, Q => Q(2),
                           QN => net645110);
   Q_reg_1_inst : DFFR_X1 port map( D => D(1), CK => clk, RN => n37, Q => Q(1),
                           QN => net645109);
   Q_reg_0_inst : DFFR_X1 port map( D => D(0), CK => clk, RN => n37, Q => Q(0),
                           QN => net645108);
   Q_reg_20_inst : DFFR_X1 port map( D => D(20), CK => clk, RN => n37, Q => 
                           Q(20), QN => net645107);
   U2 : INV_X2 port map( A => rst, ZN => n37);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity ff32_en_SIZE32_1 is

   port( D : in std_logic_vector (31 downto 0);  en, clk, rst : in std_logic;  
         Q : out std_logic_vector (31 downto 0));

end ff32_en_SIZE32_1;

architecture SYN_behavioral of ff32_en_SIZE32_1 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
      n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93
      , n94, n95, n97, net645107, net645108, net645109, net645110, net645111, 
      net645112, net645113, net645114, net645115, net645116, net645117, 
      net645118, net645119, net645120, net645121, net645122, net645123, 
      net645124, net645125, net645126, net645127, net645128, net645129, 
      net645130, net645131, net645132, net645133, net645134, net645135, 
      net645136, net645137, net645138, n35, n36, n38, n39, n40, n41, n42, n43, 
      n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58
      , n59, n60, n61, n62, n63, n64, n96, n98, n99, n100, n101 : std_logic;

begin
   
   Q_reg_31_inst : DFFR_X1 port map( D => n97, CK => clk, RN => n39, Q => Q(31)
                           , QN => net645138);
   Q_reg_30_inst : DFFR_X1 port map( D => n95, CK => clk, RN => n39, Q => Q(30)
                           , QN => net645137);
   Q_reg_29_inst : DFFR_X1 port map( D => n94, CK => clk, RN => n39, Q => Q(29)
                           , QN => net645136);
   Q_reg_28_inst : DFFR_X1 port map( D => n93, CK => clk, RN => n39, Q => Q(28)
                           , QN => net645135);
   Q_reg_27_inst : DFFR_X1 port map( D => n92, CK => clk, RN => n39, Q => Q(27)
                           , QN => net645134);
   Q_reg_26_inst : DFFR_X1 port map( D => n91, CK => clk, RN => n39, Q => Q(26)
                           , QN => net645133);
   Q_reg_25_inst : DFFR_X1 port map( D => n90, CK => clk, RN => n39, Q => Q(25)
                           , QN => net645132);
   Q_reg_24_inst : DFFR_X1 port map( D => n89, CK => clk, RN => n39, Q => Q(24)
                           , QN => net645131);
   Q_reg_23_inst : DFFR_X1 port map( D => n88, CK => clk, RN => n39, Q => Q(23)
                           , QN => net645130);
   Q_reg_22_inst : DFFR_X1 port map( D => n87, CK => clk, RN => n39, Q => Q(22)
                           , QN => net645129);
   Q_reg_21_inst : DFFR_X1 port map( D => n86, CK => clk, RN => n39, Q => Q(21)
                           , QN => net645128);
   Q_reg_19_inst : DFFR_X1 port map( D => n84, CK => clk, RN => n39, Q => Q(19)
                           , QN => net645127);
   Q_reg_18_inst : DFFR_X1 port map( D => n83, CK => clk, RN => n39, Q => Q(18)
                           , QN => net645126);
   Q_reg_17_inst : DFFR_X1 port map( D => n82, CK => clk, RN => n39, Q => Q(17)
                           , QN => net645125);
   Q_reg_16_inst : DFFR_X1 port map( D => n81, CK => clk, RN => n39, Q => Q(16)
                           , QN => net645124);
   Q_reg_15_inst : DFFR_X1 port map( D => n80, CK => clk, RN => n39, Q => Q(15)
                           , QN => net645123);
   Q_reg_14_inst : DFFR_X1 port map( D => n79, CK => clk, RN => n39, Q => Q(14)
                           , QN => net645122);
   Q_reg_13_inst : DFFR_X1 port map( D => n78, CK => clk, RN => n39, Q => Q(13)
                           , QN => net645121);
   Q_reg_12_inst : DFFR_X1 port map( D => n77, CK => clk, RN => n39, Q => Q(12)
                           , QN => net645120);
   Q_reg_11_inst : DFFR_X1 port map( D => n76, CK => clk, RN => n39, Q => Q(11)
                           , QN => net645119);
   Q_reg_10_inst : DFFR_X1 port map( D => n75, CK => clk, RN => n39, Q => Q(10)
                           , QN => net645118);
   Q_reg_9_inst : DFFR_X1 port map( D => n74, CK => clk, RN => n39, Q => Q(9), 
                           QN => net645117);
   Q_reg_8_inst : DFFR_X1 port map( D => n73, CK => clk, RN => n39, Q => Q(8), 
                           QN => net645116);
   Q_reg_7_inst : DFFR_X1 port map( D => n72, CK => clk, RN => n39, Q => Q(7), 
                           QN => net645115);
   Q_reg_6_inst : DFFR_X1 port map( D => n71, CK => clk, RN => n39, Q => Q(6), 
                           QN => net645114);
   Q_reg_5_inst : DFFR_X1 port map( D => n70, CK => clk, RN => n39, Q => Q(5), 
                           QN => net645113);
   Q_reg_4_inst : DFFR_X1 port map( D => n69, CK => clk, RN => n39, Q => Q(4), 
                           QN => net645112);
   Q_reg_3_inst : DFFR_X1 port map( D => n68, CK => clk, RN => n39, Q => Q(3), 
                           QN => net645111);
   Q_reg_2_inst : DFFR_X1 port map( D => n67, CK => clk, RN => n39, Q => Q(2), 
                           QN => net645110);
   Q_reg_1_inst : DFFR_X1 port map( D => n66, CK => clk, RN => n39, Q => Q(1), 
                           QN => net645109);
   Q_reg_0_inst : DFFR_X1 port map( D => n65, CK => clk, RN => n39, Q => Q(0), 
                           QN => net645108);
   Q_reg_20_inst : DFFR_X1 port map( D => n85, CK => clk, RN => n39, Q => Q(20)
                           , QN => net645107);
   U3 : NAND2_X1 port map( A1 => en, A2 => D(31), ZN => n101);
   U2 : OAI21_X1 port map( B1 => en, B2 => net645138, A => n101, ZN => n97);
   U19 : NAND2_X1 port map( A1 => en, A2 => D(23), ZN => n62);
   U18 : OAI21_X1 port map( B1 => en, B2 => net645130, A => n62, ZN => n88);
   U11 : NAND2_X1 port map( A1 => en, A2 => D(27), ZN => n98);
   U10 : OAI21_X1 port map( B1 => en, B2 => net645134, A => n98, ZN => n92);
   U21 : NAND2_X1 port map( A1 => en, A2 => D(22), ZN => n61);
   U20 : OAI21_X1 port map( B1 => n38, B2 => net645129, A => n61, ZN => n87);
   U13 : NAND2_X1 port map( A1 => en, A2 => D(26), ZN => n96);
   U12 : OAI21_X1 port map( B1 => en, B2 => net645133, A => n96, ZN => n91);
   U7 : NAND2_X1 port map( A1 => en, A2 => D(29), ZN => n100);
   U6 : OAI21_X1 port map( B1 => n38, B2 => net645136, A => n100, ZN => n94);
   U9 : NAND2_X1 port map( A1 => en, A2 => D(28), ZN => n99);
   U8 : OAI21_X1 port map( B1 => en, B2 => net645135, A => n99, ZN => n93);
   U15 : NAND2_X1 port map( A1 => en, A2 => D(25), ZN => n64);
   U14 : OAI21_X1 port map( B1 => en, B2 => net645132, A => n64, ZN => n90);
   U23 : NAND2_X1 port map( A1 => en, A2 => D(21), ZN => n60);
   U22 : OAI21_X1 port map( B1 => en, B2 => net645128, A => n60, ZN => n86);
   U25 : NAND2_X1 port map( A1 => en, A2 => D(20), ZN => n59);
   U24 : OAI21_X1 port map( B1 => en, B2 => net645107, A => n59, ZN => n85);
   U17 : NAND2_X1 port map( A1 => en, A2 => D(24), ZN => n63);
   U16 : OAI21_X1 port map( B1 => en, B2 => net645131, A => n63, ZN => n89);
   U27 : NAND2_X1 port map( A1 => en, A2 => D(19), ZN => n58);
   U26 : OAI21_X1 port map( B1 => en, B2 => net645127, A => n58, ZN => n84);
   U39 : NAND2_X1 port map( A1 => n38, A2 => D(13), ZN => n53);
   U38 : OAI21_X1 port map( B1 => en, B2 => net645121, A => n53, ZN => n78);
   U37 : NAND2_X1 port map( A1 => n38, A2 => D(14), ZN => n54);
   U36 : OAI21_X1 port map( B1 => n38, B2 => net645122, A => n54, ZN => n79);
   U41 : NAND2_X1 port map( A1 => en, A2 => D(12), ZN => n52);
   U40 : OAI21_X1 port map( B1 => en, B2 => net645120, A => n52, ZN => n77);
   U35 : NAND2_X1 port map( A1 => en, A2 => D(15), ZN => n55);
   U34 : OAI21_X1 port map( B1 => en, B2 => net645123, A => n55, ZN => n80);
   U51 : NAND2_X1 port map( A1 => en, A2 => D(7), ZN => n47);
   U50 : OAI21_X1 port map( B1 => en, B2 => net645115, A => n47, ZN => n72);
   U43 : NAND2_X1 port map( A1 => n38, A2 => D(11), ZN => n51);
   U42 : OAI21_X1 port map( B1 => en, B2 => net645119, A => n51, ZN => n76);
   U49 : NAND2_X1 port map( A1 => en, A2 => D(8), ZN => n48);
   U48 : OAI21_X1 port map( B1 => n38, B2 => net645116, A => n48, ZN => n73);
   U47 : NAND2_X1 port map( A1 => en, A2 => D(9), ZN => n49);
   U46 : OAI21_X1 port map( B1 => en, B2 => net645117, A => n49, ZN => n74);
   U31 : NAND2_X1 port map( A1 => en, A2 => D(17), ZN => n56);
   U30 : OAI21_X1 port map( B1 => en, B2 => net645125, A => n56, ZN => n82);
   U29 : NAND2_X1 port map( A1 => en, A2 => D(18), ZN => n57);
   U28 : OAI21_X1 port map( B1 => en, B2 => net645126, A => n57, ZN => n83);
   U45 : NAND2_X1 port map( A1 => n38, A2 => D(10), ZN => n50);
   U44 : OAI21_X1 port map( B1 => en, B2 => net645118, A => n50, ZN => n75);
   U59 : NAND2_X1 port map( A1 => en, A2 => D(3), ZN => n43);
   U58 : OAI21_X1 port map( B1 => n38, B2 => net645111, A => n43, ZN => n68);
   U53 : NAND2_X1 port map( A1 => en, A2 => D(6), ZN => n46);
   U52 : OAI21_X1 port map( B1 => n38, B2 => net645114, A => n46, ZN => n71);
   U55 : NAND2_X1 port map( A1 => en, A2 => D(5), ZN => n45);
   U54 : OAI21_X1 port map( B1 => n38, B2 => net645113, A => n45, ZN => n70);
   U57 : NAND2_X1 port map( A1 => en, A2 => D(4), ZN => n44);
   U56 : OAI21_X1 port map( B1 => n38, B2 => net645112, A => n44, ZN => n69);
   U61 : NAND2_X1 port map( A1 => en, A2 => D(2), ZN => n42);
   U60 : OAI21_X1 port map( B1 => n38, B2 => net645110, A => n42, ZN => n67);
   U63 : NAND2_X1 port map( A1 => en, A2 => D(1), ZN => n41);
   U62 : OAI21_X1 port map( B1 => n38, B2 => net645109, A => n41, ZN => n66);
   U65 : NAND2_X1 port map( A1 => en, A2 => D(0), ZN => n40);
   U64 : OAI21_X1 port map( B1 => n38, B2 => net645108, A => n40, ZN => n65);
   U4 : NAND2_X1 port map( A1 => en, A2 => D(16), ZN => n35);
   U5 : OAI21_X1 port map( B1 => en, B2 => net645124, A => n35, ZN => n81);
   U32 : NAND2_X1 port map( A1 => en, A2 => D(30), ZN => n36);
   U33 : OAI21_X1 port map( B1 => en, B2 => net645137, A => n36, ZN => n95);
   U66 : INV_X2 port map( A => rst, ZN => n39);
   U67 : BUF_X1 port map( A => en, Z => n38);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity p4add_N32_logN5_1 is

   port( A, B : in std_logic_vector (31 downto 0);  Cin, sign : in std_logic;  
         S : out std_logic_vector (31 downto 0);  Cout : out std_logic);

end p4add_N32_logN5_1;

architecture SYN_STRUCTURAL of p4add_N32_logN5_1 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component sum_gen_N32_1
      port( A, B : in std_logic_vector (31 downto 0);  Cin : in 
            std_logic_vector (8 downto 0);  S : out std_logic_vector (31 downto
            0));
   end component;
   
   component carry_tree_N32_logN5_1
      port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  
            Cout : out std_logic_vector (7 downto 0));
   end component;
   
   component xor_gen_N32_1
      port( A : in std_logic_vector (31 downto 0);  B : in std_logic;  S : out 
            std_logic_vector (31 downto 0));
   end component;
   
   signal new_B_31_port, new_B_30_port, new_B_29_port, new_B_28_port, 
      new_B_24_port, new_B_23_port, new_B_22_port, new_B_21_port, new_B_16_port
      , new_B_12_port, carry_pro_7_port, carry_pro_6_port, carry_pro_5_port, 
      carry_pro_4_port, carry_pro_3_port, carry_pro_2_port, carry_pro_1_port, 
      n1, n2, n3, n5, n6, n10, n11, n12, n13, n14, n15, n16, n17, n19, n22, n23
      , n24, n26, n27, n28, n29, n31, n32, n33, n34, n35, n36, n37, n38, n39, 
      n40, n41, n42, n43, n44, n45, n46, n47 : std_logic;

begin
   
   n26 <= '0';
   xor32 : xor_gen_N32_1 port map( A(31) => B(31), A(30) => B(30), A(29) => 
                           B(29), A(28) => B(28), A(27) => B(27), A(26) => 
                           B(26), A(25) => B(25), A(24) => B(24), A(23) => 
                           B(23), A(22) => B(22), A(21) => B(21), A(20) => 
                           B(20), A(19) => B(19), A(18) => B(18), A(17) => 
                           B(17), A(16) => B(16), A(15) => B(15), A(14) => 
                           B(14), A(13) => B(13), A(12) => B(12), A(11) => 
                           B(11), A(10) => B(10), A(9) => B(9), A(8) => B(8), 
                           A(7) => B(7), A(6) => B(6), A(5) => B(5), A(4) => 
                           B(4), A(3) => B(3), A(2) => B(2), A(1) => B(1), A(0)
                           => B(0), B => sign, S(31) => new_B_31_port, S(30) =>
                           new_B_30_port, S(29) => new_B_29_port, S(28) => 
                           new_B_28_port, S(27) => n29, S(26) => n1, S(25) => 
                           n14, S(24) => new_B_24_port, S(23) => new_B_23_port,
                           S(22) => new_B_22_port, S(21) => new_B_21_port, 
                           S(20) => n33, S(19) => n13, S(18) => n28, S(17) => 
                           n22, S(16) => new_B_16_port, S(15) => n3, S(14) => 
                           n16, S(13) => n6, S(12) => new_B_12_port, S(11) => 
                           n2, S(10) => n17, S(9) => n15, S(8) => n5, S(7) => 
                           n32, S(6) => n31, S(5) => n19, S(4) => n23, S(3) => 
                           n12, S(2) => n11, S(1) => n24, S(0) => n10);
   ct : carry_tree_N32_logN5_1 port map( A(31) => A(31), A(30) => A(30), A(29) 
                           => A(29), A(28) => A(28), A(27) => A(27), A(26) => 
                           A(26), A(25) => A(25), A(24) => A(24), A(23) => 
                           A(23), A(22) => A(22), A(21) => A(21), A(20) => 
                           A(20), A(19) => A(19), A(18) => A(18), A(17) => 
                           A(17), A(16) => A(16), A(15) => A(15), A(14) => 
                           A(14), A(13) => A(13), A(12) => A(12), A(11) => 
                           A(11), A(10) => A(10), A(9) => A(9), A(8) => A(8), 
                           A(7) => A(7), A(6) => A(6), A(5) => A(5), A(4) => 
                           A(4), A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(31) => new_B_31_port, B(30) => 
                           new_B_30_port, B(29) => new_B_29_port, B(28) => 
                           new_B_28_port, B(27) => n29, B(26) => n1, B(25) => 
                           n14, B(24) => new_B_24_port, B(23) => new_B_23_port,
                           B(22) => new_B_22_port, B(21) => new_B_21_port, 
                           B(20) => n33, B(19) => n13, B(18) => n28, B(17) => 
                           n22, B(16) => new_B_16_port, B(15) => n3, B(14) => 
                           n16, B(13) => n6, B(12) => new_B_12_port, B(11) => 
                           n2, B(10) => n17, B(9) => n15, B(8) => n5, B(7) => 
                           n32, B(6) => n31, B(5) => n19, B(4) => n23, B(3) => 
                           n12, B(2) => n11, B(1) => n24, B(0) => n10, Cin => 
                           sign, Cout(7) => Cout, Cout(6) => carry_pro_7_port, 
                           Cout(5) => carry_pro_6_port, Cout(4) => 
                           carry_pro_5_port, Cout(3) => carry_pro_4_port, 
                           Cout(2) => carry_pro_3_port, Cout(1) => 
                           carry_pro_2_port, Cout(0) => carry_pro_1_port);
   add : sum_gen_N32_1 port map( A(31) => A(31), A(30) => A(30), A(29) => A(29)
                           , A(28) => A(28), A(27) => A(27), A(26) => A(26), 
                           A(25) => A(25), A(24) => A(24), A(23) => A(23), 
                           A(22) => A(22), A(21) => A(21), A(20) => A(20), 
                           A(19) => A(19), A(18) => A(18), A(17) => A(17), 
                           A(16) => A(16), A(15) => A(15), A(14) => A(14), 
                           A(13) => A(13), A(12) => A(12), A(11) => A(11), 
                           A(10) => A(10), A(9) => A(9), A(8) => A(8), A(7) => 
                           A(7), A(6) => A(6), A(5) => A(5), A(4) => A(4), A(3)
                           => A(3), A(2) => A(2), A(1) => A(1), A(0) => A(0), 
                           B(31) => new_B_31_port, B(30) => new_B_30_port, 
                           B(29) => new_B_29_port, B(28) => new_B_28_port, 
                           B(27) => n29, B(26) => n1, B(25) => n40, B(24) => 
                           new_B_24_port, B(23) => n47, B(22) => n41, B(21) => 
                           n34, B(20) => n33, B(19) => n38, B(18) => n28, B(17)
                           => n45, B(16) => new_B_16_port, B(15) => n3, B(14) 
                           => n42, B(13) => n36, B(12) => new_B_12_port, B(11) 
                           => n37, B(10) => n39, B(9) => n27, B(8) => n5, B(7) 
                           => n32, B(6) => n43, B(5) => n19, B(4) => n23, B(3) 
                           => n35, B(2) => n46, B(1) => n24, B(0) => n44, 
                           Cin(8) => n26, Cin(7) => carry_pro_7_port, Cin(6) =>
                           carry_pro_6_port, Cin(5) => carry_pro_5_port, Cin(4)
                           => carry_pro_4_port, Cin(3) => carry_pro_3_port, 
                           Cin(2) => carry_pro_2_port, Cin(1) => 
                           carry_pro_1_port, Cin(0) => sign, S(31) => S(31), 
                           S(30) => S(30), S(29) => S(29), S(28) => S(28), 
                           S(27) => S(27), S(26) => S(26), S(25) => S(25), 
                           S(24) => S(24), S(23) => S(23), S(22) => S(22), 
                           S(21) => S(21), S(20) => S(20), S(19) => S(19), 
                           S(18) => S(18), S(17) => S(17), S(16) => S(16), 
                           S(15) => S(15), S(14) => S(14), S(13) => S(13), 
                           S(12) => S(12), S(11) => S(11), S(10) => S(10), S(9)
                           => S(9), S(8) => S(8), S(7) => S(7), S(6) => S(6), 
                           S(5) => S(5), S(4) => S(4), S(3) => S(3), S(2) => 
                           S(2), S(1) => S(1), S(0) => S(0));
   U1 : BUF_X1 port map( A => n15, Z => n27);
   U2 : BUF_X1 port map( A => n6, Z => n36);
   U3 : BUF_X1 port map( A => n12, Z => n35);
   U4 : BUF_X1 port map( A => new_B_22_port, Z => n41);
   U5 : BUF_X1 port map( A => n13, Z => n38);
   U6 : BUF_X1 port map( A => n10, Z => n44);
   U7 : BUF_X1 port map( A => n31, Z => n43);
   U8 : BUF_X1 port map( A => new_B_21_port, Z => n34);
   U9 : BUF_X1 port map( A => n14, Z => n40);
   U10 : CLKBUF_X1 port map( A => n2, Z => n37);
   U11 : CLKBUF_X1 port map( A => n17, Z => n39);
   U12 : CLKBUF_X1 port map( A => new_B_23_port, Z => n47);
   U13 : CLKBUF_X1 port map( A => n16, Z => n42);
   U14 : CLKBUF_X1 port map( A => n22, Z => n45);
   U15 : CLKBUF_X1 port map( A => n11, Z => n46);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity predictor_2_14 is

   port( clock, reset, enable, taken_i : in std_logic;  prediction_o : out 
         std_logic);

end predictor_2_14;

architecture SYN_bhe of predictor_2_14 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal prediction_o_port, next_STATE_1_port, next_STATE_0_port, N11, N12, n5
      , n6, n8, n10, n12_port, n13, n14, net684345 : std_logic;

begin
   prediction_o <= prediction_o_port;
   
   next_STATE_reg_0_inst : DLH_X1 port map( G => enable, D => N11, Q => 
                           next_STATE_0_port);
   STATE_reg_0_inst : DFFR_X1 port map( D => n6, CK => clock, RN => n12_port, Q
                           => n5, QN => n10);
   next_STATE_reg_1_inst : DLH_X1 port map( G => enable, D => N12, Q => 
                           next_STATE_1_port);
   STATE_reg_1_inst : DFFR_X1 port map( D => n8, CK => clock, RN => n12_port, Q
                           => prediction_o_port, QN => net684345);
   U8 : MUX2_X1 port map( A => prediction_o_port, B => next_STATE_1_port, S => 
                           enable, Z => n8);
   U9 : MUX2_X1 port map( A => n5, B => next_STATE_0_port, S => enable, Z => n6
                           );
   U7 : NOR2_X1 port map( A1 => prediction_o_port, A2 => taken_i, ZN => n14);
   U6 : NAND2_X1 port map( A1 => prediction_o_port, A2 => taken_i, ZN => n13);
   U3 : OAI21_X1 port map( B1 => n14, B2 => n10, A => n13, ZN => N12);
   U5 : OAI21_X1 port map( B1 => n5, B2 => n14, A => n13, ZN => N11);
   U2 : INV_X1 port map( A => reset, ZN => n12_port);

end SYN_bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity predictor_2_13 is

   port( clock, reset, enable, taken_i : in std_logic;  prediction_o : out 
         std_logic);

end predictor_2_13;

architecture SYN_bhe of predictor_2_13 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal prediction_o_port, next_STATE_1_port, next_STATE_0_port, N11, N12, n5
      , n6, n8, n10, n12_port, n13, n14, net684344 : std_logic;

begin
   prediction_o <= prediction_o_port;
   
   next_STATE_reg_0_inst : DLH_X1 port map( G => enable, D => N11, Q => 
                           next_STATE_0_port);
   STATE_reg_0_inst : DFFR_X1 port map( D => n6, CK => clock, RN => n12_port, Q
                           => n5, QN => n10);
   next_STATE_reg_1_inst : DLH_X1 port map( G => enable, D => N12, Q => 
                           next_STATE_1_port);
   STATE_reg_1_inst : DFFR_X1 port map( D => n8, CK => clock, RN => n12_port, Q
                           => prediction_o_port, QN => net684344);
   U8 : MUX2_X1 port map( A => prediction_o_port, B => next_STATE_1_port, S => 
                           enable, Z => n8);
   U9 : MUX2_X1 port map( A => n5, B => next_STATE_0_port, S => enable, Z => n6
                           );
   U7 : NOR2_X1 port map( A1 => prediction_o_port, A2 => taken_i, ZN => n14);
   U6 : NAND2_X1 port map( A1 => prediction_o_port, A2 => taken_i, ZN => n13);
   U5 : OAI21_X1 port map( B1 => n5, B2 => n14, A => n13, ZN => N11);
   U3 : OAI21_X1 port map( B1 => n14, B2 => n10, A => n13, ZN => N12);
   U2 : INV_X1 port map( A => reset, ZN => n12_port);

end SYN_bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity predictor_2_12 is

   port( clock, reset, enable, taken_i : in std_logic;  prediction_o : out 
         std_logic);

end predictor_2_12;

architecture SYN_bhe of predictor_2_12 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal prediction_o_port, next_STATE_1_port, next_STATE_0_port, N11, N12, n5
      , n6, n8, n10, n12_port, n13, n14, net684343 : std_logic;

begin
   prediction_o <= prediction_o_port;
   
   next_STATE_reg_0_inst : DLH_X1 port map( G => enable, D => N11, Q => 
                           next_STATE_0_port);
   STATE_reg_0_inst : DFFR_X1 port map( D => n6, CK => clock, RN => n12_port, Q
                           => n5, QN => n10);
   next_STATE_reg_1_inst : DLH_X1 port map( G => enable, D => N12, Q => 
                           next_STATE_1_port);
   STATE_reg_1_inst : DFFR_X1 port map( D => n8, CK => clock, RN => n12_port, Q
                           => prediction_o_port, QN => net684343);
   U8 : MUX2_X1 port map( A => prediction_o_port, B => next_STATE_1_port, S => 
                           enable, Z => n8);
   U9 : MUX2_X1 port map( A => n5, B => next_STATE_0_port, S => enable, Z => n6
                           );
   U7 : NOR2_X1 port map( A1 => prediction_o_port, A2 => taken_i, ZN => n14);
   U6 : NAND2_X1 port map( A1 => prediction_o_port, A2 => taken_i, ZN => n13);
   U5 : OAI21_X1 port map( B1 => n5, B2 => n14, A => n13, ZN => N11);
   U3 : OAI21_X1 port map( B1 => n14, B2 => n10, A => n13, ZN => N12);
   U2 : INV_X1 port map( A => reset, ZN => n12_port);

end SYN_bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity predictor_2_11 is

   port( clock, reset, enable, taken_i : in std_logic;  prediction_o : out 
         std_logic);

end predictor_2_11;

architecture SYN_bhe of predictor_2_11 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal prediction_o_port, next_STATE_1_port, next_STATE_0_port, N11, N12, n5
      , n6, n8, n10, n12_port, n13, n14, net684342 : std_logic;

begin
   prediction_o <= prediction_o_port;
   
   next_STATE_reg_0_inst : DLH_X1 port map( G => enable, D => N11, Q => 
                           next_STATE_0_port);
   STATE_reg_0_inst : DFFR_X1 port map( D => n6, CK => clock, RN => n12_port, Q
                           => n5, QN => n10);
   next_STATE_reg_1_inst : DLH_X1 port map( G => enable, D => N12, Q => 
                           next_STATE_1_port);
   STATE_reg_1_inst : DFFR_X1 port map( D => n8, CK => clock, RN => n12_port, Q
                           => prediction_o_port, QN => net684342);
   U8 : MUX2_X1 port map( A => prediction_o_port, B => next_STATE_1_port, S => 
                           enable, Z => n8);
   U9 : MUX2_X1 port map( A => n5, B => next_STATE_0_port, S => enable, Z => n6
                           );
   U7 : NOR2_X1 port map( A1 => prediction_o_port, A2 => taken_i, ZN => n14);
   U6 : NAND2_X1 port map( A1 => prediction_o_port, A2 => taken_i, ZN => n13);
   U5 : OAI21_X1 port map( B1 => n5, B2 => n14, A => n13, ZN => N11);
   U3 : OAI21_X1 port map( B1 => n14, B2 => n10, A => n13, ZN => N12);
   U2 : INV_X1 port map( A => reset, ZN => n12_port);

end SYN_bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity predictor_2_10 is

   port( clock, reset, enable, taken_i : in std_logic;  prediction_o : out 
         std_logic);

end predictor_2_10;

architecture SYN_bhe of predictor_2_10 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal prediction_o_port, next_STATE_1_port, next_STATE_0_port, N11, N12, n5
      , n6, n8, n10, n12_port, n13, n14, net684341 : std_logic;

begin
   prediction_o <= prediction_o_port;
   
   next_STATE_reg_0_inst : DLH_X1 port map( G => enable, D => N11, Q => 
                           next_STATE_0_port);
   STATE_reg_0_inst : DFFR_X1 port map( D => n6, CK => clock, RN => n12_port, Q
                           => n5, QN => n10);
   next_STATE_reg_1_inst : DLH_X1 port map( G => enable, D => N12, Q => 
                           next_STATE_1_port);
   STATE_reg_1_inst : DFFR_X1 port map( D => n8, CK => clock, RN => n12_port, Q
                           => prediction_o_port, QN => net684341);
   U8 : MUX2_X1 port map( A => prediction_o_port, B => next_STATE_1_port, S => 
                           enable, Z => n8);
   U9 : MUX2_X1 port map( A => n5, B => next_STATE_0_port, S => enable, Z => n6
                           );
   U7 : NOR2_X1 port map( A1 => prediction_o_port, A2 => taken_i, ZN => n14);
   U6 : NAND2_X1 port map( A1 => prediction_o_port, A2 => taken_i, ZN => n13);
   U3 : OAI21_X1 port map( B1 => n14, B2 => n10, A => n13, ZN => N12);
   U5 : OAI21_X1 port map( B1 => n5, B2 => n14, A => n13, ZN => N11);
   U2 : INV_X1 port map( A => reset, ZN => n12_port);

end SYN_bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity predictor_2_9 is

   port( clock, reset, enable, taken_i : in std_logic;  prediction_o : out 
         std_logic);

end predictor_2_9;

architecture SYN_bhe of predictor_2_9 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal prediction_o_port, next_STATE_1_port, next_STATE_0_port, N11, N12, n5
      , n6, n8, n10, n12_port, n13, n14, net684340 : std_logic;

begin
   prediction_o <= prediction_o_port;
   
   next_STATE_reg_0_inst : DLH_X1 port map( G => enable, D => N11, Q => 
                           next_STATE_0_port);
   STATE_reg_0_inst : DFFR_X1 port map( D => n6, CK => clock, RN => n12_port, Q
                           => n5, QN => n10);
   next_STATE_reg_1_inst : DLH_X1 port map( G => enable, D => N12, Q => 
                           next_STATE_1_port);
   STATE_reg_1_inst : DFFR_X1 port map( D => n8, CK => clock, RN => n12_port, Q
                           => prediction_o_port, QN => net684340);
   U8 : MUX2_X1 port map( A => prediction_o_port, B => next_STATE_1_port, S => 
                           enable, Z => n8);
   U9 : MUX2_X1 port map( A => n5, B => next_STATE_0_port, S => enable, Z => n6
                           );
   U7 : NOR2_X1 port map( A1 => prediction_o_port, A2 => taken_i, ZN => n14);
   U6 : NAND2_X1 port map( A1 => prediction_o_port, A2 => taken_i, ZN => n13);
   U3 : OAI21_X1 port map( B1 => n14, B2 => n10, A => n13, ZN => N12);
   U5 : OAI21_X1 port map( B1 => n5, B2 => n14, A => n13, ZN => N11);
   U2 : INV_X1 port map( A => reset, ZN => n12_port);

end SYN_bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity predictor_2_8 is

   port( clock, reset, enable, taken_i : in std_logic;  prediction_o : out 
         std_logic);

end predictor_2_8;

architecture SYN_bhe of predictor_2_8 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal prediction_o_port, next_STATE_1_port, next_STATE_0_port, N11, N12, n5
      , n6, n8, n10, n12_port, n13, n14, net684339 : std_logic;

begin
   prediction_o <= prediction_o_port;
   
   next_STATE_reg_0_inst : DLH_X1 port map( G => enable, D => N11, Q => 
                           next_STATE_0_port);
   STATE_reg_0_inst : DFFR_X1 port map( D => n6, CK => clock, RN => n12_port, Q
                           => n5, QN => n10);
   next_STATE_reg_1_inst : DLH_X1 port map( G => enable, D => N12, Q => 
                           next_STATE_1_port);
   STATE_reg_1_inst : DFFR_X1 port map( D => n8, CK => clock, RN => n12_port, Q
                           => prediction_o_port, QN => net684339);
   U8 : MUX2_X1 port map( A => prediction_o_port, B => next_STATE_1_port, S => 
                           enable, Z => n8);
   U9 : MUX2_X1 port map( A => n5, B => next_STATE_0_port, S => enable, Z => n6
                           );
   U7 : NOR2_X1 port map( A1 => prediction_o_port, A2 => taken_i, ZN => n14);
   U6 : NAND2_X1 port map( A1 => prediction_o_port, A2 => taken_i, ZN => n13);
   U3 : OAI21_X1 port map( B1 => n14, B2 => n10, A => n13, ZN => N12);
   U5 : OAI21_X1 port map( B1 => n5, B2 => n14, A => n13, ZN => N11);
   U2 : INV_X1 port map( A => reset, ZN => n12_port);

end SYN_bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity predictor_2_7 is

   port( clock, reset, enable, taken_i : in std_logic;  prediction_o : out 
         std_logic);

end predictor_2_7;

architecture SYN_bhe of predictor_2_7 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal prediction_o_port, next_STATE_1_port, next_STATE_0_port, N11, N12, n5
      , n6, n8, n10, n12_port, n13, n14, net684338 : std_logic;

begin
   prediction_o <= prediction_o_port;
   
   next_STATE_reg_0_inst : DLH_X1 port map( G => enable, D => N11, Q => 
                           next_STATE_0_port);
   STATE_reg_0_inst : DFFR_X1 port map( D => n6, CK => clock, RN => n12_port, Q
                           => n5, QN => n10);
   next_STATE_reg_1_inst : DLH_X1 port map( G => enable, D => N12, Q => 
                           next_STATE_1_port);
   STATE_reg_1_inst : DFFR_X1 port map( D => n8, CK => clock, RN => n12_port, Q
                           => prediction_o_port, QN => net684338);
   U8 : MUX2_X1 port map( A => prediction_o_port, B => next_STATE_1_port, S => 
                           enable, Z => n8);
   U9 : MUX2_X1 port map( A => n5, B => next_STATE_0_port, S => enable, Z => n6
                           );
   U7 : NOR2_X1 port map( A1 => prediction_o_port, A2 => taken_i, ZN => n14);
   U6 : NAND2_X1 port map( A1 => prediction_o_port, A2 => taken_i, ZN => n13);
   U3 : OAI21_X1 port map( B1 => n14, B2 => n10, A => n13, ZN => N12);
   U5 : OAI21_X1 port map( B1 => n5, B2 => n14, A => n13, ZN => N11);
   U2 : INV_X1 port map( A => reset, ZN => n12_port);

end SYN_bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity predictor_2_6 is

   port( clock, reset, enable, taken_i : in std_logic;  prediction_o : out 
         std_logic);

end predictor_2_6;

architecture SYN_bhe of predictor_2_6 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal prediction_o_port, next_STATE_1_port, next_STATE_0_port, N11, N12, n5
      , n6, n8, n10, n12_port, n13, n14, net684337 : std_logic;

begin
   prediction_o <= prediction_o_port;
   
   next_STATE_reg_0_inst : DLH_X1 port map( G => enable, D => N11, Q => 
                           next_STATE_0_port);
   STATE_reg_0_inst : DFFR_X1 port map( D => n6, CK => clock, RN => n12_port, Q
                           => n5, QN => n10);
   next_STATE_reg_1_inst : DLH_X1 port map( G => enable, D => N12, Q => 
                           next_STATE_1_port);
   STATE_reg_1_inst : DFFR_X1 port map( D => n8, CK => clock, RN => n12_port, Q
                           => prediction_o_port, QN => net684337);
   U8 : MUX2_X1 port map( A => prediction_o_port, B => next_STATE_1_port, S => 
                           enable, Z => n8);
   U9 : MUX2_X1 port map( A => n5, B => next_STATE_0_port, S => enable, Z => n6
                           );
   U7 : NOR2_X1 port map( A1 => prediction_o_port, A2 => taken_i, ZN => n14);
   U6 : NAND2_X1 port map( A1 => prediction_o_port, A2 => taken_i, ZN => n13);
   U3 : OAI21_X1 port map( B1 => n14, B2 => n10, A => n13, ZN => N12);
   U5 : OAI21_X1 port map( B1 => n5, B2 => n14, A => n13, ZN => N11);
   U2 : INV_X1 port map( A => reset, ZN => n12_port);

end SYN_bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity predictor_2_5 is

   port( clock, reset, enable, taken_i : in std_logic;  prediction_o : out 
         std_logic);

end predictor_2_5;

architecture SYN_bhe of predictor_2_5 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal prediction_o_port, next_STATE_1_port, next_STATE_0_port, N11, N12, n5
      , n6, n8, n10, n12_port, n13, n14, net684336 : std_logic;

begin
   prediction_o <= prediction_o_port;
   
   next_STATE_reg_0_inst : DLH_X1 port map( G => enable, D => N11, Q => 
                           next_STATE_0_port);
   STATE_reg_0_inst : DFFR_X1 port map( D => n6, CK => clock, RN => n12_port, Q
                           => n5, QN => n10);
   next_STATE_reg_1_inst : DLH_X1 port map( G => enable, D => N12, Q => 
                           next_STATE_1_port);
   STATE_reg_1_inst : DFFR_X1 port map( D => n8, CK => clock, RN => n12_port, Q
                           => prediction_o_port, QN => net684336);
   U8 : MUX2_X1 port map( A => prediction_o_port, B => next_STATE_1_port, S => 
                           enable, Z => n8);
   U9 : MUX2_X1 port map( A => n5, B => next_STATE_0_port, S => enable, Z => n6
                           );
   U7 : NOR2_X1 port map( A1 => prediction_o_port, A2 => taken_i, ZN => n14);
   U6 : NAND2_X1 port map( A1 => prediction_o_port, A2 => taken_i, ZN => n13);
   U5 : OAI21_X1 port map( B1 => n5, B2 => n14, A => n13, ZN => N11);
   U3 : OAI21_X1 port map( B1 => n14, B2 => n10, A => n13, ZN => N12);
   U2 : INV_X1 port map( A => reset, ZN => n12_port);

end SYN_bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity predictor_2_4 is

   port( clock, reset, enable, taken_i : in std_logic;  prediction_o : out 
         std_logic);

end predictor_2_4;

architecture SYN_bhe of predictor_2_4 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal prediction_o_port, next_STATE_1_port, next_STATE_0_port, N11, N12, n5
      , n6, n8, n10, n12_port, n13, n14, net684335 : std_logic;

begin
   prediction_o <= prediction_o_port;
   
   next_STATE_reg_0_inst : DLH_X1 port map( G => enable, D => N11, Q => 
                           next_STATE_0_port);
   STATE_reg_0_inst : DFFR_X1 port map( D => n6, CK => clock, RN => n12_port, Q
                           => n5, QN => n10);
   next_STATE_reg_1_inst : DLH_X1 port map( G => enable, D => N12, Q => 
                           next_STATE_1_port);
   STATE_reg_1_inst : DFFR_X1 port map( D => n8, CK => clock, RN => n12_port, Q
                           => prediction_o_port, QN => net684335);
   U8 : MUX2_X1 port map( A => prediction_o_port, B => next_STATE_1_port, S => 
                           enable, Z => n8);
   U9 : MUX2_X1 port map( A => n5, B => next_STATE_0_port, S => enable, Z => n6
                           );
   U7 : NOR2_X1 port map( A1 => prediction_o_port, A2 => taken_i, ZN => n14);
   U6 : NAND2_X1 port map( A1 => prediction_o_port, A2 => taken_i, ZN => n13);
   U3 : OAI21_X1 port map( B1 => n14, B2 => n10, A => n13, ZN => N12);
   U5 : OAI21_X1 port map( B1 => n5, B2 => n14, A => n13, ZN => N11);
   U2 : INV_X1 port map( A => reset, ZN => n12_port);

end SYN_bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity predictor_2_3 is

   port( clock, reset, enable, taken_i : in std_logic;  prediction_o : out 
         std_logic);

end predictor_2_3;

architecture SYN_bhe of predictor_2_3 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal prediction_o_port, next_STATE_1_port, next_STATE_0_port, N11, N12, n5
      , n6, n8, n10, n12_port, n13, n14, net684334 : std_logic;

begin
   prediction_o <= prediction_o_port;
   
   next_STATE_reg_0_inst : DLH_X1 port map( G => enable, D => N11, Q => 
                           next_STATE_0_port);
   STATE_reg_0_inst : DFFR_X1 port map( D => n6, CK => clock, RN => n12_port, Q
                           => n5, QN => n10);
   next_STATE_reg_1_inst : DLH_X1 port map( G => enable, D => N12, Q => 
                           next_STATE_1_port);
   STATE_reg_1_inst : DFFR_X1 port map( D => n8, CK => clock, RN => n12_port, Q
                           => prediction_o_port, QN => net684334);
   U8 : MUX2_X1 port map( A => prediction_o_port, B => next_STATE_1_port, S => 
                           enable, Z => n8);
   U9 : MUX2_X1 port map( A => n5, B => next_STATE_0_port, S => enable, Z => n6
                           );
   U7 : NOR2_X1 port map( A1 => prediction_o_port, A2 => taken_i, ZN => n14);
   U6 : NAND2_X1 port map( A1 => prediction_o_port, A2 => taken_i, ZN => n13);
   U5 : OAI21_X1 port map( B1 => n5, B2 => n14, A => n13, ZN => N11);
   U3 : OAI21_X1 port map( B1 => n14, B2 => n10, A => n13, ZN => N12);
   U2 : INV_X1 port map( A => reset, ZN => n12_port);

end SYN_bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity predictor_2_2 is

   port( clock, reset, enable, taken_i : in std_logic;  prediction_o : out 
         std_logic);

end predictor_2_2;

architecture SYN_bhe of predictor_2_2 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal prediction_o_port, next_STATE_1_port, next_STATE_0_port, N11, N12, n5
      , n6, n8, n10, n12_port, n13, n14, net684333 : std_logic;

begin
   prediction_o <= prediction_o_port;
   
   next_STATE_reg_0_inst : DLH_X1 port map( G => enable, D => N11, Q => 
                           next_STATE_0_port);
   STATE_reg_0_inst : DFFR_X1 port map( D => n6, CK => clock, RN => n12_port, Q
                           => n5, QN => n10);
   next_STATE_reg_1_inst : DLH_X1 port map( G => enable, D => N12, Q => 
                           next_STATE_1_port);
   STATE_reg_1_inst : DFFR_X1 port map( D => n8, CK => clock, RN => n12_port, Q
                           => prediction_o_port, QN => net684333);
   U8 : MUX2_X1 port map( A => prediction_o_port, B => next_STATE_1_port, S => 
                           enable, Z => n8);
   U9 : MUX2_X1 port map( A => n5, B => next_STATE_0_port, S => enable, Z => n6
                           );
   U7 : NOR2_X1 port map( A1 => prediction_o_port, A2 => taken_i, ZN => n14);
   U6 : NAND2_X1 port map( A1 => prediction_o_port, A2 => taken_i, ZN => n13);
   U5 : OAI21_X1 port map( B1 => n5, B2 => n14, A => n13, ZN => N11);
   U3 : OAI21_X1 port map( B1 => n14, B2 => n10, A => n13, ZN => N12);
   U2 : INV_X1 port map( A => reset, ZN => n12_port);

end SYN_bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity predictor_2_1 is

   port( clock, reset, enable, taken_i : in std_logic;  prediction_o : out 
         std_logic);

end predictor_2_1;

architecture SYN_bhe of predictor_2_1 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal prediction_o_port, next_STATE_1_port, next_STATE_0_port, N11, N12, n5
      , n6, n8, n10, n12_port, n13, n14, net684332 : std_logic;

begin
   prediction_o <= prediction_o_port;
   
   next_STATE_reg_0_inst : DLH_X1 port map( G => enable, D => N11, Q => 
                           next_STATE_0_port);
   STATE_reg_0_inst : DFFR_X1 port map( D => n6, CK => clock, RN => n12_port, Q
                           => n5, QN => n10);
   next_STATE_reg_1_inst : DLH_X1 port map( G => enable, D => N12, Q => 
                           next_STATE_1_port);
   STATE_reg_1_inst : DFFR_X1 port map( D => n8, CK => clock, RN => n12_port, Q
                           => prediction_o_port, QN => net684332);
   U8 : MUX2_X1 port map( A => prediction_o_port, B => next_STATE_1_port, S => 
                           enable, Z => n8);
   U9 : MUX2_X1 port map( A => n5, B => next_STATE_0_port, S => enable, Z => n6
                           );
   U7 : NOR2_X1 port map( A1 => prediction_o_port, A2 => taken_i, ZN => n14);
   U6 : NAND2_X1 port map( A1 => prediction_o_port, A2 => taken_i, ZN => n13);
   U3 : OAI21_X1 port map( B1 => n14, B2 => n10, A => n13, ZN => N12);
   U5 : OAI21_X1 port map( B1 => n5, B2 => n14, A => n13, ZN => N11);
   U2 : INV_X1 port map( A => reset, ZN => n12_port);

end SYN_bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity mux41_1 is

   port( IN0, IN1, IN2, IN3 : in std_logic_vector (31 downto 0);  CTRL : in 
         std_logic_vector (1 downto 0);  OUT1 : out std_logic_vector (31 downto
         0));

end mux41_1;

architecture SYN_bhe of mux41_1 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X3
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
      n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, 
      n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, 
      n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, 
      n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, 
      n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, 
      n153, n154, n155, n156, n157, n158 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n91, A2 => n90, ZN => OUT1(11));
   U2 : CLKBUF_X3 port map( A => n156, Z => n127);
   U3 : INV_X1 port map( A => CTRL(0), ZN => n110);
   U4 : AND2_X1 port map( A1 => CTRL(1), A2 => n110, ZN => n78);
   U5 : AND2_X1 port map( A1 => CTRL(1), A2 => CTRL(0), ZN => n158);
   U6 : CLKBUF_X3 port map( A => n157, Z => n130);
   U7 : CLKBUF_X3 port map( A => n157, Z => n129);
   U8 : CLKBUF_X3 port map( A => n157, Z => n128);
   U9 : CLKBUF_X3 port map( A => n156, Z => n125);
   U10 : CLKBUF_X3 port map( A => n156, Z => n126);
   U11 : BUF_X2 port map( A => n78, Z => n79);
   U12 : BUF_X2 port map( A => n158, Z => n133);
   U13 : BUF_X2 port map( A => n158, Z => n132);
   U14 : BUF_X2 port map( A => n78, Z => n80);
   U15 : BUF_X2 port map( A => n78, Z => n81);
   U16 : BUF_X2 port map( A => n158, Z => n131);
   U17 : AOI22_X1 port map( A1 => n131, A2 => IN3(15), B1 => n80, B2 => IN2(15)
                           , ZN => n83);
   U18 : AOI22_X1 port map( A1 => n131, A2 => IN3(18), B1 => n79, B2 => IN2(18)
                           , ZN => n103);
   U19 : AOI22_X1 port map( A1 => n132, A2 => IN3(29), B1 => n80, B2 => IN2(29)
                           , ZN => n105);
   U20 : AOI22_X1 port map( A1 => n131, A2 => IN3(16), B1 => n81, B2 => IN2(16)
                           , ZN => n112);
   U21 : AOI22_X1 port map( A1 => n132, A2 => IN3(22), B1 => n79, B2 => IN2(22)
                           , ZN => n116);
   U22 : AOI22_X1 port map( A1 => n131, A2 => IN3(19), B1 => n79, B2 => IN2(19)
                           , ZN => n118);
   U23 : AOI22_X1 port map( A1 => n131, A2 => IN3(12), B1 => n80, B2 => IN2(12)
                           , ZN => n120);
   U24 : AOI22_X1 port map( A1 => n133, A2 => IN3(4), B1 => n79, B2 => IN2(4), 
                           ZN => n124);
   U25 : AOI22_X1 port map( A1 => n133, A2 => IN3(6), B1 => n81, B2 => IN2(6), 
                           ZN => n152);
   U26 : AOI22_X1 port map( A1 => n131, A2 => IN3(1), B1 => n81, B2 => IN2(1), 
                           ZN => n138);
   U27 : AOI22_X1 port map( A1 => n133, A2 => IN3(31), B1 => n79, B2 => IN2(31)
                           , ZN => n85);
   U28 : AOI22_X1 port map( A1 => n131, A2 => IN3(10), B1 => n81, B2 => IN2(10)
                           , ZN => n93);
   U29 : AOI22_X1 port map( A1 => n132, A2 => IN3(23), B1 => n81, B2 => IN2(23)
                           , ZN => n97);
   U30 : AOI22_X1 port map( A1 => n133, A2 => IN3(3), B1 => n79, B2 => IN2(3), 
                           ZN => n107);
   U31 : AOI22_X1 port map( A1 => n132, A2 => IN3(2), B1 => n79, B2 => IN2(2), 
                           ZN => n109);
   U32 : AOI22_X1 port map( A1 => n133, A2 => IN3(5), B1 => n80, B2 => IN2(5), 
                           ZN => n114);
   U33 : AOI22_X1 port map( A1 => n131, A2 => IN3(17), B1 => n79, B2 => IN2(17)
                           , ZN => n122);
   U34 : AOI22_X1 port map( A1 => n131, A2 => IN3(13), B1 => n81, B2 => IN2(13)
                           , ZN => n136);
   U35 : AOI22_X1 port map( A1 => n132, A2 => IN3(21), B1 => n80, B2 => IN2(21)
                           , ZN => n142);
   U36 : AOI22_X1 port map( A1 => n131, A2 => IN3(0), B1 => n80, B2 => IN2(0), 
                           ZN => n134);
   U37 : AOI22_X1 port map( A1 => n133, A2 => IN3(8), B1 => n81, B2 => IN2(8), 
                           ZN => n154);
   U38 : AOI22_X1 port map( A1 => n131, A2 => IN3(14), B1 => n80, B2 => IN2(14)
                           , ZN => n87);
   U39 : AOI22_X1 port map( A1 => n133, A2 => IN3(9), B1 => n81, B2 => IN2(9), 
                           ZN => n89);
   U40 : AOI22_X1 port map( A1 => n131, A2 => IN3(11), B1 => n79, B2 => IN2(11)
                           , ZN => n91);
   U41 : AOI22_X1 port map( A1 => n133, A2 => IN3(7), B1 => n80, B2 => IN2(7), 
                           ZN => n95);
   U42 : AOI22_X1 port map( A1 => n132, A2 => IN3(26), B1 => n80, B2 => IN2(26)
                           , ZN => n99);
   U43 : AOI22_X1 port map( A1 => n132, A2 => IN3(27), B1 => n79, B2 => IN2(27)
                           , ZN => n101);
   U44 : AOI22_X1 port map( A1 => n132, A2 => IN3(28), B1 => n79, B2 => IN2(28)
                           , ZN => n148);
   U45 : AOI22_X1 port map( A1 => n132, A2 => IN3(30), B1 => n80, B2 => IN2(30)
                           , ZN => n150);
   U46 : AOI22_X1 port map( A1 => n132, A2 => IN3(25), B1 => n81, B2 => IN2(25)
                           , ZN => n146);
   U47 : AOI22_X1 port map( A1 => n132, A2 => IN3(24), B1 => n81, B2 => IN2(24)
                           , ZN => n144);
   U48 : AOI22_X1 port map( A1 => n132, A2 => IN3(20), B1 => n80, B2 => IN2(20)
                           , ZN => n140);
   U49 : NAND2_X1 port map( A1 => n121, A2 => n122, ZN => OUT1(17));
   U50 : NAND2_X1 port map( A1 => n92, A2 => n93, ZN => OUT1(10));
   U51 : NAND2_X1 port map( A1 => n86, A2 => n87, ZN => OUT1(14));
   U52 : NAND2_X1 port map( A1 => n111, A2 => n112, ZN => OUT1(16));
   U53 : NAND2_X1 port map( A1 => n102, A2 => n103, ZN => OUT1(18));
   U54 : NAND2_X1 port map( A1 => n82, A2 => n83, ZN => OUT1(15));
   U55 : NAND2_X1 port map( A1 => n84, A2 => n85, ZN => OUT1(31));
   U56 : AOI22_X1 port map( A1 => n130, A2 => IN1(15), B1 => n125, B2 => 
                           IN0(15), ZN => n82);
   U57 : AOI22_X1 port map( A1 => n130, A2 => IN1(31), B1 => n126, B2 => 
                           IN0(31), ZN => n84);
   U58 : NOR2_X1 port map( A1 => n110, A2 => CTRL(1), ZN => n157);
   U59 : AOI22_X1 port map( A1 => n128, A2 => IN1(14), B1 => n125, B2 => 
                           IN0(14), ZN => n86);
   U60 : AOI22_X1 port map( A1 => n128, A2 => IN1(9), B1 => n125, B2 => IN0(9),
                           ZN => n88);
   U61 : NAND2_X1 port map( A1 => n88, A2 => n89, ZN => OUT1(9));
   U62 : AOI22_X1 port map( A1 => n128, A2 => IN1(11), B1 => n126, B2 => 
                           IN0(11), ZN => n90);
   U63 : AOI22_X1 port map( A1 => n128, A2 => IN1(10), B1 => n125, B2 => 
                           IN0(10), ZN => n92);
   U64 : AOI22_X1 port map( A1 => n129, A2 => IN1(7), B1 => n126, B2 => IN0(7),
                           ZN => n94);
   U65 : NAND2_X1 port map( A1 => n94, A2 => n95, ZN => OUT1(7));
   U66 : AOI22_X1 port map( A1 => n129, A2 => IN1(23), B1 => n127, B2 => 
                           IN0(23), ZN => n96);
   U67 : NAND2_X1 port map( A1 => n96, A2 => n97, ZN => OUT1(23));
   U68 : AOI22_X1 port map( A1 => n128, A2 => IN1(26), B1 => n127, B2 => 
                           IN0(26), ZN => n98);
   U69 : NAND2_X1 port map( A1 => n98, A2 => n99, ZN => OUT1(26));
   U70 : AOI22_X1 port map( A1 => n129, A2 => IN1(27), B1 => n127, B2 => 
                           IN0(27), ZN => n100);
   U71 : NAND2_X1 port map( A1 => n100, A2 => n101, ZN => OUT1(27));
   U72 : AOI22_X1 port map( A1 => n129, A2 => IN1(18), B1 => n126, B2 => 
                           IN0(18), ZN => n102);
   U73 : AOI22_X1 port map( A1 => n128, A2 => IN1(29), B1 => n127, B2 => 
                           IN0(29), ZN => n104);
   U74 : NAND2_X1 port map( A1 => n104, A2 => n105, ZN => OUT1(29));
   U75 : AOI22_X1 port map( A1 => n128, A2 => IN1(3), B1 => n125, B2 => IN0(3),
                           ZN => n106);
   U76 : NAND2_X1 port map( A1 => n106, A2 => n107, ZN => OUT1(3));
   U77 : AOI22_X1 port map( A1 => n130, A2 => IN1(2), B1 => n127, B2 => IN0(2),
                           ZN => n108);
   U78 : NAND2_X1 port map( A1 => n108, A2 => n109, ZN => OUT1(2));
   U79 : AOI22_X1 port map( A1 => n129, A2 => IN1(16), B1 => n125, B2 => 
                           IN0(16), ZN => n111);
   U80 : AOI22_X1 port map( A1 => n128, A2 => IN1(5), B1 => n126, B2 => IN0(5),
                           ZN => n113);
   U81 : NAND2_X1 port map( A1 => n113, A2 => n114, ZN => OUT1(5));
   U82 : AOI22_X1 port map( A1 => n129, A2 => IN1(22), B1 => n126, B2 => 
                           IN0(22), ZN => n115);
   U83 : NAND2_X1 port map( A1 => n115, A2 => n116, ZN => OUT1(22));
   U84 : AOI22_X1 port map( A1 => n129, A2 => IN1(19), B1 => n127, B2 => 
                           IN0(19), ZN => n117);
   U85 : NAND2_X1 port map( A1 => n117, A2 => n118, ZN => OUT1(19));
   U86 : AOI22_X1 port map( A1 => n128, A2 => IN1(12), B1 => n125, B2 => 
                           IN0(12), ZN => n119);
   U87 : NAND2_X1 port map( A1 => n119, A2 => n120, ZN => OUT1(12));
   U88 : AOI22_X1 port map( A1 => n129, A2 => IN1(17), B1 => n126, B2 => 
                           IN0(17), ZN => n121);
   U89 : AOI22_X1 port map( A1 => n128, A2 => IN1(4), B1 => n127, B2 => IN0(4),
                           ZN => n123);
   U90 : NAND2_X1 port map( A1 => n123, A2 => n124, ZN => OUT1(4));
   U91 : NOR2_X1 port map( A1 => CTRL(0), A2 => CTRL(1), ZN => n156);
   U92 : NAND2_X1 port map( A1 => n151, A2 => n150, ZN => OUT1(30));
   U93 : NAND2_X1 port map( A1 => n149, A2 => n148, ZN => OUT1(28));
   U94 : NAND2_X1 port map( A1 => n153, A2 => n152, ZN => OUT1(6));
   U95 : NAND2_X1 port map( A1 => n135, A2 => n134, ZN => OUT1(0));
   U96 : NAND2_X1 port map( A1 => n139, A2 => n138, ZN => OUT1(1));
   U97 : NAND2_X1 port map( A1 => n147, A2 => n146, ZN => OUT1(25));
   U98 : NAND2_X1 port map( A1 => n141, A2 => n140, ZN => OUT1(20));
   U99 : NAND2_X1 port map( A1 => n145, A2 => n144, ZN => OUT1(24));
   U100 : NAND2_X1 port map( A1 => n143, A2 => n142, ZN => OUT1(21));
   U101 : NAND2_X1 port map( A1 => n137, A2 => n136, ZN => OUT1(13));
   U102 : NAND2_X1 port map( A1 => n155, A2 => n154, ZN => OUT1(8));
   U103 : AOI22_X1 port map( A1 => n129, A2 => IN1(6), B1 => n126, B2 => IN0(6)
                           , ZN => n153);
   U104 : AOI22_X1 port map( A1 => n129, A2 => IN1(8), B1 => n125, B2 => IN0(8)
                           , ZN => n155);
   U105 : AOI22_X1 port map( A1 => n130, A2 => IN1(28), B1 => n127, B2 => 
                           IN0(28), ZN => n149);
   U106 : AOI22_X1 port map( A1 => n130, A2 => IN1(30), B1 => n126, B2 => 
                           IN0(30), ZN => n151);
   U107 : AOI22_X1 port map( A1 => n130, A2 => IN1(20), B1 => n125, B2 => 
                           IN0(20), ZN => n141);
   U108 : AOI22_X1 port map( A1 => n130, A2 => IN1(25), B1 => n127, B2 => 
                           IN0(25), ZN => n147);
   U109 : AOI22_X1 port map( A1 => n130, A2 => IN1(24), B1 => n126, B2 => 
                           IN0(24), ZN => n145);
   U110 : AOI22_X1 port map( A1 => n130, A2 => IN1(21), B1 => n127, B2 => 
                           IN0(21), ZN => n143);
   U111 : AOI22_X1 port map( A1 => n130, A2 => IN1(0), B1 => n126, B2 => IN0(0)
                           , ZN => n135);
   U112 : AOI22_X1 port map( A1 => n129, A2 => IN1(1), B1 => n125, B2 => IN0(1)
                           , ZN => n139);
   U113 : AOI22_X1 port map( A1 => n128, A2 => IN1(13), B1 => n125, B2 => 
                           IN0(13), ZN => n137);

end SYN_bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity booth_encoder_5 is

   port( B_in : in std_logic_vector (2 downto 0);  A_out : out std_logic_vector
         (2 downto 0));

end booth_encoder_5;

architecture SYN_bhe of booth_encoder_5 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI33_X1
      port( A1, A2, A3, B1, B2, B3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n18, n19, n20, n21 : std_logic;

begin
   
   U9 : OAI33_X1 port map( A1 => B_in(0), A2 => B_in(1), A3 => n18, B1 => n21, 
                           B2 => n20, B3 => B_in(2), ZN => A_out(0));
   U6 : INV_X1 port map( A => B_in(1), ZN => n20);
   U3 : INV_X1 port map( A => B_in(2), ZN => n18);
   U4 : INV_X1 port map( A => B_in(0), ZN => n21);
   U5 : AOI21_X1 port map( B1 => B_in(0), B2 => B_in(1), A => n18, ZN => 
                           A_out(1));
   U7 : OAI221_X1 port map( B1 => B_in(1), B2 => n21, C1 => n20, C2 => B_in(2),
                           A => n19, ZN => A_out(2));
   U8 : NAND2_X1 port map( A1 => B_in(2), A2 => n21, ZN => n19);

end SYN_bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity booth_encoder_4 is

   port( B_in : in std_logic_vector (2 downto 0);  A_out : out std_logic_vector
         (2 downto 0));

end booth_encoder_4;

architecture SYN_bhe of booth_encoder_4 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI33_X1
      port( A1, A2, A3, B1, B2, B3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n18, n19, n20, n21 : std_logic;

begin
   
   U9 : OAI33_X1 port map( A1 => B_in(0), A2 => B_in(1), A3 => n18, B1 => n21, 
                           B2 => n20, B3 => B_in(2), ZN => A_out(0));
   U4 : NAND2_X1 port map( A1 => B_in(2), A2 => n21, ZN => n19);
   U8 : INV_X1 port map( A => B_in(2), ZN => n18);
   U3 : INV_X1 port map( A => B_in(0), ZN => n21);
   U5 : INV_X1 port map( A => B_in(1), ZN => n20);
   U6 : OAI221_X1 port map( B1 => B_in(1), B2 => n21, C1 => n20, C2 => B_in(2),
                           A => n19, ZN => A_out(2));
   U7 : AOI21_X1 port map( B1 => B_in(0), B2 => B_in(1), A => n18, ZN => 
                           A_out(1));

end SYN_bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity booth_encoder_3 is

   port( B_in : in std_logic_vector (2 downto 0);  A_out : out std_logic_vector
         (2 downto 0));

end booth_encoder_3;

architecture SYN_bhe of booth_encoder_3 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI33_X1
      port( A1, A2, A3, B1, B2, B3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n18, n19, n20, n21 : std_logic;

begin
   
   U9 : OAI33_X1 port map( A1 => B_in(0), A2 => B_in(1), A3 => n18, B1 => n21, 
                           B2 => n20, B3 => B_in(2), ZN => A_out(0));
   U7 : INV_X1 port map( A => B_in(0), ZN => n21);
   U3 : INV_X1 port map( A => B_in(2), ZN => n18);
   U4 : INV_X1 port map( A => B_in(1), ZN => n20);
   U5 : AOI21_X1 port map( B1 => B_in(0), B2 => B_in(1), A => n18, ZN => 
                           A_out(1));
   U6 : OAI221_X1 port map( B1 => B_in(1), B2 => n21, C1 => n20, C2 => B_in(2),
                           A => n19, ZN => A_out(2));
   U8 : NAND2_X1 port map( A1 => B_in(2), A2 => n21, ZN => n19);

end SYN_bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity booth_encoder_2 is

   port( B_in : in std_logic_vector (2 downto 0);  A_out : out std_logic_vector
         (2 downto 0));

end booth_encoder_2;

architecture SYN_bhe of booth_encoder_2 is

   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI33_X1
      port( A1, A2, A3, B1, B2, B3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n18, n19, n20, n21 : std_logic;

begin
   
   U9 : OAI33_X1 port map( A1 => B_in(0), A2 => B_in(1), A3 => n18, B1 => n21, 
                           B2 => n20, B3 => B_in(2), ZN => A_out(0));
   U4 : NAND2_X1 port map( A1 => B_in(2), A2 => n21, ZN => n19);
   U3 : INV_X1 port map( A => B_in(0), ZN => n21);
   U5 : INV_X1 port map( A => B_in(2), ZN => n18);
   U6 : INV_X1 port map( A => B_in(1), ZN => n20);
   U7 : AOI21_X1 port map( B1 => B_in(0), B2 => B_in(1), A => n18, ZN => 
                           A_out(1));
   U8 : OAI221_X1 port map( B1 => B_in(1), B2 => n21, C1 => n20, C2 => B_in(2),
                           A => n19, ZN => A_out(2));

end SYN_bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_100 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_100;

architecture SYN_BEHAVIORAL of FA_100 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n1);
   U1 : XNOR2_X1 port map( A => n1, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_110 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_110;

architecture SYN_BEHAVIORAL of FA_110 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n1);
   U1 : XNOR2_X1 port map( A => Ci, B => n1, ZN => S);
   U5 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n2);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n3);
   U3 : NAND2_X1 port map( A1 => n2, A2 => n3, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_119 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_119;

architecture SYN_BEHAVIORAL of FA_119 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_124 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_124;

architecture SYN_BEHAVIORAL of FA_124 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n1);
   U1 : XNOR2_X1 port map( A => n1, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_126 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_126;

architecture SYN_BEHAVIORAL of FA_126 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n1);
   U1 : XNOR2_X1 port map( A => Ci, B => n1, ZN => S);
   U5 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n2);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n3);
   U3 : NAND2_X1 port map( A1 => n2, A2 => n3, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_0_0 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_0_0;

architecture SYN_BEHAVIORAL of FA_0_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity RCA_N4_24 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_24;

architecture SYN_STRUCTURAL of RCA_N4_24 is

   component FA_96
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_97
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_98
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_99
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal n2, CTMP_3_port, CTMP_2_port, CTMP_1_port, net684331 : std_logic;

begin
   
   n2 <= '1';
   FAI_1 : FA_99 port map( A => A(0), B => B(0), Ci => n2, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_98 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_97 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_96 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => net684331);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity RCA_N4_25 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_25;

architecture SYN_STRUCTURAL of RCA_N4_25 is

   component FA_100
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_101
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_102
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_103
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal n2, CTMP_3_port, CTMP_2_port, CTMP_1_port, net684330 : std_logic;

begin
   
   n2 <= '0';
   FAI_1 : FA_103 port map( A => A(0), B => B(0), Ci => n2, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_102 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_101 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_100 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => net684330);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity RCA_N4_27 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_27;

architecture SYN_STRUCTURAL of RCA_N4_27 is

   component FA_108
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_109
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_110
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_111
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal n2, CTMP_3_port, CTMP_2_port, n1, net684329 : std_logic;

begin
   
   n2 <= '0';
   FAI_1 : FA_111 port map( A => A(0), B => B(0), Ci => n2, S => S(0), Co => n1
                           );
   FAI_2 : FA_110 port map( A => A(1), B => B(1), Ci => n1, S => S(1), Co => 
                           CTMP_2_port);
   FAI_3 : FA_109 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_108 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => net684329);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity mux21_SIZE4_14 is

   port( IN0, IN1 : in std_logic_vector (3 downto 0);  CTRL : in std_logic;  
         OUT1 : out std_logic_vector (3 downto 0));

end mux21_SIZE4_14;

architecture SYN_Bhe of mux21_SIZE4_14 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => IN0(3), B => IN1(3), S => CTRL, Z => OUT1(3));
   U2 : MUX2_X1 port map( A => IN0(2), B => IN1(2), S => CTRL, Z => OUT1(2));
   U3 : MUX2_X1 port map( A => IN0(1), B => IN1(1), S => CTRL, Z => OUT1(1));
   U4 : MUX2_X1 port map( A => IN0(0), B => IN1(0), S => CTRL, Z => OUT1(0));

end SYN_Bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity RCA_N4_29 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_29;

architecture SYN_STRUCTURAL of RCA_N4_29 is

   component FA_116
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_117
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_118
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_119
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal n1, CTMP_3_port, CTMP_2_port, CTMP_1_port, net684328 : std_logic;

begin
   
   n1 <= '0';
   FAI_1 : FA_119 port map( A => A(0), B => B(0), Ci => n1, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_118 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_117 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_116 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => net684328);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity mux21_SIZE4_0_0 is

   port( IN0, IN1 : in std_logic_vector (3 downto 0);  CTRL : in std_logic;  
         OUT1 : out std_logic_vector (3 downto 0));

end mux21_SIZE4_0_0;

architecture SYN_Bhe of mux21_SIZE4_0_0 is

begin
   OUT1 <= ( IN0(3), IN0(2), IN0(1), IN0(0) );

end SYN_Bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity RCA_N4_0_0 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_0_0;

architecture SYN_STRUCTURAL of RCA_N4_0_0 is

   component FA_124
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_125
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_126
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_0_0
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal n1, CTMP_3_port, CTMP_2_port, CTMP_1_port, net684327 : std_logic;

begin
   
   n1 <= '0';
   FAI_1 : FA_0_0 port map( A => A(0), B => B(0), Ci => n1, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_126 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_125 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_124 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => net684327);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity shift_thirdLevel is

   port( sel : in std_logic_vector (2 downto 0);  A : in std_logic_vector (38 
         downto 0);  Y : out std_logic_vector (31 downto 0));

end shift_thirdLevel;

architecture SYN_behav of shift_thirdLevel is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n20, n21, n23, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
      n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50
      , n51, n52, n53, n54, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, 
      n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80
      , n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, 
      n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, 
      n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, 
      n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, 
      n132, n133, n136, n137, n138, n139, n252, n253, n254, n255, n256, n257, 
      n258, n259, n260 : std_logic;

begin
   
   U138 : OAI22_X1 port map( A1 => A(3), A2 => n257, B1 => A(1), B2 => n30, ZN 
                           => n137);
   U137 : AOI21_X1 port map( B1 => n256, B2 => n38, A => n137, ZN => n136);
   U136 : OAI21_X1 port map( B1 => A(5), B2 => n40, A => n136, ZN => n98);
   U43 : OAI22_X1 port map( A1 => A(30), A2 => n30, B1 => A(34), B2 => n40, ZN 
                           => n66);
   U42 : AOI21_X1 port map( B1 => n47, B2 => n65, A => n66, ZN => n64);
   U41 : OAI21_X1 port map( B1 => A(36), B2 => n255, A => n64, ZN => n56);
   U34 : OAI22_X1 port map( A1 => A(33), A2 => n257, B1 => A(35), B2 => n40, ZN
                           => n59);
   U33 : AOI21_X1 port map( B1 => n37, B2 => n58, A => n59, ZN => n57);
   U32 : OAI21_X1 port map( B1 => A(37), B2 => n255, A => n57, ZN => n54);
   U31 : AOI22_X1 port map( A1 => n259, A2 => n56, B1 => n54, B2 => n260, ZN =>
                           Y(30));
   U56 : OAI22_X1 port map( A1 => A(27), A2 => n30, B1 => A(31), B2 => n40, ZN 
                           => n77);
   U55 : AOI21_X1 port map( B1 => n47, B2 => n69, A => n77, ZN => n76);
   U54 : OAI21_X1 port map( B1 => A(33), B2 => n255, A => n76, ZN => n71);
   U150 : NAND2_X1 port map( A1 => n139, A2 => sel(2), ZN => n29);
   U52 : OAI22_X1 port map( A1 => A(30), A2 => n29, B1 => A(32), B2 => n40, ZN 
                           => n74);
   U51 : AOI21_X1 port map( B1 => n37, B2 => n73, A => n74, ZN => n72);
   U50 : OAI21_X1 port map( B1 => A(34), B2 => n255, A => n72, ZN => n67);
   U74 : OAI22_X1 port map( A1 => A(25), A2 => n257, B1 => A(27), B2 => n40, ZN
                           => n90);
   U73 : AOI21_X1 port map( B1 => n37, B2 => n89, A => n90, ZN => n88);
   U72 : OAI21_X1 port map( B1 => A(29), B2 => n255, A => n88, ZN => n84);
   U69 : OAI22_X1 port map( A1 => A(24), A2 => n30, B1 => A(26), B2 => n257, ZN
                           => n86);
   U68 : AOI21_X1 port map( B1 => n26, B2 => n73, A => n86, ZN => n85);
   U67 : OAI21_X1 port map( B1 => A(30), B2 => n255, A => n85, ZN => n81);
   U66 : AOI22_X1 port map( A1 => n258, A2 => n84, B1 => n81, B2 => n260, ZN =>
                           Y(23));
   U60 : OAI22_X1 port map( A1 => A(26), A2 => n30, B1 => A(30), B2 => n40, ZN 
                           => n80);
   U59 : AOI21_X1 port map( B1 => n47, B2 => n73, A => n80, ZN => n79);
   U58 : OAI21_X1 port map( B1 => A(32), B2 => n255, A => n79, ZN => n75);
   U53 : AOI22_X1 port map( A1 => n258, A2 => n75, B1 => n71, B2 => n260, ZN =>
                           Y(26));
   U78 : OAI22_X1 port map( A1 => A(24), A2 => n29, B1 => A(26), B2 => n40, ZN 
                           => n94);
   U77 : AOI21_X1 port map( B1 => n37, B2 => n93, A => n94, ZN => n92);
   U76 : OAI21_X1 port map( B1 => A(28), B2 => n255, A => n92, ZN => n87);
   U71 : AOI22_X1 port map( A1 => n258, A2 => n87, B1 => n84, B2 => n260, ZN =>
                           Y(22));
   U48 : OAI22_X1 port map( A1 => A(31), A2 => n257, B1 => A(33), B2 => n40, ZN
                           => n70);
   U47 : AOI21_X1 port map( B1 => n37, B2 => n69, A => n70, ZN => n68);
   U46 : OAI21_X1 port map( B1 => A(35), B2 => n255, A => n68, ZN => n63);
   U40 : AOI22_X1 port map( A1 => n259, A2 => n63, B1 => n56, B2 => n260, ZN =>
                           Y(29));
   U45 : AOI22_X1 port map( A1 => n258, A2 => n67, B1 => n63, B2 => n260, ZN =>
                           Y(28));
   U64 : OAI22_X1 port map( A1 => A(25), A2 => n30, B1 => A(27), B2 => n29, ZN 
                           => n83);
   U63 : AOI21_X1 port map( B1 => n26, B2 => n69, A => n83, ZN => n82);
   U62 : OAI21_X1 port map( B1 => A(31), B2 => n255, A => n82, ZN => n78);
   U57 : AOI22_X1 port map( A1 => sel(0), A2 => n78, B1 => n75, B2 => n260, ZN 
                           => Y(25));
   U82 : OAI22_X1 port map( A1 => A(21), A2 => n30, B1 => A(25), B2 => n40, ZN 
                           => n97);
   U81 : AOI21_X1 port map( B1 => n47, B2 => n89, A => n97, ZN => n96);
   U80 : OAI21_X1 port map( B1 => A(27), B2 => n255, A => n96, ZN => n91);
   U75 : AOI22_X1 port map( A1 => n258, A2 => n91, B1 => n87, B2 => n260, ZN =>
                           Y(21));
   U91 : OAI22_X1 port map( A1 => A(20), A2 => n30, B1 => A(24), B2 => n40, ZN 
                           => n103);
   U90 : AOI21_X1 port map( B1 => n47, B2 => n93, A => n103, ZN => n102);
   U89 : OAI21_X1 port map( B1 => A(26), B2 => n255, A => n102, ZN => n95);
   U79 : AOI22_X1 port map( A1 => n258, A2 => n95, B1 => n91, B2 => n260, ZN =>
                           Y(20));
   U61 : AOI22_X1 port map( A1 => sel(0), A2 => n81, B1 => n78, B2 => n260, ZN 
                           => Y(24));
   U30 : AOI22_X1 port map( A1 => n47, A2 => A(34), B1 => n37, B2 => A(32), ZN 
                           => n52);
   U29 : AOI22_X1 port map( A1 => n256, A2 => A(38), B1 => n26, B2 => A(36), ZN
                           => n53);
   U28 : OAI222_X1 port map( A1 => sel(0), A2 => n52, B1 => sel(0), B2 => n53, 
                           C1 => n54, C2 => n260, ZN => Y(31));
   U95 : OAI22_X1 port map( A1 => A(19), A2 => n30, B1 => A(21), B2 => n257, ZN
                           => n106);
   U94 : AOI21_X1 port map( B1 => n26, B2 => n89, A => n106, ZN => n105);
   U93 : OAI21_X1 port map( B1 => A(25), B2 => n255, A => n105, ZN => n101);
   U88 : AOI22_X1 port map( A1 => n258, A2 => n101, B1 => n95, B2 => n260, ZN 
                           => Y(19));
   U121 : OAI22_X1 port map( A1 => A(15), A2 => n257, B1 => A(13), B2 => n30, 
                           ZN => n126);
   U120 : AOI21_X1 port map( B1 => n26, B2 => n112, A => n126, ZN => n125);
   U119 : OAI21_X1 port map( B1 => A(19), B2 => n255, A => n125, ZN => n121);
   U117 : OAI22_X1 port map( A1 => A(14), A2 => n30, B1 => A(18), B2 => n40, ZN
                           => n123);
   U116 : AOI21_X1 port map( B1 => n47, B2 => n116, A => n123, ZN => n122);
   U115 : OAI21_X1 port map( B1 => A(20), B2 => n255, A => n122, ZN => n118);
   U114 : AOI22_X1 port map( A1 => n259, A2 => n121, B1 => n118, B2 => n260, ZN
                           => Y(13));
   U113 : OAI22_X1 port map( A1 => A(15), A2 => n30, B1 => A(19), B2 => n40, ZN
                           => n120);
   U112 : AOI21_X1 port map( B1 => n47, B2 => n112, A => n120, ZN => n119);
   U111 : OAI21_X1 port map( B1 => A(21), B2 => n255, A => n119, ZN => n114);
   U110 : AOI22_X1 port map( A1 => n259, A2 => n118, B1 => n114, B2 => n260, ZN
                           => Y(14));
   U125 : OAI22_X1 port map( A1 => A(14), A2 => n29, B1 => A(12), B2 => n30, ZN
                           => n129);
   U124 : AOI21_X1 port map( B1 => n26, B2 => n116, A => n129, ZN => n128);
   U123 : OAI21_X1 port map( B1 => A(18), B2 => n255, A => n128, ZN => n124);
   U118 : AOI22_X1 port map( A1 => n259, A2 => n124, B1 => n121, B2 => n260, ZN
                           => Y(12));
   U129 : OAI22_X1 port map( A1 => A(13), A2 => n257, B1 => A(11), B2 => n30, 
                           ZN => n131);
   U128 : AOI21_X1 port map( B1 => n256, B2 => n112, A => n131, ZN => n130);
   U127 : OAI21_X1 port map( B1 => A(15), B2 => n40, A => n130, ZN => n127);
   U122 : AOI22_X1 port map( A1 => n259, A2 => n127, B1 => n124, B2 => n260, ZN
                           => Y(11));
   U109 : OAI22_X1 port map( A1 => A(18), A2 => n29, B1 => A(20), B2 => n40, ZN
                           => n117);
   U108 : AOI21_X1 port map( B1 => n37, B2 => n116, A => n117, ZN => n115);
   U107 : OAI21_X1 port map( B1 => A(22), B2 => n255, A => n115, ZN => n110);
   U106 : AOI22_X1 port map( A1 => n259, A2 => n114, B1 => n110, B2 => n260, ZN
                           => Y(15));
   U15 : OAI22_X1 port map( A1 => A(11), A2 => n40, B1 => A(9), B2 => n29, ZN 
                           => n39);
   U14 : AOI21_X1 port map( B1 => n37, B2 => n38, A => n39, ZN => n36);
   U13 : OAI21_X1 port map( B1 => A(13), B2 => n255, A => n36, ZN => n31);
   U10 : OAI22_X1 port map( A1 => A(10), A2 => n29, B1 => A(8), B2 => n30, ZN 
                           => n34);
   U9 : AOI21_X1 port map( B1 => n26, B2 => n33, A => n34, ZN => n32);
   U8 : OAI21_X1 port map( B1 => A(14), B2 => n255, A => n32, ZN => n23);
   U7 : AOI22_X1 port map( A1 => n259, A2 => n31, B1 => n23, B2 => n260, ZN => 
                           Y(7));
   U105 : OAI22_X1 port map( A1 => A(19), A2 => n257, B1 => A(21), B2 => n40, 
                           ZN => n113);
   U104 : AOI21_X1 port map( B1 => n37, B2 => n112, A => n113, ZN => n111);
   U103 : OAI21_X1 port map( B1 => A(23), B2 => n255, A => n111, ZN => n107);
   U100 : OAI22_X1 port map( A1 => A(18), A2 => n30, B1 => A(20), B2 => n29, ZN
                           => n109);
   U99 : AOI21_X1 port map( B1 => n26, B2 => n93, A => n109, ZN => n108);
   U98 : OAI21_X1 port map( B1 => A(24), B2 => n255, A => n108, ZN => n104);
   U97 : AOI22_X1 port map( A1 => n259, A2 => n107, B1 => n104, B2 => n260, ZN 
                           => Y(17));
   U133 : OAI22_X1 port map( A1 => A(12), A2 => n29, B1 => A(10), B2 => n30, ZN
                           => n133);
   U132 : AOI21_X1 port map( B1 => n256, B2 => n116, A => n133, ZN => n132);
   U131 : OAI21_X1 port map( B1 => A(14), B2 => n40, A => n132, ZN => n21);
   U126 : AOI22_X1 port map( A1 => n259, A2 => n21, B1 => n127, B2 => n260, ZN 
                           => Y(10));
   U5 : OAI22_X1 port map( A1 => A(11), A2 => n257, B1 => A(9), B2 => n30, ZN 
                           => n28);
   U4 : AOI21_X1 port map( B1 => n26, B2 => n27, A => n28, ZN => n25);
   U3 : OAI21_X1 port map( B1 => A(15), B2 => n255, A => n25, ZN => n20);
   U1 : AOI22_X1 port map( A1 => n258, A2 => n20, B1 => n21, B2 => n260, ZN => 
                           Y(9));
   U39 : OAI22_X1 port map( A1 => A(5), A2 => n29, B1 => A(3), B2 => n30, ZN =>
                           n62);
   U38 : AOI21_X1 port map( B1 => n26, B2 => n38, A => n62, ZN => n61);
   U37 : OAI21_X1 port map( B1 => A(9), B2 => n255, A => n61, ZN => n49);
   U27 : OAI22_X1 port map( A1 => A(4), A2 => n30, B1 => A(8), B2 => n40, ZN =>
                           n51);
   U26 : AOI21_X1 port map( B1 => n47, B2 => n43, A => n51, ZN => n50);
   U25 : OAI21_X1 port map( B1 => A(10), B2 => n255, A => n50, ZN => n45);
   U24 : AOI22_X1 port map( A1 => sel(0), A2 => n49, B1 => n45, B2 => n260, ZN 
                           => Y(3));
   U86 : OAI22_X1 port map( A1 => A(2), A2 => n30, B1 => A(4), B2 => n29, ZN =>
                           n100);
   U85 : AOI21_X1 port map( B1 => n26, B2 => n43, A => n100, ZN => n99);
   U84 : OAI21_X1 port map( B1 => A(8), B2 => n255, A => n99, ZN => n60);
   U83 : AOI22_X1 port map( A1 => n258, A2 => n98, B1 => n60, B2 => n260, ZN =>
                           Y(1));
   U2 : AOI22_X1 port map( A1 => n259, A2 => n23, B1 => n20, B2 => n260, ZN => 
                           Y(8));
   U92 : AOI22_X1 port map( A1 => n259, A2 => n104, B1 => n101, B2 => n260, ZN 
                           => Y(18));
   U102 : AOI22_X1 port map( A1 => n259, A2 => n110, B1 => n107, B2 => n260, ZN
                           => Y(16));
   U23 : OAI22_X1 port map( A1 => A(5), A2 => n30, B1 => A(9), B2 => n40, ZN =>
                           n48);
   U22 : AOI21_X1 port map( B1 => n47, B2 => n38, A => n48, ZN => n46);
   U21 : OAI21_X1 port map( B1 => A(11), B2 => n255, A => n46, ZN => n41);
   U19 : OAI22_X1 port map( A1 => A(10), A2 => n40, B1 => A(8), B2 => n257, ZN 
                           => n44);
   U18 : AOI21_X1 port map( B1 => n37, B2 => n43, A => n44, ZN => n42);
   U17 : OAI21_X1 port map( B1 => A(12), B2 => n255, A => n42, ZN => n35);
   U16 : AOI22_X1 port map( A1 => sel(0), A2 => n41, B1 => n35, B2 => n260, ZN 
                           => Y(5));
   U20 : AOI22_X1 port map( A1 => n258, A2 => n45, B1 => n41, B2 => n260, ZN =>
                           Y(4));
   U12 : AOI22_X1 port map( A1 => n259, A2 => n35, B1 => n31, B2 => n260, ZN =>
                           Y(6));
   U148 : INV_X1 port map( A => sel(2), ZN => n138);
   U151 : INV_X1 port map( A => sel(1), ZN => n139);
   U142 : INV_X1 port map( A => n40, ZN => n26);
   U149 : INV_X1 port map( A => n257, ZN => n47);
   U139 : INV_X1 port map( A => n37, ZN => n30);
   U35 : INV_X1 port map( A => A(31), ZN => n58);
   U44 : INV_X1 port map( A => A(32), ZN => n65);
   U101 : INV_X1 port map( A => A(22), ZN => n93);
   U65 : INV_X1 port map( A => A(29), ZN => n69);
   U96 : INV_X1 port map( A => A(23), ZN => n89);
   U70 : INV_X1 port map( A => A(28), ZN => n73);
   U6 : INV_X1 port map( A => A(13), ZN => n27);
   U87 : INV_X1 port map( A => A(6), ZN => n43);
   U130 : INV_X1 port map( A => A(17), ZN => n112);
   U134 : INV_X1 port map( A => A(16), ZN => n116);
   U11 : INV_X1 port map( A => A(12), ZN => n33);
   U36 : AOI22_X1 port map( A1 => A(4), A2 => n26, B1 => A(6), B2 => n256, ZN 
                           => n252);
   U49 : AOI22_X1 port map( A1 => A(0), A2 => n37, B1 => A(2), B2 => n47, ZN =>
                           n253);
   U135 : AND2_X1 port map( A1 => n252, A2 => n253, ZN => n254);
   U140 : OAI22_X1 port map( A1 => n260, A2 => n254, B1 => n259, B2 => n98, ZN 
                           => Y(0));
   U141 : AOI22_X1 port map( A1 => n260, A2 => n49, B1 => n60, B2 => n259, ZN 
                           => Y(2));
   U143 : INV_X1 port map( A => A(7), ZN => n38);
   U144 : AOI22_X1 port map( A1 => n260, A2 => n67, B1 => n71, B2 => n258, ZN 
                           => Y(27));
   U145 : NAND2_X2 port map( A1 => n138, A2 => sel(1), ZN => n40);
   U146 : CLKBUF_X1 port map( A => sel(0), Z => n258);
   U147 : INV_X2 port map( A => sel(0), ZN => n260);
   U152 : INV_X2 port map( A => n256, ZN => n255);
   U153 : NOR2_X1 port map( A1 => n138, A2 => n139, ZN => n37);
   U154 : AND2_X1 port map( A1 => n138, A2 => n139, ZN => n256);
   U155 : BUF_X1 port map( A => sel(0), Z => n259);
   U156 : NAND2_X1 port map( A1 => n139, A2 => sel(2), ZN => n257);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity shift_secondLevel is

   port( sel : in std_logic_vector (1 downto 0);  mask00, mask08, mask16 : in 
         std_logic_vector (38 downto 0);  Y : out std_logic_vector (38 downto 
         0));

end shift_secondLevel;

architecture SYN_behav of shift_secondLevel is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n41, n42, n43, n44, n45, n47, n48, n49, n50, n51, n52, n53, n54, n55,
      n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70
      , n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n83, n136, n137,
      n138, n139, n140 : std_logic;

begin
   
   U35 : AOI222_X1 port map( A1 => n139, A2 => mask00(2), B1 => n43, B2 => 
                           mask08(2), C1 => n138, C2 => mask16(2), ZN => n60);
   U9 : AOI222_X1 port map( A1 => n139, A2 => mask00(6), B1 => n43, B2 => 
                           mask08(6), C1 => n138, C2 => mask16(6), ZN => n47);
   U13 : AOI222_X1 port map( A1 => n139, A2 => mask00(4), B1 => n43, B2 => 
                           mask08(4), C1 => n138, C2 => mask16(4), ZN => n49);
   U11 : AOI222_X1 port map( A1 => n139, A2 => mask00(5), B1 => n43, B2 => 
                           mask08(5), C1 => n138, C2 => mask16(5), ZN => n48);
   U15 : AOI222_X1 port map( A1 => n139, A2 => mask00(3), B1 => n43, B2 => 
                           mask08(3), C1 => n138, C2 => mask16(3), ZN => n50);
   U57 : AOI222_X1 port map( A1 => n139, A2 => mask00(1), B1 => n140, B2 => 
                           mask08(1), C1 => n138, C2 => mask16(1), ZN => n71);
   U21 : AOI222_X1 port map( A1 => n139, A2 => mask00(36), B1 => n43, B2 => 
                           mask08(36), C1 => n138, C2 => mask16(36), ZN => n53)
                           ;
   U29 : AOI222_X1 port map( A1 => n139, A2 => mask00(32), B1 => n43, B2 => 
                           mask08(32), C1 => n138, C2 => mask16(32), ZN => n57)
                           ;
   U33 : AOI222_X1 port map( A1 => n139, A2 => mask00(30), B1 => n43, B2 => 
                           mask08(30), C1 => n138, C2 => mask16(30), ZN => n59)
                           ;
   U25 : AOI222_X1 port map( A1 => n139, A2 => mask00(34), B1 => n43, B2 => 
                           mask08(34), C1 => n138, C2 => mask16(34), ZN => n55)
                           ;
   U19 : AOI222_X1 port map( A1 => n139, A2 => mask00(37), B1 => n43, B2 => 
                           mask08(37), C1 => n138, C2 => mask16(37), ZN => n52)
                           ;
   U31 : AOI222_X1 port map( A1 => n139, A2 => mask00(31), B1 => n43, B2 => 
                           mask08(31), C1 => n138, C2 => mask16(31), ZN => n58)
                           ;
   U27 : AOI222_X1 port map( A1 => n139, A2 => mask00(33), B1 => n43, B2 => 
                           mask08(33), C1 => n138, C2 => mask16(33), ZN => n56)
                           ;
   U23 : AOI222_X1 port map( A1 => n139, A2 => mask00(35), B1 => n43, B2 => 
                           mask08(35), C1 => n138, C2 => mask16(35), ZN => n54)
                           ;
   U37 : AOI222_X1 port map( A1 => n139, A2 => mask00(29), B1 => n43, B2 => 
                           mask08(29), C1 => n138, C2 => mask16(29), ZN => n61)
                           ;
   U41 : AOI222_X1 port map( A1 => n139, A2 => mask00(27), B1 => n43, B2 => 
                           mask08(27), C1 => n138, C2 => mask16(27), ZN => n63)
                           ;
   U39 : AOI222_X1 port map( A1 => n139, A2 => mask00(28), B1 => n43, B2 => 
                           mask08(28), C1 => n138, C2 => mask16(28), ZN => n62)
                           ;
   U49 : AOI222_X1 port map( A1 => n139, A2 => mask00(23), B1 => n43, B2 => 
                           mask08(23), C1 => n138, C2 => mask16(23), ZN => n67)
                           ;
   U45 : AOI222_X1 port map( A1 => n139, A2 => mask00(25), B1 => n140, B2 => 
                           mask08(25), C1 => n138, C2 => mask16(25), ZN => n65)
                           ;
   U47 : AOI222_X1 port map( A1 => n139, A2 => mask00(24), B1 => n43, B2 => 
                           mask08(24), C1 => n138, C2 => mask16(24), ZN => n66)
                           ;
   U43 : AOI222_X1 port map( A1 => n139, A2 => mask00(26), B1 => n43, B2 => 
                           mask08(26), C1 => n138, C2 => mask16(26), ZN => n64)
                           ;
   U51 : AOI222_X1 port map( A1 => n139, A2 => mask00(22), B1 => n43, B2 => 
                           mask08(22), C1 => n138, C2 => mask16(22), ZN => n68)
                           ;
   U53 : AOI222_X1 port map( A1 => n139, A2 => mask00(21), B1 => n43, B2 => 
                           mask08(21), C1 => n138, C2 => mask16(21), ZN => n69)
                           ;
   U55 : AOI222_X1 port map( A1 => n139, A2 => mask00(20), B1 => n43, B2 => 
                           mask08(20), C1 => n138, C2 => mask16(20), ZN => n70)
                           ;
   U17 : AOI222_X1 port map( A1 => n139, A2 => mask00(38), B1 => n140, B2 => 
                           mask08(38), C1 => n138, C2 => mask16(38), ZN => n51)
                           ;
   U59 : AOI222_X1 port map( A1 => n139, A2 => mask00(19), B1 => n140, B2 => 
                           mask08(19), C1 => n138, C2 => mask16(19), ZN => n72)
                           ;
   U63 : AOI222_X1 port map( A1 => n139, A2 => mask00(17), B1 => n140, B2 => 
                           mask08(17), C1 => n138, C2 => mask16(17), ZN => n74)
                           ;
   U67 : AOI222_X1 port map( A1 => n139, A2 => mask00(15), B1 => n140, B2 => 
                           mask08(15), C1 => n138, C2 => mask16(15), ZN => n76)
                           ;
   U71 : AOI222_X1 port map( A1 => n139, A2 => mask00(13), B1 => n140, B2 => 
                           mask08(13), C1 => n138, C2 => mask16(13), ZN => n78)
                           ;
   U65 : AOI222_X1 port map( A1 => n139, A2 => mask00(16), B1 => n140, B2 => 
                           mask08(16), C1 => n138, C2 => mask16(16), ZN => n75)
                           ;
   U69 : AOI222_X1 port map( A1 => n139, A2 => mask00(14), B1 => n140, B2 => 
                           mask08(14), C1 => n138, C2 => mask16(14), ZN => n77)
                           ;
   U61 : AOI222_X1 port map( A1 => n139, A2 => mask00(18), B1 => n140, B2 => 
                           mask08(18), C1 => n138, C2 => mask16(18), ZN => n73)
                           ;
   U73 : AOI222_X1 port map( A1 => n139, A2 => mask00(12), B1 => n140, B2 => 
                           mask08(12), C1 => n138, C2 => mask16(12), ZN => n79)
                           ;
   U75 : AOI222_X1 port map( A1 => n139, A2 => mask00(11), B1 => n140, B2 => 
                           mask08(11), C1 => n138, C2 => mask16(11), ZN => n80)
                           ;
   U3 : AOI222_X1 port map( A1 => n139, A2 => mask00(9), B1 => n43, B2 => 
                           mask08(9), C1 => n138, C2 => mask16(9), ZN => n41);
   U77 : AOI222_X1 port map( A1 => n139, A2 => mask00(10), B1 => n140, B2 => 
                           mask08(10), C1 => n138, C2 => mask16(10), ZN => n81)
                           ;
   U5 : AOI222_X1 port map( A1 => n139, A2 => mask00(8), B1 => n43, B2 => 
                           mask08(8), C1 => n138, C2 => mask16(8), ZN => n45);
   U34 : INV_X1 port map( A => n60, ZN => Y(2));
   U58 : INV_X1 port map( A => n72, ZN => Y(19));
   U54 : INV_X1 port map( A => n70, ZN => Y(20));
   U52 : INV_X1 port map( A => n69, ZN => Y(21));
   U64 : INV_X1 port map( A => n75, ZN => Y(16));
   U10 : INV_X1 port map( A => n48, ZN => Y(5));
   U60 : INV_X1 port map( A => n73, ZN => Y(18));
   U68 : INV_X1 port map( A => n77, ZN => Y(14));
   U62 : INV_X1 port map( A => n74, ZN => Y(17));
   U56 : INV_X1 port map( A => n71, ZN => Y(1));
   U14 : INV_X1 port map( A => n50, ZN => Y(3));
   U70 : INV_X1 port map( A => n78, ZN => Y(13));
   U66 : INV_X1 port map( A => n76, ZN => Y(15));
   U12 : INV_X1 port map( A => n49, ZN => Y(4));
   U8 : INV_X1 port map( A => n47, ZN => Y(6));
   U22 : INV_X1 port map( A => n54, ZN => Y(35));
   U4 : INV_X1 port map( A => n45, ZN => Y(8));
   U76 : INV_X1 port map( A => n81, ZN => Y(10));
   U48 : INV_X1 port map( A => n67, ZN => Y(23));
   U26 : INV_X1 port map( A => n56, ZN => Y(33));
   U32 : INV_X1 port map( A => n59, ZN => Y(30));
   U46 : INV_X1 port map( A => n66, ZN => Y(24));
   U2 : INV_X1 port map( A => n41, ZN => Y(9));
   U42 : INV_X1 port map( A => n64, ZN => Y(26));
   U40 : INV_X1 port map( A => n63, ZN => Y(27));
   U20 : INV_X1 port map( A => n53, ZN => Y(36));
   U28 : INV_X1 port map( A => n57, ZN => Y(32));
   U74 : INV_X1 port map( A => n80, ZN => Y(11));
   U16 : INV_X1 port map( A => n51, ZN => Y(38));
   U24 : INV_X1 port map( A => n55, ZN => Y(34));
   U36 : INV_X1 port map( A => n61, ZN => Y(29));
   U44 : INV_X1 port map( A => n65, ZN => Y(25));
   U50 : INV_X1 port map( A => n68, ZN => Y(22));
   U18 : INV_X1 port map( A => n52, ZN => Y(37));
   U72 : INV_X1 port map( A => n79, ZN => Y(12));
   U38 : INV_X1 port map( A => n62, ZN => Y(28));
   U30 : INV_X1 port map( A => n58, ZN => Y(31));
   U6 : AOI222_X1 port map( A1 => mask00(0), A2 => n139, B1 => mask16(0), B2 =>
                           n138, C1 => mask08(0), C2 => n140, ZN => n136);
   U7 : INV_X1 port map( A => n136, ZN => Y(0));
   U78 : AOI222_X1 port map( A1 => n43, A2 => mask08(7), B1 => n138, B2 => 
                           mask16(7), C1 => mask00(7), C2 => n139, ZN => n137);
   U79 : INV_X1 port map( A => n137, ZN => Y(7));
   U80 : AND2_X2 port map( A1 => n83, A2 => sel(0), ZN => n43);
   U81 : BUF_X2 port map( A => n44, Z => n138);
   U82 : BUF_X2 port map( A => n42, Z => n139);
   U83 : INV_X1 port map( A => sel(1), ZN => n83);
   U84 : BUF_X1 port map( A => n43, Z => n140);
   U85 : NOR2_X1 port map( A1 => sel(0), A2 => n83, ZN => n44);
   U86 : NOR2_X1 port map( A1 => sel(1), A2 => sel(0), ZN => n42);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity shift_firstLevel is

   port( A : in std_logic_vector (31 downto 0);  sel : in std_logic_vector (1 
         downto 0);  mask00, mask08, mask16 : out std_logic_vector (38 downto 
         0));

end shift_firstLevel;

architecture SYN_behav of shift_firstLevel is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal mask08_38_port, mask08_37_port, mask08_36_port, mask08_35_port, 
      mask08_34_port, mask08_33_port, mask08_32_port, mask08_31_port, 
      mask08_23_port, mask08_22_port, mask08_21_port, mask08_20_port, 
      mask08_19_port, mask08_18_port, mask08_17_port, mask08_16_port, 
      mask08_15_port, mask08_7_port, mask08_6_port, mask08_5_port, 
      mask08_4_port, mask08_3_port, mask08_2_port, mask08_1_port, mask08_0_port
      , mask16_38_port, mask16_37_port, mask16_36_port, mask16_35_port, 
      mask16_34_port, mask16_33_port, mask16_32_port, mask16_31_port, 
      mask16_30_port, mask16_29_port, mask16_28_port, mask16_27_port, 
      mask16_26_port, mask16_25_port, mask16_24_port, mask16_23_port, 
      mask16_15_port, mask16_14_port, mask16_13_port, mask16_12_port, 
      mask16_11_port, mask16_10_port, mask16_9_port, mask16_8_port, 
      mask16_7_port, mask16_6_port, mask16_5_port, mask16_4_port, mask16_3_port
      , mask16_2_port, mask16_1_port, mask16_0_port, n36, n37, n38, n39, n40, 
      n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55
      , n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, 
      n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84
      , n85, n88, n89, n90, n91, n92, n93, n94, n95, n158, n159, mask16_17_port
      : std_logic;

begin
   mask08 <= ( mask08_38_port, mask08_37_port, mask08_36_port, mask08_35_port, 
      mask08_34_port, mask08_33_port, mask08_32_port, mask08_31_port, 
      mask16_38_port, mask16_37_port, mask16_36_port, mask16_35_port, 
      mask16_34_port, mask16_33_port, mask16_32_port, mask08_23_port, 
      mask08_22_port, mask08_21_port, mask08_20_port, mask08_19_port, 
      mask08_18_port, mask08_17_port, mask08_16_port, mask08_15_port, 
      mask16_6_port, mask16_5_port, mask16_4_port, mask16_3_port, mask16_2_port
      , mask16_1_port, mask16_0_port, mask08_7_port, mask08_6_port, 
      mask08_5_port, mask08_4_port, mask08_3_port, mask08_2_port, mask08_1_port
      , mask08_0_port );
   mask16 <= ( mask16_38_port, mask16_37_port, mask16_36_port, mask16_35_port, 
      mask16_34_port, mask16_33_port, mask16_32_port, mask16_31_port, 
      mask16_30_port, mask16_29_port, mask16_28_port, mask16_27_port, 
      mask16_26_port, mask16_25_port, mask16_24_port, mask16_23_port, 
      mask16_17_port, mask16_17_port, mask16_17_port, mask16_17_port, 
      mask16_17_port, mask16_17_port, mask16_17_port, mask16_15_port, 
      mask16_14_port, mask16_13_port, mask16_12_port, mask16_11_port, 
      mask16_10_port, mask16_9_port, mask16_8_port, mask16_7_port, 
      mask16_6_port, mask16_5_port, mask16_4_port, mask16_3_port, mask16_2_port
      , mask16_1_port, mask16_0_port );
   
   U155 : NAND2_X1 port map( A1 => sel(0), A2 => A(10), ZN => n81);
   U131 : NAND2_X1 port map( A1 => sel(0), A2 => A(18), ZN => n53);
   U62 : NAND2_X1 port map( A1 => sel(0), A2 => A(8), ZN => n84);
   U137 : NAND2_X1 port map( A1 => sel(0), A2 => A(16), ZN => n67);
   U143 : NAND2_X1 port map( A1 => sel(0), A2 => A(14), ZN => n69);
   U119 : NAND2_X1 port map( A1 => sel(0), A2 => A(22), ZN => n39);
   U149 : NAND2_X1 port map( A1 => sel(0), A2 => A(12), ZN => n71);
   U125 : NAND2_X1 port map( A1 => sel(0), A2 => A(20), ZN => n41);
   U146 : NAND2_X1 port map( A1 => sel(0), A2 => A(13), ZN => n70);
   U122 : NAND2_X1 port map( A1 => sel(0), A2 => A(21), ZN => n40);
   U157 : NOR2_X1 port map( A1 => sel(0), A2 => sel(1), ZN => n85);
   U67 : NAND2_X1 port map( A1 => n159, A2 => A(0), ZN => n60);
   U140 : NAND2_X1 port map( A1 => sel(0), A2 => A(15), ZN => n68);
   U116 : NAND2_X1 port map( A1 => sel(0), A2 => A(23), ZN => n38);
   U152 : NAND2_X1 port map( A1 => sel(0), A2 => A(11), ZN => n72);
   U129 : NAND2_X1 port map( A1 => sel(0), A2 => A(19), ZN => n42);
   U59 : NAND2_X1 port map( A1 => sel(0), A2 => A(9), ZN => n83);
   U134 : NAND2_X1 port map( A1 => sel(0), A2 => A(17), ZN => n61);
   U91 : NAND2_X1 port map( A1 => sel(0), A2 => A(31), ZN => n82);
   U77 : AOI21_X1 port map( B1 => A(29), B2 => n159, A => mask16_17_port, ZN =>
                           n90);
   U100 : NAND2_X1 port map( A1 => n159, A2 => A(21), ZN => n75);
   U40 : NAND2_X1 port map( A1 => n75, A2 => n44, ZN => mask08_36_port);
   U124 : NAND2_X1 port map( A1 => n159, A2 => A(13), ZN => n46);
   U11 : NAND2_X1 port map( A1 => n46, A2 => n44, ZN => mask16_36_port);
   U85 : AOI21_X1 port map( B1 => A(25), B2 => n159, A => mask16_17_port, ZN =>
                           n94);
   U112 : NAND2_X1 port map( A1 => n159, A2 => A(17), ZN => n79);
   U44 : NAND2_X1 port map( A1 => n79, A2 => n44, ZN => mask08_32_port);
   U138 : NAND2_X1 port map( A1 => n85, A2 => A(9), ZN => n50);
   U15 : NAND2_X1 port map( A1 => n50, A2 => n44, ZN => mask16_32_port);
   U94 : NAND2_X1 port map( A1 => sel(0), A2 => A(30), ZN => n62);
   U93 : NAND2_X1 port map( A1 => n159, A2 => A(23), ZN => n73);
   U92 : NAND2_X1 port map( A1 => n62, A2 => n73, ZN => mask00(30));
   U118 : NAND2_X1 port map( A1 => n159, A2 => A(15), ZN => n43);
   U9 : NAND2_X1 port map( A1 => n43, A2 => n44, ZN => mask16_38_port);
   U144 : NAND2_X1 port map( A1 => n85, A2 => A(7), ZN => n52);
   U17 : NAND2_X1 port map( A1 => n52, A2 => n44, ZN => mask16_30_port);
   U81 : AOI21_X1 port map( B1 => A(27), B2 => n159, A => mask16_17_port, ZN =>
                           n92);
   U106 : NAND2_X1 port map( A1 => n159, A2 => A(19), ZN => n77);
   U42 : NAND2_X1 port map( A1 => n77, A2 => n44, ZN => mask08_34_port);
   U132 : NAND2_X1 port map( A1 => n159, A2 => A(11), ZN => n48);
   U13 : NAND2_X1 port map( A1 => n48, A2 => n44, ZN => mask16_34_port);
   U75 : AOI21_X1 port map( B1 => A(30), B2 => n159, A => mask16_17_port, ZN =>
                           n89);
   U97 : NAND2_X1 port map( A1 => n159, A2 => A(22), ZN => n74);
   U39 : NAND2_X1 port map( A1 => n74, A2 => n44, ZN => mask08_37_port);
   U121 : NAND2_X1 port map( A1 => n159, A2 => A(14), ZN => n45);
   U10 : NAND2_X1 port map( A1 => n45, A2 => n44, ZN => mask16_37_port);
   U89 : AOI21_X1 port map( B1 => A(24), B2 => n159, A => mask16_15_port, ZN =>
                           n95);
   U115 : NAND2_X1 port map( A1 => n159, A2 => A(16), ZN => n80);
   U45 : NAND2_X1 port map( A1 => n80, A2 => n44, ZN => mask08_31_port);
   U141 : NAND2_X1 port map( A1 => n85, A2 => A(8), ZN => n51);
   U16 : NAND2_X1 port map( A1 => n51, A2 => n44, ZN => mask16_31_port);
   U83 : AOI21_X1 port map( B1 => A(26), B2 => n159, A => mask16_17_port, ZN =>
                           n93);
   U109 : NAND2_X1 port map( A1 => n159, A2 => A(18), ZN => n78);
   U43 : NAND2_X1 port map( A1 => n78, A2 => n44, ZN => mask08_33_port);
   U135 : NAND2_X1 port map( A1 => n85, A2 => A(10), ZN => n49);
   U14 : NAND2_X1 port map( A1 => n49, A2 => n44, ZN => mask16_33_port);
   U79 : AOI21_X1 port map( B1 => A(28), B2 => n159, A => mask16_17_port, ZN =>
                           n91);
   U103 : NAND2_X1 port map( A1 => n159, A2 => A(20), ZN => n76);
   U41 : NAND2_X1 port map( A1 => n76, A2 => n44, ZN => mask08_35_port);
   U128 : NAND2_X1 port map( A1 => n85, A2 => A(12), ZN => n47);
   U12 : NAND2_X1 port map( A1 => n47, A2 => n44, ZN => mask16_35_port);
   U98 : NAND2_X1 port map( A1 => sel(0), A2 => A(29), ZN => n63);
   U96 : NAND2_X1 port map( A1 => n63, A2 => n74, ZN => mask00(29));
   U147 : NAND2_X1 port map( A1 => n159, A2 => A(6), ZN => n54);
   U19 : NAND2_X1 port map( A1 => n54, A2 => n44, ZN => mask16_29_port);
   U104 : NAND2_X1 port map( A1 => sel(0), A2 => A(27), ZN => n65);
   U102 : NAND2_X1 port map( A1 => n65, A2 => n76, ZN => mask00(27));
   U153 : NAND2_X1 port map( A1 => n159, A2 => A(4), ZN => n56);
   U21 : NAND2_X1 port map( A1 => n56, A2 => n44, ZN => mask16_27_port);
   U101 : NAND2_X1 port map( A1 => sel(0), A2 => A(28), ZN => n64);
   U99 : NAND2_X1 port map( A1 => n64, A2 => n75, ZN => mask00(28));
   U150 : NAND2_X1 port map( A1 => n159, A2 => A(5), ZN => n55);
   U20 : NAND2_X1 port map( A1 => n55, A2 => n44, ZN => mask16_28_port);
   U114 : NAND2_X1 port map( A1 => n38, A2 => n80, ZN => mask00(23));
   U47 : NAND2_X1 port map( A1 => n51, A2 => n82, ZN => mask08_23_port);
   U25 : NAND2_X1 port map( A1 => n44, A2 => n60, ZN => mask16_23_port);
   U110 : NAND2_X1 port map( A1 => sel(0), A2 => A(25), ZN => n36);
   U108 : NAND2_X1 port map( A1 => n36, A2 => n78, ZN => mask00(25));
   U60 : NAND2_X1 port map( A1 => n159, A2 => A(2), ZN => n58);
   U23 : NAND2_X1 port map( A1 => n44, A2 => n58, ZN => mask16_25_port);
   U113 : NAND2_X1 port map( A1 => sel(0), A2 => A(24), ZN => n37);
   U111 : NAND2_X1 port map( A1 => n37, A2 => n79, ZN => mask00(24));
   U63 : NAND2_X1 port map( A1 => n159, A2 => A(1), ZN => n59);
   U24 : NAND2_X1 port map( A1 => n44, A2 => n59, ZN => mask16_24_port);
   U107 : NAND2_X1 port map( A1 => sel(0), A2 => A(26), ZN => n66);
   U105 : NAND2_X1 port map( A1 => n66, A2 => n77, ZN => mask00(26));
   U156 : NAND2_X1 port map( A1 => n85, A2 => A(3), ZN => n57);
   U22 : NAND2_X1 port map( A1 => n57, A2 => n44, ZN => mask16_26_port);
   U117 : NAND2_X1 port map( A1 => n39, A2 => n43, ZN => mask00(22));
   U48 : NAND2_X1 port map( A1 => n52, A2 => n62, ZN => mask08_22_port);
   U120 : NAND2_X1 port map( A1 => n40, A2 => n45, ZN => mask00(21));
   U49 : NAND2_X1 port map( A1 => n54, A2 => n63, ZN => mask08_21_port);
   U123 : NAND2_X1 port map( A1 => n41, A2 => n46, ZN => mask00(20));
   U50 : NAND2_X1 port map( A1 => n55, A2 => n64, ZN => mask08_20_port);
   U73 : AOI21_X1 port map( B1 => A(31), B2 => n159, A => mask16_17_port, ZN =>
                           n88);
   U38 : NAND2_X1 port map( A1 => n73, A2 => n44, ZN => mask08_38_port);
   U127 : NAND2_X1 port map( A1 => n42, A2 => n47, ZN => mask00(19));
   U52 : NAND2_X1 port map( A1 => n56, A2 => n65, ZN => mask08_19_port);
   U133 : NAND2_X1 port map( A1 => n49, A2 => n61, ZN => mask00(17));
   U54 : NAND2_X1 port map( A1 => n36, A2 => n58, ZN => mask08_17_port);
   U139 : NAND2_X1 port map( A1 => n51, A2 => n68, ZN => mask00(15));
   U56 : NAND2_X1 port map( A1 => n38, A2 => n60, ZN => mask08_15_port);
   U145 : NAND2_X1 port map( A1 => n54, A2 => n70, ZN => mask00(13));
   U136 : NAND2_X1 port map( A1 => n50, A2 => n67, ZN => mask00(16));
   U55 : NAND2_X1 port map( A1 => n37, A2 => n59, ZN => mask08_16_port);
   U142 : NAND2_X1 port map( A1 => n52, A2 => n69, ZN => mask00(14));
   U130 : NAND2_X1 port map( A1 => n48, A2 => n53, ZN => mask00(18));
   U53 : NAND2_X1 port map( A1 => n57, A2 => n66, ZN => mask08_18_port);
   U148 : NAND2_X1 port map( A1 => n55, A2 => n71, ZN => mask00(12));
   U151 : NAND2_X1 port map( A1 => n56, A2 => n72, ZN => mask00(11));
   U58 : NAND2_X1 port map( A1 => n58, A2 => n83, ZN => mask00(9));
   U154 : NAND2_X1 port map( A1 => n57, A2 => n81, ZN => mask00(10));
   U61 : NAND2_X1 port map( A1 => n59, A2 => n84, ZN => mask00(8));
   U69 : AND2_X1 port map( A1 => sel(0), A2 => A(5), ZN => mask00(5));
   U126 : AND2_X1 port map( A1 => sel(0), A2 => A(1), ZN => mask00(1));
   U71 : AND2_X1 port map( A1 => sel(0), A2 => A(3), ZN => mask00(3));
   U70 : AND2_X1 port map( A1 => sel(0), A2 => A(4), ZN => mask00(4));
   U68 : AND2_X1 port map( A1 => sel(0), A2 => A(6), ZN => mask00(6));
   U95 : AND2_X1 port map( A1 => sel(0), A2 => A(2), ZN => mask00(2));
   U51 : INV_X1 port map( A => n83, ZN => mask08_1_port);
   U31 : INV_X1 port map( A => n66, ZN => mask16_10_port);
   U3 : INV_X1 port map( A => n37, ZN => mask16_8_port);
   U26 : INV_X1 port map( A => n61, ZN => mask16_1_port);
   U30 : INV_X1 port map( A => n65, ZN => mask16_11_port);
   U18 : INV_X1 port map( A => n53, ZN => mask16_2_port);
   U6 : INV_X1 port map( A => n40, ZN => mask16_5_port);
   U46 : INV_X1 port map( A => n81, ZN => mask08_2_port);
   U35 : INV_X1 port map( A => n70, ZN => mask08_5_port);
   U90 : INV_X1 port map( A => n82, ZN => mask16_15_port);
   U2 : INV_X1 port map( A => n36, ZN => mask16_9_port);
   U28 : INV_X1 port map( A => n63, ZN => mask16_13_port);
   U29 : INV_X1 port map( A => n64, ZN => mask16_12_port);
   U37 : INV_X1 port map( A => n72, ZN => mask08_3_port);
   U34 : INV_X1 port map( A => n69, ZN => mask08_6_port);
   U5 : INV_X1 port map( A => n39, ZN => mask16_6_port);
   U8 : INV_X1 port map( A => n42, ZN => mask16_3_port);
   U27 : INV_X1 port map( A => n62, ZN => mask16_14_port);
   U36 : INV_X1 port map( A => n71, ZN => mask08_4_port);
   U32 : INV_X1 port map( A => n67, ZN => mask16_0_port);
   U7 : INV_X1 port map( A => n41, ZN => mask16_4_port);
   U88 : INV_X1 port map( A => n95, ZN => mask00(31));
   U74 : INV_X1 port map( A => n89, ZN => mask00(37));
   U78 : INV_X1 port map( A => n91, ZN => mask00(35));
   U76 : INV_X1 port map( A => n90, ZN => mask00(36));
   U72 : INV_X1 port map( A => n88, ZN => mask00(38));
   U82 : INV_X1 port map( A => n93, ZN => mask00(33));
   U80 : INV_X1 port map( A => n92, ZN => mask00(34));
   U84 : INV_X1 port map( A => n94, ZN => mask00(32));
   U4 : INV_X1 port map( A => n84, ZN => mask08_0_port);
   U33 : AND2_X1 port map( A1 => sel(0), A2 => A(0), ZN => mask00(0));
   U57 : INV_X1 port map( A => n38, ZN => mask16_7_port);
   U64 : INV_X1 port map( A => n68, ZN => mask08_7_port);
   U65 : NAND2_X1 port map( A1 => sel(0), A2 => A(7), ZN => n158);
   U66 : NAND2_X1 port map( A1 => n60, A2 => n158, ZN => mask00(7));
   U86 : NAND2_X1 port map( A1 => sel(1), A2 => mask16_15_port, ZN => n44);
   U87 : INV_X1 port map( A => n44, ZN => mask16_17_port);
   U158 : BUF_X1 port map( A => n85, Z => n159);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity mux21_1 is

   port( IN0, IN1 : in std_logic_vector (31 downto 0);  CTRL : in std_logic;  
         OUT1 : out std_logic_vector (31 downto 0));

end mux21_1;

architecture SYN_Bhe of mux21_1 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U3 : MUX2_X1 port map( A => IN0(9), B => IN1(9), S => CTRL, Z => OUT1(9));
   U4 : MUX2_X1 port map( A => IN0(8), B => IN1(8), S => CTRL, Z => OUT1(8));
   U5 : MUX2_X1 port map( A => IN0(7), B => IN1(7), S => CTRL, Z => OUT1(7));
   U6 : MUX2_X1 port map( A => IN0(6), B => IN1(6), S => CTRL, Z => OUT1(6));
   U7 : MUX2_X1 port map( A => IN0(5), B => IN1(5), S => CTRL, Z => OUT1(5));
   U8 : MUX2_X1 port map( A => IN0(4), B => IN1(4), S => CTRL, Z => OUT1(4));
   U10 : MUX2_X1 port map( A => IN0(31), B => IN1(31), S => CTRL, Z => OUT1(31)
                           );
   U11 : MUX2_X1 port map( A => IN0(30), B => IN1(30), S => CTRL, Z => OUT1(30)
                           );
   U12 : MUX2_X1 port map( A => IN0(2), B => IN1(2), S => CTRL, Z => OUT1(2));
   U14 : MUX2_X1 port map( A => IN0(28), B => IN1(28), S => CTRL, Z => OUT1(28)
                           );
   U15 : MUX2_X1 port map( A => IN0(27), B => IN1(27), S => CTRL, Z => OUT1(27)
                           );
   U16 : MUX2_X1 port map( A => IN0(26), B => IN1(26), S => CTRL, Z => OUT1(26)
                           );
   U17 : MUX2_X1 port map( A => IN0(25), B => IN1(25), S => CTRL, Z => OUT1(25)
                           );
   U18 : MUX2_X1 port map( A => IN0(24), B => IN1(24), S => CTRL, Z => OUT1(24)
                           );
   U19 : MUX2_X1 port map( A => IN0(23), B => IN1(23), S => CTRL, Z => OUT1(23)
                           );
   U20 : MUX2_X1 port map( A => IN0(22), B => IN1(22), S => CTRL, Z => OUT1(22)
                           );
   U21 : MUX2_X1 port map( A => IN0(21), B => IN1(21), S => CTRL, Z => OUT1(21)
                           );
   U22 : MUX2_X1 port map( A => IN0(20), B => IN1(20), S => CTRL, Z => OUT1(20)
                           );
   U23 : MUX2_X1 port map( A => IN0(1), B => IN1(1), S => CTRL, Z => OUT1(1));
   U24 : MUX2_X1 port map( A => IN0(19), B => IN1(19), S => CTRL, Z => OUT1(19)
                           );
   U25 : MUX2_X1 port map( A => IN0(18), B => IN1(18), S => CTRL, Z => OUT1(18)
                           );
   U26 : MUX2_X1 port map( A => IN0(17), B => IN1(17), S => CTRL, Z => OUT1(17)
                           );
   U28 : MUX2_X1 port map( A => IN0(15), B => IN1(15), S => CTRL, Z => OUT1(15)
                           );
   U30 : MUX2_X1 port map( A => IN0(13), B => IN1(13), S => CTRL, Z => OUT1(13)
                           );
   U31 : MUX2_X1 port map( A => IN0(12), B => IN1(12), S => CTRL, Z => OUT1(12)
                           );
   U32 : MUX2_X1 port map( A => IN0(11), B => IN1(11), S => CTRL, Z => OUT1(11)
                           );
   U33 : MUX2_X1 port map( A => IN0(10), B => IN1(10), S => CTRL, Z => OUT1(10)
                           );
   U2 : INV_X1 port map( A => IN0(0), ZN => n2);
   U1 : NOR2_X1 port map( A1 => n2, A2 => CTRL, ZN => OUT1(0));
   U9 : MUX2_X1 port map( A => IN0(3), B => IN1(3), S => CTRL, Z => OUT1(3));
   U13 : MUX2_X1 port map( A => IN0(14), B => IN1(14), S => CTRL, Z => OUT1(14)
                           );
   U27 : MUX2_X1 port map( A => IN0(16), B => IN1(16), S => CTRL, Z => OUT1(16)
                           );
   U29 : MUX2_X1 port map( A => IN0(29), B => IN1(29), S => CTRL, Z => OUT1(29)
                           );

end SYN_Bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity piso_r_2_N32 is

   port( Clock, ALOAD : in std_logic;  D : in std_logic_vector (31 downto 0);  
         SO : out std_logic_vector (31 downto 0));

end piso_r_2_N32;

architecture SYN_archi of piso_r_2_N32 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component SDFF_X1
      port( D, SI, SE, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal SO_31_port, SO_30_port, SO_29_port, SO_28_port, SO_27_port, 
      SO_26_port, SO_25_port, SO_24_port, SO_23_port, SO_22_port, SO_21_port, 
      SO_20_port, SO_19_port, SO_18_port, SO_17_port, SO_16_port, SO_15_port, 
      SO_14_port, SO_13_port, SO_12_port, SO_11_port, SO_10_port, SO_9_port, 
      SO_8_port, SO_7_port, SO_6_port, SO_5_port, SO_4_port, SO_3_port, 
      SO_2_port, SO_1_port, SO_0_port, N3, N4, N5, N6, N7, N8, N9, N10, N11, 
      N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26
      , N27, N28, N29, N30, N31, N32, net549709, net549724, n2, n7_port, 
      net645047, net645048, net645049, net645050, net645051, net645052, 
      net645053, net645054, net645055, net645056, net645057, net645058, 
      net645059, net645060, net645061, net645062, net645063, net645064, 
      net645065, net645066, net645067, net645068, net645069, net645070, 
      net645071, net645072, net645073, net645074, n1, n3_port, n4_port, n5_port
      , n6_port, n11_port, n12_port, n13_port, n16_port, n19_port, n21_port, 
      n22_port, n23_port, n24_port, n25_port, n26_port, n27_port, n28_port, 
      n29_port, n30_port : std_logic;

begin
   SO <= ( SO_31_port, SO_30_port, SO_29_port, SO_28_port, SO_27_port, 
      SO_26_port, SO_25_port, SO_24_port, SO_23_port, SO_22_port, SO_21_port, 
      SO_20_port, SO_19_port, SO_18_port, SO_17_port, SO_16_port, SO_15_port, 
      SO_14_port, SO_13_port, SO_12_port, SO_11_port, SO_10_port, SO_9_port, 
      SO_8_port, SO_7_port, SO_6_port, SO_5_port, SO_4_port, SO_3_port, 
      SO_2_port, SO_1_port, SO_0_port );
   
   tmp_reg_1_inst : DFF_X1 port map( D => N4, CK => Clock, Q => SO_1_port, QN 
                           => net645074);
   tmp_reg_3_inst : DFF_X1 port map( D => N6, CK => Clock, Q => SO_3_port, QN 
                           => net645073);
   tmp_reg_5_inst : DFF_X1 port map( D => N8, CK => Clock, Q => SO_5_port, QN 
                           => net645072);
   tmp_reg_7_inst : DFF_X1 port map( D => N10, CK => Clock, Q => SO_7_port, QN 
                           => net645071);
   tmp_reg_9_inst : DFF_X1 port map( D => N12, CK => Clock, Q => SO_9_port, QN 
                           => net645070);
   tmp_reg_11_inst : DFF_X1 port map( D => N14, CK => Clock, Q => SO_11_port, 
                           QN => net645069);
   tmp_reg_13_inst : DFF_X1 port map( D => N16, CK => Clock, Q => SO_13_port, 
                           QN => net645068);
   tmp_reg_15_inst : DFF_X1 port map( D => N18, CK => Clock, Q => SO_15_port, 
                           QN => net645067);
   tmp_reg_17_inst : DFF_X1 port map( D => N20, CK => Clock, Q => SO_17_port, 
                           QN => net645066);
   tmp_reg_19_inst : DFF_X1 port map( D => N22, CK => Clock, Q => SO_19_port, 
                           QN => net645065);
   tmp_reg_21_inst : DFF_X1 port map( D => N24, CK => Clock, Q => SO_21_port, 
                           QN => net645064);
   tmp_reg_23_inst : DFF_X1 port map( D => N26, CK => Clock, Q => SO_23_port, 
                           QN => net645063);
   tmp_reg_25_inst : DFF_X1 port map( D => N28, CK => Clock, Q => SO_25_port, 
                           QN => net645062);
   tmp_reg_27_inst : DFF_X1 port map( D => N30, CK => Clock, Q => SO_27_port, 
                           QN => net645061);
   tmp_reg_29_inst : DFF_X1 port map( D => N32, CK => Clock, Q => SO_29_port, 
                           QN => net549724);
   tmp_reg_0_inst : DFF_X1 port map( D => N3, CK => Clock, Q => SO_0_port, QN 
                           => net645060);
   tmp_reg_2_inst : DFF_X1 port map( D => N5, CK => Clock, Q => SO_2_port, QN 
                           => net645059);
   tmp_reg_4_inst : DFF_X1 port map( D => N7, CK => Clock, Q => SO_4_port, QN 
                           => net645058);
   tmp_reg_6_inst : DFF_X1 port map( D => N9, CK => Clock, Q => SO_6_port, QN 
                           => net645057);
   tmp_reg_8_inst : DFF_X1 port map( D => N11, CK => Clock, Q => SO_8_port, QN 
                           => net645056);
   tmp_reg_10_inst : DFF_X1 port map( D => N13, CK => Clock, Q => SO_10_port, 
                           QN => net645055);
   tmp_reg_12_inst : DFF_X1 port map( D => N15, CK => Clock, Q => SO_12_port, 
                           QN => net645054);
   tmp_reg_14_inst : DFF_X1 port map( D => N17, CK => Clock, Q => SO_14_port, 
                           QN => net645053);
   tmp_reg_16_inst : DFF_X1 port map( D => N19, CK => Clock, Q => SO_16_port, 
                           QN => net645052);
   tmp_reg_18_inst : DFF_X1 port map( D => N21, CK => Clock, Q => SO_18_port, 
                           QN => net645051);
   tmp_reg_20_inst : DFF_X1 port map( D => N23, CK => Clock, Q => SO_20_port, 
                           QN => net645050);
   tmp_reg_22_inst : DFF_X1 port map( D => N25, CK => Clock, Q => SO_22_port, 
                           QN => net645049);
   tmp_reg_24_inst : DFF_X1 port map( D => N27, CK => Clock, Q => SO_24_port, 
                           QN => net645048);
   tmp_reg_26_inst : DFF_X1 port map( D => N29, CK => Clock, Q => SO_26_port, 
                           QN => net645047);
   tmp_reg_28_inst : DFF_X1 port map( D => N31, CK => Clock, Q => SO_28_port, 
                           QN => net549709);
   tmp_reg_31_inst : SDFF_X1 port map( D => SO_29_port, SI => D(31), SE => 
                           ALOAD, CK => Clock, Q => SO_31_port, QN => n7_port);
   tmp_reg_30_inst : SDFF_X1 port map( D => SO_28_port, SI => D(30), SE => 
                           ALOAD, CK => Clock, Q => SO_30_port, QN => n2);
   U16 : OAI21_X1 port map( B1 => ALOAD, B2 => net645047, A => n11_port, ZN => 
                           N31);
   U22 : NAND2_X1 port map( A1 => ALOAD, A2 => D(26), ZN => n11_port);
   U21 : OAI21_X1 port map( B1 => ALOAD, B2 => net645048, A => n11_port, ZN => 
                           N29);
   U18 : OAI21_X1 port map( B1 => ALOAD, B2 => net645062, A => n12_port, ZN => 
                           N30);
   U38 : NAND2_X1 port map( A1 => ALOAD, A2 => D(18), ZN => n19_port);
   U37 : OAI21_X1 port map( B1 => ALOAD, B2 => net645052, A => n19_port, ZN => 
                           N21);
   U33 : OAI21_X1 port map( B1 => ALOAD, B2 => net645051, A => n19_port, ZN => 
                           N23);
   U32 : NAND2_X1 port map( A1 => ALOAD, A2 => D(21), ZN => n16_port);
   U31 : OAI21_X1 port map( B1 => ALOAD, B2 => net645065, A => n16_port, ZN => 
                           N24);
   U39 : OAI21_X1 port map( B1 => ALOAD, B2 => net645067, A => n16_port, ZN => 
                           N20);
   U42 : NAND2_X1 port map( A1 => ALOAD, A2 => D(16), ZN => n21_port);
   U41 : OAI21_X1 port map( B1 => ALOAD, B2 => net645053, A => n21_port, ZN => 
                           N19);
   U14 : OAI21_X1 port map( B1 => ALOAD, B2 => net645061, A => n21_port, ZN => 
                           N32);
   U24 : NAND2_X1 port map( A1 => ALOAD, A2 => D(25), ZN => n12_port);
   U23 : OAI21_X1 port map( B1 => ALOAD, B2 => net645063, A => n12_port, ZN => 
                           N28);
   U29 : OAI21_X1 port map( B1 => ALOAD, B2 => net645050, A => n13_port, ZN => 
                           N25);
   U26 : NAND2_X1 port map( A1 => ALOAD, A2 => D(24), ZN => n13_port);
   U25 : OAI21_X1 port map( B1 => ALOAD, B2 => net645049, A => n13_port, ZN => 
                           N27);
   U27 : OAI21_X1 port map( B1 => ALOAD, B2 => net645064, A => n12_port, ZN => 
                           N26);
   U35 : OAI21_X1 port map( B1 => ALOAD, B2 => net645066, A => n21_port, ZN => 
                           N22);
   U44 : NAND2_X1 port map( A1 => ALOAD, A2 => D(15), ZN => n22_port);
   U43 : OAI21_X1 port map( B1 => ALOAD, B2 => net645068, A => n22_port, ZN => 
                           N18);
   U52 : NAND2_X1 port map( A1 => ALOAD, A2 => D(11), ZN => n26_port);
   U51 : OAI21_X1 port map( B1 => ALOAD, B2 => net645070, A => n26_port, ZN => 
                           N14);
   U12 : NAND2_X1 port map( A1 => ALOAD, A2 => D(2), ZN => n6_port);
   U11 : OAI21_X1 port map( B1 => ALOAD, B2 => net645060, A => n6_port, ZN => 
                           N5);
   U54 : NAND2_X1 port map( A1 => ALOAD, A2 => D(10), ZN => n27_port);
   U53 : OAI21_X1 port map( B1 => ALOAD, B2 => net645056, A => n27_port, ZN => 
                           N13);
   U46 : NAND2_X1 port map( A1 => ALOAD, A2 => D(14), ZN => n23_port);
   U45 : OAI21_X1 port map( B1 => ALOAD, B2 => net645054, A => n23_port, ZN => 
                           N17);
   U50 : NAND2_X1 port map( A1 => ALOAD, A2 => D(12), ZN => n25_port);
   U49 : OAI21_X1 port map( B1 => ALOAD, B2 => net645055, A => n25_port, ZN => 
                           N15);
   U48 : NAND2_X1 port map( A1 => ALOAD, A2 => D(13), ZN => n24_port);
   U47 : OAI21_X1 port map( B1 => ALOAD, B2 => net645069, A => n24_port, ZN => 
                           N16);
   U58 : NAND2_X1 port map( A1 => ALOAD, A2 => D(8), ZN => n29_port);
   U57 : OAI21_X1 port map( B1 => ALOAD, B2 => net645057, A => n29_port, ZN => 
                           N11);
   U60 : NAND2_X1 port map( A1 => ALOAD, A2 => D(7), ZN => n30_port);
   U59 : OAI21_X1 port map( B1 => ALOAD, B2 => net645072, A => n30_port, ZN => 
                           N10);
   U56 : NAND2_X1 port map( A1 => ALOAD, A2 => D(9), ZN => n28_port);
   U55 : OAI21_X1 port map( B1 => ALOAD, B2 => net645071, A => n28_port, ZN => 
                           N12);
   U4 : NAND2_X1 port map( A1 => ALOAD, A2 => D(6), ZN => n1);
   U3 : OAI21_X1 port map( B1 => ALOAD, B2 => net645058, A => n1, ZN => N9);
   U8 : NAND2_X1 port map( A1 => ALOAD, A2 => D(4), ZN => n4_port);
   U7 : OAI21_X1 port map( B1 => ALOAD, B2 => net645059, A => n4_port, ZN => N7
                           );
   U10 : NAND2_X1 port map( A1 => ALOAD, A2 => D(3), ZN => n5_port);
   U9 : OAI21_X1 port map( B1 => ALOAD, B2 => net645074, A => n5_port, ZN => N6
                           );
   U6 : NAND2_X1 port map( A1 => ALOAD, A2 => D(5), ZN => n3_port);
   U5 : OAI21_X1 port map( B1 => ALOAD, B2 => net645073, A => n3_port, ZN => N8
                           );
   U13 : AND2_X1 port map( A1 => ALOAD, A2 => D(1), ZN => N4);
   U15 : AND2_X1 port map( A1 => ALOAD, A2 => D(0), ZN => N3);

end SYN_archi;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity shift_N9_1 is

   port( Clock, ALOAD : in std_logic;  D : in std_logic_vector (8 downto 0);  
         SO : out std_logic);

end shift_N9_1;

architecture SYN_archi of shift_N9_1 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component SDFF_X1
      port( D, SI, SE, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal tmp_8_port, tmp_7_port, tmp_6_port, tmp_5_port, tmp_4_port, 
      tmp_3_port, tmp_2_port, tmp_1_port, n13, n14, n15, n16, n17, n18, n19, 
      n20, n21, n22 : std_logic;

begin
   
   tmp_reg_8_inst : DFF_X1 port map( D => n22, CK => Clock, Q => tmp_8_port, QN
                           => n21);
   tmp_reg_0_inst : SDFF_X1 port map( D => tmp_1_port, SI => D(0), SE => ALOAD,
                           CK => Clock, Q => SO, QN => n20);
   tmp_reg_3_inst : SDFF_X1 port map( D => tmp_4_port, SI => D(3), SE => ALOAD,
                           CK => Clock, Q => tmp_3_port, QN => n19);
   tmp_reg_5_inst : SDFF_X1 port map( D => tmp_6_port, SI => D(5), SE => ALOAD,
                           CK => Clock, Q => tmp_5_port, QN => n18);
   tmp_reg_1_inst : SDFF_X1 port map( D => tmp_2_port, SI => D(1), SE => ALOAD,
                           CK => Clock, Q => tmp_1_port, QN => n17);
   tmp_reg_4_inst : SDFF_X1 port map( D => tmp_5_port, SI => D(4), SE => ALOAD,
                           CK => Clock, Q => tmp_4_port, QN => n16);
   tmp_reg_6_inst : SDFF_X1 port map( D => tmp_7_port, SI => D(6), SE => ALOAD,
                           CK => Clock, Q => tmp_6_port, QN => n15);
   tmp_reg_2_inst : SDFF_X1 port map( D => tmp_3_port, SI => D(2), SE => ALOAD,
                           CK => Clock, Q => tmp_2_port, QN => n14);
   tmp_reg_7_inst : SDFF_X1 port map( D => tmp_8_port, SI => D(7), SE => ALOAD,
                           CK => Clock, Q => tmp_7_port, QN => n13);
   U3 : AND2_X1 port map( A1 => ALOAD, A2 => D(8), ZN => n22);

end SYN_archi;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity shift_N9_2 is

   port( Clock, ALOAD : in std_logic;  D : in std_logic_vector (8 downto 0);  
         SO : out std_logic);

end shift_N9_2;

architecture SYN_archi of shift_N9_2 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component SDFF_X1
      port( D, SI, SE, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal tmp_8_port, tmp_7_port, tmp_6_port, tmp_5_port, tmp_4_port, 
      tmp_3_port, tmp_2_port, tmp_1_port, n13, n14, n15, n16, n17, n18, n19, 
      n20, n21, n22 : std_logic;

begin
   
   tmp_reg_8_inst : DFF_X1 port map( D => n22, CK => Clock, Q => tmp_8_port, QN
                           => n21);
   tmp_reg_0_inst : SDFF_X1 port map( D => tmp_1_port, SI => D(0), SE => ALOAD,
                           CK => Clock, Q => SO, QN => n20);
   tmp_reg_2_inst : SDFF_X1 port map( D => tmp_3_port, SI => D(2), SE => ALOAD,
                           CK => Clock, Q => tmp_2_port, QN => n19);
   tmp_reg_4_inst : SDFF_X1 port map( D => tmp_5_port, SI => D(4), SE => ALOAD,
                           CK => Clock, Q => tmp_4_port, QN => n18);
   tmp_reg_3_inst : SDFF_X1 port map( D => tmp_4_port, SI => D(3), SE => ALOAD,
                           CK => Clock, Q => tmp_3_port, QN => n17);
   tmp_reg_5_inst : SDFF_X1 port map( D => tmp_6_port, SI => D(5), SE => ALOAD,
                           CK => Clock, Q => tmp_5_port, QN => n16);
   tmp_reg_7_inst : SDFF_X1 port map( D => tmp_8_port, SI => D(7), SE => ALOAD,
                           CK => Clock, Q => tmp_7_port, QN => n15);
   tmp_reg_1_inst : SDFF_X1 port map( D => tmp_2_port, SI => D(1), SE => ALOAD,
                           CK => Clock, Q => tmp_1_port, QN => n14);
   tmp_reg_6_inst : SDFF_X1 port map( D => tmp_7_port, SI => D(6), SE => ALOAD,
                           CK => Clock, Q => tmp_6_port, QN => n13);
   U3 : AND2_X1 port map( A1 => ALOAD, A2 => D(8), ZN => n22);

end SYN_archi;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity shift_N9_0 is

   port( Clock, ALOAD : in std_logic;  D : in std_logic_vector (8 downto 0);  
         SO : out std_logic);

end shift_N9_0;

architecture SYN_archi of shift_N9_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component SDFF_X2
      port( D, SI, SE, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component SDFF_X1
      port( D, SI, SE, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal tmp_8_port, tmp_7_port, tmp_6_port, tmp_5_port, tmp_4_port, 
      tmp_3_port, tmp_2_port, tmp_1_port, n13, n14, n15, n16, n17, n18, n19, 
      n20, n21, n22 : std_logic;

begin
   
   tmp_reg_8_inst : DFF_X1 port map( D => n22, CK => Clock, Q => tmp_8_port, QN
                           => n21);
   tmp_reg_3_inst : SDFF_X1 port map( D => tmp_4_port, SI => D(3), SE => ALOAD,
                           CK => Clock, Q => tmp_3_port, QN => n20);
   tmp_reg_5_inst : SDFF_X1 port map( D => tmp_6_port, SI => D(5), SE => ALOAD,
                           CK => Clock, Q => tmp_5_port, QN => n19);
   tmp_reg_4_inst : SDFF_X1 port map( D => tmp_5_port, SI => D(4), SE => ALOAD,
                           CK => Clock, Q => tmp_4_port, QN => n18);
   tmp_reg_1_inst : SDFF_X1 port map( D => tmp_2_port, SI => D(1), SE => ALOAD,
                           CK => Clock, Q => tmp_1_port, QN => n17);
   tmp_reg_2_inst : SDFF_X1 port map( D => tmp_3_port, SI => D(2), SE => ALOAD,
                           CK => Clock, Q => tmp_2_port, QN => n16);
   tmp_reg_7_inst : SDFF_X1 port map( D => tmp_8_port, SI => D(7), SE => ALOAD,
                           CK => Clock, Q => tmp_7_port, QN => n15);
   tmp_reg_6_inst : SDFF_X1 port map( D => tmp_7_port, SI => D(6), SE => ALOAD,
                           CK => Clock, Q => tmp_6_port, QN => n14);
   tmp_reg_0_inst : SDFF_X2 port map( D => tmp_1_port, SI => D(0), SE => ALOAD,
                           CK => Clock, Q => SO, QN => n13);
   U3 : AND2_X1 port map( A1 => ALOAD, A2 => D(8), ZN => n22);

end SYN_archi;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity booth_encoder_1 is

   port( B_in : in std_logic_vector (2 downto 0);  A_out : out std_logic_vector
         (2 downto 0));

end booth_encoder_1;

architecture SYN_bhe of booth_encoder_1 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5 : std_logic;

begin
   
   U7 : NAND2_X1 port map( A1 => B_in(1), A2 => n3, ZN => n5);
   U3 : OAI221_X1 port map( B1 => B_in(0), B2 => n3, C1 => n4, C2 => B_in(1), A
                           => n5, ZN => A_out(2));
   U5 : NOR2_X1 port map( A1 => n5, A2 => n4, ZN => A_out(0));
   U8 : INV_X1 port map( A => B_in(2), ZN => n3);
   U4 : AND2_X1 port map( A1 => n4, A2 => B_in(1), ZN => A_out(1));
   U6 : INV_X1 port map( A => B_in(0), ZN => n4);

end SYN_bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity booth_encoder_6 is

   port( B_in : in std_logic_vector (2 downto 0);  A_out : out std_logic_vector
         (2 downto 0));

end booth_encoder_6;

architecture SYN_bhe of booth_encoder_6 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI33_X1
      port( A1, A2, A3, B1, B2, B3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U9 : OAI33_X1 port map( A1 => B_in(0), A2 => B_in(1), A3 => n7, B1 => n4, B2
                           => n5, B3 => B_in(2), ZN => A_out(0));
   U3 : INV_X1 port map( A => B_in(1), ZN => n5);
   U4 : INV_X1 port map( A => B_in(0), ZN => n4);
   U5 : INV_X1 port map( A => B_in(2), ZN => n7);
   U6 : NAND2_X1 port map( A1 => B_in(2), A2 => n4, ZN => n6);
   U7 : OAI221_X1 port map( B1 => B_in(1), B2 => n4, C1 => n5, C2 => B_in(2), A
                           => n6, ZN => A_out(2));
   U8 : AOI21_X1 port map( B1 => B_in(0), B2 => B_in(1), A => n7, ZN => 
                           A_out(1));

end SYN_bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity booth_encoder_7 is

   port( B_in : in std_logic_vector (2 downto 0);  A_out : out std_logic_vector
         (2 downto 0));

end booth_encoder_7;

architecture SYN_bhe of booth_encoder_7 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI33_X1
      port( A1, A2, A3, B1, B2, B3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U9 : OAI33_X1 port map( A1 => B_in(0), A2 => B_in(1), A3 => n7, B1 => n4, B2
                           => n5, B3 => B_in(2), ZN => A_out(0));
   U3 : INV_X1 port map( A => B_in(1), ZN => n5);
   U4 : INV_X1 port map( A => B_in(0), ZN => n4);
   U5 : INV_X1 port map( A => B_in(2), ZN => n7);
   U6 : AOI21_X1 port map( B1 => B_in(0), B2 => B_in(1), A => n7, ZN => 
                           A_out(1));
   U7 : OAI221_X1 port map( B1 => B_in(1), B2 => n4, C1 => n5, C2 => B_in(2), A
                           => n6, ZN => A_out(2));
   U8 : NAND2_X1 port map( A1 => B_in(2), A2 => n4, ZN => n6);

end SYN_bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity booth_encoder_8 is

   port( B_in : in std_logic_vector (2 downto 0);  A_out : out std_logic_vector
         (2 downto 0));

end booth_encoder_8;

architecture SYN_bhe of booth_encoder_8 is

   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI33_X1
      port( A1, A2, A3, B1, B2, B3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U9 : OAI33_X1 port map( A1 => B_in(0), A2 => B_in(1), A3 => n7, B1 => n4, B2
                           => n5, B3 => B_in(2), ZN => A_out(0));
   U3 : INV_X1 port map( A => B_in(2), ZN => n7);
   U4 : INV_X1 port map( A => B_in(1), ZN => n5);
   U5 : INV_X1 port map( A => B_in(0), ZN => n4);
   U6 : AOI21_X1 port map( B1 => B_in(0), B2 => B_in(1), A => n7, ZN => 
                           A_out(1));
   U7 : NAND2_X1 port map( A1 => B_in(2), A2 => n4, ZN => n6);
   U8 : OAI221_X1 port map( B1 => B_in(1), B2 => n4, C1 => n5, C2 => B_in(2), A
                           => n6, ZN => A_out(2));

end SYN_bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity booth_encoder_0 is

   port( B_in : in std_logic_vector (2 downto 0);  A_out : out std_logic_vector
         (2 downto 0));

end booth_encoder_0;

architecture SYN_bhe of booth_encoder_0 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal N53, N57, n2 : std_logic;

begin
   A_out <= ( N57, B_in(2), N53 );
   
   U3 : INV_X1 port map( A => B_in(2), ZN => n2);
   U4 : OR2_X1 port map( A1 => B_in(1), A2 => B_in(2), ZN => N57);
   U5 : NOR2_X1 port map( A1 => B_in(1), A2 => n2, ZN => N53);

end SYN_bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity carry_sel_gen_N4_11 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end carry_sel_gen_N4_11;

architecture SYN_STRUCTURAL of carry_sel_gen_N4_11 is

   component mux21_SIZE4_11
      port( IN0, IN1 : in std_logic_vector (3 downto 0);  CTRL : in std_logic; 
            OUT1 : out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_N4_22
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_23
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, nocarry_sum_to_mux_3_port, 
      nocarry_sum_to_mux_2_port, nocarry_sum_to_mux_1_port, 
      nocarry_sum_to_mux_0_port, carry_sum_to_mux_3_port, 
      carry_sum_to_mux_2_port, carry_sum_to_mux_1_port, carry_sum_to_mux_0_port
      , net684325, net684326 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   rca_nocarry : RCA_N4_23 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           nocarry_sum_to_mux_3_port, S(2) => 
                           nocarry_sum_to_mux_2_port, S(1) => 
                           nocarry_sum_to_mux_1_port, S(0) => 
                           nocarry_sum_to_mux_0_port, Co => net684326);
   rca_carry : RCA_N4_22 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           carry_sum_to_mux_3_port, S(2) => 
                           carry_sum_to_mux_2_port, S(1) => 
                           carry_sum_to_mux_1_port, S(0) => 
                           carry_sum_to_mux_0_port, Co => net684325);
   outmux : mux21_SIZE4_11 port map( IN0(3) => nocarry_sum_to_mux_3_port, 
                           IN0(2) => nocarry_sum_to_mux_2_port, IN0(1) => 
                           nocarry_sum_to_mux_1_port, IN0(0) => 
                           nocarry_sum_to_mux_0_port, IN1(3) => 
                           carry_sum_to_mux_3_port, IN1(2) => 
                           carry_sum_to_mux_2_port, IN1(1) => 
                           carry_sum_to_mux_1_port, IN1(0) => 
                           carry_sum_to_mux_0_port, CTRL => Ci, OUT1(3) => S(3)
                           , OUT1(2) => S(2), OUT1(1) => S(1), OUT1(0) => S(0))
                           ;

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity carry_sel_gen_N4_12 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end carry_sel_gen_N4_12;

architecture SYN_STRUCTURAL of carry_sel_gen_N4_12 is

   component mux21_SIZE4_12
      port( IN0, IN1 : in std_logic_vector (3 downto 0);  CTRL : in std_logic; 
            OUT1 : out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_N4_24
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_25
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, nocarry_sum_to_mux_3_port, 
      nocarry_sum_to_mux_2_port, nocarry_sum_to_mux_1_port, 
      nocarry_sum_to_mux_0_port, carry_sum_to_mux_3_port, 
      carry_sum_to_mux_2_port, carry_sum_to_mux_1_port, carry_sum_to_mux_0_port
      , net684323, net684324 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   rca_nocarry : RCA_N4_25 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           nocarry_sum_to_mux_3_port, S(2) => 
                           nocarry_sum_to_mux_2_port, S(1) => 
                           nocarry_sum_to_mux_1_port, S(0) => 
                           nocarry_sum_to_mux_0_port, Co => net684324);
   rca_carry : RCA_N4_24 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           carry_sum_to_mux_3_port, S(2) => 
                           carry_sum_to_mux_2_port, S(1) => 
                           carry_sum_to_mux_1_port, S(0) => 
                           carry_sum_to_mux_0_port, Co => net684323);
   outmux : mux21_SIZE4_12 port map( IN0(3) => nocarry_sum_to_mux_3_port, 
                           IN0(2) => nocarry_sum_to_mux_2_port, IN0(1) => 
                           nocarry_sum_to_mux_1_port, IN0(0) => 
                           nocarry_sum_to_mux_0_port, IN1(3) => 
                           carry_sum_to_mux_3_port, IN1(2) => 
                           carry_sum_to_mux_2_port, IN1(1) => 
                           carry_sum_to_mux_1_port, IN1(0) => 
                           carry_sum_to_mux_0_port, CTRL => Ci, OUT1(3) => S(3)
                           , OUT1(2) => S(2), OUT1(1) => S(1), OUT1(0) => S(0))
                           ;

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity carry_sel_gen_N4_13 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end carry_sel_gen_N4_13;

architecture SYN_STRUCTURAL of carry_sel_gen_N4_13 is

   component mux21_SIZE4_13
      port( IN0, IN1 : in std_logic_vector (3 downto 0);  CTRL : in std_logic; 
            OUT1 : out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_N4_26
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_27
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, nocarry_sum_to_mux_3_port, 
      nocarry_sum_to_mux_2_port, nocarry_sum_to_mux_1_port, 
      nocarry_sum_to_mux_0_port, carry_sum_to_mux_3_port, 
      carry_sum_to_mux_2_port, carry_sum_to_mux_1_port, carry_sum_to_mux_0_port
      , net684321, net684322 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   rca_nocarry : RCA_N4_27 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           nocarry_sum_to_mux_3_port, S(2) => 
                           nocarry_sum_to_mux_2_port, S(1) => 
                           nocarry_sum_to_mux_1_port, S(0) => 
                           nocarry_sum_to_mux_0_port, Co => net684322);
   rca_carry : RCA_N4_26 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           carry_sum_to_mux_3_port, S(2) => 
                           carry_sum_to_mux_2_port, S(1) => 
                           carry_sum_to_mux_1_port, S(0) => 
                           carry_sum_to_mux_0_port, Co => net684321);
   outmux : mux21_SIZE4_13 port map( IN0(3) => nocarry_sum_to_mux_3_port, 
                           IN0(2) => nocarry_sum_to_mux_2_port, IN0(1) => 
                           nocarry_sum_to_mux_1_port, IN0(0) => 
                           nocarry_sum_to_mux_0_port, IN1(3) => 
                           carry_sum_to_mux_3_port, IN1(2) => 
                           carry_sum_to_mux_2_port, IN1(1) => 
                           carry_sum_to_mux_1_port, IN1(0) => 
                           carry_sum_to_mux_0_port, CTRL => Ci, OUT1(3) => S(3)
                           , OUT1(2) => S(2), OUT1(1) => S(1), OUT1(0) => S(0))
                           ;

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity carry_sel_gen_N4_14 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end carry_sel_gen_N4_14;

architecture SYN_STRUCTURAL of carry_sel_gen_N4_14 is

   component mux21_SIZE4_14
      port( IN0, IN1 : in std_logic_vector (3 downto 0);  CTRL : in std_logic; 
            OUT1 : out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_N4_28
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_29
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, nocarry_sum_to_mux_3_port, 
      nocarry_sum_to_mux_2_port, nocarry_sum_to_mux_1_port, 
      nocarry_sum_to_mux_0_port, carry_sum_to_mux_3_port, 
      carry_sum_to_mux_2_port, carry_sum_to_mux_1_port, carry_sum_to_mux_0_port
      , net684319, net684320 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   rca_nocarry : RCA_N4_29 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           nocarry_sum_to_mux_3_port, S(2) => 
                           nocarry_sum_to_mux_2_port, S(1) => 
                           nocarry_sum_to_mux_1_port, S(0) => 
                           nocarry_sum_to_mux_0_port, Co => net684320);
   rca_carry : RCA_N4_28 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           carry_sum_to_mux_3_port, S(2) => 
                           carry_sum_to_mux_2_port, S(1) => 
                           carry_sum_to_mux_1_port, S(0) => 
                           carry_sum_to_mux_0_port, Co => net684319);
   outmux : mux21_SIZE4_14 port map( IN0(3) => nocarry_sum_to_mux_3_port, 
                           IN0(2) => nocarry_sum_to_mux_2_port, IN0(1) => 
                           nocarry_sum_to_mux_1_port, IN0(0) => 
                           nocarry_sum_to_mux_0_port, IN1(3) => 
                           carry_sum_to_mux_3_port, IN1(2) => 
                           carry_sum_to_mux_2_port, IN1(1) => 
                           carry_sum_to_mux_1_port, IN1(0) => 
                           carry_sum_to_mux_0_port, CTRL => Ci, OUT1(3) => S(3)
                           , OUT1(2) => S(2), OUT1(1) => S(1), OUT1(0) => S(0))
                           ;

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity carry_sel_gen_N4_0_0 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end carry_sel_gen_N4_0_0;

architecture SYN_STRUCTURAL of carry_sel_gen_N4_0_0 is

   component mux21_SIZE4_0_0
      port( IN0, IN1 : in std_logic_vector (3 downto 0);  CTRL : in std_logic; 
            OUT1 : out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_N4_0_0
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic0_port, n5, nocarry_sum_to_mux_3_port, 
      nocarry_sum_to_mux_2_port, nocarry_sum_to_mux_1_port, 
      nocarry_sum_to_mux_0_port, n1, n2, n3, n4, net684318 : std_logic;

begin
   
   X_Logic0_port <= '0';
   rca_nocarry : RCA_N4_0_0 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1),
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           nocarry_sum_to_mux_3_port, S(2) => 
                           nocarry_sum_to_mux_2_port, S(1) => 
                           nocarry_sum_to_mux_1_port, S(0) => 
                           nocarry_sum_to_mux_0_port, Co => net684318);
   outmux : mux21_SIZE4_0_0 port map( IN0(3) => nocarry_sum_to_mux_3_port, 
                           IN0(2) => nocarry_sum_to_mux_2_port, IN0(1) => 
                           nocarry_sum_to_mux_1_port, IN0(0) => 
                           nocarry_sum_to_mux_0_port, IN1(3) => n1, IN1(2) => 
                           n2, IN1(1) => n3, IN1(0) => n4, CTRL => n5, OUT1(3) 
                           => S(3), OUT1(2) => S(2), OUT1(1) => S(1), OUT1(0) 
                           => S(0));
   n1 <= '0';
   n2 <= '0';
   n3 <= '0';
   n4 <= '0';
   n5 <= '0';

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_37 is

   port( p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic;  
         g_BAR : in std_logic);

end pg_37;

architecture SYN_beh of pg_37 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U3 : NAND2_X1 port map( A1 => p, A2 => g_prec, ZN => n1);
   U2 : NAND2_X1 port map( A1 => g_BAR, A2 => n1, ZN => g_out);
   U1 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_38 is

   port( p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic;  
         g_BAR : in std_logic);

end pg_38;

architecture SYN_beh of pg_38 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U3 : NAND2_X1 port map( A1 => p, A2 => g_prec, ZN => n1);
   U2 : NAND2_X1 port map( A1 => g_BAR, A2 => n1, ZN => g_out);
   U1 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity g_17 is

   port( g, p, g_prec : in std_logic;  g_out : out std_logic);

end g_17;

architecture SYN_beh of g_17 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U2 : AOI21_X1 port map( B1 => p, B2 => g_prec, A => g, ZN => n2);
   U1 : INV_X1 port map( A => n2, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_46 is

   port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic);

end pg_46;

architecture SYN_beh of pg_46 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n6, n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => g, ZN => n7);
   U2 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);
   U3 : NAND2_X1 port map( A1 => p, A2 => g_prec, ZN => n6);
   U4 : NAND2_X1 port map( A1 => n6, A2 => n7, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_51 is

   port( g, p, g_prec, p_prec : in std_logic;  p_out, g_out_BAR : out std_logic
         );

end pg_51;

architecture SYN_beh of pg_51 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U2 : AOI21_X1 port map( B1 => g_prec, B2 => p, A => g, ZN => g_out_BAR);
   U1 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_52 is

   port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic);

end pg_52;

architecture SYN_beh of pg_52 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U3 : AOI21_X1 port map( B1 => g_prec, B2 => p, A => g, ZN => n2);
   U1 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);
   U2 : INV_X1 port map( A => n2, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_0_0 is

   port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic);

end pg_0_0;

architecture SYN_beh of pg_0_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U3 : AOI21_X1 port map( B1 => g_prec, B2 => p, A => g, ZN => n2);
   U1 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);
   U2 : INV_X1 port map( A => n2, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity g_18 is

   port( g, p, g_prec : in std_logic;  g_out : out std_logic);

end g_18;

architecture SYN_beh of g_18 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U2 : AOI21_X1 port map( B1 => p, B2 => g_prec, A => g, ZN => n2);
   U1 : INV_X1 port map( A => n2, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity g_0_0 is

   port( g, p, g_prec : in std_logic;  g_out : out std_logic);

end g_0_0;

architecture SYN_beh of g_0_0 is

begin
   g_out <= g;

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_49 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_49;

architecture SYN_beh of pg_net_49 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_62 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_62;

architecture SYN_beh of pg_net_62 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_0_0 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_0_0;

architecture SYN_beh of pg_net_0_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity logic_unit_SIZE32 is

   port( IN1, IN2 : in std_logic_vector (31 downto 0);  CTRL : in 
         std_logic_vector (1 downto 0);  OUT1 : out std_logic_vector (31 downto
         0));

end logic_unit_SIZE32;

architecture SYN_Bhe of logic_unit_SIZE32 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n22, n23, n24, n25, n28, n29, n30, n31, n32, n33, n34, 
      n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49
      , n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, 
      n64, n65, n268, n269, n270, n271, n272, n273 : std_logic;

begin
   
   U98 : XOR2_X1 port map( A => n273, B => CTRL(0), Z => n3);
   U95 : OAI21_X1 port map( B1 => n273, B2 => n64, A => n65, ZN => OUT1(0));
   U28 : NAND2_X1 port map( A1 => IN2(30), A2 => IN1(30), ZN => n18);
   U27 : OAI211_X1 port map( C1 => IN2(30), C2 => IN1(30), A => n272, B => n18,
                           ZN => n19);
   U26 : OAI21_X1 port map( B1 => CTRL(1), B2 => n18, A => n19, ZN => OUT1(30))
                           ;
   U52 : NAND2_X1 port map( A1 => IN2(23), A2 => IN1(23), ZN => n34);
   U51 : OAI211_X1 port map( C1 => IN2(23), C2 => IN1(23), A => n272, B => n34,
                           ZN => n35);
   U50 : OAI21_X1 port map( B1 => CTRL(1), B2 => n34, A => n35, ZN => OUT1(23))
                           ;
   U43 : NAND2_X1 port map( A1 => IN2(26), A2 => IN1(26), ZN => n28);
   U42 : OAI211_X1 port map( C1 => IN2(26), C2 => IN1(26), A => n272, B => n28,
                           ZN => n29);
   U41 : OAI21_X1 port map( B1 => CTRL(1), B2 => n28, A => n29, ZN => OUT1(26))
                           ;
   U55 : NAND2_X1 port map( A1 => IN2(22), A2 => IN1(22), ZN => n36);
   U54 : OAI211_X1 port map( C1 => IN2(22), C2 => IN1(22), A => n272, B => n36,
                           ZN => n37);
   U53 : OAI21_X1 port map( B1 => CTRL(1), B2 => n36, A => n37, ZN => OUT1(22))
                           ;
   U34 : NAND2_X1 port map( A1 => IN2(29), A2 => IN1(29), ZN => n22);
   U33 : OAI211_X1 port map( C1 => IN2(29), C2 => IN1(29), A => n272, B => n22,
                           ZN => n23);
   U32 : OAI21_X1 port map( B1 => n273, B2 => n22, A => n23, ZN => OUT1(29));
   U37 : NAND2_X1 port map( A1 => IN2(28), A2 => IN1(28), ZN => n24);
   U36 : OAI211_X1 port map( C1 => IN2(28), C2 => IN1(28), A => n272, B => n24,
                           ZN => n25);
   U35 : OAI21_X1 port map( B1 => n273, B2 => n24, A => n25, ZN => OUT1(28));
   U46 : NAND2_X1 port map( A1 => IN2(25), A2 => IN1(25), ZN => n30);
   U45 : OAI211_X1 port map( C1 => IN2(25), C2 => IN1(25), A => n272, B => n30,
                           ZN => n31);
   U44 : OAI21_X1 port map( B1 => CTRL(1), B2 => n30, A => n31, ZN => OUT1(25))
                           ;
   U58 : NAND2_X1 port map( A1 => IN2(21), A2 => IN1(21), ZN => n38);
   U57 : OAI211_X1 port map( C1 => IN2(21), C2 => IN1(21), A => n272, B => n38,
                           ZN => n39);
   U56 : OAI21_X1 port map( B1 => n273, B2 => n38, A => n39, ZN => OUT1(21));
   U61 : NAND2_X1 port map( A1 => IN2(20), A2 => IN1(20), ZN => n40);
   U60 : OAI211_X1 port map( C1 => IN2(20), C2 => IN1(20), A => n272, B => n40,
                           ZN => n41);
   U59 : OAI21_X1 port map( B1 => n273, B2 => n40, A => n41, ZN => OUT1(20));
   U49 : NAND2_X1 port map( A1 => IN2(24), A2 => IN1(24), ZN => n32);
   U48 : OAI211_X1 port map( C1 => IN2(24), C2 => IN1(24), A => n272, B => n32,
                           ZN => n33);
   U47 : OAI21_X1 port map( B1 => n273, B2 => n32, A => n33, ZN => OUT1(24));
   U25 : NAND2_X1 port map( A1 => IN2(31), A2 => IN1(31), ZN => n16);
   U24 : OAI211_X1 port map( C1 => IN2(31), C2 => IN1(31), A => n272, B => n16,
                           ZN => n17);
   U23 : OAI21_X1 port map( B1 => n273, B2 => n16, A => n17, ZN => OUT1(31));
   U67 : NAND2_X1 port map( A1 => IN2(19), A2 => IN1(19), ZN => n44);
   U66 : OAI211_X1 port map( C1 => IN2(19), C2 => IN1(19), A => n272, B => n44,
                           ZN => n45);
   U65 : OAI21_X1 port map( B1 => n273, B2 => n44, A => n45, ZN => OUT1(19));
   U83 : OAI21_X1 port map( B1 => CTRL(1), B2 => n56, A => n57, ZN => OUT1(13))
                           ;
   U80 : OAI21_X1 port map( B1 => CTRL(1), B2 => n54, A => n55, ZN => OUT1(14))
                           ;
   U86 : OAI21_X1 port map( B1 => CTRL(1), B2 => n58, A => n59, ZN => OUT1(12))
                           ;
   U91 : NAND2_X1 port map( A1 => IN2(11), A2 => IN1(11), ZN => n60);
   U90 : OAI211_X1 port map( C1 => IN2(11), C2 => IN1(11), A => n272, B => n60,
                           ZN => n61);
   U89 : OAI21_X1 port map( B1 => n273, B2 => n60, A => n61, ZN => OUT1(11));
   U79 : NAND2_X1 port map( A1 => IN2(15), A2 => IN1(15), ZN => n52);
   U78 : OAI211_X1 port map( C1 => IN2(15), C2 => IN1(15), A => n272, B => n52,
                           ZN => n53);
   U77 : OAI21_X1 port map( B1 => CTRL(1), B2 => n52, A => n53, ZN => OUT1(15))
                           ;
   U8 : OAI21_X1 port map( B1 => n273, B2 => n6, A => n7, ZN => OUT1(7));
   U71 : OAI21_X1 port map( B1 => CTRL(1), B2 => n48, A => n49, ZN => OUT1(17))
                           ;
   U92 : OAI21_X1 port map( B1 => CTRL(1), B2 => n62, A => n63, ZN => OUT1(10))
                           ;
   U2 : OAI21_X1 port map( B1 => n273, B2 => n1, A => n2, ZN => OUT1(9));
   U20 : OAI21_X1 port map( B1 => n273, B2 => n14, A => n15, ZN => OUT1(3));
   U62 : OAI21_X1 port map( B1 => CTRL(1), B2 => n42, A => n43, ZN => OUT1(1));
   U7 : NAND2_X1 port map( A1 => IN2(8), A2 => IN1(8), ZN => n4);
   U6 : OAI211_X1 port map( C1 => IN2(8), C2 => IN1(8), A => n3, B => n4, ZN =>
                           n5);
   U5 : OAI21_X1 port map( B1 => n273, B2 => n4, A => n5, ZN => OUT1(8));
   U70 : NAND2_X1 port map( A1 => IN2(18), A2 => IN1(18), ZN => n46);
   U69 : OAI211_X1 port map( C1 => IN2(18), C2 => IN1(18), A => n272, B => n46,
                           ZN => n47);
   U68 : OAI21_X1 port map( B1 => n273, B2 => n46, A => n47, ZN => OUT1(18));
   U76 : NAND2_X1 port map( A1 => IN2(16), A2 => IN1(16), ZN => n50);
   U75 : OAI211_X1 port map( C1 => IN2(16), C2 => IN1(16), A => n272, B => n50,
                           ZN => n51);
   U74 : OAI21_X1 port map( B1 => CTRL(1), B2 => n50, A => n51, ZN => OUT1(16))
                           ;
   U14 : OAI21_X1 port map( B1 => n273, B2 => n10, A => n11, ZN => OUT1(5));
   U17 : OAI21_X1 port map( B1 => n273, B2 => n12, A => n13, ZN => OUT1(4));
   U11 : OAI21_X1 port map( B1 => n273, B2 => n8, A => n9, ZN => OUT1(6));
   U3 : NAND2_X1 port map( A1 => IN2(2), A2 => IN1(2), ZN => n268);
   U4 : OAI211_X1 port map( C1 => IN2(2), C2 => IN1(2), A => n272, B => n268, 
                           ZN => n269);
   U9 : OAI21_X1 port map( B1 => CTRL(1), B2 => n268, A => n269, ZN => OUT1(2))
                           ;
   U10 : NAND2_X1 port map( A1 => IN2(27), A2 => IN1(27), ZN => n270);
   U12 : OAI211_X1 port map( C1 => IN2(27), C2 => IN1(27), A => n272, B => n270
                           , ZN => n271);
   U13 : OAI21_X1 port map( B1 => CTRL(1), B2 => n270, A => n271, ZN => 
                           OUT1(27));
   U15 : BUF_X2 port map( A => n3, Z => n272);
   U16 : BUF_X1 port map( A => CTRL(1), Z => n273);
   U18 : OAI211_X1 port map( C1 => IN2(10), C2 => IN1(10), A => n272, B => n62,
                           ZN => n63);
   U19 : NAND2_X1 port map( A1 => IN2(10), A2 => IN1(10), ZN => n62);
   U21 : OAI211_X1 port map( C1 => IN2(12), C2 => IN1(12), A => n272, B => n58,
                           ZN => n59);
   U22 : NAND2_X1 port map( A1 => IN2(12), A2 => IN1(12), ZN => n58);
   U29 : OAI211_X1 port map( C1 => IN2(4), C2 => IN1(4), A => n272, B => n12, 
                           ZN => n13);
   U30 : NAND2_X1 port map( A1 => IN2(4), A2 => IN1(4), ZN => n12);
   U31 : OAI211_X1 port map( C1 => IN2(17), C2 => IN1(17), A => n272, B => n48,
                           ZN => n49);
   U38 : NAND2_X1 port map( A1 => IN2(17), A2 => IN1(17), ZN => n48);
   U39 : OAI211_X1 port map( C1 => IN2(1), C2 => IN1(1), A => n272, B => n42, 
                           ZN => n43);
   U40 : NAND2_X1 port map( A1 => IN2(1), A2 => IN1(1), ZN => n42);
   U63 : OAI211_X1 port map( C1 => IN2(13), C2 => IN1(13), A => n272, B => n56,
                           ZN => n57);
   U64 : NAND2_X1 port map( A1 => IN2(13), A2 => IN1(13), ZN => n56);
   U72 : OAI211_X1 port map( C1 => IN2(7), C2 => IN1(7), A => n272, B => n6, ZN
                           => n7);
   U73 : NAND2_X1 port map( A1 => IN2(7), A2 => IN1(7), ZN => n6);
   U81 : OAI211_X1 port map( C1 => IN2(3), C2 => IN1(3), A => n272, B => n14, 
                           ZN => n15);
   U82 : NAND2_X1 port map( A1 => IN2(3), A2 => IN1(3), ZN => n14);
   U84 : OAI211_X1 port map( C1 => IN2(14), C2 => IN1(14), A => n272, B => n54,
                           ZN => n55);
   U85 : NAND2_X1 port map( A1 => IN2(14), A2 => IN1(14), ZN => n54);
   U87 : OAI211_X1 port map( C1 => IN2(6), C2 => IN1(6), A => n3, B => n8, ZN 
                           => n9);
   U88 : NAND2_X1 port map( A1 => IN2(6), A2 => IN1(6), ZN => n8);
   U93 : OAI211_X1 port map( C1 => IN2(0), C2 => IN1(0), A => n272, B => n64, 
                           ZN => n65);
   U94 : NAND2_X1 port map( A1 => IN2(0), A2 => IN1(0), ZN => n64);
   U96 : OAI211_X1 port map( C1 => IN2(9), C2 => IN1(9), A => n272, B => n1, ZN
                           => n2);
   U97 : NAND2_X1 port map( A1 => IN2(9), A2 => IN1(9), ZN => n1);
   U99 : OAI211_X1 port map( C1 => IN2(5), C2 => IN1(5), A => n3, B => n10, ZN 
                           => n11);
   U100 : NAND2_X1 port map( A1 => IN2(5), A2 => IN1(5), ZN => n10);

end SYN_Bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity shifter is

   port( A : in std_logic_vector (31 downto 0);  B : in std_logic_vector (4 
         downto 0);  LOGIC_ARITH, LEFT_RIGHT : in std_logic;  OUTPUT : out 
         std_logic_vector (31 downto 0));

end shifter;

architecture SYN_struct of shifter is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component shift_thirdLevel
      port( sel : in std_logic_vector (2 downto 0);  A : in std_logic_vector 
            (38 downto 0);  Y : out std_logic_vector (31 downto 0));
   end component;
   
   component shift_secondLevel
      port( sel : in std_logic_vector (1 downto 0);  mask00, mask08, mask16 : 
            in std_logic_vector (38 downto 0);  Y : out std_logic_vector (38 
            downto 0));
   end component;
   
   component shift_firstLevel
      port( A : in std_logic_vector (31 downto 0);  sel : in std_logic_vector 
            (1 downto 0);  mask00, mask08, mask16 : out std_logic_vector (38 
            downto 0));
   end component;
   
   signal s3_2_port, s3_1_port, s3_0_port, m0_38_port, m0_37_port, m0_36_port, 
      m0_35_port, m0_34_port, m0_33_port, m0_32_port, m0_31_port, m0_30_port, 
      m0_29_port, m0_28_port, m0_27_port, m0_26_port, m0_25_port, m0_24_port, 
      m0_23_port, m0_22_port, m0_21_port, m0_20_port, m0_19_port, m0_18_port, 
      m0_17_port, m0_16_port, m0_15_port, m0_14_port, m0_13_port, m0_12_port, 
      m0_11_port, m0_10_port, m0_9_port, m0_8_port, m0_7_port, m0_6_port, 
      m0_5_port, m0_4_port, m0_3_port, m0_2_port, m0_1_port, m0_0_port, 
      m8_38_port, m8_37_port, m8_36_port, m8_35_port, m8_34_port, m8_33_port, 
      m8_32_port, m8_31_port, m8_30_port, m8_29_port, m8_28_port, m8_27_port, 
      m8_26_port, m8_25_port, m8_24_port, m8_23_port, m8_22_port, m8_21_port, 
      m8_20_port, m8_19_port, m8_18_port, m8_17_port, m8_16_port, m8_15_port, 
      m8_14_port, m8_13_port, m8_12_port, m8_11_port, m8_10_port, m8_9_port, 
      m8_8_port, m8_7_port, m8_6_port, m8_5_port, m8_4_port, m8_3_port, 
      m8_2_port, m8_1_port, m8_0_port, m16_38_port, m16_37_port, m16_36_port, 
      m16_35_port, m16_34_port, m16_33_port, m16_32_port, m16_31_port, 
      m16_30_port, m16_29_port, m16_28_port, m16_27_port, m16_26_port, 
      m16_25_port, m16_24_port, m16_23_port, m16_15_port, m16_14_port, 
      m16_13_port, m16_12_port, m16_11_port, m16_10_port, m16_9_port, 
      m16_8_port, m16_7_port, m16_6_port, m16_5_port, m16_4_port, m16_3_port, 
      m16_2_port, m16_1_port, m16_0_port, y_38_port, y_37_port, y_36_port, 
      y_35_port, y_34_port, y_33_port, y_32_port, y_31_port, y_30_port, 
      y_29_port, y_28_port, y_27_port, y_26_port, y_25_port, y_24_port, 
      y_23_port, y_22_port, y_21_port, y_20_port, y_19_port, y_18_port, 
      y_17_port, y_16_port, y_15_port, y_14_port, y_13_port, y_12_port, 
      y_11_port, y_10_port, y_9_port, y_8_port, y_7_port, y_6_port, y_5_port, 
      y_4_port, y_3_port, y_2_port, y_1_port, y_0_port, n2, n3, n4, n6, n10, 
      n11, n12, n9, n14, n15, n16, n17 : std_logic;

begin
   
   IL : shift_firstLevel port map( A(31) => A(31), A(30) => A(30), A(29) => 
                           A(29), A(28) => A(28), A(27) => A(27), A(26) => 
                           A(26), A(25) => A(25), A(24) => A(24), A(23) => 
                           A(23), A(22) => A(22), A(21) => A(21), A(20) => 
                           A(20), A(19) => A(19), A(18) => A(18), A(17) => 
                           A(17), A(16) => A(16), A(15) => A(15), A(14) => 
                           A(14), A(13) => A(13), A(12) => A(12), A(11) => 
                           A(11), A(10) => A(10), A(9) => A(9), A(8) => A(8), 
                           A(7) => A(7), A(6) => A(6), A(5) => A(5), A(4) => 
                           A(4), A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), sel(1) => LOGIC_ARITH, sel(0) => LEFT_RIGHT
                           , mask00(38) => m0_38_port, mask00(37) => m0_37_port
                           , mask00(36) => m0_36_port, mask00(35) => m0_35_port
                           , mask00(34) => m0_34_port, mask00(33) => m0_33_port
                           , mask00(32) => m0_32_port, mask00(31) => m0_31_port
                           , mask00(30) => m0_30_port, mask00(29) => m0_29_port
                           , mask00(28) => m0_28_port, mask00(27) => m0_27_port
                           , mask00(26) => m0_26_port, mask00(25) => m0_25_port
                           , mask00(24) => m0_24_port, mask00(23) => m0_23_port
                           , mask00(22) => m0_22_port, mask00(21) => m0_21_port
                           , mask00(20) => m0_20_port, mask00(19) => m0_19_port
                           , mask00(18) => m0_18_port, mask00(17) => m0_17_port
                           , mask00(16) => m0_16_port, mask00(15) => m0_15_port
                           , mask00(14) => m0_14_port, mask00(13) => m0_13_port
                           , mask00(12) => m0_12_port, mask00(11) => m0_11_port
                           , mask00(10) => m0_10_port, mask00(9) => m0_9_port, 
                           mask00(8) => m0_8_port, mask00(7) => m0_7_port, 
                           mask00(6) => m0_6_port, mask00(5) => m0_5_port, 
                           mask00(4) => m0_4_port, mask00(3) => m0_3_port, 
                           mask00(2) => m0_2_port, mask00(1) => m0_1_port, 
                           mask00(0) => m0_0_port, mask08(38) => m8_38_port, 
                           mask08(37) => m8_37_port, mask08(36) => m8_36_port, 
                           mask08(35) => m8_35_port, mask08(34) => m8_34_port, 
                           mask08(33) => m8_33_port, mask08(32) => m8_32_port, 
                           mask08(31) => m8_31_port, mask08(30) => m8_30_port, 
                           mask08(29) => m8_29_port, mask08(28) => m8_28_port, 
                           mask08(27) => m8_27_port, mask08(26) => m8_26_port, 
                           mask08(25) => m8_25_port, mask08(24) => m8_24_port, 
                           mask08(23) => m8_23_port, mask08(22) => m8_22_port, 
                           mask08(21) => m8_21_port, mask08(20) => m8_20_port, 
                           mask08(19) => m8_19_port, mask08(18) => m8_18_port, 
                           mask08(17) => m8_17_port, mask08(16) => m8_16_port, 
                           mask08(15) => m8_15_port, mask08(14) => m8_14_port, 
                           mask08(13) => m8_13_port, mask08(12) => m8_12_port, 
                           mask08(11) => m8_11_port, mask08(10) => m8_10_port, 
                           mask08(9) => m8_9_port, mask08(8) => m8_8_port, 
                           mask08(7) => m8_7_port, mask08(6) => m8_6_port, 
                           mask08(5) => m8_5_port, mask08(4) => m8_4_port, 
                           mask08(3) => m8_3_port, mask08(2) => m8_2_port, 
                           mask08(1) => m8_1_port, mask08(0) => m8_0_port, 
                           mask16(38) => m16_38_port, mask16(37) => m16_37_port
                           , mask16(36) => m16_36_port, mask16(35) => 
                           m16_35_port, mask16(34) => m16_34_port, mask16(33) 
                           => m16_33_port, mask16(32) => m16_32_port, 
                           mask16(31) => m16_31_port, mask16(30) => m16_30_port
                           , mask16(29) => m16_29_port, mask16(28) => 
                           m16_28_port, mask16(27) => m16_27_port, mask16(26) 
                           => m16_26_port, mask16(25) => m16_25_port, 
                           mask16(24) => m16_24_port, mask16(23) => m16_23_port
                           , mask16(22) => n3, mask16(21) => n11, mask16(20) =>
                           n6, mask16(19) => n2, mask16(18) => n12, mask16(17) 
                           => n4, mask16(16) => n10, mask16(15) => m16_15_port,
                           mask16(14) => m16_14_port, mask16(13) => m16_13_port
                           , mask16(12) => m16_12_port, mask16(11) => 
                           m16_11_port, mask16(10) => m16_10_port, mask16(9) =>
                           m16_9_port, mask16(8) => m16_8_port, mask16(7) => 
                           m16_7_port, mask16(6) => m16_6_port, mask16(5) => 
                           m16_5_port, mask16(4) => m16_4_port, mask16(3) => 
                           m16_3_port, mask16(2) => m16_2_port, mask16(1) => 
                           m16_1_port, mask16(0) => m16_0_port);
   IIL : shift_secondLevel port map( sel(1) => B(4), sel(0) => B(3), mask00(38)
                           => m0_38_port, mask00(37) => m0_37_port, mask00(36) 
                           => m0_36_port, mask00(35) => m0_35_port, mask00(34) 
                           => m0_34_port, mask00(33) => m0_33_port, mask00(32) 
                           => m0_32_port, mask00(31) => m0_31_port, mask00(30) 
                           => m0_30_port, mask00(29) => m0_29_port, mask00(28) 
                           => m0_28_port, mask00(27) => m0_27_port, mask00(26) 
                           => m0_26_port, mask00(25) => m0_25_port, mask00(24) 
                           => m0_24_port, mask00(23) => m0_23_port, mask00(22) 
                           => m0_22_port, mask00(21) => m0_21_port, mask00(20) 
                           => m0_20_port, mask00(19) => m0_19_port, mask00(18) 
                           => m0_18_port, mask00(17) => m0_17_port, mask00(16) 
                           => m0_16_port, mask00(15) => m0_15_port, mask00(14) 
                           => m0_14_port, mask00(13) => m0_13_port, mask00(12) 
                           => m0_12_port, mask00(11) => m0_11_port, mask00(10) 
                           => m0_10_port, mask00(9) => m0_9_port, mask00(8) => 
                           m0_8_port, mask00(7) => m0_7_port, mask00(6) => 
                           m0_6_port, mask00(5) => m0_5_port, mask00(4) => 
                           m0_4_port, mask00(3) => m0_3_port, mask00(2) => 
                           m0_2_port, mask00(1) => m0_1_port, mask00(0) => 
                           m0_0_port, mask08(38) => m8_38_port, mask08(37) => 
                           m8_37_port, mask08(36) => m8_36_port, mask08(35) => 
                           m8_35_port, mask08(34) => m8_34_port, mask08(33) => 
                           m8_33_port, mask08(32) => m8_32_port, mask08(31) => 
                           m8_31_port, mask08(30) => m8_30_port, mask08(29) => 
                           m8_29_port, mask08(28) => m8_28_port, mask08(27) => 
                           m8_27_port, mask08(26) => m8_26_port, mask08(25) => 
                           m8_25_port, mask08(24) => m8_24_port, mask08(23) => 
                           m8_23_port, mask08(22) => m8_22_port, mask08(21) => 
                           m8_21_port, mask08(20) => m8_20_port, mask08(19) => 
                           m8_19_port, mask08(18) => m8_18_port, mask08(17) => 
                           m8_17_port, mask08(16) => m8_16_port, mask08(15) => 
                           m8_15_port, mask08(14) => m8_14_port, mask08(13) => 
                           m8_13_port, mask08(12) => m8_12_port, mask08(11) => 
                           m8_11_port, mask08(10) => m8_10_port, mask08(9) => 
                           m8_9_port, mask08(8) => m8_8_port, mask08(7) => 
                           m8_7_port, mask08(6) => m8_6_port, mask08(5) => 
                           m8_5_port, mask08(4) => m8_4_port, mask08(3) => 
                           m8_3_port, mask08(2) => m8_2_port, mask08(1) => 
                           m8_1_port, mask08(0) => m8_0_port, mask16(38) => 
                           m16_38_port, mask16(37) => m16_37_port, mask16(36) 
                           => m16_36_port, mask16(35) => m16_35_port, 
                           mask16(34) => m16_34_port, mask16(33) => m16_33_port
                           , mask16(32) => m16_32_port, mask16(31) => 
                           m16_31_port, mask16(30) => m16_30_port, mask16(29) 
                           => m16_29_port, mask16(28) => m16_28_port, 
                           mask16(27) => m16_27_port, mask16(26) => m16_26_port
                           , mask16(25) => m16_25_port, mask16(24) => 
                           m16_24_port, mask16(23) => m16_23_port, mask16(22) 
                           => n3, mask16(21) => n11, mask16(20) => n6, 
                           mask16(19) => n2, mask16(18) => n12, mask16(17) => 
                           n4, mask16(16) => n10, mask16(15) => m16_15_port, 
                           mask16(14) => m16_14_port, mask16(13) => m16_13_port
                           , mask16(12) => m16_12_port, mask16(11) => 
                           m16_11_port, mask16(10) => m16_10_port, mask16(9) =>
                           m16_9_port, mask16(8) => m16_8_port, mask16(7) => 
                           m16_7_port, mask16(6) => m16_6_port, mask16(5) => 
                           m16_5_port, mask16(4) => m16_4_port, mask16(3) => 
                           m16_3_port, mask16(2) => m16_2_port, mask16(1) => 
                           m16_1_port, mask16(0) => m16_0_port, Y(38) => 
                           y_38_port, Y(37) => y_37_port, Y(36) => y_36_port, 
                           Y(35) => y_35_port, Y(34) => y_34_port, Y(33) => 
                           y_33_port, Y(32) => y_32_port, Y(31) => y_31_port, 
                           Y(30) => y_30_port, Y(29) => y_29_port, Y(28) => 
                           y_28_port, Y(27) => y_27_port, Y(26) => y_26_port, 
                           Y(25) => y_25_port, Y(24) => y_24_port, Y(23) => 
                           y_23_port, Y(22) => y_22_port, Y(21) => y_21_port, 
                           Y(20) => y_20_port, Y(19) => y_19_port, Y(18) => 
                           y_18_port, Y(17) => y_17_port, Y(16) => y_16_port, 
                           Y(15) => y_15_port, Y(14) => y_14_port, Y(13) => 
                           y_13_port, Y(12) => y_12_port, Y(11) => y_11_port, 
                           Y(10) => y_10_port, Y(9) => y_9_port, Y(8) => 
                           y_8_port, Y(7) => y_7_port, Y(6) => y_6_port, Y(5) 
                           => y_5_port, Y(4) => y_4_port, Y(3) => y_3_port, 
                           Y(2) => y_2_port, Y(1) => y_1_port, Y(0) => y_0_port
                           );
   IIIL : shift_thirdLevel port map( sel(2) => s3_2_port, sel(1) => s3_1_port, 
                           sel(0) => s3_0_port, A(38) => y_38_port, A(37) => 
                           y_37_port, A(36) => y_36_port, A(35) => y_35_port, 
                           A(34) => y_34_port, A(33) => y_33_port, A(32) => 
                           y_32_port, A(31) => y_31_port, A(30) => y_30_port, 
                           A(29) => y_29_port, A(28) => y_28_port, A(27) => 
                           y_27_port, A(26) => y_26_port, A(25) => y_25_port, 
                           A(24) => y_24_port, A(23) => y_23_port, A(22) => 
                           y_22_port, A(21) => y_21_port, A(20) => y_20_port, 
                           A(19) => y_19_port, A(18) => y_18_port, A(17) => 
                           y_17_port, A(16) => y_16_port, A(15) => y_15_port, 
                           A(14) => y_14_port, A(13) => y_13_port, A(12) => 
                           y_12_port, A(11) => y_11_port, A(10) => y_10_port, 
                           A(9) => y_9_port, A(8) => y_8_port, A(7) => y_7_port
                           , A(6) => y_6_port, A(5) => y_5_port, A(4) => 
                           y_4_port, A(3) => y_3_port, A(2) => y_2_port, A(1) 
                           => y_1_port, A(0) => y_0_port, Y(31) => OUTPUT(31), 
                           Y(30) => OUTPUT(30), Y(29) => OUTPUT(29), Y(28) => 
                           OUTPUT(28), Y(27) => OUTPUT(27), Y(26) => OUTPUT(26)
                           , Y(25) => OUTPUT(25), Y(24) => OUTPUT(24), Y(23) =>
                           OUTPUT(23), Y(22) => OUTPUT(22), Y(21) => OUTPUT(21)
                           , Y(20) => OUTPUT(20), Y(19) => OUTPUT(19), Y(18) =>
                           OUTPUT(18), Y(17) => OUTPUT(17), Y(16) => OUTPUT(16)
                           , Y(15) => OUTPUT(15), Y(14) => OUTPUT(14), Y(13) =>
                           OUTPUT(13), Y(12) => OUTPUT(12), Y(11) => OUTPUT(11)
                           , Y(10) => OUTPUT(10), Y(9) => OUTPUT(9), Y(8) => 
                           OUTPUT(8), Y(7) => OUTPUT(7), Y(6) => OUTPUT(6), 
                           Y(5) => OUTPUT(5), Y(4) => OUTPUT(4), Y(3) => 
                           OUTPUT(3), Y(2) => OUTPUT(2), Y(1) => OUTPUT(1), 
                           Y(0) => OUTPUT(0));
   U8 : OR2_X1 port map( A1 => LOGIC_ARITH, A2 => LEFT_RIGHT, ZN => n9);
   U1 : INV_X1 port map( A => LEFT_RIGHT, ZN => n17);
   U2 : INV_X1 port map( A => B(0), ZN => n16);
   U3 : INV_X1 port map( A => B(2), ZN => n14);
   U4 : INV_X1 port map( A => B(1), ZN => n15);
   U5 : AOI22_X1 port map( A1 => B(0), A2 => n9, B1 => n17, B2 => n16, ZN => 
                           s3_0_port);
   U6 : AOI22_X1 port map( A1 => B(2), A2 => n9, B1 => n17, B2 => n14, ZN => 
                           s3_2_port);
   U7 : AOI22_X1 port map( A1 => B(1), A2 => n9, B1 => n17, B2 => n15, ZN => 
                           s3_1_port);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity comparator_M32 is

   port( C, V : in std_logic;  SUM : in std_logic_vector (31 downto 0);  sel : 
         in std_logic_vector (2 downto 0);  sign : in std_logic;  S : out 
         std_logic);

end comparator_M32;

architecture SYN_BEHAVIORAL of comparator_M32 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   signal n6, n24, n23, n22, n21, n20, n19, n18, n17, n66, n67, n68, n69, n70, 
      n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83 : 
      std_logic;

begin
   
   U14 : NOR4_X1 port map( A1 => SUM(9), A2 => SUM(8), A3 => SUM(7), A4 => 
                           SUM(6), ZN => n18);
   U17 : NOR4_X1 port map( A1 => SUM(16), A2 => SUM(15), A3 => SUM(14), A4 => 
                           SUM(13), ZN => n24);
   U18 : NOR4_X1 port map( A1 => SUM(12), A2 => SUM(11), A3 => SUM(10), A4 => 
                           SUM(0), ZN => n23);
   U20 : NOR4_X1 port map( A1 => SUM(1), A2 => SUM(19), A3 => SUM(18), A4 => 
                           SUM(17), ZN => n21);
   U1 : XNOR2_X1 port map( A => n83, B => V, ZN => n66);
   U2 : MUX2_X1 port map( A => C, B => n66, S => sign, Z => n6);
   U3 : INV_X1 port map( A => sel(0), ZN => n77);
   U4 : INV_X1 port map( A => sel(1), ZN => n80);
   U5 : INV_X1 port map( A => sel(2), ZN => n79);
   U6 : AND3_X1 port map( A1 => n21, A2 => n68, A3 => n22, ZN => n69);
   U7 : AND2_X1 port map( A1 => n24, A2 => n23, ZN => n68);
   U8 : CLKBUF_X1 port map( A => SUM(31), Z => n83);
   U9 : AND2_X1 port map( A1 => n67, A2 => n69, ZN => n71);
   U10 : AND2_X1 port map( A1 => n67, A2 => n69, ZN => n70);
   U11 : AND4_X1 port map( A1 => n17, A2 => n18, A3 => n19, A4 => n20, ZN => 
                           n67);
   U12 : NOR2_X1 port map( A1 => sel(0), A2 => sel(1), ZN => n76);
   U13 : NAND2_X1 port map( A1 => n79, A2 => n80, ZN => n78);
   U15 : AOI21_X1 port map( B1 => n71, B2 => n77, A => n78, ZN => n74);
   U16 : XNOR2_X1 port map( A => n70, B => n76, ZN => n75);
   U19 : NAND2_X1 port map( A1 => n71, A2 => sel(0), ZN => n82);
   U21 : NAND2_X1 port map( A1 => n73, A2 => n72, ZN => S);
   U22 : NOR4_X1 port map( A1 => SUM(23), A2 => SUM(22), A3 => SUM(21), A4 => 
                           SUM(20), ZN => n22);
   U23 : NOR4_X1 port map( A1 => SUM(30), A2 => SUM(28), A3 => SUM(29), A4 => 
                           SUM(2), ZN => n20);
   U24 : NOR4_X1 port map( A1 => SUM(27), A2 => SUM(26), A3 => SUM(25), A4 => 
                           SUM(24), ZN => n19);
   U25 : NOR4_X1 port map( A1 => SUM(31), A2 => SUM(5), A3 => SUM(3), A4 => 
                           SUM(4), ZN => n17);
   U26 : NAND3_X1 port map( A1 => n81, A2 => n79, A3 => sel(1), ZN => n72);
   U27 : NAND2_X1 port map( A1 => n6, A2 => n82, ZN => n81);
   U28 : AOI22_X1 port map( A1 => n6, A2 => n74, B1 => n75, B2 => sel(2), ZN =>
                           n73);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity simple_booth_add_ext_N16 is

   port( Clock, Reset, sign, enable : in std_logic;  valid : out std_logic;  A,
         B : in std_logic_vector (15 downto 0);  A_to_add, B_to_add : out 
         std_logic_vector (31 downto 0);  sign_to_add : out std_logic;  
         final_out : out std_logic_vector (31 downto 0);  ACC_from_add : in 
         std_logic_vector (31 downto 0));

end simple_booth_add_ext_N16;

architecture SYN_struct of simple_booth_add_ext_N16 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X8
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component ff32_en_SIZE32_1
      port( D : in std_logic_vector (31 downto 0);  en, clk, rst : in std_logic
            ;  Q : out std_logic_vector (31 downto 0));
   end component;
   
   component mux21_1
      port( IN0, IN1 : in std_logic_vector (31 downto 0);  CTRL : in std_logic;
            OUT1 : out std_logic_vector (31 downto 0));
   end component;
   
   component piso_r_2_N32
      port( Clock, ALOAD : in std_logic;  D : in std_logic_vector (31 downto 0)
            ;  SO : out std_logic_vector (31 downto 0));
   end component;
   
   component shift_N9_1
      port( Clock, ALOAD : in std_logic;  D : in std_logic_vector (8 downto 0);
            SO : out std_logic);
   end component;
   
   component shift_N9_2
      port( Clock, ALOAD : in std_logic;  D : in std_logic_vector (8 downto 0);
            SO : out std_logic);
   end component;
   
   component shift_N9_0
      port( Clock, ALOAD : in std_logic;  D : in std_logic_vector (8 downto 0);
            SO : out std_logic);
   end component;
   
   component booth_encoder_1
      port( B_in : in std_logic_vector (2 downto 0);  A_out : out 
            std_logic_vector (2 downto 0));
   end component;
   
   component booth_encoder_2
      port( B_in : in std_logic_vector (2 downto 0);  A_out : out 
            std_logic_vector (2 downto 0));
   end component;
   
   component booth_encoder_3
      port( B_in : in std_logic_vector (2 downto 0);  A_out : out 
            std_logic_vector (2 downto 0));
   end component;
   
   component booth_encoder_4
      port( B_in : in std_logic_vector (2 downto 0);  A_out : out 
            std_logic_vector (2 downto 0));
   end component;
   
   component booth_encoder_5
      port( B_in : in std_logic_vector (2 downto 0);  A_out : out 
            std_logic_vector (2 downto 0));
   end component;
   
   component booth_encoder_6
      port( B_in : in std_logic_vector (2 downto 0);  A_out : out 
            std_logic_vector (2 downto 0));
   end component;
   
   component booth_encoder_7
      port( B_in : in std_logic_vector (2 downto 0);  A_out : out 
            std_logic_vector (2 downto 0));
   end component;
   
   component booth_encoder_8
      port( B_in : in std_logic_vector (2 downto 0);  A_out : out 
            std_logic_vector (2 downto 0));
   end component;
   
   component booth_encoder_0
      port( B_in : in std_logic_vector (2 downto 0);  A_out : out 
            std_logic_vector (2 downto 0));
   end component;
   
   component DFFS_X1
      port( D, CK, SN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal X_Logic0_port, valid_port, A_to_add_31_port, A_to_add_30_port, 
      A_to_add_29_port, A_to_add_28_port, A_to_add_27_port, A_to_add_26_port, 
      A_to_add_25_port, A_to_add_24_port, A_to_add_23_port, A_to_add_22_port, 
      A_to_add_21_port, A_to_add_20_port, A_to_add_19_port, A_to_add_18_port, 
      A_to_add_17_port, A_to_add_16_port, A_to_add_15_port, A_to_add_14_port, 
      A_to_add_13_port, A_to_add_12_port, A_to_add_11_port, A_to_add_10_port, 
      A_to_add_9_port, A_to_add_8_port, A_to_add_7_port, A_to_add_6_port, 
      A_to_add_5_port, A_to_add_4_port, A_to_add_3_port, A_to_add_2_port, 
      A_to_add_1_port, A_to_add_0_port, enc_N2_in_2_port, piso_0_in_8_port, 
      piso_0_in_7_port, piso_0_in_6_port, piso_0_in_5_port, piso_0_in_4_port, 
      piso_0_in_3_port, piso_0_in_2_port, piso_0_in_1_port, piso_0_in_0_port, 
      piso_1_in_8_port, piso_1_in_7_port, piso_1_in_6_port, piso_1_in_5_port, 
      piso_1_in_4_port, piso_1_in_3_port, piso_1_in_2_port, piso_1_in_1_port, 
      piso_1_in_0_port, piso_2_in_8_port, piso_2_in_7_port, piso_2_in_6_port, 
      piso_2_in_5_port, piso_2_in_4_port, piso_2_in_3_port, piso_2_in_2_port, 
      piso_2_in_1_port, piso_2_in_0_port, extend_vector_15_port, 
      A_to_mux_31_port, A_to_mux_30_port, A_to_mux_29_port, A_to_mux_28_port, 
      A_to_mux_27_port, A_to_mux_26_port, A_to_mux_25_port, A_to_mux_24_port, 
      A_to_mux_23_port, A_to_mux_22_port, A_to_mux_21_port, A_to_mux_20_port, 
      A_to_mux_19_port, A_to_mux_18_port, A_to_mux_17_port, A_to_mux_16_port, 
      A_to_mux_15_port, A_to_mux_14_port, A_to_mux_13_port, A_to_mux_12_port, 
      A_to_mux_11_port, A_to_mux_10_port, A_to_mux_9_port, A_to_mux_8_port, 
      A_to_mux_7_port, A_to_mux_6_port, A_to_mux_5_port, A_to_mux_4_port, 
      A_to_mux_3_port, A_to_mux_2_port, A_to_mux_1_port, A_to_mux_0_port, 
      input_mux_sel_2_port, input_mux_sel_0, next_accumulate_31_port, 
      next_accumulate_30_port, next_accumulate_29_port, next_accumulate_28_port
      , next_accumulate_27_port, next_accumulate_26_port, 
      next_accumulate_25_port, next_accumulate_24_port, next_accumulate_23_port
      , next_accumulate_22_port, next_accumulate_21_port, 
      next_accumulate_20_port, next_accumulate_19_port, next_accumulate_18_port
      , next_accumulate_17_port, next_accumulate_16_port, 
      next_accumulate_15_port, next_accumulate_14_port, next_accumulate_13_port
      , next_accumulate_12_port, next_accumulate_11_port, 
      next_accumulate_10_port, next_accumulate_9_port, next_accumulate_8_port, 
      next_accumulate_7_port, next_accumulate_6_port, next_accumulate_5_port, 
      next_accumulate_4_port, next_accumulate_3_port, next_accumulate_2_port, 
      next_accumulate_1_port, next_accumulate_0_port, reg_enable, n50, n51, n52
      , n54, n22, n37, n40, net645046, n49, n53, n55, n56, n57, n58, n59, n60, 
      n61, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76
      , n77, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n90, n91, n92, 
      n93, n41, n42, n46, n47, n48, n62, n78, net684315, net684316, net684317 :
      std_logic;

begin
   valid <= valid_port;
   A_to_add <= ( A_to_add_31_port, A_to_add_30_port, A_to_add_29_port, 
      A_to_add_28_port, A_to_add_27_port, A_to_add_26_port, A_to_add_25_port, 
      A_to_add_24_port, A_to_add_23_port, A_to_add_22_port, A_to_add_21_port, 
      A_to_add_20_port, A_to_add_19_port, A_to_add_18_port, A_to_add_17_port, 
      A_to_add_16_port, A_to_add_15_port, A_to_add_14_port, A_to_add_13_port, 
      A_to_add_12_port, A_to_add_11_port, A_to_add_10_port, A_to_add_9_port, 
      A_to_add_8_port, A_to_add_7_port, A_to_add_6_port, A_to_add_5_port, 
      A_to_add_4_port, A_to_add_3_port, A_to_add_2_port, A_to_add_1_port, 
      A_to_add_0_port );
   
   X_Logic0_port <= '0';
   count_reg_1_inst : DFFR_X1 port map( D => n51, CK => Clock, RN => n78, Q => 
                           n48, QN => net645046);
   count_reg_2_inst : DFFR_X1 port map( D => n50, CK => Clock, RN => n78, Q => 
                           net684317, QN => n37);
   count_reg_0_inst : DFFS_X1 port map( D => n54, CK => Clock, SN => n78, Q => 
                           net684316, QN => n40);
   count_reg_3_inst : DFFS_X1 port map( D => n52, CK => Clock, SN => n78, Q => 
                           net684315, QN => n47);
   U85 : MUX2_X1 port map( A => n49, B => n48, S => n86, Z => n51);
   U87 : MUX2_X1 port map( A => A_to_add_9_port, B => ACC_from_add(9), S => n62
                           , Z => final_out(9));
   U88 : MUX2_X1 port map( A => A_to_add_8_port, B => ACC_from_add(8), S => 
                           input_mux_sel_2_port, Z => final_out(8));
   U89 : MUX2_X1 port map( A => A_to_add_7_port, B => ACC_from_add(7), S => 
                           input_mux_sel_2_port, Z => final_out(7));
   U90 : MUX2_X1 port map( A => A_to_add_6_port, B => ACC_from_add(6), S => n62
                           , Z => final_out(6));
   U91 : MUX2_X1 port map( A => A_to_add_5_port, B => ACC_from_add(5), S => 
                           input_mux_sel_2_port, Z => final_out(5));
   U92 : MUX2_X1 port map( A => A_to_add_4_port, B => ACC_from_add(4), S => 
                           input_mux_sel_2_port, Z => final_out(4));
   U93 : MUX2_X1 port map( A => A_to_add_3_port, B => ACC_from_add(3), S => 
                           input_mux_sel_2_port, Z => final_out(3));
   U94 : MUX2_X1 port map( A => A_to_add_31_port, B => ACC_from_add(31), S => 
                           input_mux_sel_2_port, Z => final_out(31));
   U95 : MUX2_X1 port map( A => A_to_add_30_port, B => ACC_from_add(30), S => 
                           input_mux_sel_2_port, Z => final_out(30));
   U97 : MUX2_X1 port map( A => A_to_add_29_port, B => ACC_from_add(29), S => 
                           input_mux_sel_2_port, Z => final_out(29));
   U98 : MUX2_X1 port map( A => A_to_add_28_port, B => ACC_from_add(28), S => 
                           input_mux_sel_2_port, Z => final_out(28));
   U100 : MUX2_X1 port map( A => A_to_add_26_port, B => ACC_from_add(26), S => 
                           input_mux_sel_2_port, Z => final_out(26));
   U101 : MUX2_X1 port map( A => A_to_add_25_port, B => ACC_from_add(25), S => 
                           input_mux_sel_2_port, Z => final_out(25));
   U102 : MUX2_X1 port map( A => A_to_add_24_port, B => ACC_from_add(24), S => 
                           input_mux_sel_2_port, Z => final_out(24));
   U103 : MUX2_X1 port map( A => A_to_add_23_port, B => ACC_from_add(23), S => 
                           input_mux_sel_2_port, Z => final_out(23));
   U104 : MUX2_X1 port map( A => A_to_add_22_port, B => ACC_from_add(22), S => 
                           input_mux_sel_2_port, Z => final_out(22));
   U105 : MUX2_X1 port map( A => A_to_add_21_port, B => ACC_from_add(21), S => 
                           input_mux_sel_2_port, Z => final_out(21));
   U106 : MUX2_X1 port map( A => A_to_add_20_port, B => ACC_from_add(20), S => 
                           input_mux_sel_2_port, Z => final_out(20));
   U107 : MUX2_X1 port map( A => A_to_add_1_port, B => ACC_from_add(1), S => 
                           n62, Z => final_out(1));
   U108 : MUX2_X1 port map( A => A_to_add_19_port, B => ACC_from_add(19), S => 
                           n62, Z => final_out(19));
   U109 : MUX2_X1 port map( A => A_to_add_18_port, B => ACC_from_add(18), S => 
                           n62, Z => final_out(18));
   U110 : MUX2_X1 port map( A => A_to_add_17_port, B => ACC_from_add(17), S => 
                           n62, Z => final_out(17));
   U111 : MUX2_X1 port map( A => A_to_add_16_port, B => ACC_from_add(16), S => 
                           n62, Z => final_out(16));
   U112 : MUX2_X1 port map( A => A_to_add_15_port, B => ACC_from_add(15), S => 
                           n62, Z => final_out(15));
   U113 : MUX2_X1 port map( A => A_to_add_14_port, B => ACC_from_add(14), S => 
                           n62, Z => final_out(14));
   U114 : MUX2_X1 port map( A => A_to_add_13_port, B => ACC_from_add(13), S => 
                           n62, Z => final_out(13));
   U115 : MUX2_X1 port map( A => A_to_add_12_port, B => ACC_from_add(12), S => 
                           n62, Z => final_out(12));
   U116 : MUX2_X1 port map( A => A_to_add_11_port, B => ACC_from_add(11), S => 
                           n62, Z => final_out(11));
   U117 : MUX2_X1 port map( A => A_to_add_10_port, B => ACC_from_add(10), S => 
                           n62, Z => final_out(10));
   encod_0_0 : booth_encoder_0 port map( B_in(2) => B(1), B_in(1) => B(0), 
                           B_in(0) => X_Logic0_port, A_out(2) => 
                           piso_2_in_0_port, A_out(1) => piso_1_in_0_port, 
                           A_out(0) => piso_0_in_0_port);
   encod_i_1 : booth_encoder_8 port map( B_in(2) => B(3), B_in(1) => B(2), 
                           B_in(0) => B(1), A_out(2) => piso_2_in_1_port, 
                           A_out(1) => piso_1_in_1_port, A_out(0) => 
                           piso_0_in_1_port);
   encod_i_2 : booth_encoder_7 port map( B_in(2) => B(5), B_in(1) => B(4), 
                           B_in(0) => B(3), A_out(2) => piso_2_in_2_port, 
                           A_out(1) => piso_1_in_2_port, A_out(0) => 
                           piso_0_in_2_port);
   encod_i_3 : booth_encoder_6 port map( B_in(2) => B(7), B_in(1) => B(6), 
                           B_in(0) => B(5), A_out(2) => piso_2_in_3_port, 
                           A_out(1) => piso_1_in_3_port, A_out(0) => 
                           piso_0_in_3_port);
   encod_i_4 : booth_encoder_5 port map( B_in(2) => B(9), B_in(1) => B(8), 
                           B_in(0) => B(7), A_out(2) => piso_2_in_4_port, 
                           A_out(1) => piso_1_in_4_port, A_out(0) => 
                           piso_0_in_4_port);
   encod_i_5 : booth_encoder_4 port map( B_in(2) => B(11), B_in(1) => B(10), 
                           B_in(0) => B(9), A_out(2) => piso_2_in_5_port, 
                           A_out(1) => piso_1_in_5_port, A_out(0) => 
                           piso_0_in_5_port);
   encod_i_6 : booth_encoder_3 port map( B_in(2) => B(13), B_in(1) => B(12), 
                           B_in(0) => B(11), A_out(2) => piso_2_in_6_port, 
                           A_out(1) => piso_1_in_6_port, A_out(0) => 
                           piso_0_in_6_port);
   encod_i_7 : booth_encoder_2 port map( B_in(2) => B(15), B_in(1) => B(14), 
                           B_in(0) => B(13), A_out(2) => piso_2_in_7_port, 
                           A_out(1) => piso_1_in_7_port, A_out(0) => 
                           piso_0_in_7_port);
   encod_i_8 : booth_encoder_1 port map( B_in(2) => enc_N2_in_2_port, B_in(1) 
                           => enc_N2_in_2_port, B_in(0) => B(15), A_out(2) => 
                           piso_2_in_8_port, A_out(1) => piso_1_in_8_port, 
                           A_out(0) => piso_0_in_8_port);
   piso_0 : shift_N9_0 port map( Clock => Clock, ALOAD => n46, D(8) => 
                           piso_0_in_8_port, D(7) => piso_0_in_7_port, D(6) => 
                           piso_0_in_6_port, D(5) => piso_0_in_5_port, D(4) => 
                           piso_0_in_4_port, D(3) => piso_0_in_3_port, D(2) => 
                           piso_0_in_2_port, D(1) => piso_0_in_1_port, D(0) => 
                           piso_0_in_0_port, SO => input_mux_sel_0);
   piso_1 : shift_N9_2 port map( Clock => Clock, ALOAD => n46, D(8) => 
                           piso_1_in_8_port, D(7) => piso_1_in_7_port, D(6) => 
                           piso_1_in_6_port, D(5) => piso_1_in_5_port, D(4) => 
                           piso_1_in_4_port, D(3) => piso_1_in_3_port, D(2) => 
                           piso_1_in_2_port, D(1) => piso_1_in_1_port, D(0) => 
                           piso_1_in_0_port, SO => sign_to_add);
   piso_2 : shift_N9_1 port map( Clock => Clock, ALOAD => n46, D(8) => 
                           piso_2_in_8_port, D(7) => piso_2_in_7_port, D(6) => 
                           piso_2_in_6_port, D(5) => piso_2_in_5_port, D(4) => 
                           piso_2_in_4_port, D(3) => piso_2_in_3_port, D(2) => 
                           piso_2_in_2_port, D(1) => piso_2_in_1_port, D(0) => 
                           piso_2_in_0_port, SO => input_mux_sel_2_port);
   A_reg : piso_r_2_N32 port map( Clock => Clock, ALOAD => n46, D(31) => 
                           extend_vector_15_port, D(30) => 
                           extend_vector_15_port, D(29) => 
                           extend_vector_15_port, D(28) => 
                           extend_vector_15_port, D(27) => 
                           extend_vector_15_port, D(26) => 
                           extend_vector_15_port, D(25) => 
                           extend_vector_15_port, D(24) => 
                           extend_vector_15_port, D(23) => 
                           extend_vector_15_port, D(22) => 
                           extend_vector_15_port, D(21) => 
                           extend_vector_15_port, D(20) => 
                           extend_vector_15_port, D(19) => 
                           extend_vector_15_port, D(18) => 
                           extend_vector_15_port, D(17) => 
                           extend_vector_15_port, D(16) => 
                           extend_vector_15_port, D(15) => A(15), D(14) => 
                           A(14), D(13) => A(13), D(12) => A(12), D(11) => 
                           A(11), D(10) => A(10), D(9) => A(9), D(8) => A(8), 
                           D(7) => A(7), D(6) => A(6), D(5) => A(5), D(4) => 
                           A(4), D(3) => A(3), D(2) => A(2), D(1) => A(1), D(0)
                           => A(0), SO(31) => A_to_mux_31_port, SO(30) => 
                           A_to_mux_30_port, SO(29) => A_to_mux_29_port, SO(28)
                           => A_to_mux_28_port, SO(27) => A_to_mux_27_port, 
                           SO(26) => A_to_mux_26_port, SO(25) => 
                           A_to_mux_25_port, SO(24) => A_to_mux_24_port, SO(23)
                           => A_to_mux_23_port, SO(22) => A_to_mux_22_port, 
                           SO(21) => A_to_mux_21_port, SO(20) => 
                           A_to_mux_20_port, SO(19) => A_to_mux_19_port, SO(18)
                           => A_to_mux_18_port, SO(17) => A_to_mux_17_port, 
                           SO(16) => A_to_mux_16_port, SO(15) => 
                           A_to_mux_15_port, SO(14) => A_to_mux_14_port, SO(13)
                           => A_to_mux_13_port, SO(12) => A_to_mux_12_port, 
                           SO(11) => A_to_mux_11_port, SO(10) => 
                           A_to_mux_10_port, SO(9) => A_to_mux_9_port, SO(8) =>
                           A_to_mux_8_port, SO(7) => A_to_mux_7_port, SO(6) => 
                           A_to_mux_6_port, SO(5) => A_to_mux_5_port, SO(4) => 
                           A_to_mux_4_port, SO(3) => A_to_mux_3_port, SO(2) => 
                           A_to_mux_2_port, SO(1) => A_to_mux_1_port, SO(0) => 
                           A_to_mux_0_port);
   INPUTMUX : mux21_1 port map( IN0(31) => A_to_mux_31_port, IN0(30) => 
                           A_to_mux_30_port, IN0(29) => A_to_mux_29_port, 
                           IN0(28) => A_to_mux_28_port, IN0(27) => 
                           A_to_mux_27_port, IN0(26) => A_to_mux_26_port, 
                           IN0(25) => A_to_mux_25_port, IN0(24) => 
                           A_to_mux_24_port, IN0(23) => A_to_mux_23_port, 
                           IN0(22) => A_to_mux_22_port, IN0(21) => 
                           A_to_mux_21_port, IN0(20) => A_to_mux_20_port, 
                           IN0(19) => A_to_mux_19_port, IN0(18) => 
                           A_to_mux_18_port, IN0(17) => A_to_mux_17_port, 
                           IN0(16) => A_to_mux_16_port, IN0(15) => 
                           A_to_mux_15_port, IN0(14) => A_to_mux_14_port, 
                           IN0(13) => A_to_mux_13_port, IN0(12) => 
                           A_to_mux_12_port, IN0(11) => A_to_mux_11_port, 
                           IN0(10) => A_to_mux_10_port, IN0(9) => 
                           A_to_mux_9_port, IN0(8) => A_to_mux_8_port, IN0(7) 
                           => A_to_mux_7_port, IN0(6) => A_to_mux_6_port, 
                           IN0(5) => A_to_mux_5_port, IN0(4) => A_to_mux_4_port
                           , IN0(3) => A_to_mux_3_port, IN0(2) => 
                           A_to_mux_2_port, IN0(1) => A_to_mux_1_port, IN0(0) 
                           => A_to_mux_0_port, IN1(31) => A_to_mux_30_port, 
                           IN1(30) => A_to_mux_29_port, IN1(29) => 
                           A_to_mux_28_port, IN1(28) => A_to_mux_27_port, 
                           IN1(27) => A_to_mux_26_port, IN1(26) => 
                           A_to_mux_25_port, IN1(25) => A_to_mux_24_port, 
                           IN1(24) => A_to_mux_23_port, IN1(23) => 
                           A_to_mux_22_port, IN1(22) => A_to_mux_21_port, 
                           IN1(21) => A_to_mux_20_port, IN1(20) => 
                           A_to_mux_19_port, IN1(19) => A_to_mux_18_port, 
                           IN1(18) => A_to_mux_17_port, IN1(17) => 
                           A_to_mux_16_port, IN1(16) => A_to_mux_15_port, 
                           IN1(15) => A_to_mux_14_port, IN1(14) => 
                           A_to_mux_13_port, IN1(13) => A_to_mux_12_port, 
                           IN1(12) => A_to_mux_11_port, IN1(11) => 
                           A_to_mux_10_port, IN1(10) => A_to_mux_9_port, IN1(9)
                           => A_to_mux_8_port, IN1(8) => A_to_mux_7_port, 
                           IN1(7) => A_to_mux_6_port, IN1(6) => A_to_mux_5_port
                           , IN1(5) => A_to_mux_4_port, IN1(4) => 
                           A_to_mux_3_port, IN1(3) => A_to_mux_2_port, IN1(2) 
                           => A_to_mux_1_port, IN1(1) => A_to_mux_0_port, 
                           IN1(0) => X_Logic0_port, CTRL => input_mux_sel_0, 
                           OUT1(31) => B_to_add(31), OUT1(30) => B_to_add(30), 
                           OUT1(29) => B_to_add(29), OUT1(28) => B_to_add(28), 
                           OUT1(27) => B_to_add(27), OUT1(26) => B_to_add(26), 
                           OUT1(25) => B_to_add(25), OUT1(24) => B_to_add(24), 
                           OUT1(23) => B_to_add(23), OUT1(22) => B_to_add(22), 
                           OUT1(21) => B_to_add(21), OUT1(20) => B_to_add(20), 
                           OUT1(19) => B_to_add(19), OUT1(18) => B_to_add(18), 
                           OUT1(17) => B_to_add(17), OUT1(16) => B_to_add(16), 
                           OUT1(15) => B_to_add(15), OUT1(14) => B_to_add(14), 
                           OUT1(13) => B_to_add(13), OUT1(12) => B_to_add(12), 
                           OUT1(11) => B_to_add(11), OUT1(10) => B_to_add(10), 
                           OUT1(9) => B_to_add(9), OUT1(8) => B_to_add(8), 
                           OUT1(7) => B_to_add(7), OUT1(6) => B_to_add(6), 
                           OUT1(5) => B_to_add(5), OUT1(4) => B_to_add(4), 
                           OUT1(3) => B_to_add(3), OUT1(2) => B_to_add(2), 
                           OUT1(1) => B_to_add(1), OUT1(0) => B_to_add(0));
   ACCUMULATOR : ff32_en_SIZE32_1 port map( D(31) => next_accumulate_31_port, 
                           D(30) => next_accumulate_30_port, D(29) => 
                           next_accumulate_29_port, D(28) => 
                           next_accumulate_28_port, D(27) => 
                           next_accumulate_27_port, D(26) => 
                           next_accumulate_26_port, D(25) => 
                           next_accumulate_25_port, D(24) => 
                           next_accumulate_24_port, D(23) => 
                           next_accumulate_23_port, D(22) => 
                           next_accumulate_22_port, D(21) => 
                           next_accumulate_21_port, D(20) => 
                           next_accumulate_20_port, D(19) => 
                           next_accumulate_19_port, D(18) => 
                           next_accumulate_18_port, D(17) => 
                           next_accumulate_17_port, D(16) => 
                           next_accumulate_16_port, D(15) => 
                           next_accumulate_15_port, D(14) => 
                           next_accumulate_14_port, D(13) => 
                           next_accumulate_13_port, D(12) => 
                           next_accumulate_12_port, D(11) => 
                           next_accumulate_11_port, D(10) => 
                           next_accumulate_10_port, D(9) => 
                           next_accumulate_9_port, D(8) => 
                           next_accumulate_8_port, D(7) => 
                           next_accumulate_7_port, D(6) => 
                           next_accumulate_6_port, D(5) => 
                           next_accumulate_5_port, D(4) => 
                           next_accumulate_4_port, D(3) => 
                           next_accumulate_3_port, D(2) => 
                           next_accumulate_2_port, D(1) => 
                           next_accumulate_1_port, D(0) => 
                           next_accumulate_0_port, en => reg_enable, clk => 
                           Clock, rst => Reset, Q(31) => A_to_add_31_port, 
                           Q(30) => A_to_add_30_port, Q(29) => A_to_add_29_port
                           , Q(28) => A_to_add_28_port, Q(27) => 
                           A_to_add_27_port, Q(26) => A_to_add_26_port, Q(25) 
                           => A_to_add_25_port, Q(24) => A_to_add_24_port, 
                           Q(23) => A_to_add_23_port, Q(22) => A_to_add_22_port
                           , Q(21) => A_to_add_21_port, Q(20) => 
                           A_to_add_20_port, Q(19) => A_to_add_19_port, Q(18) 
                           => A_to_add_18_port, Q(17) => A_to_add_17_port, 
                           Q(16) => A_to_add_16_port, Q(15) => A_to_add_15_port
                           , Q(14) => A_to_add_14_port, Q(13) => 
                           A_to_add_13_port, Q(12) => A_to_add_12_port, Q(11) 
                           => A_to_add_11_port, Q(10) => A_to_add_10_port, Q(9)
                           => A_to_add_9_port, Q(8) => A_to_add_8_port, Q(7) =>
                           A_to_add_7_port, Q(6) => A_to_add_6_port, Q(5) => 
                           A_to_add_5_port, Q(4) => A_to_add_4_port, Q(3) => 
                           A_to_add_3_port, Q(2) => A_to_add_2_port, Q(1) => 
                           A_to_add_1_port, Q(0) => A_to_add_0_port);
   U20 : NOR2_X1 port map( A1 => n46, A2 => n61, ZN => next_accumulate_31_port)
                           ;
   U38 : NOR2_X1 port map( A1 => n46, A2 => n70, ZN => next_accumulate_23_port)
                           ;
   U30 : NOR2_X1 port map( A1 => n46, A2 => n66, ZN => next_accumulate_27_port)
                           ;
   U40 : NOR2_X1 port map( A1 => n46, A2 => n71, ZN => next_accumulate_22_port)
                           ;
   U32 : NOR2_X1 port map( A1 => n46, A2 => n67, ZN => next_accumulate_26_port)
                           ;
   U26 : NOR2_X1 port map( A1 => n46, A2 => n64, ZN => next_accumulate_29_port)
                           ;
   U28 : NOR2_X1 port map( A1 => n46, A2 => n65, ZN => next_accumulate_28_port)
                           ;
   U34 : NOR2_X1 port map( A1 => n46, A2 => n68, ZN => next_accumulate_25_port)
                           ;
   U42 : NOR2_X1 port map( A1 => n46, A2 => n72, ZN => next_accumulate_21_port)
                           ;
   U44 : NOR2_X1 port map( A1 => n46, A2 => n73, ZN => next_accumulate_20_port)
                           ;
   U36 : NOR2_X1 port map( A1 => n46, A2 => n69, ZN => next_accumulate_24_port)
                           ;
   U48 : NOR2_X1 port map( A1 => n46, A2 => n75, ZN => next_accumulate_19_port)
                           ;
   U60 : NOR2_X1 port map( A1 => n46, A2 => n81, ZN => next_accumulate_13_port)
                           ;
   U58 : NOR2_X1 port map( A1 => n46, A2 => n80, ZN => next_accumulate_14_port)
                           ;
   U62 : NOR2_X1 port map( A1 => n46, A2 => n82, ZN => next_accumulate_12_port)
                           ;
   U56 : NOR2_X1 port map( A1 => n46, A2 => n79, ZN => next_accumulate_15_port)
                           ;
   U10 : NOR2_X1 port map( A1 => n46, A2 => n56, ZN => next_accumulate_7_port);
   U64 : NOR2_X1 port map( A1 => n46, A2 => n83, ZN => next_accumulate_11_port)
                           ;
   U8 : NOR2_X1 port map( A1 => n46, A2 => n55, ZN => next_accumulate_8_port);
   U6 : NOR2_X1 port map( A1 => n46, A2 => n53, ZN => next_accumulate_9_port);
   U52 : NOR2_X1 port map( A1 => n46, A2 => n77, ZN => next_accumulate_17_port)
                           ;
   U50 : NOR2_X1 port map( A1 => n46, A2 => n76, ZN => next_accumulate_18_port)
                           ;
   U66 : NOR2_X1 port map( A1 => n46, A2 => n84, ZN => next_accumulate_10_port)
                           ;
   U18 : NOR2_X1 port map( A1 => n46, A2 => n60, ZN => next_accumulate_3_port);
   U12 : NOR2_X1 port map( A1 => n46, A2 => n57, ZN => next_accumulate_6_port);
   U14 : NOR2_X1 port map( A1 => n46, A2 => n58, ZN => next_accumulate_5_port);
   U16 : NOR2_X1 port map( A1 => n46, A2 => n59, ZN => next_accumulate_4_port);
   U24 : NOR2_X1 port map( A1 => n46, A2 => n63, ZN => next_accumulate_2_port);
   U46 : NOR2_X1 port map( A1 => n46, A2 => n74, ZN => next_accumulate_1_port);
   U68 : NOR2_X1 port map( A1 => n46, A2 => n85, ZN => next_accumulate_0_port);
   U4 : NOR2_X1 port map( A1 => valid_port, A2 => n48, ZN => n49);
   U78 : NAND2_X1 port map( A1 => n40, A2 => enable, ZN => n86);
   U76 : NOR2_X1 port map( A1 => n93, A2 => n86, ZN => n88);
   U74 : NAND2_X1 port map( A1 => n88, A2 => n87, ZN => n91);
   U73 : OAI221_X1 port map( B1 => n37, B2 => net645046, C1 => n37, C2 => n90, 
                           A => n91, ZN => n50);
   U70 : OAI211_X1 port map( C1 => n40, C2 => enable, A => n86, B => n87, ZN =>
                           n54);
   U71 : OAI21_X1 port map( B1 => n88, B2 => n47, A => n87, ZN => n52);
   U80 : NOR3_X1 port map( A1 => n40, A2 => n47, A3 => n93, ZN => n22);
   U81 : NAND2_X1 port map( A1 => n37, A2 => net645046, ZN => n93);
   U86 : NAND3_X1 port map( A1 => n47, A2 => n92, A3 => n40, ZN => n87);
   U77 : INV_X1 port map( A => n86, ZN => n90);
   U75 : INV_X1 port map( A => n93, ZN => n92);
   U72 : INV_X1 port map( A => n87, ZN => valid_port);
   U69 : INV_X1 port map( A => ACC_from_add(0), ZN => n85);
   U47 : INV_X1 port map( A => ACC_from_add(1), ZN => n74);
   U25 : INV_X1 port map( A => ACC_from_add(2), ZN => n63);
   U15 : INV_X1 port map( A => ACC_from_add(5), ZN => n58);
   U19 : INV_X1 port map( A => ACC_from_add(3), ZN => n60);
   U13 : INV_X1 port map( A => ACC_from_add(6), ZN => n57);
   U17 : INV_X1 port map( A => ACC_from_add(4), ZN => n59);
   U11 : INV_X1 port map( A => ACC_from_add(7), ZN => n56);
   U65 : INV_X1 port map( A => ACC_from_add(11), ZN => n83);
   U67 : INV_X1 port map( A => ACC_from_add(10), ZN => n84);
   U7 : INV_X1 port map( A => ACC_from_add(9), ZN => n53);
   U9 : INV_X1 port map( A => ACC_from_add(8), ZN => n55);
   U53 : INV_X1 port map( A => ACC_from_add(17), ZN => n77);
   U49 : INV_X1 port map( A => ACC_from_add(19), ZN => n75);
   U63 : INV_X1 port map( A => ACC_from_add(12), ZN => n82);
   U51 : INV_X1 port map( A => ACC_from_add(18), ZN => n76);
   U31 : INV_X1 port map( A => ACC_from_add(27), ZN => n66);
   U39 : INV_X1 port map( A => ACC_from_add(23), ZN => n70);
   U41 : INV_X1 port map( A => ACC_from_add(22), ZN => n71);
   U3 : MUX2_X1 port map( A => A_to_add_0_port, B => ACC_from_add(0), S => n62,
                           Z => final_out(0));
   U5 : MUX2_X1 port map( A => A_to_add_2_port, B => ACC_from_add(2), S => 
                           input_mux_sel_2_port, Z => final_out(2));
   U21 : MUX2_X1 port map( A => A_to_add_27_port, B => ACC_from_add(27), S => 
                           input_mux_sel_2_port, Z => final_out(27));
   U22 : INV_X1 port map( A => ACC_from_add(16), ZN => n41);
   U23 : NOR2_X1 port map( A1 => n46, A2 => n41, ZN => next_accumulate_16_port)
                           ;
   U27 : INV_X1 port map( A => ACC_from_add(30), ZN => n42);
   U29 : NOR2_X1 port map( A1 => n46, A2 => n42, ZN => next_accumulate_30_port)
                           ;
   U33 : OR2_X2 port map( A1 => n46, A2 => input_mux_sel_2_port, ZN => 
                           reg_enable);
   U35 : AND2_X1 port map( A1 => sign, A2 => A(15), ZN => extend_vector_15_port
                           );
   U37 : BUF_X8 port map( A => n22, Z => n46);
   U43 : INV_X1 port map( A => Reset, ZN => n78);
   U45 : INV_X1 port map( A => ACC_from_add(14), ZN => n80);
   U54 : INV_X1 port map( A => ACC_from_add(21), ZN => n72);
   U55 : INV_X1 port map( A => ACC_from_add(26), ZN => n67);
   U57 : INV_X1 port map( A => ACC_from_add(20), ZN => n73);
   U59 : INV_X1 port map( A => ACC_from_add(15), ZN => n79);
   U61 : INV_X1 port map( A => ACC_from_add(13), ZN => n81);
   U79 : INV_X1 port map( A => ACC_from_add(29), ZN => n64);
   U82 : INV_X1 port map( A => ACC_from_add(25), ZN => n68);
   U83 : AND2_X1 port map( A1 => sign, A2 => B(15), ZN => enc_N2_in_2_port);
   U84 : INV_X1 port map( A => ACC_from_add(31), ZN => n61);
   U96 : INV_X1 port map( A => ACC_from_add(24), ZN => n69);
   U99 : INV_X1 port map( A => ACC_from_add(28), ZN => n65);
   U118 : BUF_X1 port map( A => input_mux_sel_2_port, Z => n62);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity sum_gen_N32_0 is

   port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic_vector 
         (8 downto 0);  S : out std_logic_vector (31 downto 0));

end sum_gen_N32_0;

architecture SYN_STRUCTURAL of sum_gen_N32_0 is

   component carry_sel_gen_N4_8
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component carry_sel_gen_N4_9
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component carry_sel_gen_N4_10
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component carry_sel_gen_N4_11
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component carry_sel_gen_N4_12
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component carry_sel_gen_N4_13
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component carry_sel_gen_N4_14
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component carry_sel_gen_N4_0_0
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal n4, net684307, net684308, net684309, net684310, net684311, net684312,
      net684313, net684314 : std_logic;

begin
   
   csel_N_0 : carry_sel_gen_N4_0_0 port map( A(3) => A(3), A(2) => A(2), A(1) 
                           => A(1), A(0) => A(0), B(3) => B(3), B(2) => B(2), 
                           B(1) => B(1), B(0) => B(0), Ci => n4, S(3) => S(3), 
                           S(2) => S(2), S(1) => S(1), S(0) => S(0), Co => 
                           net684314);
   csel_N_1 : carry_sel_gen_N4_14 port map( A(3) => A(7), A(2) => A(6), A(1) =>
                           A(5), A(0) => A(4), B(3) => B(7), B(2) => B(6), B(1)
                           => B(5), B(0) => B(4), Ci => Cin(1), S(3) => S(7), 
                           S(2) => S(6), S(1) => S(5), S(0) => S(4), Co => 
                           net684313);
   csel_N_2 : carry_sel_gen_N4_13 port map( A(3) => A(11), A(2) => A(10), A(1) 
                           => A(9), A(0) => A(8), B(3) => B(11), B(2) => B(10),
                           B(1) => B(9), B(0) => B(8), Ci => Cin(2), S(3) => 
                           S(11), S(2) => S(10), S(1) => S(9), S(0) => S(8), Co
                           => net684312);
   csel_N_3 : carry_sel_gen_N4_12 port map( A(3) => A(15), A(2) => A(14), A(1) 
                           => A(13), A(0) => A(12), B(3) => B(15), B(2) => 
                           B(14), B(1) => B(13), B(0) => B(12), Ci => Cin(3), 
                           S(3) => S(15), S(2) => S(14), S(1) => S(13), S(0) =>
                           S(12), Co => net684311);
   csel_N_4 : carry_sel_gen_N4_11 port map( A(3) => A(19), A(2) => A(18), A(1) 
                           => A(17), A(0) => A(16), B(3) => B(19), B(2) => 
                           B(18), B(1) => B(17), B(0) => B(16), Ci => Cin(4), 
                           S(3) => S(19), S(2) => S(18), S(1) => S(17), S(0) =>
                           S(16), Co => net684310);
   csel_N_5 : carry_sel_gen_N4_10 port map( A(3) => A(23), A(2) => A(22), A(1) 
                           => A(21), A(0) => A(20), B(3) => B(23), B(2) => 
                           B(22), B(1) => B(21), B(0) => B(20), Ci => Cin(5), 
                           S(3) => S(23), S(2) => S(22), S(1) => S(21), S(0) =>
                           S(20), Co => net684309);
   csel_N_6 : carry_sel_gen_N4_9 port map( A(3) => A(27), A(2) => A(26), A(1) 
                           => A(25), A(0) => A(24), B(3) => B(27), B(2) => 
                           B(26), B(1) => B(25), B(0) => B(24), Ci => Cin(6), 
                           S(3) => S(27), S(2) => S(26), S(1) => S(25), S(0) =>
                           S(24), Co => net684308);
   csel_N_7 : carry_sel_gen_N4_8 port map( A(3) => A(31), A(2) => A(30), A(1) 
                           => A(29), A(0) => A(28), B(3) => B(31), B(2) => 
                           B(30), B(1) => B(29), B(0) => B(28), Ci => Cin(7), 
                           S(3) => S(31), S(2) => S(30), S(1) => S(29), S(0) =>
                           S(28), Co => net684307);
   n4 <= '0';

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity carry_tree_N32_logN5_0 is

   port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  Cout :
         out std_logic_vector (7 downto 0));

end carry_tree_N32_logN5_0;

architecture SYN_arch of carry_tree_N32_logN5_0 is

   component pg_28
      port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic
            );
   end component;
   
   component pg_30
      port( p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic;  
            g_BAR : in std_logic);
   end component;
   
   component pg_31
      port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic
            );
   end component;
   
   component g_11
      port( g, p, g_prec : in std_logic;  g_out : out std_logic);
   end component;
   
   component g_12
      port( g, p, g_prec : in std_logic;  g_out : out std_logic);
   end component;
   
   component g_13
      port( g, p, g_prec : in std_logic;  g_out : out std_logic);
   end component;
   
   component g_14
      port( g, p, g_prec : in std_logic;  g_out : out std_logic);
   end component;
   
   component g_15
      port( g, p, g_prec : in std_logic;  g_out : out std_logic);
   end component;
   
   component g_16
      port( g, p, g_prec : in std_logic;  g_out : out std_logic);
   end component;
   
   component pg_33
      port( p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic;  
            g_BAR : in std_logic);
   end component;
   
   component pg_34
      port( g, p, g_prec, p_prec : in std_logic;  p_out, g_out_BAR : out 
            std_logic);
   end component;
   
   component pg_35
      port( p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic;  
            g_BAR : in std_logic);
   end component;
   
   component pg_36
      port( p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic;  
            g_BAR : in std_logic);
   end component;
   
   component pg_37
      port( p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic;  
            g_BAR : in std_logic);
   end component;
   
   component pg_38
      port( p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic;  
            g_BAR : in std_logic);
   end component;
   
   component g_17
      port( g, p, g_prec : in std_logic;  g_out : out std_logic);
   end component;
   
   component pg_41
      port( g, p, g_prec, p_prec : in std_logic;  p_out, g_out_BAR : out 
            std_logic);
   end component;
   
   component pg_42
      port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic
            );
   end component;
   
   component pg_43
      port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic
            );
   end component;
   
   component pg_44
      port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic
            );
   end component;
   
   component pg_45
      port( g, p, g_prec, p_prec : in std_logic;  p_out, g_out_BAR : out 
            std_logic);
   end component;
   
   component pg_46
      port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic
            );
   end component;
   
   component pg_47
      port( g, p, g_prec, p_prec : in std_logic;  p_out, g_out_BAR : out 
            std_logic);
   end component;
   
   component pg_48
      port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic
            );
   end component;
   
   component pg_49
      port( g, p, g_prec, p_prec : in std_logic;  p_out, g_out_BAR : out 
            std_logic);
   end component;
   
   component pg_50
      port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic
            );
   end component;
   
   component pg_51
      port( g, p, g_prec, p_prec : in std_logic;  p_out, g_out_BAR : out 
            std_logic);
   end component;
   
   component pg_52
      port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic
            );
   end component;
   
   component pg_0_0
      port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic
            );
   end component;
   
   component g_18
      port( g, p, g_prec : in std_logic;  g_out : out std_logic);
   end component;
   
   component g_0_0
      port( g, p, g_prec : in std_logic;  g_out : out std_logic);
   end component;
   
   component pg_net_32
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_37
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_38
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_39
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_40
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_41
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_42
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_43
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_44
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_45
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_46
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_47
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_48
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_49
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_50
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_51
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_52
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_53
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_54
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_55
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_56
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_57
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_58
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_59
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_60
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_61
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_62
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_0_0
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   signal n14, Cout_6_port, Cout_5_port, Cout_4_port, Cout_2_port, 
      p_net_27_port, p_net_26_port, p_net_25_port, p_net_24_port, p_net_23_port
      , p_net_22_port, p_net_21_port, p_net_20_port, p_net_19_port, 
      p_net_18_port, p_net_17_port, p_net_16_port, p_net_15_port, p_net_14_port
      , p_net_13_port, p_net_12_port, p_net_11_port, p_net_10_port, 
      p_net_9_port, p_net_8_port, p_net_7_port, p_net_6_port, p_net_5_port, 
      p_net_4_port, p_net_3_port, p_net_2_port, p_net_1_port, g_net_27_port, 
      g_net_26_port, g_net_25_port, g_net_24_port, g_net_23_port, g_net_22_port
      , g_net_21_port, g_net_20_port, g_net_19_port, g_net_18_port, 
      g_net_17_port, g_net_16_port, g_net_15_port, g_net_14_port, g_net_13_port
      , g_net_12_port, g_net_11_port, g_net_10_port, g_net_9_port, g_net_8_port
      , g_net_7_port, g_net_6_port, g_net_5_port, g_net_4_port, g_net_3_port, 
      g_net_2_port, g_net_1_port, g_net_0_port, magic_pro_0_port, 
      pg_1_13_1_port, pg_1_13_0_port, pg_1_12_1_port, pg_1_12_0_port, 
      pg_1_11_1_port, pg_1_11_0_port, pg_1_10_1_port, pg_1_10_0_port, 
      pg_1_9_1_port, pg_1_9_0_port, pg_1_8_1_port, pg_1_8_0_port, pg_1_7_1_port
      , pg_1_7_0_port, pg_1_6_1_port, pg_1_6_0_port, pg_1_5_1_port, 
      pg_1_5_0_port, pg_1_4_1_port, pg_1_4_0_port, pg_1_3_1_port, pg_1_3_0_port
      , pg_1_2_1_port, pg_1_2_0_port, pg_1_1_1_port, pg_1_1_0_port, 
      pg_1_0_0_port, pg_n_4_6_1_port, pg_n_4_6_0_port, pg_n_3_5_1_port, 
      pg_n_3_3_1_port, pg_n_3_3_0_port, pg_n_2_6_1_port, pg_n_2_6_0_port, 
      pg_n_2_5_1_port, pg_n_2_5_0_port, pg_n_2_4_1_port, pg_n_2_3_1_port, 
      pg_n_2_3_0_port, pg_n_2_2_1_port, pg_n_2_2_0_port, pg_n_2_1_1_port, 
      pg_n_2_1_0_port, n1, n5, Cout_0_port, n7, n8, n13, net684306, n_1175 : 
      std_logic;

begin
   Cout <= ( n_1175, Cout_6_port, Cout_5_port, Cout_4_port, n1, Cout_2_port, n8
      , Cout_0_port );
   
   pg_net_x_1 : pg_net_0_0 port map( a => A(1), b => B(1), g_out => 
                           g_net_1_port, p_out => p_net_1_port);
   pg_net_x_2 : pg_net_62 port map( a => A(2), b => B(2), g_out => g_net_2_port
                           , p_out => p_net_2_port);
   pg_net_x_3 : pg_net_61 port map( a => A(3), b => B(3), g_out => g_net_3_port
                           , p_out => p_net_3_port);
   pg_net_x_4 : pg_net_60 port map( a => A(4), b => B(4), g_out => g_net_4_port
                           , p_out => p_net_4_port);
   pg_net_x_5 : pg_net_59 port map( a => A(5), b => B(5), g_out => g_net_5_port
                           , p_out => p_net_5_port);
   pg_net_x_6 : pg_net_58 port map( a => A(6), b => B(6), g_out => g_net_6_port
                           , p_out => p_net_6_port);
   pg_net_x_7 : pg_net_57 port map( a => A(7), b => B(7), g_out => g_net_7_port
                           , p_out => p_net_7_port);
   pg_net_x_8 : pg_net_56 port map( a => A(8), b => B(8), g_out => g_net_8_port
                           , p_out => p_net_8_port);
   pg_net_x_9 : pg_net_55 port map( a => A(9), b => B(9), g_out => g_net_9_port
                           , p_out => p_net_9_port);
   pg_net_x_10 : pg_net_54 port map( a => A(10), b => B(10), g_out => 
                           g_net_10_port, p_out => p_net_10_port);
   pg_net_x_11 : pg_net_53 port map( a => A(11), b => B(11), g_out => 
                           g_net_11_port, p_out => p_net_11_port);
   pg_net_x_12 : pg_net_52 port map( a => A(12), b => B(12), g_out => 
                           g_net_12_port, p_out => p_net_12_port);
   pg_net_x_13 : pg_net_51 port map( a => A(13), b => B(13), g_out => 
                           g_net_13_port, p_out => p_net_13_port);
   pg_net_x_14 : pg_net_50 port map( a => A(14), b => B(14), g_out => 
                           g_net_14_port, p_out => p_net_14_port);
   pg_net_x_15 : pg_net_49 port map( a => A(15), b => B(15), g_out => 
                           g_net_15_port, p_out => p_net_15_port);
   pg_net_x_16 : pg_net_48 port map( a => A(16), b => B(16), g_out => 
                           g_net_16_port, p_out => p_net_16_port);
   pg_net_x_17 : pg_net_47 port map( a => A(17), b => B(17), g_out => 
                           g_net_17_port, p_out => p_net_17_port);
   pg_net_x_18 : pg_net_46 port map( a => A(18), b => B(18), g_out => 
                           g_net_18_port, p_out => p_net_18_port);
   pg_net_x_19 : pg_net_45 port map( a => A(19), b => B(19), g_out => 
                           g_net_19_port, p_out => p_net_19_port);
   pg_net_x_20 : pg_net_44 port map( a => A(20), b => B(20), g_out => 
                           g_net_20_port, p_out => p_net_20_port);
   pg_net_x_21 : pg_net_43 port map( a => A(21), b => B(21), g_out => 
                           g_net_21_port, p_out => p_net_21_port);
   pg_net_x_22 : pg_net_42 port map( a => A(22), b => B(22), g_out => 
                           g_net_22_port, p_out => p_net_22_port);
   pg_net_x_23 : pg_net_41 port map( a => A(23), b => B(23), g_out => 
                           g_net_23_port, p_out => p_net_23_port);
   pg_net_x_24 : pg_net_40 port map( a => A(24), b => B(24), g_out => 
                           g_net_24_port, p_out => p_net_24_port);
   pg_net_x_25 : pg_net_39 port map( a => A(25), b => B(25), g_out => 
                           g_net_25_port, p_out => p_net_25_port);
   pg_net_x_26 : pg_net_38 port map( a => A(26), b => B(26), g_out => 
                           g_net_26_port, p_out => p_net_26_port);
   pg_net_x_27 : pg_net_37 port map( a => A(27), b => B(27), g_out => 
                           g_net_27_port, p_out => p_net_27_port);
   pg_net_0_MAGIC : pg_net_32 port map( a => A(0), b => B(0), g_out => 
                           magic_pro_0_port, p_out => net684306);
   xG_0_0_MAGIC : g_0_0 port map( g => magic_pro_0_port, p => n13, g_prec => 
                           n14, g_out => g_net_0_port);
   xG_1_0 : g_18 port map( g => g_net_1_port, p => p_net_1_port, g_prec => 
                           g_net_0_port, g_out => pg_1_0_0_port);
   xPG_1_1 : pg_0_0 port map( g => g_net_3_port, p => p_net_3_port, g_prec => 
                           g_net_2_port, p_prec => p_net_2_port, g_out => 
                           pg_1_1_0_port, p_out => pg_1_1_1_port);
   xPG_1_2 : pg_52 port map( g => g_net_5_port, p => p_net_5_port, g_prec => 
                           g_net_4_port, p_prec => p_net_4_port, g_out => 
                           pg_1_2_0_port, p_out => pg_1_2_1_port);
   xPG_1_3 : pg_51 port map( g => g_net_7_port, p => p_net_7_port, g_prec => 
                           g_net_6_port, p_prec => p_net_6_port, p_out => 
                           pg_1_3_1_port, g_out_BAR => pg_1_3_0_port);
   xPG_1_4 : pg_50 port map( g => g_net_9_port, p => p_net_9_port, g_prec => 
                           g_net_8_port, p_prec => p_net_8_port, g_out => 
                           pg_1_4_0_port, p_out => pg_1_4_1_port);
   xPG_1_5 : pg_49 port map( g => g_net_11_port, p => p_net_11_port, g_prec => 
                           g_net_10_port, p_prec => p_net_10_port, p_out => 
                           pg_1_5_1_port, g_out_BAR => pg_1_5_0_port);
   xPG_1_6 : pg_48 port map( g => g_net_13_port, p => p_net_13_port, g_prec => 
                           g_net_12_port, p_prec => p_net_12_port, g_out => 
                           pg_1_6_0_port, p_out => pg_1_6_1_port);
   xPG_1_7 : pg_47 port map( g => g_net_15_port, p => p_net_15_port, g_prec => 
                           g_net_14_port, p_prec => p_net_14_port, p_out => 
                           pg_1_7_1_port, g_out_BAR => pg_1_7_0_port);
   xPG_1_8 : pg_46 port map( g => g_net_17_port, p => p_net_17_port, g_prec => 
                           g_net_16_port, p_prec => p_net_16_port, g_out => 
                           pg_1_8_0_port, p_out => pg_1_8_1_port);
   xPG_1_9 : pg_45 port map( g => g_net_19_port, p => p_net_19_port, g_prec => 
                           g_net_18_port, p_prec => p_net_18_port, p_out => 
                           pg_1_9_1_port, g_out_BAR => pg_1_9_0_port);
   xPG_1_10 : pg_44 port map( g => g_net_21_port, p => p_net_21_port, g_prec =>
                           g_net_20_port, p_prec => p_net_20_port, g_out => 
                           pg_1_10_0_port, p_out => pg_1_10_1_port);
   xPG_1_11 : pg_43 port map( g => g_net_23_port, p => p_net_23_port, g_prec =>
                           g_net_22_port, p_prec => p_net_22_port, g_out => 
                           pg_1_11_0_port, p_out => pg_1_11_1_port);
   xPG_1_12 : pg_42 port map( g => g_net_25_port, p => p_net_25_port, g_prec =>
                           g_net_24_port, p_prec => p_net_24_port, g_out => 
                           pg_1_12_0_port, p_out => pg_1_12_1_port);
   xPG_1_13 : pg_41 port map( g => g_net_27_port, p => p_net_27_port, g_prec =>
                           g_net_26_port, p_prec => p_net_26_port, p_out => 
                           pg_1_13_1_port, g_out_BAR => pg_1_13_0_port);
   xG_2_0 : g_17 port map( g => pg_1_1_0_port, p => pg_1_1_1_port, g_prec => 
                           pg_1_0_0_port, g_out => Cout_0_port);
   xPG_2_1 : pg_38 port map( p => pg_1_3_1_port, g_prec => pg_1_2_0_port, 
                           p_prec => pg_1_2_1_port, g_out => pg_n_2_1_0_port, 
                           p_out => pg_n_2_1_1_port, g_BAR => pg_1_3_0_port);
   xPG_2_2 : pg_37 port map( p => pg_1_5_1_port, g_prec => pg_1_4_0_port, 
                           p_prec => pg_1_4_1_port, g_out => pg_n_2_2_0_port, 
                           p_out => pg_n_2_2_1_port, g_BAR => pg_1_5_0_port);
   xPG_2_3 : pg_36 port map( p => pg_1_7_1_port, g_prec => pg_1_6_0_port, 
                           p_prec => pg_1_6_1_port, g_out => pg_n_2_3_0_port, 
                           p_out => pg_n_2_3_1_port, g_BAR => pg_1_7_0_port);
   xPG_2_4 : pg_35 port map( p => pg_1_9_1_port, g_prec => pg_1_8_0_port, 
                           p_prec => pg_1_8_1_port, g_out => n5, p_out => 
                           pg_n_2_4_1_port, g_BAR => pg_1_9_0_port);
   xPG_2_5 : pg_34 port map( g => pg_1_11_0_port, p => pg_1_11_1_port, g_prec 
                           => pg_1_10_0_port, p_prec => pg_1_10_1_port, p_out 
                           => pg_n_2_5_1_port, g_out_BAR => pg_n_2_5_0_port);
   xPG_2_6 : pg_33 port map( p => pg_1_13_1_port, g_prec => pg_1_12_0_port, 
                           p_prec => pg_1_12_1_port, g_out => pg_n_2_6_0_port, 
                           p_out => pg_n_2_6_1_port, g_BAR => pg_1_13_0_port);
   xG_3_1 : g_16 port map( g => pg_n_2_1_0_port, p => pg_n_2_1_1_port, g_prec 
                           => Cout_0_port, g_out => n8);
   xG_4_2 : g_15 port map( g => pg_n_2_2_0_port, p => pg_n_2_2_1_port, g_prec 
                           => n8, g_out => Cout_2_port);
   xG_4_3 : g_14 port map( g => pg_n_3_3_0_port, p => pg_n_3_3_1_port, g_prec 
                           => n8, g_out => n1);
   xG_5_4 : g_13 port map( g => n5, p => pg_n_2_4_1_port, g_prec => n1, g_out 
                           => Cout_4_port);
   xG_5_5 : g_12 port map( g => n7, p => pg_n_3_5_1_port, g_prec => n1, g_out 
                           => Cout_5_port);
   xG_5_6 : g_11 port map( g => pg_n_4_6_0_port, p => pg_n_4_6_1_port, g_prec 
                           => n1, g_out => Cout_6_port);
   xPG_3_3 : pg_31 port map( g => pg_n_2_3_0_port, p => pg_n_2_3_1_port, g_prec
                           => pg_n_2_2_0_port, p_prec => pg_n_2_2_1_port, g_out
                           => pg_n_3_3_0_port, p_out => pg_n_3_3_1_port);
   xPG_3_5 : pg_30 port map( p => pg_n_2_5_1_port, g_prec => n5, p_prec => 
                           pg_n_2_4_1_port, g_out => n7, p_out => 
                           pg_n_3_5_1_port, g_BAR => pg_n_2_5_0_port);
   xPG_4_6 : pg_28 port map( g => pg_n_2_6_0_port, p => pg_n_2_6_1_port, g_prec
                           => n7, p_prec => pg_n_3_5_1_port, g_out => 
                           pg_n_4_6_0_port, p_out => pg_n_4_6_1_port);
   n13 <= '0';
   n14 <= '0';

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity xor_gen_N32_0 is

   port( A : in std_logic_vector (31 downto 0);  B : in std_logic;  S : out 
         std_logic_vector (31 downto 0));

end xor_gen_N32_0;

architecture SYN_bhe of xor_gen_N32_0 is

begin
   S <= ( A(31), A(30), A(29), A(28), A(27), A(26), A(25), A(24), A(23), A(22),
      A(21), A(20), A(19), A(18), A(17), A(16), A(15), A(14), A(13), A(12), 
      A(11), A(10), A(9), A(8), A(7), A(6), A(5), A(4), A(3), A(2), A(1), A(0) 
      );

end SYN_bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity ff32_SIZE5 is

   port( D : in std_logic_vector (4 downto 0);  clk, rst : in std_logic;  Q : 
         out std_logic_vector (4 downto 0));

end ff32_SIZE5;

architecture SYN_behavioral of ff32_SIZE5 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n4, n6, n8, n10, net684301, net684302, net684303, net684304, 
      net684305 : std_logic;

begin
   
   Q_reg_4_inst : DFFR_X1 port map( D => D(4), CK => clk, RN => n10, Q => Q(4),
                           QN => net684305);
   Q_reg_3_inst : DFFR_X1 port map( D => D(3), CK => clk, RN => n10, Q => 
                           net684304, QN => n4);
   Q_reg_2_inst : DFFR_X1 port map( D => D(2), CK => clk, RN => n10, Q => 
                           net684303, QN => n6);
   Q_reg_1_inst : DFFR_X1 port map( D => D(1), CK => clk, RN => n10, Q => 
                           net684302, QN => n1);
   Q_reg_0_inst : DFFR_X1 port map( D => D(0), CK => clk, RN => n10, Q => 
                           net684301, QN => n8);
   U3 : INV_X1 port map( A => n1, ZN => Q(1));
   U4 : INV_X1 port map( A => n4, ZN => Q(3));
   U5 : INV_X1 port map( A => n6, ZN => Q(2));
   U6 : INV_X1 port map( A => rst, ZN => n10);
   U7 : INV_X1 port map( A => n8, ZN => Q(0));

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity ff32_SIZE32 is

   port( D : in std_logic_vector (31 downto 0);  clk, rst : in std_logic;  Q : 
         out std_logic_vector (31 downto 0));

end ff32_SIZE32;

architecture SYN_behavioral of ff32_SIZE32 is

   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n33, n32 : std_logic;

begin
   
   Q_reg_31_inst : DFFR_X1 port map( D => D(31), CK => clk, RN => n32, Q => 
                           Q(31), QN => n33);
   Q_reg_30_inst : DFFR_X1 port map( D => D(30), CK => clk, RN => n32, Q => 
                           Q(30), QN => n31);
   Q_reg_29_inst : DFFR_X1 port map( D => D(29), CK => clk, RN => n32, Q => 
                           Q(29), QN => n30);
   Q_reg_28_inst : DFFR_X1 port map( D => D(28), CK => clk, RN => n32, Q => 
                           Q(28), QN => n29);
   Q_reg_27_inst : DFFR_X1 port map( D => D(27), CK => clk, RN => n32, Q => 
                           Q(27), QN => n28);
   Q_reg_26_inst : DFFR_X1 port map( D => D(26), CK => clk, RN => n32, Q => 
                           Q(26), QN => n27);
   Q_reg_25_inst : DFFR_X1 port map( D => D(25), CK => clk, RN => n32, Q => 
                           Q(25), QN => n26);
   Q_reg_24_inst : DFFR_X1 port map( D => D(24), CK => clk, RN => n32, Q => 
                           Q(24), QN => n25);
   Q_reg_23_inst : DFFR_X1 port map( D => D(23), CK => clk, RN => n32, Q => 
                           Q(23), QN => n24);
   Q_reg_22_inst : DFFR_X1 port map( D => D(22), CK => clk, RN => n32, Q => 
                           Q(22), QN => n23);
   Q_reg_21_inst : DFFR_X1 port map( D => D(21), CK => clk, RN => n32, Q => 
                           Q(21), QN => n22);
   Q_reg_20_inst : DFFR_X1 port map( D => D(20), CK => clk, RN => n32, Q => 
                           Q(20), QN => n21);
   Q_reg_19_inst : DFFR_X1 port map( D => D(19), CK => clk, RN => n32, Q => 
                           Q(19), QN => n20);
   Q_reg_18_inst : DFFR_X1 port map( D => D(18), CK => clk, RN => n32, Q => 
                           Q(18), QN => n19);
   Q_reg_17_inst : DFFR_X1 port map( D => D(17), CK => clk, RN => n32, Q => 
                           Q(17), QN => n18);
   Q_reg_16_inst : DFFR_X1 port map( D => D(16), CK => clk, RN => n32, Q => 
                           Q(16), QN => n17);
   Q_reg_15_inst : DFFR_X1 port map( D => D(15), CK => clk, RN => n32, Q => 
                           Q(15), QN => n16);
   Q_reg_14_inst : DFFR_X1 port map( D => D(14), CK => clk, RN => n32, Q => 
                           Q(14), QN => n15);
   Q_reg_13_inst : DFFR_X1 port map( D => D(13), CK => clk, RN => n32, Q => 
                           Q(13), QN => n14);
   Q_reg_12_inst : DFFR_X1 port map( D => D(12), CK => clk, RN => n32, Q => 
                           Q(12), QN => n13);
   Q_reg_11_inst : DFFR_X1 port map( D => D(11), CK => clk, RN => n32, Q => 
                           Q(11), QN => n12);
   Q_reg_10_inst : DFFR_X1 port map( D => D(10), CK => clk, RN => n32, Q => 
                           Q(10), QN => n11);
   Q_reg_9_inst : DFFR_X1 port map( D => D(9), CK => clk, RN => n32, Q => Q(9),
                           QN => n10);
   Q_reg_8_inst : DFFR_X1 port map( D => D(8), CK => clk, RN => n32, Q => Q(8),
                           QN => n9);
   Q_reg_7_inst : DFFR_X1 port map( D => D(7), CK => clk, RN => n32, Q => Q(7),
                           QN => n8);
   Q_reg_6_inst : DFFR_X1 port map( D => D(6), CK => clk, RN => n32, Q => Q(6),
                           QN => n7);
   Q_reg_5_inst : DFFR_X1 port map( D => D(5), CK => clk, RN => n32, Q => Q(5),
                           QN => n6);
   Q_reg_4_inst : DFFR_X1 port map( D => D(4), CK => clk, RN => n32, Q => Q(4),
                           QN => n5);
   Q_reg_3_inst : DFFR_X1 port map( D => D(3), CK => clk, RN => n32, Q => Q(3),
                           QN => n4);
   Q_reg_2_inst : DFFR_X1 port map( D => D(2), CK => clk, RN => n32, Q => Q(2),
                           QN => n3);
   Q_reg_1_inst : DFFR_X1 port map( D => D(1), CK => clk, RN => n32, Q => Q(1),
                           QN => n2);
   Q_reg_0_inst : DFFR_X1 port map( D => D(0), CK => clk, RN => n32, Q => Q(0),
                           QN => n1);
   U3 : INV_X2 port map( A => rst, ZN => n32);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity mux41_MUX_SIZE32_1 is

   port( IN0, IN1, IN2, IN3 : in std_logic_vector (31 downto 0);  CTRL : in 
         std_logic_vector (1 downto 0);  OUT1 : out std_logic_vector (31 downto
         0));

end mux41_MUX_SIZE32_1;

architecture SYN_bhe of mux41_MUX_SIZE32_1 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n35, n36, n38, n39, n40, n42, n44, n45, n47, n48, n49, n50, n51, n52,
      n53, n54, n55, n56, n58, n61, n65, n66, n67, n37, n69, n186, n187, n188, 
      n189, n190, n191, n192, n194, n195, n196, n197, n199, n202, n203, n204, 
      n205, n206, n207, n210, n211, n212, n213, n214, n215, n216, n217, n218, 
      n220, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, 
      n234, n235, n236 : std_logic;

begin
   
   U23 : INV_X1 port map( A => n48, ZN => OUT1(28));
   U31 : INV_X1 port map( A => n52, ZN => OUT1(24));
   U25 : INV_X1 port map( A => n49, ZN => OUT1(27));
   U21 : INV_X1 port map( A => n47, ZN => OUT1(29));
   U15 : INV_X1 port map( A => n44, ZN => OUT1(31));
   U17 : INV_X1 port map( A => n45, ZN => OUT1(30));
   U39 : INV_X1 port map( A => n56, ZN => OUT1(20));
   U1 : BUF_X2 port map( A => n35, Z => n234);
   U2 : BUF_X2 port map( A => n36, Z => n233);
   U3 : BUF_X2 port map( A => n36, Z => n231);
   U4 : OR3_X1 port map( A1 => n205, A2 => n206, A3 => n207, ZN => OUT1(2));
   U5 : OR3_X1 port map( A1 => n225, A2 => n224, A3 => n223, ZN => OUT1(13));
   U6 : NAND2_X1 port map( A1 => IN1(3), A2 => n233, ZN => n186);
   U7 : AOI21_X1 port map( B1 => n236, B2 => IN0(3), A => n220, ZN => n187);
   U8 : NAND2_X1 port map( A1 => n186, A2 => n187, ZN => OUT1(3));
   U9 : NAND2_X1 port map( A1 => IN2(15), A2 => n229, ZN => n188);
   U10 : AOI21_X1 port map( B1 => n234, B2 => IN0(15), A => n194, ZN => n189);
   U11 : NAND2_X1 port map( A1 => n188, A2 => n189, ZN => OUT1(15));
   U12 : NAND2_X1 port map( A1 => IN1(17), A2 => n231, ZN => n190);
   U13 : AOI21_X1 port map( B1 => n234, B2 => IN0(17), A => n199, ZN => n191);
   U14 : NAND2_X1 port map( A1 => n190, A2 => n191, ZN => OUT1(17));
   U16 : NAND2_X1 port map( A1 => IN0(18), A2 => n234, ZN => n192);
   U18 : NAND3_X1 port map( A1 => n192, A2 => n196, A3 => n197, ZN => OUT1(18))
                           ;
   U19 : BUF_X2 port map( A => n36, Z => n232);
   U20 : BUF_X2 port map( A => n37, Z => n230);
   U22 : AND2_X1 port map( A1 => n231, A2 => IN1(15), ZN => n194);
   U24 : BUF_X2 port map( A => n37, Z => n195);
   U26 : NAND2_X1 port map( A1 => n231, A2 => IN1(18), ZN => n196);
   U27 : NAND2_X1 port map( A1 => n195, A2 => IN2(18), ZN => n197);
   U28 : BUF_X1 port map( A => n37, Z => n229);
   U29 : BUF_X1 port map( A => n37, Z => n210);
   U30 : AND2_X1 port map( A1 => n210, A2 => IN2(17), ZN => n199);
   U32 : NAND3_X1 port map( A1 => n202, A2 => n203, A3 => n204, ZN => OUT1(14))
                           ;
   U33 : BUF_X1 port map( A => n35, Z => n235);
   U34 : INV_X1 port map( A => n50, ZN => OUT1(26));
   U35 : AND2_X1 port map( A1 => n234, A2 => IN0(13), ZN => n223);
   U36 : BUF_X1 port map( A => n35, Z => n236);
   U37 : INV_X1 port map( A => n61, ZN => OUT1(16));
   U38 : INV_X1 port map( A => n55, ZN => OUT1(21));
   U40 : INV_X1 port map( A => n53, ZN => OUT1(23));
   U41 : INV_X1 port map( A => n58, ZN => OUT1(19));
   U42 : INV_X1 port map( A => n54, ZN => OUT1(22));
   U43 : INV_X1 port map( A => n66, ZN => OUT1(11));
   U44 : AND2_X1 port map( A1 => n233, A2 => IN1(13), ZN => n224);
   U45 : NAND2_X1 port map( A1 => n234, A2 => IN0(14), ZN => n202);
   U46 : NAND2_X1 port map( A1 => n233, A2 => IN1(14), ZN => n203);
   U47 : NAND2_X1 port map( A1 => n230, A2 => IN2(14), ZN => n204);
   U48 : AND2_X1 port map( A1 => n235, A2 => IN0(2), ZN => n205);
   U49 : AND2_X1 port map( A1 => n232, A2 => IN1(2), ZN => n206);
   U50 : AND2_X1 port map( A1 => n229, A2 => IN2(2), ZN => n207);
   U51 : INV_X1 port map( A => n39, ZN => OUT1(7));
   U52 : INV_X1 port map( A => n51, ZN => OUT1(25));
   U53 : AND2_X1 port map( A1 => n69, A2 => CTRL(0), ZN => n36);
   U54 : INV_X1 port map( A => n38, ZN => OUT1(8));
   U55 : INV_X1 port map( A => n65, ZN => OUT1(12));
   U56 : INV_X1 port map( A => n67, ZN => OUT1(10));
   U57 : NOR2_X1 port map( A1 => n69, A2 => CTRL(0), ZN => n37);
   U58 : INV_X1 port map( A => n40, ZN => OUT1(6));
   U59 : INV_X1 port map( A => n42, ZN => OUT1(4));
   U60 : AND2_X1 port map( A1 => n210, A2 => IN2(13), ZN => n225);
   U61 : AND2_X1 port map( A1 => n210, A2 => IN2(3), ZN => n220);
   U62 : NAND3_X1 port map( A1 => n227, A2 => n226, A3 => n228, ZN => OUT1(9));
   U63 : INV_X1 port map( A => CTRL(1), ZN => n69);
   U64 : NAND2_X1 port map( A1 => n230, A2 => IN2(5), ZN => n211);
   U65 : NAND2_X1 port map( A1 => n195, A2 => IN2(0), ZN => n216);
   U66 : AOI222_X1 port map( A1 => n235, A2 => IN0(30), B1 => n233, B2 => 
                           IN1(30), C1 => n210, C2 => IN2(30), ZN => n45);
   U67 : AOI222_X1 port map( A1 => n235, A2 => IN0(22), B1 => n233, B2 => 
                           IN1(22), C1 => n210, C2 => IN2(22), ZN => n54);
   U68 : AOI222_X1 port map( A1 => n234, A2 => IN0(16), B1 => n233, B2 => 
                           IN1(16), C1 => n210, C2 => IN2(16), ZN => n61);
   U69 : AOI222_X1 port map( A1 => n235, A2 => IN0(26), B1 => n231, B2 => 
                           IN1(26), C1 => n195, C2 => IN2(26), ZN => n50);
   U70 : NAND2_X1 port map( A1 => n230, A2 => IN2(9), ZN => n228);
   U71 : AOI222_X1 port map( A1 => n235, A2 => IN0(25), B1 => n231, B2 => 
                           IN1(25), C1 => n230, C2 => IN2(25), ZN => n51);
   U72 : AOI222_X1 port map( A1 => n236, A2 => IN0(6), B1 => n232, B2 => IN1(6)
                           , C1 => n210, C2 => IN2(6), ZN => n40);
   U73 : AOI222_X1 port map( A1 => n236, A2 => IN0(7), B1 => n232, B2 => IN1(7)
                           , C1 => n195, C2 => IN2(7), ZN => n39);
   U74 : NAND3_X1 port map( A1 => n216, A2 => n215, A3 => n214, ZN => OUT1(0));
   U75 : NAND3_X1 port map( A1 => n212, A2 => n211, A3 => n213, ZN => OUT1(5));
   U76 : NAND2_X1 port map( A1 => n232, A2 => IN1(5), ZN => n212);
   U77 : NAND2_X1 port map( A1 => n236, A2 => IN0(5), ZN => n213);
   U78 : NAND2_X1 port map( A1 => n234, A2 => IN0(0), ZN => n214);
   U79 : NAND2_X1 port map( A1 => n232, A2 => IN1(0), ZN => n215);
   U80 : NAND2_X1 port map( A1 => n195, A2 => IN2(1), ZN => n217);
   U81 : NAND2_X1 port map( A1 => n217, A2 => n218, ZN => OUT1(1));
   U82 : AOI22_X1 port map( A1 => n231, A2 => IN1(1), B1 => n234, B2 => IN0(1),
                           ZN => n218);
   U83 : AOI222_X1 port map( A1 => n236, A2 => IN0(31), B1 => n231, B2 => 
                           IN1(31), C1 => n230, C2 => IN2(31), ZN => n44);
   U84 : AOI222_X1 port map( A1 => n236, A2 => IN0(4), B1 => n232, B2 => IN1(4)
                           , C1 => n230, C2 => IN2(4), ZN => n42);
   U85 : AOI222_X1 port map( A1 => n236, A2 => IN0(8), B1 => n233, B2 => IN1(8)
                           , C1 => n229, C2 => IN2(8), ZN => n38);
   U86 : AOI222_X1 port map( A1 => n235, A2 => IN0(24), B1 => n232, B2 => 
                           IN1(24), C1 => n230, C2 => IN2(24), ZN => n52);
   U87 : NAND2_X1 port map( A1 => n236, A2 => IN0(9), ZN => n226);
   U88 : NAND2_X1 port map( A1 => n233, A2 => IN1(9), ZN => n227);
   U89 : AOI222_X1 port map( A1 => n235, A2 => IN0(20), B1 => n232, B2 => 
                           IN1(20), C1 => n229, C2 => IN2(20), ZN => n56);
   U90 : AOI222_X1 port map( A1 => n235, A2 => IN0(28), B1 => n233, B2 => 
                           IN1(28), C1 => n210, C2 => IN2(28), ZN => n48);
   U91 : AOI222_X1 port map( A1 => n235, A2 => IN0(29), B1 => n232, B2 => 
                           IN1(29), C1 => n195, C2 => IN2(29), ZN => n47);
   U92 : AOI222_X1 port map( A1 => n235, A2 => IN0(23), B1 => n231, B2 => 
                           IN1(23), C1 => n230, C2 => IN2(23), ZN => n53);
   U93 : AOI222_X1 port map( A1 => n235, A2 => IN0(27), B1 => n232, B2 => 
                           IN1(27), C1 => n229, C2 => IN2(27), ZN => n49);
   U94 : AOI222_X1 port map( A1 => n235, A2 => IN0(21), B1 => n231, B2 => 
                           IN1(21), C1 => n210, C2 => IN2(21), ZN => n55);
   U95 : AOI222_X1 port map( A1 => n234, A2 => IN0(19), B1 => n233, B2 => 
                           IN1(19), C1 => n230, C2 => IN2(19), ZN => n58);
   U96 : AOI222_X1 port map( A1 => n234, A2 => IN0(12), B1 => n231, B2 => 
                           IN1(12), C1 => n229, C2 => IN2(12), ZN => n65);
   U97 : AOI222_X1 port map( A1 => n234, A2 => IN0(11), B1 => n233, B2 => 
                           IN1(11), C1 => n230, C2 => IN2(11), ZN => n66);
   U98 : AOI222_X1 port map( A1 => n234, A2 => IN0(10), B1 => n231, B2 => 
                           IN1(10), C1 => n230, C2 => IN2(10), ZN => n67);
   U99 : NOR2_X1 port map( A1 => CTRL(0), A2 => CTRL(1), ZN => n35);

end SYN_bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity mux41_MUX_SIZE32_0 is

   port( IN0, IN1, IN2, IN3 : in std_logic_vector (31 downto 0);  CTRL : in 
         std_logic_vector (1 downto 0);  OUT1 : out std_logic_vector (31 downto
         0));

end mux41_MUX_SIZE32_0;

architecture SYN_bhe of mux41_MUX_SIZE32_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
      n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62
      , n63, n64, n65, n66, n67, n69, n114, n116, n117, n118, n119, n120, n121,
      n122, n123 : std_logic;

begin
   
   U18 : AOI222_X1 port map( A1 => n122, A2 => IN2(30), B1 => n114, B2 => 
                           IN0(30), C1 => n120, C2 => IN1(30), ZN => n45);
   U22 : AOI222_X1 port map( A1 => n122, A2 => IN2(29), B1 => n114, B2 => 
                           IN0(29), C1 => n120, C2 => IN1(29), ZN => n47);
   U24 : AOI222_X1 port map( A1 => n123, A2 => IN2(28), B1 => n114, B2 => 
                           IN0(28), C1 => n120, C2 => IN1(28), ZN => n48);
   U16 : AOI222_X1 port map( A1 => n123, A2 => IN2(31), B1 => n114, B2 => 
                           IN0(31), C1 => n119, C2 => IN1(31), ZN => n44);
   U42 : AOI222_X1 port map( A1 => n35, A2 => IN2(1), B1 => n121, B2 => IN0(1),
                           C1 => n119, C2 => IN1(1), ZN => n57);
   U20 : AOI222_X1 port map( A1 => n35, A2 => IN2(2), B1 => n114, B2 => IN0(2),
                           C1 => n119, C2 => IN1(2), ZN => n46);
   U14 : AOI222_X1 port map( A1 => n122, A2 => IN2(3), B1 => n114, B2 => IN0(3)
                           , C1 => n120, C2 => IN1(3), ZN => n43);
   U8 : AOI222_X1 port map( A1 => n123, A2 => IN2(6), B1 => n114, B2 => IN0(6),
                           C1 => n119, C2 => IN1(6), ZN => n40);
   U6 : AOI222_X1 port map( A1 => n122, A2 => IN2(7), B1 => n114, B2 => IN0(7),
                           C1 => n120, C2 => IN1(7), ZN => n39);
   U10 : AOI222_X1 port map( A1 => n123, A2 => IN2(5), B1 => n114, B2 => IN0(5)
                           , C1 => n119, C2 => IN1(5), ZN => n41);
   U12 : AOI222_X1 port map( A1 => n122, A2 => IN2(4), B1 => n114, B2 => IN0(4)
                           , C1 => n120, C2 => IN1(4), ZN => n42);
   U56 : AOI222_X1 port map( A1 => n122, A2 => IN2(13), B1 => n121, B2 => 
                           IN0(13), C1 => n119, C2 => IN1(13), ZN => n64);
   U62 : AOI222_X1 port map( A1 => n122, A2 => IN2(10), B1 => n121, B2 => 
                           IN0(10), C1 => n119, C2 => IN1(10), ZN => n67);
   U2 : AOI222_X1 port map( A1 => n123, A2 => IN2(9), B1 => n114, B2 => IN0(9),
                           C1 => n119, C2 => IN1(9), ZN => n34);
   U4 : AOI222_X1 port map( A1 => n123, A2 => IN2(8), B1 => n114, B2 => IN0(8),
                           C1 => n120, C2 => IN1(8), ZN => n38);
   U26 : AOI222_X1 port map( A1 => n123, A2 => IN2(27), B1 => n114, B2 => 
                           IN0(27), C1 => n120, C2 => IN1(27), ZN => n49);
   U28 : AOI222_X1 port map( A1 => n122, A2 => IN2(26), B1 => n114, B2 => 
                           IN0(26), C1 => n120, C2 => IN1(26), ZN => n50);
   U30 : AOI222_X1 port map( A1 => n122, A2 => IN2(25), B1 => n114, B2 => 
                           IN0(25), C1 => n120, C2 => IN1(25), ZN => n51);
   U32 : AOI222_X1 port map( A1 => n123, A2 => IN2(24), B1 => n114, B2 => 
                           IN0(24), C1 => n119, C2 => IN1(24), ZN => n52);
   U38 : AOI222_X1 port map( A1 => n122, A2 => IN2(21), B1 => n114, B2 => 
                           IN0(21), C1 => n120, C2 => IN1(21), ZN => n55);
   U40 : AOI222_X1 port map( A1 => n123, A2 => IN2(20), B1 => n114, B2 => 
                           IN0(20), C1 => n119, C2 => IN1(20), ZN => n56);
   U34 : AOI222_X1 port map( A1 => n123, A2 => IN2(23), B1 => n114, B2 => 
                           IN0(23), C1 => n120, C2 => IN1(23), ZN => n53);
   U36 : AOI222_X1 port map( A1 => n122, A2 => IN2(22), B1 => n114, B2 => 
                           IN0(22), C1 => n120, C2 => IN1(22), ZN => n54);
   U46 : AOI222_X1 port map( A1 => n123, A2 => IN2(18), B1 => n121, B2 => 
                           IN0(18), C1 => n120, C2 => IN1(18), ZN => n59);
   U48 : AOI222_X1 port map( A1 => n123, A2 => IN2(17), B1 => n121, B2 => 
                           IN0(17), C1 => n120, C2 => IN1(17), ZN => n60);
   U67 : AND2_X1 port map( A1 => CTRL(1), A2 => n69, ZN => n35);
   U57 : INV_X1 port map( A => n65, ZN => OUT1(12));
   U49 : INV_X1 port map( A => n61, ZN => OUT1(16));
   U53 : INV_X1 port map( A => n63, ZN => OUT1(14));
   U47 : INV_X1 port map( A => n60, ZN => OUT1(17));
   U51 : INV_X1 port map( A => n62, ZN => OUT1(15));
   U45 : INV_X1 port map( A => n59, ZN => OUT1(18));
   U55 : INV_X1 port map( A => n64, ZN => OUT1(13));
   U11 : INV_X1 port map( A => n42, ZN => OUT1(4));
   U15 : INV_X1 port map( A => n44, ZN => OUT1(31));
   U17 : INV_X1 port map( A => n45, ZN => OUT1(30));
   U21 : INV_X1 port map( A => n47, ZN => OUT1(29));
   U23 : INV_X1 port map( A => n48, ZN => OUT1(28));
   U5 : INV_X1 port map( A => n39, ZN => OUT1(7));
   U25 : INV_X1 port map( A => n49, ZN => OUT1(27));
   U3 : INV_X1 port map( A => n38, ZN => OUT1(8));
   U27 : INV_X1 port map( A => n50, ZN => OUT1(26));
   U1 : INV_X1 port map( A => n34, ZN => OUT1(9));
   U29 : INV_X1 port map( A => n51, ZN => OUT1(25));
   U31 : INV_X1 port map( A => n52, ZN => OUT1(24));
   U33 : INV_X1 port map( A => n53, ZN => OUT1(23));
   U35 : INV_X1 port map( A => n54, ZN => OUT1(22));
   U37 : INV_X1 port map( A => n55, ZN => OUT1(21));
   U7 : INV_X1 port map( A => n40, ZN => OUT1(6));
   U39 : INV_X1 port map( A => n56, ZN => OUT1(20));
   U43 : INV_X1 port map( A => n58, ZN => OUT1(19));
   U61 : INV_X1 port map( A => n67, ZN => OUT1(10));
   U59 : INV_X1 port map( A => n66, ZN => OUT1(11));
   U9 : BUF_X2 port map( A => n37, Z => n120);
   U13 : BUF_X2 port map( A => n37, Z => n119);
   U19 : BUF_X2 port map( A => n35, Z => n123);
   U41 : BUF_X1 port map( A => n35, Z => n122);
   U44 : BUF_X1 port map( A => n36, Z => n121);
   U50 : BUF_X2 port map( A => n36, Z => n114);
   U52 : AND2_X1 port map( A1 => n119, A2 => IN1(0), ZN => n117);
   U54 : INV_X1 port map( A => n43, ZN => OUT1(3));
   U58 : INV_X1 port map( A => n57, ZN => OUT1(1));
   U60 : INV_X1 port map( A => n46, ZN => OUT1(2));
   U63 : INV_X1 port map( A => n41, ZN => OUT1(5));
   U64 : AOI222_X1 port map( A1 => n123, A2 => IN2(11), B1 => n121, B2 => 
                           IN0(11), C1 => n120, C2 => IN1(11), ZN => n66);
   U65 : AOI222_X1 port map( A1 => n123, A2 => IN2(12), B1 => n121, B2 => 
                           IN0(12), C1 => n120, C2 => IN1(12), ZN => n65);
   U66 : AOI222_X1 port map( A1 => n123, A2 => IN2(19), B1 => n121, B2 => 
                           IN0(19), C1 => n120, C2 => IN1(19), ZN => n58);
   U68 : AOI222_X1 port map( A1 => n122, A2 => IN2(14), B1 => n121, B2 => 
                           IN0(14), C1 => n120, C2 => IN1(14), ZN => n63);
   U69 : AOI222_X1 port map( A1 => n122, A2 => IN2(15), B1 => n121, B2 => 
                           IN0(15), C1 => n120, C2 => IN1(15), ZN => n62);
   U70 : AOI222_X1 port map( A1 => n122, A2 => IN2(16), B1 => n121, B2 => 
                           IN0(16), C1 => n120, C2 => IN1(16), ZN => n61);
   U71 : AND2_X1 port map( A1 => n121, A2 => IN0(0), ZN => n118);
   U72 : AND2_X1 port map( A1 => n35, A2 => IN2(0), ZN => n116);
   U73 : OR3_X2 port map( A1 => n118, A2 => n117, A3 => n116, ZN => OUT1(0));
   U74 : NOR2_X1 port map( A1 => CTRL(1), A2 => CTRL(0), ZN => n36);
   U75 : NOR2_X1 port map( A1 => CTRL(1), A2 => n69, ZN => n37);
   U76 : INV_X1 port map( A => CTRL(0), ZN => n69);

end SYN_bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity mux41_MUX_SIZE5 is

   port( IN0, IN1, IN2, IN3 : in std_logic_vector (4 downto 0);  CTRL : in 
         std_logic_vector (1 downto 0);  OUT1 : out std_logic_vector (4 downto 
         0));

end mux41_MUX_SIZE5;

architecture SYN_bhe of mux41_MUX_SIZE5 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6 : std_logic;

begin
   
   U6 : AOI22_X1 port map( A1 => CTRL(0), A2 => IN1(2), B1 => CTRL(1), B2 => 
                           IN2(2), ZN => n4);
   U8 : AOI22_X1 port map( A1 => CTRL(0), A2 => IN1(1), B1 => CTRL(1), B2 => 
                           IN2(1), ZN => n5);
   U4 : AOI22_X1 port map( A1 => CTRL(0), A2 => IN1(3), B1 => CTRL(1), B2 => 
                           IN2(3), ZN => n3);
   U2 : AOI22_X1 port map( A1 => CTRL(0), A2 => IN1(4), B1 => CTRL(1), B2 => 
                           IN2(4), ZN => n1);
   U11 : AOI22_X1 port map( A1 => CTRL(0), A2 => IN1(0), B1 => CTRL(1), B2 => 
                           IN2(0), ZN => n6);
   U9 : NAND2_X1 port map( A1 => n6, A2 => n2, ZN => OUT1(0));
   U3 : NAND2_X1 port map( A1 => n3, A2 => n2, ZN => OUT1(3));
   U1 : NAND2_X1 port map( A1 => n1, A2 => n2, ZN => OUT1(4));
   U5 : NAND2_X1 port map( A1 => n4, A2 => n2, ZN => OUT1(2));
   U7 : NAND2_X1 port map( A1 => n5, A2 => n2, ZN => OUT1(1));
   U10 : NAND2_X1 port map( A1 => CTRL(0), A2 => CTRL(1), ZN => n2);

end SYN_bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity real_alu_DATA_SIZE32 is

   port( IN1, IN2 : in std_logic_vector (31 downto 0);  ALUW_i : in 
         std_logic_vector (12 downto 0);  DOUT : out std_logic_vector (31 
         downto 0);  stall_o : out std_logic;  Clock, Reset : in std_logic);

end real_alu_DATA_SIZE32;

architecture SYN_Bhe of real_alu_DATA_SIZE32 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X2
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X3
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component logic_unit_SIZE32
      port( IN1, IN2 : in std_logic_vector (31 downto 0);  CTRL : in 
            std_logic_vector (1 downto 0);  OUT1 : out std_logic_vector (31 
            downto 0));
   end component;
   
   component shifter
      port( A : in std_logic_vector (31 downto 0);  B : in std_logic_vector (4 
            downto 0);  LOGIC_ARITH, LEFT_RIGHT : in std_logic;  OUTPUT : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component comparator_M32
      port( C, V : in std_logic;  SUM : in std_logic_vector (31 downto 0);  sel
            : in std_logic_vector (2 downto 0);  sign : in std_logic;  S : out 
            std_logic);
   end component;
   
   component p4add_N32_logN5_1
      port( A, B : in std_logic_vector (31 downto 0);  Cin, sign : in std_logic
            ;  S : out std_logic_vector (31 downto 0);  Cout : out std_logic);
   end component;
   
   component simple_booth_add_ext_N16
      port( Clock, Reset, sign, enable : in std_logic;  valid : out std_logic; 
            A, B : in std_logic_vector (15 downto 0);  A_to_add, B_to_add : out
            std_logic_vector (31 downto 0);  sign_to_add : out std_logic;  
            final_out : out std_logic_vector (31 downto 0);  ACC_from_add : in 
            std_logic_vector (31 downto 0));
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal X_Logic0_port, mux_A_31_port, mux_A_30_port, mux_A_29_port, 
      mux_A_28_port, mux_A_27_port, mux_A_26_port, mux_A_25_port, mux_A_24_port
      , mux_A_23_port, mux_A_22_port, mux_A_21_port, mux_A_20_port, 
      mux_A_19_port, mux_A_18_port, mux_A_17_port, mux_A_16_port, mux_A_15_port
      , mux_A_14_port, mux_A_13_port, mux_A_12_port, mux_A_11_port, 
      mux_A_10_port, mux_A_9_port, mux_A_8_port, mux_A_7_port, mux_A_6_port, 
      mux_A_5_port, mux_A_4_port, mux_A_3_port, mux_A_2_port, mux_A_1_port, 
      mux_A_0_port, A_booth_to_add_31_port, A_booth_to_add_30_port, 
      A_booth_to_add_29_port, A_booth_to_add_28_port, A_booth_to_add_27_port, 
      A_booth_to_add_26_port, A_booth_to_add_25_port, A_booth_to_add_24_port, 
      A_booth_to_add_23_port, A_booth_to_add_22_port, A_booth_to_add_21_port, 
      A_booth_to_add_20_port, A_booth_to_add_19_port, A_booth_to_add_18_port, 
      A_booth_to_add_17_port, A_booth_to_add_16_port, A_booth_to_add_15_port, 
      A_booth_to_add_14_port, A_booth_to_add_13_port, A_booth_to_add_12_port, 
      A_booth_to_add_11_port, A_booth_to_add_10_port, A_booth_to_add_9_port, 
      A_booth_to_add_8_port, A_booth_to_add_7_port, A_booth_to_add_6_port, 
      A_booth_to_add_5_port, A_booth_to_add_4_port, A_booth_to_add_3_port, 
      A_booth_to_add_2_port, A_booth_to_add_1_port, A_booth_to_add_0_port, 
      mux_B_31_port, mux_B_30_port, mux_B_29_port, mux_B_28_port, mux_B_27_port
      , mux_B_26_port, mux_B_25_port, mux_B_24_port, mux_B_23_port, 
      mux_B_22_port, mux_B_21_port, mux_B_20_port, mux_B_19_port, mux_B_18_port
      , mux_B_17_port, mux_B_16_port, mux_B_15_port, mux_B_14_port, 
      mux_B_13_port, mux_B_12_port, mux_B_11_port, mux_B_10_port, mux_B_9_port,
      mux_B_8_port, mux_B_7_port, mux_B_6_port, mux_B_5_port, mux_B_4_port, 
      mux_B_3_port, mux_B_2_port, mux_B_1_port, mux_B_0_port, 
      B_booth_to_add_31_port, B_booth_to_add_30_port, B_booth_to_add_29_port, 
      B_booth_to_add_28_port, B_booth_to_add_27_port, B_booth_to_add_26_port, 
      B_booth_to_add_25_port, B_booth_to_add_24_port, B_booth_to_add_23_port, 
      B_booth_to_add_22_port, B_booth_to_add_21_port, B_booth_to_add_20_port, 
      B_booth_to_add_19_port, B_booth_to_add_18_port, B_booth_to_add_17_port, 
      B_booth_to_add_16_port, B_booth_to_add_15_port, B_booth_to_add_14_port, 
      B_booth_to_add_13_port, B_booth_to_add_12_port, B_booth_to_add_11_port, 
      B_booth_to_add_10_port, B_booth_to_add_9_port, B_booth_to_add_8_port, 
      B_booth_to_add_7_port, B_booth_to_add_6_port, B_booth_to_add_5_port, 
      B_booth_to_add_4_port, B_booth_to_add_3_port, B_booth_to_add_2_port, 
      B_booth_to_add_1_port, B_booth_to_add_0_port, mux_sign, sign_booth_to_add
      , valid_from_booth, mult_out_31_port, mult_out_30_port, mult_out_29_port,
      mult_out_28_port, mult_out_27_port, mult_out_26_port, mult_out_25_port, 
      mult_out_24_port, mult_out_23_port, mult_out_22_port, mult_out_21_port, 
      mult_out_20_port, mult_out_19_port, mult_out_18_port, mult_out_17_port, 
      mult_out_16_port, mult_out_15_port, mult_out_14_port, mult_out_13_port, 
      mult_out_12_port, mult_out_11_port, mult_out_10_port, mult_out_9_port, 
      mult_out_8_port, mult_out_7_port, mult_out_6_port, mult_out_5_port, 
      mult_out_4_port, mult_out_3_port, mult_out_2_port, mult_out_1_port, 
      mult_out_0_port, sum_out_30_port, sum_out_27_port, sum_out_26_port, 
      sum_out_23_port, sum_out_18_port, sum_out_17_port, sum_out_16_port, 
      sum_out_15_port, sum_out_14_port, sum_out_13_port, sum_out_12_port, 
      sum_out_11_port, sum_out_10_port, sum_out_9_port, sum_out_8_port, 
      sum_out_7_port, sum_out_6_port, sum_out_5_port, sum_out_4_port, 
      sum_out_3_port, sum_out_2_port, sum_out_1_port, sum_out_0_port, 
      carry_from_adder, overflow, comp_out, shift_out_31_port, 
      shift_out_30_port, shift_out_29_port, shift_out_28_port, 
      shift_out_27_port, shift_out_26_port, shift_out_25_port, 
      shift_out_24_port, shift_out_23_port, shift_out_22_port, 
      shift_out_21_port, shift_out_20_port, shift_out_19_port, 
      shift_out_18_port, shift_out_17_port, shift_out_16_port, 
      shift_out_15_port, shift_out_14_port, shift_out_13_port, 
      shift_out_12_port, shift_out_11_port, shift_out_10_port, shift_out_9_port
      , shift_out_8_port, shift_out_7_port, shift_out_6_port, shift_out_5_port,
      shift_out_4_port, shift_out_3_port, shift_out_2_port, shift_out_1_port, 
      shift_out_0_port, lu_out_31_port, lu_out_30_port, lu_out_29_port, 
      lu_out_28_port, lu_out_27_port, lu_out_26_port, lu_out_25_port, 
      lu_out_24_port, lu_out_23_port, lu_out_22_port, lu_out_21_port, 
      lu_out_20_port, lu_out_19_port, lu_out_18_port, lu_out_17_port, 
      lu_out_16_port, lu_out_15_port, lu_out_14_port, lu_out_13_port, 
      lu_out_12_port, lu_out_11_port, lu_out_10_port, lu_out_9_port, 
      lu_out_8_port, lu_out_7_port, lu_out_6_port, lu_out_5_port, lu_out_4_port
      , lu_out_3_port, lu_out_2_port, lu_out_1_port, lu_out_0_port, n120, n149,
      n150, n168, n169, n172, n174, n179, n185, n8, n10, n12, n13, n14, n15, 
      n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30
      , n31, n32, n33, n34, n35, n38, n39, n40, n41, n44, n45, n46, n47, n48, 
      n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63
      , n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, 
      n78, n79, n80, n84, n267, n268, n269, n270, n271, n272, n273, n274, n275,
      n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, 
      n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, 
      n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, 
      n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, 
      n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, 
      n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, 
      n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, 
      n360, n361, n362, n363, n364 : std_logic;

begin
   
   X_Logic0_port <= '0';
   U120 : MUX2_X1 port map( A => B_booth_to_add_31_port, B => IN2(31), S => n8,
                           Z => mux_B_31_port);
   U121 : MUX2_X1 port map( A => B_booth_to_add_30_port, B => IN2(30), S => n8,
                           Z => mux_B_30_port);
   U124 : MUX2_X1 port map( A => B_booth_to_add_28_port, B => IN2(28), S => n8,
                           Z => mux_B_28_port);
   U126 : MUX2_X1 port map( A => B_booth_to_add_26_port, B => IN2(26), S => n8,
                           Z => mux_B_26_port);
   U127 : MUX2_X1 port map( A => B_booth_to_add_25_port, B => IN2(25), S => n8,
                           Z => mux_B_25_port);
   U128 : MUX2_X1 port map( A => B_booth_to_add_24_port, B => IN2(24), S => n8,
                           Z => mux_B_24_port);
   U129 : MUX2_X1 port map( A => B_booth_to_add_23_port, B => IN2(23), S => n8,
                           Z => mux_B_23_port);
   U130 : MUX2_X1 port map( A => B_booth_to_add_22_port, B => IN2(22), S => n8,
                           Z => mux_B_22_port);
   U132 : MUX2_X1 port map( A => B_booth_to_add_20_port, B => IN2(20), S => n8,
                           Z => mux_B_20_port);
   U145 : MUX2_X1 port map( A => A_booth_to_add_9_port, B => IN1(9), S => n282,
                           Z => mux_A_9_port);
   U146 : MUX2_X1 port map( A => A_booth_to_add_8_port, B => IN1(8), S => n282,
                           Z => mux_A_8_port);
   U147 : MUX2_X1 port map( A => A_booth_to_add_7_port, B => IN1(7), S => n282,
                           Z => mux_A_7_port);
   U150 : MUX2_X1 port map( A => A_booth_to_add_4_port, B => IN1(4), S => n282,
                           Z => mux_A_4_port);
   U151 : MUX2_X1 port map( A => A_booth_to_add_3_port, B => IN1(3), S => n282,
                           Z => mux_A_3_port);
   U152 : MUX2_X1 port map( A => A_booth_to_add_31_port, B => IN1(31), S => 
                           n282, Z => mux_A_31_port);
   U153 : MUX2_X1 port map( A => A_booth_to_add_30_port, B => IN1(30), S => 
                           n282, Z => mux_A_30_port);
   U155 : MUX2_X1 port map( A => A_booth_to_add_29_port, B => IN1(29), S => 
                           n282, Z => mux_A_29_port);
   U156 : MUX2_X1 port map( A => A_booth_to_add_28_port, B => IN1(28), S => 
                           n282, Z => mux_A_28_port);
   U157 : MUX2_X1 port map( A => A_booth_to_add_27_port, B => IN1(27), S => 
                           n282, Z => mux_A_27_port);
   U158 : MUX2_X1 port map( A => A_booth_to_add_26_port, B => IN1(26), S => 
                           n282, Z => mux_A_26_port);
   U159 : MUX2_X1 port map( A => A_booth_to_add_25_port, B => IN1(25), S => 
                           n282, Z => mux_A_25_port);
   U160 : MUX2_X1 port map( A => A_booth_to_add_24_port, B => IN1(24), S => 
                           n282, Z => mux_A_24_port);
   U161 : MUX2_X1 port map( A => A_booth_to_add_23_port, B => IN1(23), S => 
                           n282, Z => mux_A_23_port);
   U162 : MUX2_X1 port map( A => A_booth_to_add_22_port, B => IN1(22), S => 
                           n282, Z => mux_A_22_port);
   U163 : MUX2_X1 port map( A => A_booth_to_add_21_port, B => IN1(21), S => 
                           n282, Z => mux_A_21_port);
   U164 : MUX2_X1 port map( A => A_booth_to_add_20_port, B => IN1(20), S => 
                           n282, Z => mux_A_20_port);
   U165 : MUX2_X1 port map( A => A_booth_to_add_1_port, B => IN1(1), S => n282,
                           Z => mux_A_1_port);
   U166 : MUX2_X1 port map( A => A_booth_to_add_19_port, B => IN1(19), S => 
                           n282, Z => mux_A_19_port);
   U167 : MUX2_X1 port map( A => A_booth_to_add_18_port, B => IN1(18), S => 
                           n282, Z => mux_A_18_port);
   U168 : MUX2_X1 port map( A => A_booth_to_add_17_port, B => IN1(17), S => 
                           n282, Z => mux_A_17_port);
   U169 : MUX2_X1 port map( A => A_booth_to_add_16_port, B => IN1(16), S => 
                           n282, Z => mux_A_16_port);
   U170 : MUX2_X1 port map( A => A_booth_to_add_15_port, B => IN1(15), S => 
                           n282, Z => mux_A_15_port);
   U171 : MUX2_X1 port map( A => A_booth_to_add_14_port, B => IN1(14), S => 
                           n282, Z => mux_A_14_port);
   U172 : MUX2_X1 port map( A => A_booth_to_add_13_port, B => IN1(13), S => 
                           n282, Z => mux_A_13_port);
   U173 : MUX2_X1 port map( A => A_booth_to_add_12_port, B => IN1(12), S => 
                           n282, Z => mux_A_12_port);
   U174 : MUX2_X1 port map( A => A_booth_to_add_11_port, B => IN1(11), S => 
                           n282, Z => mux_A_11_port);
   U175 : MUX2_X1 port map( A => A_booth_to_add_10_port, B => IN1(10), S => 
                           n282, Z => mux_A_10_port);
   U178 : NAND3_X1 port map( A1 => n84, A2 => n80, A3 => ALUW_i(12), ZN => n31)
                           ;
   MULT : simple_booth_add_ext_N16 port map( Clock => Clock, Reset => Reset, 
                           sign => ALUW_i(0), enable => ALUW_i(1), valid => 
                           valid_from_booth, A(15) => IN1(15), A(14) => IN1(14)
                           , A(13) => IN1(13), A(12) => IN1(12), A(11) => 
                           IN1(11), A(10) => IN1(10), A(9) => IN1(9), A(8) => 
                           IN1(8), A(7) => IN1(7), A(6) => IN1(6), A(5) => 
                           IN1(5), A(4) => IN1(4), A(3) => IN1(3), A(2) => 
                           IN1(2), A(1) => IN1(1), A(0) => IN1(0), B(15) => 
                           n286, B(14) => IN2(14), B(13) => n288, B(12) => n287
                           , B(11) => n363, B(10) => n300, B(9) => n362, B(8) 
                           => n291, B(7) => n289, B(6) => n285, B(5) => n299, 
                           B(4) => n293, B(3) => n297, B(2) => IN2(2), B(1) => 
                           n298, B(0) => n292, A_to_add(31) => 
                           A_booth_to_add_31_port, A_to_add(30) => 
                           A_booth_to_add_30_port, A_to_add(29) => 
                           A_booth_to_add_29_port, A_to_add(28) => 
                           A_booth_to_add_28_port, A_to_add(27) => 
                           A_booth_to_add_27_port, A_to_add(26) => 
                           A_booth_to_add_26_port, A_to_add(25) => 
                           A_booth_to_add_25_port, A_to_add(24) => 
                           A_booth_to_add_24_port, A_to_add(23) => 
                           A_booth_to_add_23_port, A_to_add(22) => 
                           A_booth_to_add_22_port, A_to_add(21) => 
                           A_booth_to_add_21_port, A_to_add(20) => 
                           A_booth_to_add_20_port, A_to_add(19) => 
                           A_booth_to_add_19_port, A_to_add(18) => 
                           A_booth_to_add_18_port, A_to_add(17) => 
                           A_booth_to_add_17_port, A_to_add(16) => 
                           A_booth_to_add_16_port, A_to_add(15) => 
                           A_booth_to_add_15_port, A_to_add(14) => 
                           A_booth_to_add_14_port, A_to_add(13) => 
                           A_booth_to_add_13_port, A_to_add(12) => 
                           A_booth_to_add_12_port, A_to_add(11) => 
                           A_booth_to_add_11_port, A_to_add(10) => 
                           A_booth_to_add_10_port, A_to_add(9) => 
                           A_booth_to_add_9_port, A_to_add(8) => 
                           A_booth_to_add_8_port, A_to_add(7) => 
                           A_booth_to_add_7_port, A_to_add(6) => 
                           A_booth_to_add_6_port, A_to_add(5) => 
                           A_booth_to_add_5_port, A_to_add(4) => 
                           A_booth_to_add_4_port, A_to_add(3) => 
                           A_booth_to_add_3_port, A_to_add(2) => 
                           A_booth_to_add_2_port, A_to_add(1) => 
                           A_booth_to_add_1_port, A_to_add(0) => 
                           A_booth_to_add_0_port, B_to_add(31) => 
                           B_booth_to_add_31_port, B_to_add(30) => 
                           B_booth_to_add_30_port, B_to_add(29) => 
                           B_booth_to_add_29_port, B_to_add(28) => 
                           B_booth_to_add_28_port, B_to_add(27) => 
                           B_booth_to_add_27_port, B_to_add(26) => 
                           B_booth_to_add_26_port, B_to_add(25) => 
                           B_booth_to_add_25_port, B_to_add(24) => 
                           B_booth_to_add_24_port, B_to_add(23) => 
                           B_booth_to_add_23_port, B_to_add(22) => 
                           B_booth_to_add_22_port, B_to_add(21) => 
                           B_booth_to_add_21_port, B_to_add(20) => 
                           B_booth_to_add_20_port, B_to_add(19) => 
                           B_booth_to_add_19_port, B_to_add(18) => 
                           B_booth_to_add_18_port, B_to_add(17) => 
                           B_booth_to_add_17_port, B_to_add(16) => 
                           B_booth_to_add_16_port, B_to_add(15) => 
                           B_booth_to_add_15_port, B_to_add(14) => 
                           B_booth_to_add_14_port, B_to_add(13) => 
                           B_booth_to_add_13_port, B_to_add(12) => 
                           B_booth_to_add_12_port, B_to_add(11) => 
                           B_booth_to_add_11_port, B_to_add(10) => 
                           B_booth_to_add_10_port, B_to_add(9) => 
                           B_booth_to_add_9_port, B_to_add(8) => 
                           B_booth_to_add_8_port, B_to_add(7) => 
                           B_booth_to_add_7_port, B_to_add(6) => 
                           B_booth_to_add_6_port, B_to_add(5) => 
                           B_booth_to_add_5_port, B_to_add(4) => 
                           B_booth_to_add_4_port, B_to_add(3) => 
                           B_booth_to_add_3_port, B_to_add(2) => 
                           B_booth_to_add_2_port, B_to_add(1) => 
                           B_booth_to_add_1_port, B_to_add(0) => 
                           B_booth_to_add_0_port, sign_to_add => 
                           sign_booth_to_add, final_out(31) => mult_out_31_port
                           , final_out(30) => mult_out_30_port, final_out(29) 
                           => mult_out_29_port, final_out(28) => 
                           mult_out_28_port, final_out(27) => mult_out_27_port,
                           final_out(26) => mult_out_26_port, final_out(25) => 
                           mult_out_25_port, final_out(24) => mult_out_24_port,
                           final_out(23) => mult_out_23_port, final_out(22) => 
                           mult_out_22_port, final_out(21) => mult_out_21_port,
                           final_out(20) => mult_out_20_port, final_out(19) => 
                           mult_out_19_port, final_out(18) => mult_out_18_port,
                           final_out(17) => mult_out_17_port, final_out(16) => 
                           mult_out_16_port, final_out(15) => mult_out_15_port,
                           final_out(14) => mult_out_14_port, final_out(13) => 
                           mult_out_13_port, final_out(12) => mult_out_12_port,
                           final_out(11) => mult_out_11_port, final_out(10) => 
                           mult_out_10_port, final_out(9) => mult_out_9_port, 
                           final_out(8) => mult_out_8_port, final_out(7) => 
                           mult_out_7_port, final_out(6) => mult_out_6_port, 
                           final_out(5) => mult_out_5_port, final_out(4) => 
                           mult_out_4_port, final_out(3) => mult_out_3_port, 
                           final_out(2) => mult_out_2_port, final_out(1) => 
                           mult_out_1_port, final_out(0) => mult_out_0_port, 
                           ACC_from_add(31) => n185, ACC_from_add(30) => 
                           sum_out_30_port, ACC_from_add(29) => n296, 
                           ACC_from_add(28) => n290, ACC_from_add(27) => 
                           sum_out_27_port, ACC_from_add(26) => sum_out_26_port
                           , ACC_from_add(25) => n294, ACC_from_add(24) => n295
                           , ACC_from_add(23) => sum_out_23_port, 
                           ACC_from_add(22) => n169, ACC_from_add(21) => n174, 
                           ACC_from_add(20) => n179, ACC_from_add(19) => n120, 
                           ACC_from_add(18) => sum_out_18_port, 
                           ACC_from_add(17) => sum_out_17_port, 
                           ACC_from_add(16) => sum_out_16_port, 
                           ACC_from_add(15) => sum_out_15_port, 
                           ACC_from_add(14) => sum_out_14_port, 
                           ACC_from_add(13) => n283, ACC_from_add(12) => 
                           sum_out_12_port, ACC_from_add(11) => sum_out_11_port
                           , ACC_from_add(10) => sum_out_10_port, 
                           ACC_from_add(9) => sum_out_9_port, ACC_from_add(8) 
                           => sum_out_8_port, ACC_from_add(7) => sum_out_7_port
                           , ACC_from_add(6) => sum_out_6_port, ACC_from_add(5)
                           => sum_out_5_port, ACC_from_add(4) => sum_out_4_port
                           , ACC_from_add(3) => sum_out_3_port, ACC_from_add(2)
                           => sum_out_2_port, ACC_from_add(1) => sum_out_1_port
                           , ACC_from_add(0) => sum_out_0_port);
   ADDER : p4add_N32_logN5_1 port map( A(31) => mux_A_31_port, A(30) => 
                           mux_A_30_port, A(29) => mux_A_29_port, A(28) => 
                           mux_A_28_port, A(27) => mux_A_27_port, A(26) => 
                           mux_A_26_port, A(25) => mux_A_25_port, A(24) => 
                           mux_A_24_port, A(23) => mux_A_23_port, A(22) => 
                           mux_A_22_port, A(21) => mux_A_21_port, A(20) => 
                           mux_A_20_port, A(19) => mux_A_19_port, A(18) => 
                           mux_A_18_port, A(17) => mux_A_17_port, A(16) => 
                           mux_A_16_port, A(15) => mux_A_15_port, A(14) => 
                           mux_A_14_port, A(13) => mux_A_13_port, A(12) => 
                           mux_A_12_port, A(11) => mux_A_11_port, A(10) => 
                           mux_A_10_port, A(9) => mux_A_9_port, A(8) => 
                           mux_A_8_port, A(7) => mux_A_7_port, A(6) => 
                           mux_A_6_port, A(5) => mux_A_5_port, A(4) => 
                           mux_A_4_port, A(3) => mux_A_3_port, A(2) => 
                           mux_A_2_port, A(1) => mux_A_1_port, A(0) => 
                           mux_A_0_port, B(31) => mux_B_31_port, B(30) => 
                           mux_B_30_port, B(29) => mux_B_29_port, B(28) => 
                           mux_B_28_port, B(27) => mux_B_27_port, B(26) => 
                           mux_B_26_port, B(25) => mux_B_25_port, B(24) => 
                           mux_B_24_port, B(23) => mux_B_23_port, B(22) => 
                           mux_B_22_port, B(21) => mux_B_21_port, B(20) => 
                           mux_B_20_port, B(19) => mux_B_19_port, B(18) => 
                           mux_B_18_port, B(17) => mux_B_17_port, B(16) => 
                           mux_B_16_port, B(15) => mux_B_15_port, B(14) => 
                           mux_B_14_port, B(13) => mux_B_13_port, B(12) => 
                           mux_B_12_port, B(11) => mux_B_11_port, B(10) => 
                           mux_B_10_port, B(9) => mux_B_9_port, B(8) => 
                           mux_B_8_port, B(7) => mux_B_7_port, B(6) => 
                           mux_B_6_port, B(5) => mux_B_5_port, B(4) => 
                           mux_B_4_port, B(3) => mux_B_3_port, B(2) => 
                           mux_B_2_port, B(1) => mux_B_1_port, B(0) => 
                           mux_B_0_port, Cin => X_Logic0_port, sign => mux_sign
                           , S(31) => n185, S(30) => sum_out_30_port, S(29) => 
                           n168, S(28) => n172, S(27) => sum_out_27_port, S(26)
                           => sum_out_26_port, S(25) => n149, S(24) => n150, 
                           S(23) => sum_out_23_port, S(22) => n169, S(21) => 
                           n174, S(20) => n179, S(19) => n120, S(18) => 
                           sum_out_18_port, S(17) => sum_out_17_port, S(16) => 
                           sum_out_16_port, S(15) => sum_out_15_port, S(14) => 
                           sum_out_14_port, S(13) => sum_out_13_port, S(12) => 
                           sum_out_12_port, S(11) => sum_out_11_port, S(10) => 
                           sum_out_10_port, S(9) => sum_out_9_port, S(8) => 
                           sum_out_8_port, S(7) => sum_out_7_port, S(6) => 
                           sum_out_6_port, S(5) => sum_out_5_port, S(4) => 
                           sum_out_4_port, S(3) => sum_out_3_port, S(2) => 
                           sum_out_2_port, S(1) => sum_out_1_port, S(0) => 
                           sum_out_0_port, Cout => carry_from_adder);
   COMP : comparator_M32 port map( C => carry_from_adder, V => overflow, 
                           SUM(31) => n185, SUM(30) => sum_out_30_port, SUM(29)
                           => n168, SUM(28) => n172, SUM(27) => sum_out_27_port
                           , SUM(26) => sum_out_26_port, SUM(25) => n149, 
                           SUM(24) => n150, SUM(23) => sum_out_23_port, SUM(22)
                           => n169, SUM(21) => n174, SUM(20) => n179, SUM(19) 
                           => n120, SUM(18) => sum_out_18_port, SUM(17) => 
                           sum_out_17_port, SUM(16) => sum_out_16_port, SUM(15)
                           => sum_out_15_port, SUM(14) => sum_out_14_port, 
                           SUM(13) => sum_out_13_port, SUM(12) => 
                           sum_out_12_port, SUM(11) => sum_out_11_port, SUM(10)
                           => sum_out_10_port, SUM(9) => sum_out_9_port, SUM(8)
                           => sum_out_8_port, SUM(7) => sum_out_7_port, SUM(6) 
                           => sum_out_6_port, SUM(5) => sum_out_5_port, SUM(4) 
                           => sum_out_4_port, SUM(3) => sum_out_3_port, SUM(2) 
                           => sum_out_2_port, SUM(1) => sum_out_1_port, SUM(0) 
                           => sum_out_0_port, sel(2) => ALUW_i(4), sel(1) => 
                           ALUW_i(3), sel(0) => ALUW_i(2), sign => ALUW_i(0), S
                           => comp_out);
   SHIFT : shifter port map( A(31) => IN1(31), A(30) => IN1(30), A(29) => 
                           IN1(29), A(28) => IN1(28), A(27) => IN1(27), A(26) 
                           => IN1(26), A(25) => IN1(25), A(24) => IN1(24), 
                           A(23) => IN1(23), A(22) => IN1(22), A(21) => IN1(21)
                           , A(20) => IN1(20), A(19) => IN1(19), A(18) => 
                           IN1(18), A(17) => IN1(17), A(16) => IN1(16), A(15) 
                           => IN1(15), A(14) => IN1(14), A(13) => IN1(13), 
                           A(12) => IN1(12), A(11) => IN1(11), A(10) => IN1(10)
                           , A(9) => IN1(9), A(8) => IN1(8), A(7) => IN1(7), 
                           A(6) => IN1(6), A(5) => IN1(5), A(4) => IN1(4), A(3)
                           => IN1(3), A(2) => IN1(2), A(1) => IN1(1), A(0) => 
                           IN1(0), B(4) => n293, B(3) => n297, B(2) => IN2(2), 
                           B(1) => n298, B(0) => n292, LOGIC_ARITH => ALUW_i(8)
                           , LEFT_RIGHT => ALUW_i(9), OUTPUT(31) => 
                           shift_out_31_port, OUTPUT(30) => shift_out_30_port, 
                           OUTPUT(29) => shift_out_29_port, OUTPUT(28) => 
                           shift_out_28_port, OUTPUT(27) => shift_out_27_port, 
                           OUTPUT(26) => shift_out_26_port, OUTPUT(25) => 
                           shift_out_25_port, OUTPUT(24) => shift_out_24_port, 
                           OUTPUT(23) => shift_out_23_port, OUTPUT(22) => 
                           shift_out_22_port, OUTPUT(21) => shift_out_21_port, 
                           OUTPUT(20) => shift_out_20_port, OUTPUT(19) => 
                           shift_out_19_port, OUTPUT(18) => shift_out_18_port, 
                           OUTPUT(17) => shift_out_17_port, OUTPUT(16) => 
                           shift_out_16_port, OUTPUT(15) => shift_out_15_port, 
                           OUTPUT(14) => shift_out_14_port, OUTPUT(13) => 
                           shift_out_13_port, OUTPUT(12) => shift_out_12_port, 
                           OUTPUT(11) => shift_out_11_port, OUTPUT(10) => 
                           shift_out_10_port, OUTPUT(9) => shift_out_9_port, 
                           OUTPUT(8) => shift_out_8_port, OUTPUT(7) => 
                           shift_out_7_port, OUTPUT(6) => shift_out_6_port, 
                           OUTPUT(5) => shift_out_5_port, OUTPUT(4) => 
                           shift_out_4_port, OUTPUT(3) => shift_out_3_port, 
                           OUTPUT(2) => shift_out_2_port, OUTPUT(1) => 
                           shift_out_1_port, OUTPUT(0) => shift_out_0_port);
   LU : logic_unit_SIZE32 port map( IN1(31) => IN1(31), IN1(30) => IN1(30), 
                           IN1(29) => IN1(29), IN1(28) => IN1(28), IN1(27) => 
                           IN1(27), IN1(26) => IN1(26), IN1(25) => IN1(25), 
                           IN1(24) => IN1(24), IN1(23) => IN1(23), IN1(22) => 
                           IN1(22), IN1(21) => IN1(21), IN1(20) => IN1(20), 
                           IN1(19) => IN1(19), IN1(18) => IN1(18), IN1(17) => 
                           IN1(17), IN1(16) => IN1(16), IN1(15) => IN1(15), 
                           IN1(14) => IN1(14), IN1(13) => IN1(13), IN1(12) => 
                           IN1(12), IN1(11) => IN1(11), IN1(10) => IN1(10), 
                           IN1(9) => IN1(9), IN1(8) => IN1(8), IN1(7) => IN1(7)
                           , IN1(6) => IN1(6), IN1(5) => IN1(5), IN1(4) => 
                           IN1(4), IN1(3) => IN1(3), IN1(2) => IN1(2), IN1(1) 
                           => IN1(1), IN1(0) => IN1(0), IN2(31) => IN2(31), 
                           IN2(30) => IN2(30), IN2(29) => IN2(29), IN2(28) => 
                           IN2(28), IN2(27) => IN2(27), IN2(26) => IN2(26), 
                           IN2(25) => IN2(25), IN2(24) => IN2(24), IN2(23) => 
                           IN2(23), IN2(22) => IN2(22), IN2(21) => IN2(21), 
                           IN2(20) => IN2(20), IN2(19) => IN2(19), IN2(18) => 
                           IN2(18), IN2(17) => n284, IN2(16) => IN2(16), 
                           IN2(15) => n286, IN2(14) => IN2(14), IN2(13) => n288
                           , IN2(12) => n287, IN2(11) => n363, IN2(10) => n300,
                           IN2(9) => n362, IN2(8) => n291, IN2(7) => n289, 
                           IN2(6) => IN2(6), IN2(5) => n299, IN2(4) => n293, 
                           IN2(3) => n297, IN2(2) => IN2(2), IN2(1) => n298, 
                           IN2(0) => n292, CTRL(1) => ALUW_i(6), CTRL(0) => 
                           ALUW_i(5), OUT1(31) => lu_out_31_port, OUT1(30) => 
                           lu_out_30_port, OUT1(29) => lu_out_29_port, OUT1(28)
                           => lu_out_28_port, OUT1(27) => lu_out_27_port, 
                           OUT1(26) => lu_out_26_port, OUT1(25) => 
                           lu_out_25_port, OUT1(24) => lu_out_24_port, OUT1(23)
                           => lu_out_23_port, OUT1(22) => lu_out_22_port, 
                           OUT1(21) => lu_out_21_port, OUT1(20) => 
                           lu_out_20_port, OUT1(19) => lu_out_19_port, OUT1(18)
                           => lu_out_18_port, OUT1(17) => lu_out_17_port, 
                           OUT1(16) => lu_out_16_port, OUT1(15) => 
                           lu_out_15_port, OUT1(14) => lu_out_14_port, OUT1(13)
                           => lu_out_13_port, OUT1(12) => lu_out_12_port, 
                           OUT1(11) => lu_out_11_port, OUT1(10) => 
                           lu_out_10_port, OUT1(9) => lu_out_9_port, OUT1(8) =>
                           lu_out_8_port, OUT1(7) => lu_out_7_port, OUT1(6) => 
                           lu_out_6_port, OUT1(5) => lu_out_5_port, OUT1(4) => 
                           lu_out_4_port, OUT1(3) => lu_out_3_port, OUT1(2) => 
                           lu_out_2_port, OUT1(1) => lu_out_1_port, OUT1(0) => 
                           lu_out_0_port);
   U134 : MUX2_X1 port map( A => B_booth_to_add_19_port, B => IN2(19), S => n8,
                           Z => mux_B_19_port);
   U33 : AOI222_X1 port map( A1 => IN2(30), A2 => n16, B1 => n17, B2 => 
                           mult_out_30_port, C1 => n280, C2 => 
                           shift_out_30_port, ZN => n34);
   U32 : AOI22_X1 port map( A1 => n281, A2 => lu_out_30_port, B1 => n15, B2 => 
                           sum_out_30_port, ZN => n35);
   U31 : NAND2_X1 port map( A1 => n34, A2 => n35, ZN => DOUT(30));
   U57 : AOI222_X1 port map( A1 => IN2(23), A2 => n16, B1 => n17, B2 => 
                           mult_out_23_port, C1 => n280, C2 => 
                           shift_out_23_port, ZN => n50);
   U56 : AOI22_X1 port map( A1 => n281, A2 => lu_out_23_port, B1 => n364, B2 =>
                           sum_out_23_port, ZN => n51);
   U55 : NAND2_X1 port map( A1 => n50, A2 => n51, ZN => DOUT(23));
   U48 : AOI222_X1 port map( A1 => IN2(26), A2 => n16, B1 => n17, B2 => 
                           mult_out_26_port, C1 => n280, C2 => 
                           shift_out_26_port, ZN => n44);
   U47 : AOI22_X1 port map( A1 => n281, A2 => lu_out_26_port, B1 => 
                           sum_out_26_port, B2 => n15, ZN => n45);
   U46 : NAND2_X1 port map( A1 => n44, A2 => n45, ZN => DOUT(26));
   U60 : AOI222_X1 port map( A1 => IN2(22), A2 => n16, B1 => n17, B2 => 
                           mult_out_22_port, C1 => n280, C2 => 
                           shift_out_22_port, ZN => n52);
   U59 : AOI22_X1 port map( A1 => n281, A2 => lu_out_22_port, B1 => n364, B2 =>
                           n169, ZN => n53);
   U58 : NAND2_X1 port map( A1 => n52, A2 => n53, ZN => DOUT(22));
   U39 : AOI222_X1 port map( A1 => IN2(29), A2 => n16, B1 => n17, B2 => 
                           mult_out_29_port, C1 => n280, C2 => 
                           shift_out_29_port, ZN => n38);
   U37 : NAND2_X1 port map( A1 => n38, A2 => n39, ZN => DOUT(29));
   U42 : AOI222_X1 port map( A1 => IN2(28), A2 => n16, B1 => n17, B2 => 
                           mult_out_28_port, C1 => n280, C2 => 
                           shift_out_28_port, ZN => n40);
   U40 : NAND2_X1 port map( A1 => n40, A2 => n41, ZN => DOUT(28));
   U49 : NAND2_X1 port map( A1 => n46, A2 => n47, ZN => DOUT(25));
   U63 : AOI222_X1 port map( A1 => IN2(21), A2 => n16, B1 => n17, B2 => 
                           mult_out_21_port, C1 => n280, C2 => 
                           shift_out_21_port, ZN => n54);
   U61 : NAND2_X1 port map( A1 => n54, A2 => n55, ZN => DOUT(21));
   U66 : AOI222_X1 port map( A1 => IN2(20), A2 => n16, B1 => n17, B2 => 
                           mult_out_20_port, C1 => n280, C2 => 
                           shift_out_20_port, ZN => n56);
   U64 : NAND2_X1 port map( A1 => n56, A2 => n57, ZN => DOUT(20));
   U54 : AOI222_X1 port map( A1 => IN2(24), A2 => n16, B1 => n17, B2 => 
                           mult_out_24_port, C1 => n280, C2 => 
                           shift_out_24_port, ZN => n48);
   U52 : NAND2_X1 port map( A1 => n48, A2 => n49, ZN => DOUT(24));
   U28 : AOI22_X1 port map( A1 => n17, A2 => mult_out_31_port, B1 => n280, B2 
                           => shift_out_31_port, ZN => n33);
   U27 : OAI211_X1 port map( C1 => n31, C2 => n10, A => n32, B => n33, ZN => 
                           DOUT(31));
   U72 : AOI222_X1 port map( A1 => IN2(19), A2 => n16, B1 => n17, B2 => 
                           mult_out_19_port, C1 => n280, C2 => 
                           shift_out_19_port, ZN => n60);
   U71 : AOI22_X1 port map( A1 => n281, A2 => lu_out_19_port, B1 => n364, B2 =>
                           n120, ZN => n61);
   U70 : NAND2_X1 port map( A1 => n60, A2 => n61, ZN => DOUT(19));
   U89 : AOI22_X1 port map( A1 => n281, A2 => lu_out_13_port, B1 => n364, B2 =>
                           n283, ZN => n73);
   U88 : NAND2_X1 port map( A1 => n72, A2 => n73, ZN => DOUT(13));
   U86 : AOI22_X1 port map( A1 => n281, A2 => lu_out_14_port, B1 => n364, B2 =>
                           sum_out_14_port, ZN => n71);
   U85 : NAND2_X1 port map( A1 => n70, A2 => n71, ZN => DOUT(14));
   U92 : AOI22_X1 port map( A1 => n281, A2 => lu_out_12_port, B1 => n364, B2 =>
                           sum_out_12_port, ZN => n75);
   U91 : NAND2_X1 port map( A1 => n74, A2 => n75, ZN => DOUT(12));
   U96 : AOI222_X1 port map( A1 => n363, A2 => n16, B1 => n17, B2 => 
                           mult_out_11_port, C1 => n280, C2 => 
                           shift_out_11_port, ZN => n76);
   U95 : AOI22_X1 port map( A1 => n281, A2 => lu_out_11_port, B1 => n364, B2 =>
                           sum_out_11_port, ZN => n77);
   U94 : NAND2_X1 port map( A1 => n76, A2 => n77, ZN => DOUT(11));
   U84 : AOI222_X1 port map( A1 => n286, A2 => n16, B1 => n17, B2 => 
                           mult_out_15_port, C1 => n18, C2 => shift_out_15_port
                           , ZN => n68);
   U83 : AOI22_X1 port map( A1 => n281, A2 => lu_out_15_port, B1 => n364, B2 =>
                           sum_out_15_port, ZN => n69);
   U82 : NAND2_X1 port map( A1 => n68, A2 => n69, ZN => DOUT(15));
   U13 : AOI22_X1 port map( A1 => n281, A2 => lu_out_7_port, B1 => n15, B2 => 
                           sum_out_7_port, ZN => n22);
   U12 : NAND2_X1 port map( A1 => n21, A2 => n22, ZN => DOUT(7));
   U77 : AOI22_X1 port map( A1 => n281, A2 => lu_out_17_port, B1 => n364, B2 =>
                           sum_out_17_port, ZN => n65);
   U76 : NAND2_X1 port map( A1 => n64, A2 => n65, ZN => DOUT(17));
   U98 : AOI22_X1 port map( A1 => n281, A2 => lu_out_10_port, B1 => n364, B2 =>
                           sum_out_10_port, ZN => n79);
   U97 : NAND2_X1 port map( A1 => n78, A2 => n79, ZN => DOUT(10));
   U7 : AOI22_X1 port map( A1 => n281, A2 => lu_out_9_port, B1 => n364, B2 => 
                           sum_out_9_port, ZN => n13);
   U6 : NAND2_X1 port map( A1 => n12, A2 => n13, ZN => DOUT(9));
   U25 : AOI22_X1 port map( A1 => n14, A2 => lu_out_3_port, B1 => n364, B2 => 
                           sum_out_3_port, ZN => n30);
   U24 : NAND2_X1 port map( A1 => n29, A2 => n30, ZN => DOUT(3));
   U68 : AOI22_X1 port map( A1 => n281, A2 => lu_out_1_port, B1 => n364, B2 => 
                           sum_out_1_port, ZN => n59);
   U67 : NAND2_X1 port map( A1 => n58, A2 => n59, ZN => DOUT(1));
   U11 : AOI222_X1 port map( A1 => n291, A2 => n16, B1 => n17, B2 => 
                           mult_out_8_port, C1 => n280, C2 => shift_out_8_port,
                           ZN => n19);
   U10 : AOI22_X1 port map( A1 => n281, A2 => lu_out_8_port, B1 => n364, B2 => 
                           sum_out_8_port, ZN => n20);
   U9 : NAND2_X1 port map( A1 => n19, A2 => n20, ZN => DOUT(8));
   U75 : AOI222_X1 port map( A1 => IN2(18), A2 => n16, B1 => n17, B2 => 
                           mult_out_18_port, C1 => n280, C2 => 
                           shift_out_18_port, ZN => n62);
   U74 : AOI22_X1 port map( A1 => n281, A2 => lu_out_18_port, B1 => n364, B2 =>
                           sum_out_18_port, ZN => n63);
   U73 : NAND2_X1 port map( A1 => n62, A2 => n63, ZN => DOUT(18));
   U81 : AOI222_X1 port map( A1 => IN2(16), A2 => n16, B1 => n17, B2 => 
                           mult_out_16_port, C1 => n18, C2 => shift_out_16_port
                           , ZN => n66);
   U80 : AOI22_X1 port map( A1 => n281, A2 => lu_out_16_port, B1 => n364, B2 =>
                           sum_out_16_port, ZN => n67);
   U79 : NAND2_X1 port map( A1 => n66, A2 => n67, ZN => DOUT(16));
   U19 : AOI22_X1 port map( A1 => n281, A2 => lu_out_5_port, B1 => n364, B2 => 
                           sum_out_5_port, ZN => n26);
   U18 : NAND2_X1 port map( A1 => n25, A2 => n26, ZN => DOUT(5));
   U22 : AOI22_X1 port map( A1 => n281, A2 => lu_out_4_port, B1 => n364, B2 => 
                           sum_out_4_port, ZN => n28);
   U21 : NAND2_X1 port map( A1 => n27, A2 => n28, ZN => DOUT(4));
   U16 : AOI22_X1 port map( A1 => n281, A2 => lu_out_6_port, B1 => n364, B2 => 
                           sum_out_6_port, ZN => n24);
   U15 : NAND2_X1 port map( A1 => n23, A2 => n24, ZN => DOUT(6));
   U154 : MUX2_X1 port map( A => A_booth_to_add_2_port, B => IN1(2), S => n282,
                           Z => mux_A_2_port);
   U149 : MUX2_X1 port map( A => A_booth_to_add_5_port, B => IN1(5), S => n282,
                           Z => mux_A_5_port);
   U148 : MUX2_X1 port map( A => A_booth_to_add_6_port, B => IN1(6), S => n282,
                           Z => mux_A_6_port);
   U109 : INV_X1 port map( A => ALUW_i(10), ZN => n80);
   U2 : NOR2_X1 port map( A1 => valid_from_booth, A2 => n282, ZN => stall_o);
   U3 : NAND2_X1 port map( A1 => n329, A2 => n317, ZN => mux_A_0_port);
   U4 : MUX2_X1 port map( A => B_booth_to_add_0_port, B => IN2(0), S => n282, Z
                           => mux_B_0_port);
   U5 : NAND2_X1 port map( A1 => n315, A2 => n349, ZN => mux_B_3_port);
   U8 : AOI22_X1 port map( A1 => sum_out_0_port, A2 => n364, B1 => n280, B2 => 
                           shift_out_0_port, ZN => n267);
   U14 : AOI22_X1 port map( A1 => n16, A2 => n292, B1 => n17, B2 => 
                           mult_out_0_port, ZN => n268);
   U17 : AND2_X1 port map( A1 => n267, A2 => n268, ZN => n359);
   U20 : MUX2_X1 port map( A => B_booth_to_add_5_port, B => IN2(5), S => n282, 
                           Z => mux_B_5_port);
   U23 : OAI21_X1 port map( B1 => n282, B2 => n319, A => n318, ZN => 
                           mux_B_9_port);
   U26 : INV_X1 port map( A => IN2(2), ZN => n269);
   U29 : INV_X1 port map( A => n16, ZN => n270);
   U30 : AOI22_X1 port map( A1 => shift_out_2_port, A2 => n280, B1 => 
                           mult_out_2_port, B2 => n17, ZN => n271);
   U34 : AOI22_X1 port map( A1 => sum_out_2_port, A2 => n364, B1 => 
                           lu_out_2_port, B2 => n281, ZN => n272);
   U35 : OAI211_X1 port map( C1 => n269, C2 => n270, A => n271, B => n272, ZN 
                           => DOUT(2));
   U36 : INV_X1 port map( A => n282, ZN => n273);
   U38 : NAND2_X1 port map( A1 => B_booth_to_add_3_port, A2 => n273, ZN => n315
                           );
   U41 : MUX2_X1 port map( A => B_booth_to_add_14_port, B => IN2(14), S => n8, 
                           Z => mux_B_14_port);
   U43 : MUX2_X1 port map( A => B_booth_to_add_21_port, B => IN2(21), S => n8, 
                           Z => mux_B_21_port);
   U44 : INV_X1 port map( A => n8, ZN => n274);
   U45 : NAND2_X1 port map( A1 => B_booth_to_add_16_port, A2 => n274, ZN => 
                           n304);
   U50 : MUX2_X1 port map( A => B_booth_to_add_29_port, B => IN2(29), S => n8, 
                           Z => mux_B_29_port);
   U51 : INV_X1 port map( A => IN2(27), ZN => n275);
   U53 : INV_X1 port map( A => n16, ZN => n276);
   U62 : AOI22_X1 port map( A1 => shift_out_27_port, A2 => n280, B1 => 
                           mult_out_27_port, B2 => n17, ZN => n277);
   U65 : AOI22_X1 port map( A1 => sum_out_27_port, A2 => n364, B1 => 
                           lu_out_27_port, B2 => n281, ZN => n278);
   U69 : OAI211_X1 port map( C1 => n275, C2 => n276, A => n277, B => n278, ZN 
                           => DOUT(27));
   U78 : CLKBUF_X1 port map( A => IN2(15), Z => n279);
   U87 : CLKBUF_X1 port map( A => IN2(12), Z => n287);
   U90 : AOI222_X1 port map( A1 => IN2(25), A2 => n16, B1 => n17, B2 => 
                           mult_out_25_port, C1 => n280, C2 => 
                           shift_out_25_port, ZN => n46);
   U93 : BUF_X1 port map( A => n149, Z => n294);
   U99 : AOI222_X1 port map( A1 => n284, A2 => n16, B1 => n17, B2 => 
                           mult_out_17_port, C1 => n280, C2 => 
                           shift_out_17_port, ZN => n64);
   U100 : AOI222_X1 port map( A1 => n300, A2 => n16, B1 => n17, B2 => 
                           mult_out_10_port, C1 => n280, C2 => 
                           shift_out_10_port, ZN => n78);
   U101 : AOI222_X1 port map( A1 => n299, A2 => n16, B1 => n17, B2 => 
                           mult_out_5_port, C1 => n280, C2 => shift_out_5_port,
                           ZN => n25);
   U102 : AOI222_X1 port map( A1 => n289, A2 => n16, B1 => n17, B2 => 
                           mult_out_7_port, C1 => n280, C2 => shift_out_7_port,
                           ZN => n21);
   U103 : AOI222_X1 port map( A1 => n298, A2 => n16, B1 => n17, B2 => 
                           mult_out_1_port, C1 => n280, C2 => shift_out_1_port,
                           ZN => n58);
   U104 : BUF_X1 port map( A => IN2(0), Z => n292);
   U105 : BUF_X1 port map( A => IN2(10), Z => n300);
   U106 : BUF_X1 port map( A => IN2(1), Z => n298);
   U107 : BUF_X1 port map( A => IN2(17), Z => n284);
   U108 : OR2_X1 port map( A1 => n282, A2 => n330, ZN => n317);
   U110 : OR2_X1 port map( A1 => n282, A2 => n332, ZN => n311);
   U111 : OR2_X1 port map( A1 => n282, A2 => n342, ZN => n312);
   U112 : OR2_X1 port map( A1 => n282, A2 => n340, ZN => n316);
   U113 : OR2_X1 port map( A1 => n282, A2 => n346, ZN => n313);
   U114 : OR2_X1 port map( A1 => n282, A2 => n328, ZN => n310);
   U115 : OR2_X1 port map( A1 => n282, A2 => n348, ZN => n314);
   U116 : AND2_X2 port map( A1 => n31, A2 => ALUW_i(12), ZN => n17);
   U117 : CLKBUF_X3 port map( A => n8, Z => n282);
   U118 : INV_X2 port map( A => ALUW_i(1), ZN => n8);
   U119 : AOI222_X1 port map( A1 => IN2(14), A2 => n16, B1 => n17, B2 => 
                           mult_out_14_port, C1 => n18, C2 => shift_out_14_port
                           , ZN => n70);
   U122 : BUF_X1 port map( A => n172, Z => n290);
   U123 : INV_X1 port map( A => n359, ZN => n358);
   U125 : INV_X1 port map( A => n360, ZN => n357);
   U131 : BUF_X1 port map( A => IN2(6), Z => n285);
   U133 : BUF_X1 port map( A => IN2(7), Z => n289);
   U135 : INV_X1 port map( A => IN2(31), ZN => n10);
   U136 : BUF_X1 port map( A => IN2(4), Z => n293);
   U137 : BUF_X1 port map( A => IN2(8), Z => n291);
   U138 : OR2_X1 port map( A1 => n8, A2 => n336, ZN => n306);
   U139 : OR2_X1 port map( A1 => n8, A2 => n338, ZN => n307);
   U140 : OR2_X1 port map( A1 => n8, A2 => n323, ZN => n302);
   U141 : OR2_X1 port map( A1 => n8, A2 => n344, ZN => n308);
   U142 : OR2_X1 port map( A1 => n8, A2 => n325, ZN => n303);
   U143 : OR2_X1 port map( A1 => n8, A2 => n321, ZN => n301);
   U144 : OR2_X1 port map( A1 => n8, A2 => n334, ZN => n305);
   U176 : OR2_X1 port map( A1 => n8, A2 => n351, ZN => n309);
   U177 : INV_X1 port map( A => B_booth_to_add_9_port, ZN => n319);
   U179 : INV_X1 port map( A => B_booth_to_add_4_port, ZN => n346);
   U180 : INV_X1 port map( A => B_booth_to_add_8_port, ZN => n342);
   U181 : INV_X1 port map( A => B_booth_to_add_6_port, ZN => n328);
   U182 : INV_X1 port map( A => B_booth_to_add_7_port, ZN => n348);
   U183 : BUF_X2 port map( A => n15, Z => n364);
   U184 : INV_X1 port map( A => B_booth_to_add_13_port, ZN => n338);
   U185 : INV_X1 port map( A => B_booth_to_add_12_port, ZN => n323);
   U186 : BUF_X2 port map( A => n18, Z => n280);
   U187 : INV_X1 port map( A => B_booth_to_add_11_port, ZN => n334);
   U188 : INV_X1 port map( A => B_booth_to_add_1_port, ZN => n351);
   U189 : INV_X1 port map( A => B_booth_to_add_10_port, ZN => n340);
   U190 : INV_X1 port map( A => B_booth_to_add_15_port, ZN => n336);
   U191 : INV_X1 port map( A => B_booth_to_add_2_port, ZN => n332);
   U192 : INV_X1 port map( A => B_booth_to_add_17_port, ZN => n344);
   U193 : BUF_X2 port map( A => n14, Z => n281);
   U194 : INV_X1 port map( A => B_booth_to_add_27_port, ZN => n321);
   U195 : INV_X1 port map( A => B_booth_to_add_18_port, ZN => n325);
   U196 : INV_X1 port map( A => ALUW_i(11), ZN => n84);
   U197 : INV_X1 port map( A => A_booth_to_add_0_port, ZN => n330);
   U198 : BUF_X1 port map( A => sum_out_13_port, Z => n283);
   U199 : CLKBUF_X1 port map( A => IN2(9), Z => n362);
   U200 : BUF_X1 port map( A => n279, Z => n286);
   U201 : CLKBUF_X1 port map( A => IN2(13), Z => n288);
   U202 : CLKBUF_X1 port map( A => n150, Z => n295);
   U203 : CLKBUF_X1 port map( A => n168, Z => n296);
   U204 : BUF_X1 port map( A => IN2(3), Z => n297);
   U205 : BUF_X1 port map( A => IN2(5), Z => n299);
   U206 : AOI222_X1 port map( A1 => n285, A2 => n16, B1 => n17, B2 => 
                           mult_out_6_port, C1 => n280, C2 => shift_out_6_port,
                           ZN => n23);
   U207 : INV_X1 port map( A => n355, ZN => DOUT(0));
   U208 : NOR3_X1 port map( A1 => ALUW_i(12), A2 => ALUW_i(11), A3 => 
                           ALUW_i(10), ZN => n15);
   U209 : NOR3_X1 port map( A1 => ALUW_i(12), A2 => ALUW_i(10), A3 => n84, ZN 
                           => n18);
   U210 : BUF_X1 port map( A => IN2(11), Z => n363);
   U211 : INV_X2 port map( A => n31, ZN => n16);
   U212 : MUX2_X2 port map( A => sign_booth_to_add, B => ALUW_i(7), S => n8, Z 
                           => mux_sign);
   U213 : AOI222_X1 port map( A1 => n293, A2 => n16, B1 => n17, B2 => 
                           mult_out_4_port, C1 => n280, C2 => shift_out_4_port,
                           ZN => n27);
   U214 : AOI222_X1 port map( A1 => n297, A2 => n16, B1 => n17, B2 => 
                           mult_out_3_port, C1 => n280, C2 => shift_out_3_port,
                           ZN => n29);
   U215 : AOI222_X1 port map( A1 => n362, A2 => n16, B1 => n17, B2 => 
                           mult_out_9_port, C1 => n280, C2 => shift_out_9_port,
                           ZN => n12);
   U216 : AOI222_X1 port map( A1 => n287, A2 => n16, B1 => n17, B2 => 
                           mult_out_12_port, C1 => n18, C2 => shift_out_12_port
                           , ZN => n74);
   U217 : AOI222_X1 port map( A1 => n288, A2 => n16, B1 => n17, B2 => 
                           mult_out_13_port, C1 => n280, C2 => 
                           shift_out_13_port, ZN => n72);
   U218 : OAI21_X1 port map( B1 => lu_out_0_port, B2 => ALUW_i(11), A => n361, 
                           ZN => n360);
   U219 : NOR2_X1 port map( A1 => n80, A2 => ALUW_i(12), ZN => n361);
   U220 : NAND2_X1 port map( A1 => n359, A2 => ALUW_i(11), ZN => n356);
   U221 : NOR2_X1 port map( A1 => n10, A2 => IN1(31), ZN => n354);
   U222 : NAND2_X1 port map( A1 => n10, A2 => IN1(31), ZN => n352);
   U223 : NOR3_X1 port map( A1 => ALUW_i(12), A2 => ALUW_i(11), A3 => n80, ZN 
                           => n14);
   U224 : NAND2_X1 port map( A1 => IN2(9), A2 => n282, ZN => n318);
   U225 : NAND2_X1 port map( A1 => IN2(27), A2 => n8, ZN => n320);
   U226 : NAND2_X1 port map( A1 => n320, A2 => n301, ZN => mux_B_27_port);
   U227 : NAND2_X1 port map( A1 => IN2(12), A2 => n8, ZN => n322);
   U228 : NAND2_X1 port map( A1 => n322, A2 => n302, ZN => mux_B_12_port);
   U229 : NAND2_X1 port map( A1 => IN2(18), A2 => n8, ZN => n324);
   U230 : NAND2_X1 port map( A1 => n324, A2 => n303, ZN => mux_B_18_port);
   U231 : NAND2_X1 port map( A1 => IN2(16), A2 => n8, ZN => n326);
   U232 : NAND2_X1 port map( A1 => n326, A2 => n304, ZN => mux_B_16_port);
   U233 : NAND2_X1 port map( A1 => IN2(6), A2 => n282, ZN => n327);
   U234 : NAND2_X1 port map( A1 => n327, A2 => n310, ZN => mux_B_6_port);
   U235 : NAND2_X1 port map( A1 => IN1(0), A2 => n282, ZN => n329);
   U236 : NAND2_X1 port map( A1 => IN2(2), A2 => n282, ZN => n331);
   U237 : NAND2_X1 port map( A1 => n331, A2 => n311, ZN => mux_B_2_port);
   U238 : NAND2_X1 port map( A1 => IN2(11), A2 => n8, ZN => n333);
   U239 : NAND2_X1 port map( A1 => n333, A2 => n305, ZN => mux_B_11_port);
   U240 : NAND2_X1 port map( A1 => IN2(15), A2 => n8, ZN => n335);
   U241 : NAND2_X1 port map( A1 => n335, A2 => n306, ZN => mux_B_15_port);
   U242 : NAND2_X1 port map( A1 => IN2(13), A2 => n8, ZN => n337);
   U243 : NAND2_X1 port map( A1 => n337, A2 => n307, ZN => mux_B_13_port);
   U244 : NAND2_X1 port map( A1 => IN2(10), A2 => n282, ZN => n339);
   U245 : NAND2_X1 port map( A1 => n339, A2 => n316, ZN => mux_B_10_port);
   U246 : NAND2_X1 port map( A1 => IN2(8), A2 => n282, ZN => n341);
   U247 : NAND2_X1 port map( A1 => n341, A2 => n312, ZN => mux_B_8_port);
   U248 : NAND2_X1 port map( A1 => IN2(17), A2 => n8, ZN => n343);
   U249 : NAND2_X1 port map( A1 => n343, A2 => n308, ZN => mux_B_17_port);
   U250 : NAND2_X1 port map( A1 => IN2(4), A2 => n282, ZN => n345);
   U251 : NAND2_X1 port map( A1 => n345, A2 => n313, ZN => mux_B_4_port);
   U252 : NAND2_X1 port map( A1 => IN2(7), A2 => n282, ZN => n347);
   U253 : NAND2_X1 port map( A1 => n347, A2 => n314, ZN => mux_B_7_port);
   U254 : NAND2_X1 port map( A1 => IN2(3), A2 => n282, ZN => n349);
   U255 : NAND2_X1 port map( A1 => IN2(1), A2 => n8, ZN => n350);
   U256 : NAND2_X1 port map( A1 => n350, A2 => n309, ZN => mux_B_1_port);
   U257 : NAND2_X1 port map( A1 => n185, A2 => n354, ZN => n353);
   U258 : OAI21_X1 port map( B1 => n185, B2 => n352, A => n353, ZN => overflow)
                           ;
   U259 : OAI22_X1 port map( A1 => comp_out, A2 => n356, B1 => n357, B2 => n358
                           , ZN => n355);
   U260 : AOI22_X1 port map( A1 => n281, A2 => lu_out_25_port, B1 => n15, B2 =>
                           n294, ZN => n47);
   U261 : AOI22_X1 port map( A1 => n281, A2 => lu_out_21_port, B1 => n364, B2 
                           => n174, ZN => n55);
   U262 : AOI22_X1 port map( A1 => n281, A2 => lu_out_29_port, B1 => n364, B2 
                           => n296, ZN => n39);
   U263 : AOI22_X1 port map( A1 => n281, A2 => lu_out_28_port, B1 => n364, B2 
                           => n290, ZN => n41);
   U264 : AOI22_X1 port map( A1 => n281, A2 => lu_out_24_port, B1 => n364, B2 
                           => n295, ZN => n49);
   U265 : AOI22_X1 port map( A1 => n281, A2 => lu_out_20_port, B1 => n364, B2 
                           => n179, ZN => n57);
   U266 : AOI22_X1 port map( A1 => n281, A2 => lu_out_31_port, B1 => n185, B2 
                           => n364, ZN => n32);

end SYN_Bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity mux21_0 is

   port( IN0, IN1 : in std_logic_vector (31 downto 0);  CTRL : in std_logic;  
         OUT1 : out std_logic_vector (31 downto 0));

end mux21_0;

architecture SYN_Bhe of mux21_0 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X2
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n15, n16, n17, n18, n19, n20, n21 : std_logic;

begin
   
   U8 : MUX2_X1 port map( A => IN0(31), B => IN1(31), S => CTRL, Z => OUT1(31))
                           ;
   U9 : MUX2_X1 port map( A => IN0(30), B => IN1(30), S => CTRL, Z => OUT1(30))
                           ;
   U11 : MUX2_X1 port map( A => IN0(29), B => IN1(29), S => CTRL, Z => OUT1(29)
                           );
   U12 : MUX2_X1 port map( A => IN0(28), B => IN1(28), S => CTRL, Z => OUT1(28)
                           );
   U14 : MUX2_X1 port map( A => IN0(26), B => IN1(26), S => CTRL, Z => OUT1(26)
                           );
   U16 : MUX2_X1 port map( A => IN0(24), B => IN1(24), S => CTRL, Z => OUT1(24)
                           );
   U18 : MUX2_X1 port map( A => IN0(22), B => IN1(22), S => CTRL, Z => OUT1(22)
                           );
   U19 : MUX2_X1 port map( A => IN0(21), B => IN1(21), S => CTRL, Z => OUT1(21)
                           );
   U20 : MUX2_X1 port map( A => IN0(20), B => IN1(20), S => CTRL, Z => OUT1(20)
                           );
   U22 : MUX2_X1 port map( A => IN0(19), B => IN1(19), S => CTRL, Z => OUT1(19)
                           );
   U1 : MUX2_X1 port map( A => IN0(13), B => IN1(13), S => CTRL, Z => OUT1(13))
                           ;
   U2 : MUX2_X1 port map( A => IN0(17), B => IN1(17), S => CTRL, Z => OUT1(17))
                           ;
   U3 : MUX2_X1 port map( A => IN0(12), B => IN1(12), S => CTRL, Z => OUT1(12))
                           ;
   U4 : MUX2_X1 port map( A => IN0(18), B => IN1(18), S => CTRL, Z => OUT1(18))
                           ;
   U5 : MUX2_X1 port map( A => IN0(14), B => IN1(14), S => CTRL, Z => OUT1(14))
                           ;
   U6 : MUX2_X1 port map( A => IN0(15), B => IN1(15), S => CTRL, Z => OUT1(15))
                           ;
   U7 : MUX2_X2 port map( A => IN0(27), B => IN1(27), S => CTRL, Z => OUT1(27))
                           ;
   U10 : MUX2_X2 port map( A => IN0(16), B => IN1(16), S => CTRL, Z => OUT1(16)
                           );
   U13 : MUX2_X1 port map( A => IN0(8), B => IN1(8), S => CTRL, Z => OUT1(8));
   U15 : MUX2_X1 port map( A => IN0(10), B => IN1(10), S => CTRL, Z => OUT1(10)
                           );
   U17 : MUX2_X1 port map( A => IN0(4), B => IN1(4), S => CTRL, Z => OUT1(4));
   U21 : MUX2_X2 port map( A => IN0(23), B => IN1(23), S => CTRL, Z => OUT1(23)
                           );
   U23 : NAND2_X1 port map( A1 => n16, A2 => n17, ZN => OUT1(6));
   U24 : NAND2_X1 port map( A1 => n20, A2 => n21, ZN => OUT1(7));
   U25 : NAND2_X1 port map( A1 => n18, A2 => n19, ZN => OUT1(0));
   U26 : MUX2_X1 port map( A => IN0(3), B => IN1(3), S => CTRL, Z => OUT1(3));
   U27 : NAND2_X1 port map( A1 => IN0(6), A2 => n15, ZN => n16);
   U28 : NAND2_X1 port map( A1 => IN1(6), A2 => CTRL, ZN => n17);
   U29 : INV_X1 port map( A => CTRL, ZN => n15);
   U30 : MUX2_X2 port map( A => IN0(2), B => IN1(2), S => CTRL, Z => OUT1(2));
   U31 : MUX2_X1 port map( A => IN0(1), B => IN1(1), S => CTRL, Z => OUT1(1));
   U32 : MUX2_X1 port map( A => IN0(5), B => IN1(5), S => CTRL, Z => OUT1(5));
   U33 : MUX2_X1 port map( A => IN0(25), B => IN1(25), S => CTRL, Z => OUT1(25)
                           );
   U34 : MUX2_X1 port map( A => IN0(11), B => IN1(11), S => CTRL, Z => OUT1(11)
                           );
   U35 : NAND2_X1 port map( A1 => CTRL, A2 => IN1(7), ZN => n21);
   U36 : NAND2_X1 port map( A1 => IN1(0), A2 => CTRL, ZN => n19);
   U37 : NAND2_X1 port map( A1 => IN0(0), A2 => n15, ZN => n18);
   U38 : NAND2_X1 port map( A1 => IN0(7), A2 => n15, ZN => n20);
   U39 : MUX2_X1 port map( A => IN0(9), B => IN1(9), S => CTRL, Z => OUT1(9));

end SYN_Bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity ff32_en_SIZE13 is

   port( D : in std_logic_vector (12 downto 0);  en, clk, rst : in std_logic;  
         Q : out std_logic_vector (12 downto 0));

end ff32_en_SIZE13;

architecture SYN_behavioral of ff32_en_SIZE13 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X2
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   signal Q_12_port, Q_11_port, Q_10_port, Q_9_port, Q_8_port, Q_7_port, 
      Q_6_port, Q_5_port, Q_4_port, Q_3_port, Q_2_port, Q_0_port, n27, n28, n29
      , n30, n31, n32, n33, n34, n35, n36, n37, n38, n40, n1, n2, Q_1_port, 
      net645036, net645037, net645038, net645039, net645040, net645041, 
      net645042, net645043, net645044, net645045, n5, n6, n7, n8, n9, n10, n11,
      n12, n13, n14, n15, n16, n18, net684300 : std_logic;

begin
   Q <= ( Q_12_port, Q_11_port, Q_10_port, Q_9_port, Q_8_port, Q_7_port, 
      Q_6_port, Q_5_port, Q_4_port, Q_3_port, Q_2_port, Q_1_port, Q_0_port );
   
   Q_reg_12_inst : DFFR_X1 port map( D => n40, CK => clk, RN => n18, Q => 
                           Q_12_port, QN => net645045);
   Q_reg_11_inst : DFFR_X1 port map( D => n38, CK => clk, RN => n18, Q => 
                           Q_11_port, QN => net645044);
   Q_reg_10_inst : DFFR_X1 port map( D => n37, CK => clk, RN => n18, Q => 
                           Q_10_port, QN => net645043);
   Q_reg_8_inst : DFFR_X1 port map( D => n35, CK => clk, RN => n18, Q => 
                           Q_8_port, QN => net645042);
   Q_reg_7_inst : DFFR_X1 port map( D => n34, CK => clk, RN => n18, Q => 
                           Q_7_port, QN => net645041);
   Q_reg_5_inst : DFFR_X1 port map( D => n32, CK => clk, RN => n18, Q => 
                           Q_5_port, QN => net645040);
   Q_reg_4_inst : DFFR_X1 port map( D => n31, CK => clk, RN => n18, Q => 
                           Q_4_port, QN => net645039);
   Q_reg_3_inst : DFFR_X1 port map( D => n30, CK => clk, RN => n18, Q => 
                           Q_3_port, QN => net645038);
   Q_reg_2_inst : DFFR_X1 port map( D => n29, CK => clk, RN => n18, Q => 
                           Q_2_port, QN => net645037);
   Q_reg_1_inst : DFFR_X1 port map( D => n28, CK => clk, RN => n18, Q => 
                           Q_1_port, QN => net684300);
   Q_reg_0_inst : DFFR_X1 port map( D => n27, CK => clk, RN => n18, Q => 
                           Q_0_port, QN => net645036);
   U27 : MUX2_X1 port map( A => Q_1_port, B => D(1), S => en, Z => n28);
   Q_reg_6_inst : DFFR_X1 port map( D => n33, CK => clk, RN => n18, Q => 
                           Q_6_port, QN => n1);
   U8 : NAND2_X1 port map( A1 => en, A2 => D(10), ZN => n7);
   U7 : OAI21_X1 port map( B1 => en, B2 => net645043, A => n7, ZN => n37);
   U6 : NAND2_X1 port map( A1 => en, A2 => D(11), ZN => n6);
   U5 : OAI21_X1 port map( B1 => en, B2 => net645044, A => n6, ZN => n38);
   U3 : NAND2_X1 port map( A1 => en, A2 => D(12), ZN => n5);
   U2 : OAI21_X1 port map( B1 => en, B2 => net645045, A => n5, ZN => n40);
   U12 : NAND2_X1 port map( A1 => en, A2 => D(8), ZN => n9);
   U11 : OAI21_X1 port map( B1 => en, B2 => net645042, A => n9, ZN => n35);
   U10 : NAND2_X1 port map( A1 => en, A2 => D(9), ZN => n8);
   U9 : OAI21_X1 port map( B1 => en, B2 => n2, A => n8, ZN => n36);
   U24 : NAND2_X1 port map( A1 => en, A2 => D(2), ZN => n15);
   U23 : OAI21_X1 port map( B1 => en, B2 => net645037, A => n15, ZN => n29);
   U22 : NAND2_X1 port map( A1 => en, A2 => D(3), ZN => n14);
   U21 : OAI21_X1 port map( B1 => en, B2 => net645038, A => n14, ZN => n30);
   U16 : NAND2_X1 port map( A1 => en, A2 => D(6), ZN => n11);
   U15 : OAI21_X1 port map( B1 => en, B2 => n1, A => n11, ZN => n33);
   U14 : NAND2_X1 port map( A1 => en, A2 => D(7), ZN => n10);
   U13 : OAI21_X1 port map( B1 => en, B2 => net645041, A => n10, ZN => n34);
   U18 : NAND2_X1 port map( A1 => en, A2 => D(5), ZN => n12);
   U17 : OAI21_X1 port map( B1 => en, B2 => net645040, A => n12, ZN => n32);
   U26 : NAND2_X1 port map( A1 => en, A2 => D(0), ZN => n16);
   U25 : OAI21_X1 port map( B1 => en, B2 => net645036, A => n16, ZN => n27);
   U20 : NAND2_X1 port map( A1 => en, A2 => D(4), ZN => n13);
   U19 : OAI21_X1 port map( B1 => en, B2 => net645039, A => n13, ZN => n31);
   Q_reg_9_inst : DFFR_X2 port map( D => n36, CK => clk, RN => n18, Q => 
                           Q_9_port, QN => n2);
   U4 : INV_X1 port map( A => rst, ZN => n18);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity ff32_en_SIZE5_3 is

   port( D : in std_logic_vector (4 downto 0);  en, clk, rst : in std_logic;  Q
         : out std_logic_vector (4 downto 0));

end ff32_en_SIZE5_3;

architecture SYN_behavioral of ff32_en_SIZE5_3 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n3, n4, n5, n6, net645267, net645268, net645269, net645270, 
      net645271, n8, n9, n10, n11, n12, n13 : std_logic;

begin
   
   Q_reg_4_inst : DFFR_X1 port map( D => n1, CK => clk, RN => n13, Q => Q(4), 
                           QN => net645271);
   Q_reg_3_inst : DFFR_X1 port map( D => n3, CK => clk, RN => n13, Q => Q(3), 
                           QN => net645270);
   Q_reg_2_inst : DFFR_X1 port map( D => n4, CK => clk, RN => n13, Q => Q(2), 
                           QN => net645269);
   Q_reg_0_inst : DFFR_X1 port map( D => n6, CK => clk, RN => n13, Q => Q(0), 
                           QN => net645267);
   Q_reg_1_inst : DFFR_X1 port map( D => n5, CK => clk, RN => n13, Q => Q(1), 
                           QN => net645268);
   U7 : NAND2_X1 port map( A1 => en, A2 => D(2), ZN => n10);
   U6 : OAI21_X1 port map( B1 => en, B2 => net645269, A => n10, ZN => n4);
   U9 : NAND2_X1 port map( A1 => en, A2 => D(3), ZN => n11);
   U8 : OAI21_X1 port map( B1 => en, B2 => net645270, A => n11, ZN => n3);
   U12 : NAND2_X1 port map( A1 => en, A2 => D(4), ZN => n12);
   U11 : OAI21_X1 port map( B1 => en, B2 => net645271, A => n12, ZN => n1);
   U5 : NAND2_X1 port map( A1 => en, A2 => D(1), ZN => n9);
   U4 : OAI21_X1 port map( B1 => en, B2 => net645268, A => n9, ZN => n5);
   U3 : NAND2_X1 port map( A1 => en, A2 => D(0), ZN => n8);
   U2 : OAI21_X1 port map( B1 => en, B2 => net645267, A => n8, ZN => n6);
   U10 : INV_X1 port map( A => rst, ZN => n13);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity ff32_en_SIZE5_0 is

   port( D : in std_logic_vector (4 downto 0);  en, clk, rst : in std_logic;  Q
         : out std_logic_vector (4 downto 0));

end ff32_en_SIZE5_0;

architecture SYN_behavioral of ff32_en_SIZE5_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n11, n12, n13, n14, n16, net645031, net645032, net645033, net645034, 
      net645035, n2, n3, n4, n5, n6, n7 : std_logic;

begin
   
   Q_reg_4_inst : DFFR_X1 port map( D => n16, CK => clk, RN => n7, Q => Q(4), 
                           QN => net645035);
   Q_reg_3_inst : DFFR_X1 port map( D => n14, CK => clk, RN => n7, Q => Q(3), 
                           QN => net645034);
   Q_reg_2_inst : DFFR_X1 port map( D => n13, CK => clk, RN => n7, Q => Q(2), 
                           QN => net645033);
   Q_reg_1_inst : DFFR_X1 port map( D => n12, CK => clk, RN => n7, Q => Q(1), 
                           QN => net645032);
   Q_reg_0_inst : DFFR_X1 port map( D => n11, CK => clk, RN => n7, Q => Q(0), 
                           QN => net645031);
   U10 : NAND2_X1 port map( A1 => en, A2 => D(1), ZN => n5);
   U9 : OAI21_X1 port map( B1 => en, B2 => net645032, A => n5, ZN => n12);
   U8 : NAND2_X1 port map( A1 => en, A2 => D(2), ZN => n4);
   U7 : OAI21_X1 port map( B1 => en, B2 => net645033, A => n4, ZN => n13);
   U6 : NAND2_X1 port map( A1 => en, A2 => D(3), ZN => n3);
   U5 : OAI21_X1 port map( B1 => en, B2 => net645034, A => n3, ZN => n14);
   U12 : NAND2_X1 port map( A1 => en, A2 => D(0), ZN => n6);
   U11 : OAI21_X1 port map( B1 => en, B2 => net645031, A => n6, ZN => n11);
   U3 : NAND2_X1 port map( A1 => en, A2 => D(4), ZN => n2);
   U2 : OAI21_X1 port map( B1 => en, B2 => net645035, A => n2, ZN => n16);
   U4 : INV_X1 port map( A => rst, ZN => n7);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity ff32_en_SIZE32_0 is

   port( D : in std_logic_vector (31 downto 0);  en, clk, rst : in std_logic;  
         Q : out std_logic_vector (31 downto 0));

end ff32_en_SIZE32_0;

architecture SYN_behavioral of ff32_en_SIZE32_0 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
      n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93
      , n94, n95, n97, net645107, net645108, net645109, net645110, net645111, 
      net645112, net645113, net645114, net645115, net645116, net645117, 
      net645118, net645119, net645120, net645121, net645122, net645123, 
      net645124, net645125, net645126, net645127, net645128, net645129, 
      net645130, net645131, net645132, net645133, net645134, net645135, 
      net645136, net645137, net645138, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11
      , n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, 
      n26, n27, n28, n29, n30, n31, n32, n33, n36, n37, n38 : std_logic;

begin
   
   Q_reg_31_inst : DFFR_X1 port map( D => n97, CK => clk, RN => n38, Q => Q(31)
                           , QN => net645138);
   Q_reg_30_inst : DFFR_X1 port map( D => n95, CK => clk, RN => n38, Q => Q(30)
                           , QN => net645137);
   Q_reg_29_inst : DFFR_X1 port map( D => n94, CK => clk, RN => n38, Q => Q(29)
                           , QN => net645136);
   Q_reg_28_inst : DFFR_X1 port map( D => n93, CK => clk, RN => n38, Q => Q(28)
                           , QN => net645135);
   Q_reg_27_inst : DFFR_X1 port map( D => n92, CK => clk, RN => n38, Q => Q(27)
                           , QN => net645134);
   Q_reg_26_inst : DFFR_X1 port map( D => n91, CK => clk, RN => n38, Q => Q(26)
                           , QN => net645133);
   Q_reg_25_inst : DFFR_X1 port map( D => n90, CK => clk, RN => n38, Q => Q(25)
                           , QN => net645132);
   Q_reg_24_inst : DFFR_X1 port map( D => n89, CK => clk, RN => n38, Q => Q(24)
                           , QN => net645131);
   Q_reg_23_inst : DFFR_X1 port map( D => n88, CK => clk, RN => n38, Q => Q(23)
                           , QN => net645130);
   Q_reg_22_inst : DFFR_X1 port map( D => n87, CK => clk, RN => n38, Q => Q(22)
                           , QN => net645129);
   Q_reg_21_inst : DFFR_X1 port map( D => n86, CK => clk, RN => n38, Q => Q(21)
                           , QN => net645128);
   Q_reg_19_inst : DFFR_X1 port map( D => n84, CK => clk, RN => n38, Q => Q(19)
                           , QN => net645127);
   Q_reg_18_inst : DFFR_X1 port map( D => n83, CK => clk, RN => n38, Q => Q(18)
                           , QN => net645126);
   Q_reg_17_inst : DFFR_X1 port map( D => n82, CK => clk, RN => n38, Q => Q(17)
                           , QN => net645125);
   Q_reg_16_inst : DFFR_X1 port map( D => n81, CK => clk, RN => n38, Q => Q(16)
                           , QN => net645124);
   Q_reg_15_inst : DFFR_X1 port map( D => n80, CK => clk, RN => n38, Q => Q(15)
                           , QN => net645123);
   Q_reg_14_inst : DFFR_X1 port map( D => n79, CK => clk, RN => n38, Q => Q(14)
                           , QN => net645122);
   Q_reg_13_inst : DFFR_X1 port map( D => n78, CK => clk, RN => n38, Q => Q(13)
                           , QN => net645121);
   Q_reg_12_inst : DFFR_X1 port map( D => n77, CK => clk, RN => n38, Q => Q(12)
                           , QN => net645120);
   Q_reg_11_inst : DFFR_X1 port map( D => n76, CK => clk, RN => n38, Q => Q(11)
                           , QN => net645119);
   Q_reg_10_inst : DFFR_X1 port map( D => n75, CK => clk, RN => n38, Q => Q(10)
                           , QN => net645118);
   Q_reg_9_inst : DFFR_X1 port map( D => n74, CK => clk, RN => n38, Q => Q(9), 
                           QN => net645117);
   Q_reg_8_inst : DFFR_X1 port map( D => n73, CK => clk, RN => n38, Q => Q(8), 
                           QN => net645116);
   Q_reg_7_inst : DFFR_X1 port map( D => n72, CK => clk, RN => n38, Q => Q(7), 
                           QN => net645115);
   Q_reg_6_inst : DFFR_X1 port map( D => n71, CK => clk, RN => n38, Q => Q(6), 
                           QN => net645114);
   Q_reg_5_inst : DFFR_X1 port map( D => n70, CK => clk, RN => n38, Q => Q(5), 
                           QN => net645113);
   Q_reg_4_inst : DFFR_X1 port map( D => n69, CK => clk, RN => n38, Q => Q(4), 
                           QN => net645112);
   Q_reg_3_inst : DFFR_X1 port map( D => n68, CK => clk, RN => n38, Q => Q(3), 
                           QN => net645111);
   Q_reg_2_inst : DFFR_X1 port map( D => n67, CK => clk, RN => n38, Q => Q(2), 
                           QN => net645110);
   Q_reg_1_inst : DFFR_X1 port map( D => n66, CK => clk, RN => n38, Q => Q(1), 
                           QN => net645109);
   Q_reg_0_inst : DFFR_X1 port map( D => n65, CK => clk, RN => n38, Q => Q(0), 
                           QN => net645108);
   Q_reg_20_inst : DFFR_X1 port map( D => n85, CK => clk, RN => n38, Q => Q(20)
                           , QN => net645107);
   U39 : NAND2_X1 port map( A1 => n36, A2 => D(13), ZN => n20);
   U38 : OAI21_X1 port map( B1 => en, B2 => net645121, A => n20, ZN => n78);
   U37 : NAND2_X1 port map( A1 => n36, A2 => D(14), ZN => n19);
   U36 : OAI21_X1 port map( B1 => en, B2 => net645122, A => n19, ZN => n79);
   U45 : NAND2_X1 port map( A1 => n36, A2 => D(10), ZN => n23);
   U44 : OAI21_X1 port map( B1 => en, B2 => net645118, A => n23, ZN => n75);
   U43 : NAND2_X1 port map( A1 => n36, A2 => D(11), ZN => n22);
   U42 : OAI21_X1 port map( B1 => en, B2 => net645119, A => n22, ZN => n76);
   U59 : NAND2_X1 port map( A1 => n37, A2 => D(3), ZN => n30);
   U58 : OAI21_X1 port map( B1 => n36, B2 => net645111, A => n30, ZN => n68);
   U23 : NAND2_X1 port map( A1 => n37, A2 => D(21), ZN => n12);
   U22 : OAI21_X1 port map( B1 => n36, B2 => net645128, A => n12, ZN => n86);
   U57 : NAND2_X1 port map( A1 => n37, A2 => D(4), ZN => n29);
   U56 : OAI21_X1 port map( B1 => n36, B2 => net645112, A => n29, ZN => n69);
   U55 : NAND2_X1 port map( A1 => en, A2 => D(5), ZN => n28);
   U54 : OAI21_X1 port map( B1 => n36, B2 => net645113, A => n28, ZN => n70);
   U61 : NAND2_X1 port map( A1 => n37, A2 => D(2), ZN => n31);
   U60 : OAI21_X1 port map( B1 => n36, B2 => net645110, A => n31, ZN => n67);
   U49 : NAND2_X1 port map( A1 => en, A2 => D(8), ZN => n25);
   U48 : OAI21_X1 port map( B1 => n36, B2 => net645116, A => n25, ZN => n73);
   U53 : NAND2_X1 port map( A1 => n37, A2 => D(6), ZN => n27);
   U52 : OAI21_X1 port map( B1 => n36, B2 => net645114, A => n27, ZN => n71);
   U25 : NAND2_X1 port map( A1 => en, A2 => D(20), ZN => n13);
   U24 : OAI21_X1 port map( B1 => n37, B2 => net645107, A => n13, ZN => n85);
   U27 : NAND2_X1 port map( A1 => en, A2 => D(19), ZN => n14);
   U26 : OAI21_X1 port map( B1 => en, B2 => net645127, A => n14, ZN => n84);
   U47 : NAND2_X1 port map( A1 => en, A2 => D(9), ZN => n24);
   U46 : OAI21_X1 port map( B1 => en, B2 => net645117, A => n24, ZN => n74);
   U51 : NAND2_X1 port map( A1 => en, A2 => D(7), ZN => n26);
   U50 : OAI21_X1 port map( B1 => en, B2 => net645115, A => n26, ZN => n72);
   U19 : NAND2_X1 port map( A1 => n37, A2 => D(23), ZN => n10);
   U18 : OAI21_X1 port map( B1 => en, B2 => net645130, A => n10, ZN => n88);
   U9 : NAND2_X1 port map( A1 => n37, A2 => D(28), ZN => n5);
   U8 : OAI21_X1 port map( B1 => en, B2 => net645135, A => n5, ZN => n93);
   U7 : NAND2_X1 port map( A1 => n37, A2 => D(29), ZN => n4);
   U6 : OAI21_X1 port map( B1 => en, B2 => net645136, A => n4, ZN => n94);
   U41 : NAND2_X1 port map( A1 => en, A2 => D(12), ZN => n21);
   U40 : OAI21_X1 port map( B1 => en, B2 => net645120, A => n21, ZN => n77);
   U21 : NAND2_X1 port map( A1 => en, A2 => D(22), ZN => n11);
   U20 : OAI21_X1 port map( B1 => en, B2 => net645129, A => n11, ZN => n87);
   U29 : NAND2_X1 port map( A1 => en, A2 => D(18), ZN => n15);
   U28 : OAI21_X1 port map( B1 => en, B2 => net645126, A => n15, ZN => n83);
   U11 : NAND2_X1 port map( A1 => n37, A2 => D(27), ZN => n6);
   U10 : OAI21_X1 port map( B1 => en, B2 => net645134, A => n6, ZN => n92);
   U31 : NAND2_X1 port map( A1 => en, A2 => D(17), ZN => n16);
   U30 : OAI21_X1 port map( B1 => en, B2 => net645125, A => n16, ZN => n82);
   U35 : NAND2_X1 port map( A1 => en, A2 => D(15), ZN => n18);
   U34 : OAI21_X1 port map( B1 => en, B2 => net645123, A => n18, ZN => n80);
   U33 : NAND2_X1 port map( A1 => en, A2 => D(16), ZN => n17);
   U32 : OAI21_X1 port map( B1 => en, B2 => net645124, A => n17, ZN => n81);
   U15 : NAND2_X1 port map( A1 => n37, A2 => D(25), ZN => n8);
   U14 : OAI21_X1 port map( B1 => en, B2 => net645132, A => n8, ZN => n90);
   U13 : NAND2_X1 port map( A1 => n37, A2 => D(26), ZN => n7);
   U12 : OAI21_X1 port map( B1 => en, B2 => net645133, A => n7, ZN => n91);
   U17 : NAND2_X1 port map( A1 => n37, A2 => D(24), ZN => n9);
   U16 : OAI21_X1 port map( B1 => en, B2 => net645131, A => n9, ZN => n89);
   U63 : NAND2_X1 port map( A1 => en, A2 => D(1), ZN => n32);
   U62 : OAI21_X1 port map( B1 => n36, B2 => net645109, A => n32, ZN => n66);
   U65 : NAND2_X1 port map( A1 => en, A2 => D(0), ZN => n33);
   U64 : OAI21_X1 port map( B1 => n36, B2 => net645108, A => n33, ZN => n65);
   U5 : NAND2_X1 port map( A1 => en, A2 => D(30), ZN => n3);
   U4 : OAI21_X1 port map( B1 => en, B2 => net645137, A => n3, ZN => n95);
   U3 : NAND2_X1 port map( A1 => en, A2 => D(31), ZN => n2);
   U2 : OAI21_X1 port map( B1 => en, B2 => net645138, A => n2, ZN => n97);
   U66 : INV_X2 port map( A => rst, ZN => n38);
   U67 : BUF_X1 port map( A => en, Z => n37);
   U68 : BUF_X1 port map( A => en, Z => n36);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity alu_ctrl is

   port( OP : in std_logic_vector (0 to 4);  ALU_WORD : out std_logic_vector 
         (12 downto 0));

end alu_ctrl;

architecture SYN_bhe of alu_ctrl is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI33_X1
      port( A1, A2, A3, B1, B2, B3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal ALU_WORD_12_port, ALU_WORD_11_port, ALU_WORD_10_port, ALU_WORD_9_port
      , ALU_WORD_8_port, ALU_WORD_7_port, ALU_WORD_6_port, ALU_WORD_5_port, 
      ALU_WORD_4_port, ALU_WORD_3_port, ALU_WORD_2_port, ALU_WORD_1_port, 
      ALU_WORD_0_port, N20, N21, N22, N23, N24, N25, N26, N27, N29, N30, N31, 
      N32, N33, n37, n12, n13, n14, n15, n16, n17, n18, n19, n20_port, n21_port
      , n22_port, n23_port, n24_port, n25_port, n26_port, n27_port, n28, 
      n29_port, n30_port, n31_port, n32_port, n33_port, n34, n35, n36, n38, n39
      , n40 : std_logic;

begin
   ALU_WORD <= ( ALU_WORD_12_port, ALU_WORD_11_port, ALU_WORD_10_port, 
      ALU_WORD_9_port, ALU_WORD_8_port, ALU_WORD_7_port, ALU_WORD_6_port, 
      ALU_WORD_5_port, ALU_WORD_4_port, ALU_WORD_3_port, ALU_WORD_2_port, 
      ALU_WORD_1_port, ALU_WORD_0_port );
   
   comp_sel_reg_2_inst : DLH_X1 port map( G => N32, D => N33, Q => 
                           ALU_WORD_4_port);
   comp_sel_reg_1_inst : DLH_X1 port map( G => N32, D => N31, Q => 
                           ALU_WORD_3_port);
   comp_sel_reg_0_inst : DLH_X1 port map( G => N32, D => N30, Q => 
                           ALU_WORD_2_port);
   sign_to_booth_reg : DLH_X1 port map( G => N20, D => N21, Q => 
                           ALU_WORD_0_port);
   left_right_reg : DLH_X1 port map( G => N23, D => N22, Q => ALU_WORD_9_port);
   logic_arith_reg : DLH_X1 port map( G => N23, D => N24, Q => ALU_WORD_8_port)
                           ;
   sign_to_adder_reg : DLH_X1 port map( G => N25, D => N26, Q => 
                           ALU_WORD_7_port);
   lu_ctrl_reg_1_inst : DLL_X1 port map( D => N29, GN => n37, Q => 
                           ALU_WORD_6_port);
   lu_ctrl_reg_0_inst : DLL_X1 port map( D => N27, GN => n37, Q => 
                           ALU_WORD_5_port);
   U43 : NAND3_X1 port map( A1 => n21_port, A2 => n37, A3 => n27_port, ZN => 
                           ALU_WORD_10_port);
   U44 : NAND3_X1 port map( A1 => n17, A2 => n29_port, A3 => OP(2), ZN => n13);
   U45 : OAI33_X1 port map( A1 => n14, A2 => n17, A3 => n19, B1 => n26_port, B2
                           => n30_port, B3 => OP(1), ZN => n25_port);
   U46 : NAND3_X1 port map( A1 => n15, A2 => OP(4), A3 => OP(3), ZN => n12);
   U47 : NAND3_X1 port map( A1 => OP(3), A2 => n17, A3 => n15, ZN => n35);
   U42 : NAND2_X1 port map( A1 => OP(0), A2 => OP(1), ZN => n16);
   U36 : NOR2_X1 port map( A1 => OP(2), A2 => OP(3), ZN => n33_port);
   U35 : NAND2_X1 port map( A1 => OP(4), A2 => n33_port, ZN => n18);
   U34 : NOR2_X1 port map( A1 => n18, A2 => n16, ZN => n39);
   U32 : NAND2_X1 port map( A1 => OP(2), A2 => OP(3), ZN => n19);
   U31 : NAND2_X1 port map( A1 => n33_port, A2 => n17, ZN => n26_port);
   U28 : AOI221_X1 port map( B1 => n13, B2 => n30_port, C1 => n13, C2 => n12, A
                           => n31_port, ZN => n40);
   U26 : AOI211_X1 port map( C1 => n38, C2 => n34, A => n39, B => N30, ZN => 
                           n36);
   U25 : OAI221_X1 port map( B1 => n17, B2 => n29_port, C1 => OP(4), C2 => 
                           OP(3), A => OP(2), ZN => n32_port);
   U23 : OAI211_X1 port map( C1 => n16, C2 => n35, A => n36, B => n23_port, ZN 
                           => N32);
   U21 : NOR2_X1 port map( A1 => n14, A2 => n35, ZN => N29);
   U20 : AOI21_X1 port map( B1 => n33_port, B2 => n34, A => N29, ZN => n37);
   U19 : NOR2_X1 port map( A1 => n16, A2 => n32_port, ZN => ALU_WORD_1_port);
   U16 : NOR3_X1 port map( A1 => OP(2), A2 => n29_port, A3 => n20_port, ZN => 
                           N22);
   U14 : OAI21_X1 port map( B1 => n18, B2 => n20_port, A => n28, ZN => N23);
   U12 : OAI21_X1 port map( B1 => n26_port, B2 => n20_port, A => n27_port, ZN 
                           => ALU_WORD_12_port);
   U4 : NOR2_X1 port map( A1 => n14, A2 => n18, ZN => N27);
   U7 : NOR2_X1 port map( A1 => n12, A2 => n20_port, ZN => N24);
   U5 : OAI21_X1 port map( B1 => n19, B2 => n20_port, A => n21_port, ZN => N26)
                           ;
   U2 : AOI21_X1 port map( B1 => n12, B2 => n13, A => n14, ZN => N33);
   U8 : OAI211_X1 port map( C1 => n19, C2 => n22_port, A => n23_port, B => 
                           n24_port, ZN => N21);
   U3 : AOI221_X1 port map( B1 => OP(2), B2 => n14, C1 => n15, C2 => n16, A => 
                           n17, ZN => N31);
   U6 : OAI21_X1 port map( B1 => n15, B2 => n20_port, A => n21_port, ZN => N25)
                           ;
   U37 : NOR2_X1 port map( A1 => n31_port, A2 => OP(0), ZN => n34);
   U17 : NAND2_X1 port map( A1 => n30_port, A2 => n31_port, ZN => n20_port);
   U29 : INV_X1 port map( A => OP(3), ZN => n29_port);
   U41 : INV_X1 port map( A => OP(4), ZN => n17);
   U40 : INV_X1 port map( A => OP(2), ZN => n15);
   U30 : INV_X1 port map( A => OP(0), ZN => n30_port);
   U38 : INV_X1 port map( A => OP(1), ZN => n31_port);
   U10 : OR2_X1 port map( A1 => OP(4), A2 => n16, ZN => n22_port);
   U39 : INV_X1 port map( A => n12, ZN => n38);
   U33 : INV_X1 port map( A => n34, ZN => n14);
   U18 : INV_X1 port map( A => ALU_WORD_1_port, ZN => n27_port);
   U24 : OR2_X1 port map( A1 => n14, A2 => n32_port, ZN => n23_port);
   U15 : INV_X1 port map( A => N22, ZN => n28);
   U9 : INV_X1 port map( A => n25_port, ZN => n24_port);
   U27 : OR2_X1 port map( A1 => n25_port, A2 => n40, ZN => N30);
   U13 : OR2_X1 port map( A1 => N32, A2 => N23, ZN => ALU_WORD_11_port);
   U11 : OR2_X1 port map( A1 => N32, A2 => ALU_WORD_12_port, ZN => N20);
   U22 : INV_X1 port map( A => N32, ZN => n21_port);

end SYN_bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity cw_mem_MICROCODE_MEM_SIZE64_OP_CODE_SIZE6_CW_SIZE13 is

   port( OPCODE_IN : in std_logic_vector (5 downto 0);  CW_OUT : out 
         std_logic_vector (12 downto 0));

end cw_mem_MICROCODE_MEM_SIZE64_OP_CODE_SIZE6_CW_SIZE13;

architecture SYN_bhe of cw_mem_MICROCODE_MEM_SIZE64_OP_CODE_SIZE6_CW_SIZE13 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal CW_OUT_12_port, CW_OUT_11_port, CW_OUT_10_port, CW_OUT_9_port, 
      CW_OUT_8_port, CW_OUT_7_port, CW_OUT_6_port, CW_OUT_4, CW_OUT_3, CW_OUT_2
      , CW_OUT_1, CW_OUT_0, n9, n10, n11, n12, n13, n14, n15, n16, n19, n20, 
      n21, n22, n23, n24, n25, n26, n27, n28, n29, n17, n30, n31, n32, n33, n34
      , n35, n36, n37, n_1187 : std_logic;

begin
   CW_OUT <= ( CW_OUT_12_port, CW_OUT_11_port, CW_OUT_10_port, CW_OUT_9_port, 
      CW_OUT_8_port, CW_OUT_7_port, CW_OUT_6_port, n_1187, CW_OUT_4, CW_OUT_3, 
      CW_OUT_2, CW_OUT_1, CW_OUT_0 );
   
   U29 : NAND2_X1 port map( A1 => n29, A2 => n28, ZN => n14);
   U11 : AOI21_X1 port map( B1 => n20, B2 => n26, A => CW_OUT_7_port, ZN => n25
                           );
   U19 : INV_X1 port map( A => OPCODE_IN(0), ZN => n12);
   U2 : OR3_X1 port map( A1 => CW_OUT_1, A2 => CW_OUT_4, A3 => n13, ZN => 
                           CW_OUT_0);
   U9 : OR2_X1 port map( A1 => CW_OUT_3, A2 => n13, ZN => CW_OUT_6_port);
   U1 : OAI21_X1 port map( B1 => n14, B2 => n30, A => n35, ZN => CW_OUT_11_port
                           );
   U3 : OR2_X1 port map( A1 => n22, A2 => n27, ZN => n30);
   U4 : OAI221_X1 port map( B1 => n22, B2 => n23, C1 => n22, C2 => n24, A => 
                           n25, ZN => n13);
   U5 : NAND2_X1 port map( A1 => n16, A2 => n21, ZN => CW_OUT_12_port);
   U6 : CLKBUF_X1 port map( A => n21, Z => n35);
   U7 : OR2_X1 port map( A1 => n33, A2 => CW_OUT_12_port, ZN => CW_OUT_9_port);
   U8 : NOR2_X1 port map( A1 => n11, A2 => n31, ZN => CW_OUT_10_port);
   U10 : NOR2_X1 port map( A1 => n10, A2 => OPCODE_IN(5), ZN => n20);
   U12 : INV_X1 port map( A => OPCODE_IN(1), ZN => n27);
   U13 : NAND2_X1 port map( A1 => OPCODE_IN(1), A2 => n19, ZN => n11);
   U14 : INV_X1 port map( A => OPCODE_IN(4), ZN => n22);
   U15 : NOR2_X1 port map( A1 => OPCODE_IN(4), A2 => OPCODE_IN(2), ZN => n19);
   U16 : INV_X1 port map( A => OPCODE_IN(3), ZN => n10);
   U17 : INV_X1 port map( A => OPCODE_IN(2), ZN => n28);
   U18 : OR2_X1 port map( A1 => OPCODE_IN(3), A2 => OPCODE_IN(5), ZN => n37);
   U20 : INV_X1 port map( A => CW_OUT_10_port, ZN => n16);
   U21 : BUF_X1 port map( A => n11, Z => n36);
   U22 : OR3_X2 port map( A1 => n15, A2 => n28, A3 => n37, ZN => n21);
   U23 : OR2_X1 port map( A1 => OPCODE_IN(5), A2 => OPCODE_IN(3), ZN => n31);
   U24 : NOR2_X1 port map( A1 => OPCODE_IN(2), A2 => OPCODE_IN(4), ZN => n32);
   U25 : NAND2_X1 port map( A1 => n32, A2 => n20, ZN => n17);
   U26 : NOR2_X1 port map( A1 => OPCODE_IN(0), A2 => n17, ZN => n33);
   U27 : NAND2_X1 port map( A1 => n22, A2 => n27, ZN => n34);
   U28 : OAI22_X1 port map( A1 => n14, A2 => n34, B1 => n16, B2 => n12, ZN => 
                           CW_OUT_4);
   U30 : INV_X1 port map( A => OPCODE_IN(5), ZN => n9);
   U31 : NOR2_X1 port map( A1 => OPCODE_IN(5), A2 => OPCODE_IN(3), ZN => n29);
   U32 : NOR4_X1 port map( A1 => n9, A2 => n10, A3 => n36, A4 => n12, ZN => 
                           CW_OUT_2);
   U33 : NOR3_X1 port map( A1 => n9, A2 => n36, A3 => n12, ZN => CW_OUT_3);
   U34 : NOR4_X1 port map( A1 => OPCODE_IN(3), A2 => n9, A3 => n36, A4 => n12, 
                           ZN => CW_OUT_1);
   U35 : NOR2_X1 port map( A1 => n12, A2 => n35, ZN => CW_OUT_8_port);
   U36 : OAI221_X1 port map( B1 => OPCODE_IN(2), B2 => OPCODE_IN(1), C1 => n28,
                           C2 => n27, A => OPCODE_IN(3), ZN => n24);
   U37 : OAI211_X1 port map( C1 => OPCODE_IN(1), C2 => n12, A => n29, B => 
                           OPCODE_IN(2), ZN => n23);
   U38 : OAI211_X1 port map( C1 => OPCODE_IN(4), C2 => OPCODE_IN(0), A => 
                           OPCODE_IN(2), B => OPCODE_IN(1), ZN => n26);
   U39 : NOR3_X1 port map( A1 => n14, A2 => n27, A3 => n12, ZN => CW_OUT_7_port
                           );
   U40 : NAND2_X1 port map( A1 => n22, A2 => n27, ZN => n15);

end SYN_bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity stall_logic_FUNC_SIZE11_OP_CODE_SIZE6 is

   port( OPCODE_i : in std_logic_vector (5 downto 0);  FUNC_i : in 
         std_logic_vector (10 downto 0);  rA_i, rB_i, D1_i, D2_i : in 
         std_logic_vector (4 downto 0);  S_mem_LOAD_i, S_exe_LOAD_i : in 
         std_logic;  S_MUX_PC_BUS_i : in std_logic_vector (1 downto 0);  
         mispredict_i : in std_logic;  bubble_dec_o, bubble_exe_o, stall_exe_o,
         stall_dec_o, stall_btb_o, stall_fetch_o : out std_logic;  
         S_exe_WRITE_i_BAR : in std_logic);

end stall_logic_FUNC_SIZE11_OP_CODE_SIZE6;

architecture SYN_stall_logic_hw of stall_logic_FUNC_SIZE11_OP_CODE_SIZE6 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI33_X1
      port( A1, A2, A3, B1, B2, B3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal stall_fetch_o_port, n16, n27, n28, n29, n30, n31, n32, n33, n34, n41,
      n43, n44, n45, n46, n47, n48, n50, n51, n52, n53, n54, n55, n56, n42, n49
      , n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, 
      n71, n72, n73 : std_logic;

begin
   stall_fetch_o <= stall_fetch_o_port;
   
   U38 : OAI22_X1 port map( A1 => n54, A2 => D1_i(2), B1 => n55, B2 => D1_i(1),
                           ZN => n56);
   U37 : AOI221_X1 port map( B1 => n54, B2 => D1_i(2), C1 => D1_i(1), C2 => n55
                           , A => n56, ZN => n50);
   U34 : OAI22_X1 port map( A1 => n44, A2 => D1_i(3), B1 => n46, B2 => D1_i(4),
                           ZN => n53);
   U33 : AOI221_X1 port map( B1 => n44, B2 => D1_i(3), C1 => D1_i(4), C2 => n46
                           , A => n53, ZN => n51);
   U32 : XNOR2_X1 port map( A => rA_i(0), B => D1_i(0), ZN => n52);
   U12 : OAI22_X1 port map( A1 => n33, A2 => rB_i(2), B1 => n32, B2 => rB_i(1),
                           ZN => n34);
   U11 : AOI221_X1 port map( B1 => rB_i(1), B2 => n32, C1 => n33, C2 => rB_i(2)
                           , A => n34, ZN => n27);
   U8 : OAI22_X1 port map( A1 => n30, A2 => rB_i(3), B1 => n29, B2 => rB_i(4), 
                           ZN => n31);
   U7 : AOI221_X1 port map( B1 => rB_i(4), B2 => n29, C1 => n30, C2 => rB_i(3),
                           A => n31, ZN => n28);
   U2 : NOR2_X1 port map( A1 => stall_fetch_o_port, A2 => n16, ZN => 
                           bubble_dec_o);
   U40 : INV_X1 port map( A => rA_i(2), ZN => n54);
   U39 : INV_X1 port map( A => rA_i(1), ZN => n55);
   U36 : INV_X1 port map( A => rA_i(3), ZN => n44);
   U22 : INV_X1 port map( A => D2_i(2), ZN => n43);
   U9 : INV_X1 port map( A => D1_i(3), ZN => n30);
   U10 : INV_X1 port map( A => D1_i(4), ZN => n29);
   U13 : INV_X1 port map( A => D1_i(2), ZN => n33);
   U14 : INV_X1 port map( A => D1_i(1), ZN => n32);
   U35 : INV_X1 port map( A => rA_i(4), ZN => n46);
   U3 : INV_X1 port map( A => S_exe_LOAD_i, ZN => n42);
   U4 : NOR2_X1 port map( A1 => OPCODE_i(4), A2 => OPCODE_i(1), ZN => n49);
   U5 : INV_X1 port map( A => OPCODE_i(2), ZN => n57);
   U6 : NAND2_X1 port map( A1 => OPCODE_i(4), A2 => OPCODE_i(1), ZN => n58);
   U15 : OAI221_X1 port map( B1 => n57, B2 => OPCODE_i(0), C1 => n57, C2 => 
                           OPCODE_i(4), A => n58, ZN => n59);
   U16 : NOR4_X1 port map( A1 => n49, A2 => OPCODE_i(5), A3 => OPCODE_i(3), A4 
                           => n59, ZN => n60);
   U17 : NAND3_X1 port map( A1 => n50, A2 => n52, A3 => n51, ZN => n61);
   U18 : INV_X1 port map( A => n49, ZN => n62);
   U19 : AOI22_X1 port map( A1 => OPCODE_i(2), A2 => n62, B1 => n58, B2 => n57,
                           ZN => n63);
   U20 : INV_X1 port map( A => rA_i(1), ZN => n64);
   U21 : AOI22_X1 port map( A1 => n47, A2 => D2_i(0), B1 => n46, B2 => D2_i(4),
                           ZN => n65);
   U23 : OAI21_X1 port map( B1 => n64, B2 => D2_i(1), A => n65, ZN => n66);
   U24 : AOI211_X1 port map( C1 => n64, C2 => D2_i(1), A => n48, B => n66, ZN 
                           => n67);
   U25 : NAND3_X1 port map( A1 => n41, A2 => S_mem_LOAD_i, A3 => n67, ZN => n68
                           );
   U26 : OAI21_X1 port map( B1 => S_exe_WRITE_i_BAR, B2 => n61, A => n68, ZN =>
                           n69);
   U27 : XOR2_X1 port map( A => D1_i(0), B => rB_i(0), Z => n70);
   U28 : NAND4_X1 port map( A1 => S_exe_LOAD_i, A2 => n49, A3 => n28, A4 => n27
                           , ZN => n71);
   U29 : NOR4_X1 port map( A1 => OPCODE_i(0), A2 => OPCODE_i(2), A3 => n70, A4 
                           => n71, ZN => n72);
   U30 : AOI21_X1 port map( B1 => n63, B2 => n69, A => n72, ZN => n73);
   U31 : OAI33_X1 port map( A1 => n42, A2 => n60, A3 => n61, B1 => OPCODE_i(5),
                           B2 => n73, B3 => OPCODE_i(3), ZN => 
                           stall_fetch_o_port);
   U41 : INV_X1 port map( A => mispredict_i, ZN => n16);
   U42 : INV_X1 port map( A => rA_i(0), ZN => n47);
   U43 : AOI221_X1 port map( B1 => rA_i(2), B2 => n43, C1 => n44, C2 => D2_i(3)
                           , A => n45, ZN => n41);
   U44 : OAI22_X1 port map( A1 => n47, A2 => D2_i(0), B1 => n46, B2 => D2_i(4),
                           ZN => n48);
   U45 : OAI22_X1 port map( A1 => n44, A2 => D2_i(3), B1 => n43, B2 => rA_i(2),
                           ZN => n45);

end SYN_stall_logic_hw;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity mux41_MUX_SIZE32 is

   port( IN0, IN1, IN2, IN3 : in std_logic_vector (31 downto 0);  CTRL : in 
         std_logic_vector (1 downto 0);  OUT1 : out std_logic_vector (31 downto
         0));

end mux41_MUX_SIZE32;

architecture SYN_bhe of mux41_MUX_SIZE32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n5, n6, n7, n8, n9, n10, n11, n12, n13, n16, n17, n18, n19, 
      n20, n21, n24, n25, n28, n29, n30, n31, n34, n35, n36, n37, n44, n45, n46
      , n47, n60, n61, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, 
      n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91
      , n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, 
      n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, 
      n117, n118, n119, n120, n121, n122, n123, n124, n125, n126 : std_logic;

begin
   
   U61 : NAND2_X1 port map( A1 => n46, A2 => n47, ZN => OUT1(1));
   U1 : BUF_X1 port map( A => n6, Z => n71);
   U2 : BUF_X1 port map( A => n6, Z => n73);
   U3 : BUF_X2 port map( A => n6, Z => n72);
   U4 : AND2_X2 port map( A1 => n70, A2 => CTRL(0), ZN => n6);
   U5 : BUF_X1 port map( A => n7, Z => n119);
   U6 : BUF_X2 port map( A => n5, Z => n125);
   U7 : BUF_X2 port map( A => n7, Z => n121);
   U8 : BUF_X2 port map( A => n7, Z => n120);
   U9 : BUF_X2 port map( A => n6, Z => n123);
   U10 : NOR2_X1 port map( A1 => CTRL(0), A2 => n70, ZN => n5);
   U11 : NOR2_X1 port map( A1 => CTRL(0), A2 => n118, ZN => n7);
   U12 : BUF_X2 port map( A => n6, Z => n122);
   U13 : BUF_X2 port map( A => n5, Z => n126);
   U14 : BUF_X2 port map( A => n5, Z => n124);
   U15 : BUF_X1 port map( A => CTRL(1), Z => n118);
   U16 : NAND2_X1 port map( A1 => n126, A2 => IN2(28), ZN => n29);
   U17 : NAND2_X1 port map( A1 => n125, A2 => IN2(24), ZN => n37);
   U18 : NAND2_X1 port map( A1 => n126, A2 => IN2(20), ZN => n45);
   U19 : NAND3_X1 port map( A1 => n75, A2 => n74, A3 => n76, ZN => OUT1(12));
   U20 : NAND2_X1 port map( A1 => n6, A2 => IN1(12), ZN => n75);
   U21 : NAND2_X1 port map( A1 => n119, A2 => IN0(12), ZN => n76);
   U22 : NAND2_X1 port map( A1 => n125, A2 => IN2(12), ZN => n74);
   U23 : NAND3_X1 port map( A1 => n79, A2 => n78, A3 => n77, ZN => OUT1(29));
   U24 : NAND2_X1 port map( A1 => n123, A2 => IN1(29), ZN => n79);
   U25 : NAND2_X1 port map( A1 => n120, A2 => IN0(29), ZN => n78);
   U26 : NAND2_X1 port map( A1 => n125, A2 => IN2(29), ZN => n77);
   U27 : NAND3_X1 port map( A1 => n82, A2 => n81, A3 => n80, ZN => OUT1(26));
   U28 : NAND2_X1 port map( A1 => n72, A2 => IN1(26), ZN => n82);
   U29 : NAND2_X1 port map( A1 => n120, A2 => IN0(26), ZN => n81);
   U30 : NAND2_X1 port map( A1 => n126, A2 => IN2(26), ZN => n80);
   U31 : NAND3_X1 port map( A1 => n84, A2 => n83, A3 => n85, ZN => OUT1(14));
   U32 : NAND2_X1 port map( A1 => n72, A2 => IN1(14), ZN => n84);
   U33 : NAND2_X1 port map( A1 => n119, A2 => IN0(14), ZN => n85);
   U34 : NAND2_X1 port map( A1 => n124, A2 => IN2(14), ZN => n83);
   U35 : NAND3_X1 port map( A1 => n88, A2 => n87, A3 => n86, ZN => OUT1(18));
   U36 : NAND2_X1 port map( A1 => n123, A2 => IN1(18), ZN => n88);
   U37 : NAND2_X1 port map( A1 => n120, A2 => IN0(18), ZN => n87);
   U38 : NAND2_X1 port map( A1 => n124, A2 => IN2(18), ZN => n86);
   U39 : AOI22_X1 port map( A1 => n120, A2 => IN0(5), B1 => n73, B2 => IN1(5), 
                           ZN => n90);
   U40 : NAND2_X1 port map( A1 => n90, A2 => n89, ZN => OUT1(5));
   U41 : NAND2_X1 port map( A1 => n125, A2 => IN2(5), ZN => n89);
   U42 : NAND3_X1 port map( A1 => n93, A2 => n92, A3 => n91, ZN => OUT1(22));
   U43 : NAND2_X1 port map( A1 => n72, A2 => IN1(22), ZN => n93);
   U44 : NAND2_X1 port map( A1 => n120, A2 => IN0(22), ZN => n92);
   U45 : NAND2_X1 port map( A1 => n124, A2 => IN2(22), ZN => n91);
   U46 : NAND3_X1 port map( A1 => n95, A2 => n94, A3 => n96, ZN => OUT1(30));
   U47 : NAND2_X1 port map( A1 => n122, A2 => IN1(30), ZN => n95);
   U48 : NAND2_X1 port map( A1 => n120, A2 => IN0(30), ZN => n96);
   U49 : NAND2_X1 port map( A1 => n124, A2 => IN2(30), ZN => n94);
   U50 : NAND3_X1 port map( A1 => n98, A2 => n97, A3 => n99, ZN => OUT1(19));
   U51 : NAND2_X1 port map( A1 => n71, A2 => IN1(19), ZN => n98);
   U52 : NAND2_X1 port map( A1 => n120, A2 => IN0(19), ZN => n99);
   U53 : NAND2_X1 port map( A1 => n124, A2 => IN2(19), ZN => n97);
   U54 : NAND3_X1 port map( A1 => n101, A2 => n100, A3 => n102, ZN => OUT1(11))
                           ;
   U55 : NAND2_X1 port map( A1 => n71, A2 => IN1(11), ZN => n101);
   U56 : NAND2_X1 port map( A1 => n120, A2 => IN0(11), ZN => n102);
   U57 : NAND2_X1 port map( A1 => n125, A2 => IN2(11), ZN => n100);
   U58 : NAND3_X1 port map( A1 => n105, A2 => n104, A3 => n103, ZN => OUT1(17))
                           ;
   U59 : NAND2_X1 port map( A1 => n122, A2 => IN1(17), ZN => n105);
   U60 : NAND2_X1 port map( A1 => n120, A2 => IN0(17), ZN => n104);
   U62 : NAND2_X1 port map( A1 => n124, A2 => IN2(17), ZN => n103);
   U63 : NAND3_X1 port map( A1 => n107, A2 => n106, A3 => n108, ZN => OUT1(15))
                           ;
   U64 : NAND2_X1 port map( A1 => n122, A2 => IN1(15), ZN => n107);
   U65 : NAND2_X1 port map( A1 => n119, A2 => IN0(15), ZN => n108);
   U66 : NAND2_X1 port map( A1 => n125, A2 => IN2(15), ZN => n106);
   U67 : NAND3_X1 port map( A1 => n110, A2 => n109, A3 => n111, ZN => OUT1(21))
                           ;
   U68 : NAND2_X1 port map( A1 => n72, A2 => IN1(21), ZN => n110);
   U69 : NAND2_X1 port map( A1 => n119, A2 => IN0(21), ZN => n111);
   U70 : NAND2_X1 port map( A1 => n124, A2 => IN2(21), ZN => n109);
   U71 : NAND3_X1 port map( A1 => n114, A2 => n113, A3 => n112, ZN => OUT1(23))
                           ;
   U72 : NAND2_X1 port map( A1 => n123, A2 => IN1(23), ZN => n114);
   U73 : NAND2_X1 port map( A1 => n119, A2 => IN0(23), ZN => n113);
   U74 : NAND2_X1 port map( A1 => n125, A2 => IN2(23), ZN => n112);
   U75 : NAND3_X1 port map( A1 => n117, A2 => n116, A3 => n115, ZN => OUT1(16))
                           ;
   U76 : NAND2_X1 port map( A1 => n122, A2 => IN1(16), ZN => n117);
   U77 : NAND2_X1 port map( A1 => n120, A2 => IN0(16), ZN => n116);
   U78 : NAND2_X1 port map( A1 => n126, A2 => IN2(16), ZN => n115);
   U79 : NAND2_X1 port map( A1 => n66, A2 => n67, ZN => OUT1(10));
   U80 : NAND2_X1 port map( A1 => n60, A2 => n61, ZN => OUT1(13));
   U81 : AOI22_X1 port map( A1 => n71, A2 => IN1(9), B1 => n121, B2 => IN0(9), 
                           ZN => n2);
   U82 : AOI22_X1 port map( A1 => n123, A2 => IN1(4), B1 => n121, B2 => IN0(4),
                           ZN => n16);
   U83 : AOI22_X1 port map( A1 => n73, A2 => IN1(8), B1 => n121, B2 => IN0(8), 
                           ZN => n8);
   U84 : AOI22_X1 port map( A1 => n123, A2 => IN1(3), B1 => n120, B2 => IN0(3),
                           ZN => n18);
   U85 : AOI22_X1 port map( A1 => n72, A2 => IN1(7), B1 => n119, B2 => IN0(7), 
                           ZN => n10);
   U86 : NAND2_X1 port map( A1 => n68, A2 => n69, ZN => OUT1(0));
   U87 : NAND2_X1 port map( A1 => n126, A2 => IN2(27), ZN => n31);
   U88 : NAND2_X1 port map( A1 => n126, A2 => IN2(2), ZN => n25);
   U89 : NAND2_X1 port map( A1 => n126, A2 => IN2(25), ZN => n35);
   U90 : NAND2_X1 port map( A1 => n12, A2 => n13, ZN => OUT1(6));
   U91 : NAND2_X1 port map( A1 => n2, A2 => n3, ZN => OUT1(9));
   U92 : AOI22_X1 port map( A1 => n123, A2 => IN1(27), B1 => n121, B2 => 
                           IN0(27), ZN => n30);
   U93 : AOI22_X1 port map( A1 => n122, A2 => IN1(2), B1 => n120, B2 => IN0(2),
                           ZN => n24);
   U94 : AOI22_X1 port map( A1 => n123, A2 => IN1(25), B1 => n121, B2 => 
                           IN0(25), ZN => n34);
   U95 : AOI22_X1 port map( A1 => n73, A2 => IN1(28), B1 => n121, B2 => IN0(28)
                           , ZN => n28);
   U96 : AOI22_X1 port map( A1 => n72, A2 => IN1(20), B1 => n121, B2 => IN0(20)
                           , ZN => n44);
   U97 : AOI22_X1 port map( A1 => n72, A2 => IN1(24), B1 => n121, B2 => IN0(24)
                           , ZN => n36);
   U98 : NAND2_X1 port map( A1 => n30, A2 => n31, ZN => OUT1(27));
   U99 : NAND2_X1 port map( A1 => n125, A2 => IN2(1), ZN => n47);
   U100 : NAND2_X1 port map( A1 => n125, A2 => IN2(10), ZN => n67);
   U101 : AOI22_X1 port map( A1 => n122, A2 => IN1(6), B1 => n121, B2 => IN0(6)
                           , ZN => n12);
   U102 : NAND2_X1 port map( A1 => n10, A2 => n11, ZN => OUT1(7));
   U103 : NAND2_X1 port map( A1 => n8, A2 => n9, ZN => OUT1(8));
   U104 : AOI22_X1 port map( A1 => n71, A2 => IN1(1), B1 => n119, B2 => IN0(1),
                           ZN => n46);
   U105 : AOI22_X1 port map( A1 => n71, A2 => IN1(10), B1 => n121, B2 => 
                           IN0(10), ZN => n66);
   U106 : AOI22_X1 port map( A1 => n71, A2 => IN1(0), B1 => n119, B2 => IN0(0),
                           ZN => n68);
   U107 : AOI22_X1 port map( A1 => n122, A2 => IN1(13), B1 => n120, B2 => 
                           IN0(13), ZN => n60);
   U108 : AOI22_X1 port map( A1 => n73, A2 => IN1(31), B1 => n121, B2 => 
                           IN0(31), ZN => n20);
   U109 : NAND2_X1 port map( A1 => n125, A2 => IN2(31), ZN => n21);
   U110 : NAND2_X1 port map( A1 => n18, A2 => n19, ZN => OUT1(3));
   U111 : NAND2_X1 port map( A1 => n34, A2 => n35, ZN => OUT1(25));
   U112 : NAND2_X1 port map( A1 => n20, A2 => n21, ZN => OUT1(31));
   U113 : NAND2_X1 port map( A1 => n16, A2 => n17, ZN => OUT1(4));
   U114 : NAND2_X1 port map( A1 => n28, A2 => n29, ZN => OUT1(28));
   U115 : NAND2_X1 port map( A1 => n24, A2 => n25, ZN => OUT1(2));
   U116 : NAND2_X1 port map( A1 => n36, A2 => n37, ZN => OUT1(24));
   U117 : NAND2_X1 port map( A1 => n44, A2 => n45, ZN => OUT1(20));
   U118 : NAND2_X1 port map( A1 => n125, A2 => IN2(9), ZN => n3);
   U119 : NAND2_X1 port map( A1 => n125, A2 => IN2(4), ZN => n17);
   U120 : NAND2_X1 port map( A1 => n126, A2 => IN2(8), ZN => n9);
   U121 : NAND2_X1 port map( A1 => n126, A2 => IN2(3), ZN => n19);
   U122 : NAND2_X1 port map( A1 => n126, A2 => IN2(7), ZN => n11);
   U123 : NAND2_X1 port map( A1 => n126, A2 => IN2(6), ZN => n13);
   U124 : NAND2_X1 port map( A1 => n126, A2 => IN2(0), ZN => n69);
   U125 : NAND2_X1 port map( A1 => n126, A2 => IN2(13), ZN => n61);
   U126 : INV_X1 port map( A => CTRL(1), ZN => n70);

end SYN_bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity zerocheck is

   port( IN0 : in std_logic_vector (31 downto 0);  CTRL : in std_logic;  OUT1 :
         out std_logic);

end zerocheck;

architecture SYN_Bhe of zerocheck is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
      n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42
      : std_logic;

begin
   
   U1 : INV_X1 port map( A => IN0(7), ZN => n32);
   U2 : INV_X1 port map( A => IN0(13), ZN => n28);
   U3 : INV_X1 port map( A => IN0(12), ZN => n21);
   U4 : INV_X1 port map( A => IN0(1), ZN => n20);
   U5 : NOR2_X1 port map( A1 => n25, A2 => n26, ZN => n15);
   U6 : AND3_X1 port map( A1 => n14, A2 => n16, A3 => n15, ZN => n42);
   U7 : XNOR2_X1 port map( A => n42, B => CTRL, ZN => OUT1);
   U8 : INV_X1 port map( A => IN0(3), ZN => n31);
   U9 : INV_X1 port map( A => IN0(0), ZN => n29);
   U10 : NAND3_X1 port map( A1 => n19, A2 => n20, A3 => n21, ZN => n18);
   U11 : NAND3_X1 port map( A1 => n23, A2 => n24, A3 => n22, ZN => n17);
   U12 : NAND3_X1 port map( A1 => n27, A2 => n28, A3 => n29, ZN => n26);
   U13 : NAND3_X1 port map( A1 => n30, A2 => n31, A3 => n32, ZN => n25);
   U14 : NAND3_X1 port map( A1 => n35, A2 => n36, A3 => n37, ZN => n34);
   U15 : NOR2_X1 port map( A1 => IN0(31), A2 => IN0(14), ZN => n38);
   U16 : NAND4_X1 port map( A1 => n38, A2 => n39, A3 => n40, A4 => n41, ZN => 
                           n33);
   U17 : NOR2_X1 port map( A1 => IN0(18), A2 => IN0(19), ZN => n39);
   U18 : NOR2_X1 port map( A1 => IN0(22), A2 => IN0(17), ZN => n40);
   U19 : NOR2_X1 port map( A1 => IN0(30), A2 => IN0(21), ZN => n41);
   U20 : NOR2_X1 port map( A1 => IN0(20), A2 => IN0(15), ZN => n35);
   U21 : NOR2_X1 port map( A1 => IN0(27), A2 => IN0(29), ZN => n36);
   U22 : NOR2_X1 port map( A1 => IN0(25), A2 => IN0(26), ZN => n37);
   U23 : NOR2_X1 port map( A1 => IN0(11), A2 => IN0(23), ZN => n19);
   U24 : NOR2_X1 port map( A1 => IN0(5), A2 => IN0(16), ZN => n27);
   U25 : NOR2_X1 port map( A1 => IN0(10), A2 => IN0(6), ZN => n30);
   U26 : NOR2_X1 port map( A1 => IN0(24), A2 => IN0(28), ZN => n22);
   U27 : NOR2_X1 port map( A1 => IN0(4), A2 => IN0(9), ZN => n23);
   U28 : NOR2_X1 port map( A1 => IN0(2), A2 => IN0(8), ZN => n24);
   U29 : NOR2_X1 port map( A1 => n17, A2 => n18, ZN => n16);
   U30 : NOR2_X1 port map( A1 => n33, A2 => n34, ZN => n14);

end SYN_Bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity mux21_2 is

   port( IN0, IN1 : in std_logic_vector (31 downto 0);  CTRL : in std_logic;  
         OUT1 : out std_logic_vector (31 downto 0));

end mux21_2;

architecture SYN_Bhe of mux21_2 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X3
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8 : std_logic;

begin
   
   U1 : MUX2_X1 port map( A => IN0(9), B => IN1(9), S => n8, Z => OUT1(9));
   U3 : MUX2_X1 port map( A => IN0(7), B => IN1(7), S => n8, Z => OUT1(7));
   U5 : MUX2_X1 port map( A => IN0(5), B => IN1(5), S => n8, Z => OUT1(5));
   U10 : MUX2_X1 port map( A => IN0(2), B => IN1(2), S => n3, Z => OUT1(2));
   U17 : MUX2_X1 port map( A => IN0(23), B => IN1(23), S => n3, Z => OUT1(23));
   U20 : MUX2_X1 port map( A => IN0(20), B => IN1(20), S => n7, Z => OUT1(20));
   U22 : MUX2_X1 port map( A => IN0(19), B => IN1(19), S => n7, Z => OUT1(19));
   U23 : MUX2_X1 port map( A => IN0(18), B => IN1(18), S => n8, Z => OUT1(18));
   U24 : MUX2_X1 port map( A => IN0(17), B => IN1(17), S => n7, Z => OUT1(17));
   U25 : MUX2_X1 port map( A => IN0(16), B => IN1(16), S => n7, Z => OUT1(16));
   U26 : MUX2_X1 port map( A => IN0(15), B => IN1(15), S => n8, Z => OUT1(15));
   U28 : MUX2_X1 port map( A => IN0(13), B => IN1(13), S => n3, Z => OUT1(13));
   U29 : MUX2_X1 port map( A => IN0(12), B => IN1(12), S => n3, Z => OUT1(12));
   U14 : MUX2_X1 port map( A => IN0(26), B => IN1(26), S => n7, Z => OUT1(26));
   U4 : MUX2_X1 port map( A => IN0(6), B => IN1(6), S => n3, Z => OUT1(6));
   U6 : MUX2_X1 port map( A => IN0(4), B => IN1(4), S => n3, Z => OUT1(4));
   U7 : MUX2_X1 port map( A => IN0(3), B => IN1(3), S => n7, Z => OUT1(3));
   U9 : MUX2_X1 port map( A => IN0(30), B => IN1(30), S => n7, Z => OUT1(30));
   U32 : MUX2_X1 port map( A => IN0(0), B => IN1(0), S => n3, Z => OUT1(0));
   U13 : MUX2_X1 port map( A => IN0(27), B => IN1(27), S => n3, Z => OUT1(27));
   U19 : MUX2_X1 port map( A => IN0(21), B => IN1(21), S => n3, Z => OUT1(21));
   U21 : MUX2_X1 port map( A => IN0(1), B => IN1(1), S => n7, Z => OUT1(1));
   U16 : MUX2_X1 port map( A => IN0(24), B => IN1(24), S => n7, Z => OUT1(24));
   U30 : MUX2_X1 port map( A => IN0(11), B => IN1(11), S => n8, Z => OUT1(11));
   U2 : MUX2_X1 port map( A => IN0(10), B => IN1(10), S => n7, Z => OUT1(10));
   U8 : MUX2_X1 port map( A => IN0(8), B => IN1(8), S => n7, Z => OUT1(8));
   U11 : MUX2_X1 port map( A => IN0(14), B => IN1(14), S => n7, Z => OUT1(14));
   U12 : MUX2_X1 port map( A => IN0(25), B => IN1(25), S => n3, Z => OUT1(25));
   U15 : MUX2_X1 port map( A => IN0(22), B => IN1(22), S => n7, Z => OUT1(22));
   U18 : CLKBUF_X2 port map( A => CTRL, Z => n8);
   U27 : CLKBUF_X3 port map( A => CTRL, Z => n3);
   U31 : CLKBUF_X3 port map( A => CTRL, Z => n7);
   U33 : INV_X1 port map( A => n7, ZN => n4);
   U34 : NAND2_X1 port map( A1 => n3, A2 => IN1(31), ZN => n2);
   U35 : NAND2_X1 port map( A1 => IN0(31), A2 => n4, ZN => n1);
   U36 : NAND2_X1 port map( A1 => n1, A2 => n2, ZN => OUT1(31));
   U37 : NAND2_X1 port map( A1 => IN1(28), A2 => n3, ZN => n6);
   U38 : NAND2_X1 port map( A1 => IN0(28), A2 => n4, ZN => n5);
   U39 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => OUT1(28));
   U40 : MUX2_X1 port map( A => IN0(29), B => IN1(29), S => n3, Z => OUT1(29));

end SYN_Bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity p4add_N32_logN5_0 is

   port( A, B : in std_logic_vector (31 downto 0);  Cin, sign : in std_logic;  
         S : out std_logic_vector (31 downto 0);  Cout : out std_logic);

end p4add_N32_logN5_0;

architecture SYN_STRUCTURAL of p4add_N32_logN5_0 is

   component sum_gen_N32_0
      port( A, B : in std_logic_vector (31 downto 0);  Cin : in 
            std_logic_vector (8 downto 0);  S : out std_logic_vector (31 downto
            0));
   end component;
   
   component carry_tree_N32_logN5_0
      port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  
            Cout : out std_logic_vector (7 downto 0));
   end component;
   
   component xor_gen_N32_0
      port( A : in std_logic_vector (31 downto 0);  B : in std_logic;  S : out 
            std_logic_vector (31 downto 0));
   end component;
   
   signal new_B_31_port, new_B_30_port, new_B_29_port, new_B_28_port, 
      new_B_27_port, new_B_24_port, new_B_23_port, new_B_22_port, new_B_21_port
      , new_B_20_port, new_B_16_port, new_B_12_port, new_B_6_port, 
      carry_pro_7_port, carry_pro_6_port, carry_pro_5_port, carry_pro_4_port, 
      carry_pro_3_port, carry_pro_2_port, carry_pro_1_port, n1, n2, n3, n5, n6,
      n8, n10, n11, n12, n14, n15, n16, n17, n19, n20, n22, n23, n24, n25, n26,
      n27, n29, n30, n31, n32, n33, n34, n35, n36, net684299 : std_logic;

begin
   
   n26 <= '0';
   xor32 : xor_gen_N32_0 port map( A(31) => B(31), A(30) => B(30), A(29) => 
                           B(29), A(28) => B(28), A(27) => B(27), A(26) => 
                           B(26), A(25) => B(25), A(24) => B(24), A(23) => 
                           B(23), A(22) => B(22), A(21) => B(21), A(20) => 
                           B(20), A(19) => B(19), A(18) => B(18), A(17) => 
                           B(17), A(16) => B(16), A(15) => B(15), A(14) => 
                           B(14), A(13) => B(13), A(12) => B(12), A(11) => 
                           B(11), A(10) => B(10), A(9) => B(9), A(8) => B(8), 
                           A(7) => B(7), A(6) => B(6), A(5) => B(5), A(4) => 
                           B(4), A(3) => B(3), A(2) => B(2), A(1) => B(1), A(0)
                           => B(0), B => n20, S(31) => new_B_31_port, S(30) => 
                           new_B_30_port, S(29) => new_B_29_port, S(28) => 
                           new_B_28_port, S(27) => new_B_27_port, S(26) => n1, 
                           S(25) => n14, S(24) => new_B_24_port, S(23) => 
                           new_B_23_port, S(22) => new_B_22_port, S(21) => 
                           new_B_21_port, S(20) => new_B_20_port, S(19) => n27,
                           S(18) => n8, S(17) => n22, S(16) => new_B_16_port, 
                           S(15) => n3, S(14) => n16, S(13) => n6, S(12) => 
                           new_B_12_port, S(11) => n2, S(10) => n17, S(9) => 
                           n15, S(8) => n5, S(7) => n25, S(6) => new_B_6_port, 
                           S(5) => n19, S(4) => n23, S(3) => n12, S(2) => n11, 
                           S(1) => n24, S(0) => n10);
   ct : carry_tree_N32_logN5_0 port map( A(31) => n29, A(30) => n30, A(29) => 
                           n31, A(28) => n32, A(27) => A(27), A(26) => A(26), 
                           A(25) => A(25), A(24) => A(24), A(23) => A(23), 
                           A(22) => A(22), A(21) => A(21), A(20) => A(20), 
                           A(19) => A(19), A(18) => A(18), A(17) => A(17), 
                           A(16) => A(16), A(15) => A(15), A(14) => A(14), 
                           A(13) => A(13), A(12) => A(12), A(11) => A(11), 
                           A(10) => A(10), A(9) => A(9), A(8) => A(8), A(7) => 
                           A(7), A(6) => A(6), A(5) => A(5), A(4) => A(4), A(3)
                           => A(3), A(2) => A(2), A(1) => A(1), A(0) => A(0), 
                           B(31) => n33, B(30) => n34, B(29) => n35, B(28) => 
                           n36, B(27) => new_B_27_port, B(26) => n1, B(25) => 
                           n14, B(24) => new_B_24_port, B(23) => new_B_23_port,
                           B(22) => new_B_22_port, B(21) => new_B_21_port, 
                           B(20) => new_B_20_port, B(19) => n27, B(18) => n8, 
                           B(17) => n22, B(16) => new_B_16_port, B(15) => n3, 
                           B(14) => n16, B(13) => n6, B(12) => new_B_12_port, 
                           B(11) => n2, B(10) => n17, B(9) => n15, B(8) => n5, 
                           B(7) => n25, B(6) => new_B_6_port, B(5) => n19, B(4)
                           => n23, B(3) => n12, B(2) => n11, B(1) => n24, B(0) 
                           => n10, Cin => n20, Cout(7) => net684299, Cout(6) =>
                           carry_pro_7_port, Cout(5) => carry_pro_6_port, 
                           Cout(4) => carry_pro_5_port, Cout(3) => 
                           carry_pro_4_port, Cout(2) => carry_pro_3_port, 
                           Cout(1) => carry_pro_2_port, Cout(0) => 
                           carry_pro_1_port);
   add : sum_gen_N32_0 port map( A(31) => A(31), A(30) => A(30), A(29) => A(29)
                           , A(28) => A(28), A(27) => A(27), A(26) => A(26), 
                           A(25) => A(25), A(24) => A(24), A(23) => A(23), 
                           A(22) => A(22), A(21) => A(21), A(20) => A(20), 
                           A(19) => A(19), A(18) => A(18), A(17) => A(17), 
                           A(16) => A(16), A(15) => A(15), A(14) => A(14), 
                           A(13) => A(13), A(12) => A(12), A(11) => A(11), 
                           A(10) => A(10), A(9) => A(9), A(8) => A(8), A(7) => 
                           A(7), A(6) => A(6), A(5) => A(5), A(4) => A(4), A(3)
                           => A(3), A(2) => A(2), A(1) => A(1), A(0) => A(0), 
                           B(31) => new_B_31_port, B(30) => new_B_30_port, 
                           B(29) => new_B_29_port, B(28) => new_B_28_port, 
                           B(27) => new_B_27_port, B(26) => n1, B(25) => n14, 
                           B(24) => new_B_24_port, B(23) => new_B_23_port, 
                           B(22) => new_B_22_port, B(21) => new_B_21_port, 
                           B(20) => new_B_20_port, B(19) => n27, B(18) => n8, 
                           B(17) => n22, B(16) => new_B_16_port, B(15) => n3, 
                           B(14) => n16, B(13) => n6, B(12) => new_B_12_port, 
                           B(11) => n2, B(10) => n17, B(9) => n15, B(8) => n5, 
                           B(7) => n25, B(6) => new_B_6_port, B(5) => n19, B(4)
                           => n23, B(3) => n12, B(2) => n11, B(1) => n24, B(0) 
                           => n10, Cin(8) => n26, Cin(7) => carry_pro_7_port, 
                           Cin(6) => carry_pro_6_port, Cin(5) => 
                           carry_pro_5_port, Cin(4) => carry_pro_4_port, Cin(3)
                           => carry_pro_3_port, Cin(2) => carry_pro_2_port, 
                           Cin(1) => carry_pro_1_port, Cin(0) => n20, S(31) => 
                           S(31), S(30) => S(30), S(29) => S(29), S(28) => 
                           S(28), S(27) => S(27), S(26) => S(26), S(25) => 
                           S(25), S(24) => S(24), S(23) => S(23), S(22) => 
                           S(22), S(21) => S(21), S(20) => S(20), S(19) => 
                           S(19), S(18) => S(18), S(17) => S(17), S(16) => 
                           S(16), S(15) => S(15), S(14) => S(14), S(13) => 
                           S(13), S(12) => S(12), S(11) => S(11), S(10) => 
                           S(10), S(9) => S(9), S(8) => S(8), S(7) => S(7), 
                           S(6) => S(6), S(5) => S(5), S(4) => S(4), S(3) => 
                           S(3), S(2) => S(2), S(1) => S(1), S(0) => S(0));
   n20 <= '0';
   n29 <= '0';
   n30 <= '0';
   n31 <= '0';
   n32 <= '0';
   n33 <= '0';
   n34 <= '0';
   n35 <= '0';
   n36 <= '0';

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity extender_32 is

   port( IN1 : in std_logic_vector (31 downto 0);  CTRL, SIGN : in std_logic;  
         OUT1 : out std_logic_vector (31 downto 0));

end extender_32;

architecture SYN_Bhe of extender_32 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal OUT1_25_port, OUT1_24_port, OUT1_23_port, OUT1_22_port, OUT1_21_port,
      OUT1_20_port, OUT1_19_port, OUT1_18_port, OUT1_17_port, OUT1_16_port, n2,
      n3, n4, n5, n7, n8, n9, n10, n12, n11, n13, n14, n15, n16, OUT1_28_port, 
      OUT1_27_port, OUT1_26_port : std_logic;

begin
   OUT1 <= ( OUT1_26_port, OUT1_28_port, OUT1_28_port, OUT1_28_port, 
      OUT1_27_port, OUT1_26_port, OUT1_27_port, OUT1_24_port, OUT1_23_port, 
      OUT1_22_port, OUT1_21_port, OUT1_20_port, OUT1_19_port, OUT1_18_port, 
      OUT1_17_port, OUT1_16_port, IN1(15), IN1(14), IN1(13), IN1(12), IN1(11), 
      IN1(10), IN1(9), IN1(8), IN1(7), IN1(6), IN1(5), IN1(4), IN1(3), IN1(2), 
      IN1(1), IN1(0) );
   
   U2 : BUF_X2 port map( A => OUT1_25_port, Z => OUT1_28_port);
   U3 : NAND2_X1 port map( A1 => IN1(22), A2 => CTRL, ZN => n14);
   U4 : NAND2_X1 port map( A1 => n15, A2 => n14, ZN => OUT1_22_port);
   U5 : INV_X1 port map( A => CTRL, ZN => n13);
   U6 : NAND3_X1 port map( A1 => SIGN, A2 => IN1(15), A3 => n13, ZN => n16);
   U7 : NAND3_X1 port map( A1 => SIGN, A2 => IN1(15), A3 => n13, ZN => n15);
   U8 : NAND3_X1 port map( A1 => SIGN, A2 => IN1(15), A3 => n13, ZN => n2);
   U9 : NAND2_X1 port map( A1 => n2, A2 => n10, ZN => OUT1_18_port);
   U10 : NAND2_X1 port map( A1 => n2, A2 => n11, ZN => OUT1_17_port);
   U11 : NAND2_X1 port map( A1 => n2, A2 => n3, ZN => OUT1_25_port);
   U12 : BUF_X2 port map( A => OUT1_25_port, Z => OUT1_27_port);
   U13 : CLKBUF_X2 port map( A => OUT1_25_port, Z => OUT1_26_port);
   U14 : NAND2_X1 port map( A1 => n16, A2 => n7, ZN => OUT1_21_port);
   U15 : NAND2_X1 port map( A1 => CTRL, A2 => IN1(17), ZN => n11);
   U16 : NAND2_X1 port map( A1 => CTRL, A2 => IN1(24), ZN => n4);
   U17 : NAND2_X1 port map( A1 => CTRL, A2 => IN1(20), ZN => n8);
   U18 : NAND2_X1 port map( A1 => CTRL, A2 => IN1(16), ZN => n12);
   U19 : NAND2_X1 port map( A1 => CTRL, A2 => IN1(23), ZN => n5);
   U20 : NAND2_X1 port map( A1 => CTRL, A2 => IN1(19), ZN => n9);
   U21 : NAND2_X1 port map( A1 => CTRL, A2 => IN1(21), ZN => n7);
   U22 : NAND2_X1 port map( A1 => CTRL, A2 => IN1(18), ZN => n10);
   U23 : NAND2_X1 port map( A1 => CTRL, A2 => IN1(25), ZN => n3);
   U24 : NAND2_X1 port map( A1 => n15, A2 => n4, ZN => OUT1_24_port);
   U25 : NAND2_X1 port map( A1 => n15, A2 => n8, ZN => OUT1_20_port);
   U26 : NAND2_X1 port map( A1 => n15, A2 => n5, ZN => OUT1_23_port);
   U27 : NAND2_X1 port map( A1 => n16, A2 => n9, ZN => OUT1_19_port);
   U28 : NAND2_X1 port map( A1 => n16, A2 => n12, ZN => OUT1_16_port);

end SYN_Bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity ff32_en_IR is

   port( D : in std_logic_vector (31 downto 0);  en, clk, rst : in std_logic;  
         Q : out std_logic_vector (31 downto 0));

end ff32_en_IR;

architecture SYN_behavioral of ff32_en_IR is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFS_X2
      port( D, CK, SN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFS_X1
      port( D, CK, SN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFR_X2
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
      n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93
      , n94, n95, n97, net644967, net644968, net644969, net644970, net644971, 
      net644972, net644973, net644974, net644975, net644976, net644977, 
      net644978, net644979, net644980, net644981, net644982, net644983, 
      net644984, net644985, net644986, net644987, net644988, net644989, 
      net644990, net644991, net644992, net644993, net644994, net644995, 
      net644996, net644997, net644998, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11
      , n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, 
      n26, n27, n28, n29, n30, n31, n32, n33, n34, n35 : std_logic;

begin
   
   Q_reg_24_inst : DFFR_X1 port map( D => n89, CK => clk, RN => n35, Q => Q(24)
                           , QN => net644991);
   Q_reg_23_inst : DFFR_X1 port map( D => n88, CK => clk, RN => n35, Q => Q(23)
                           , QN => net644990);
   Q_reg_22_inst : DFFR_X1 port map( D => n87, CK => clk, RN => n35, Q => Q(22)
                           , QN => net644989);
   Q_reg_20_inst : DFFR_X1 port map( D => n85, CK => clk, RN => n35, Q => Q(20)
                           , QN => net644987);
   Q_reg_19_inst : DFFR_X1 port map( D => n84, CK => clk, RN => n35, Q => Q(19)
                           , QN => net644986);
   Q_reg_18_inst : DFFR_X1 port map( D => n83, CK => clk, RN => n35, Q => Q(18)
                           , QN => net644985);
   Q_reg_17_inst : DFFR_X1 port map( D => n82, CK => clk, RN => n35, Q => Q(17)
                           , QN => net644984);
   Q_reg_16_inst : DFFR_X1 port map( D => n81, CK => clk, RN => n35, Q => Q(16)
                           , QN => net644983);
   Q_reg_15_inst : DFFR_X1 port map( D => n80, CK => clk, RN => n35, Q => Q(15)
                           , QN => net644982);
   Q_reg_14_inst : DFFR_X1 port map( D => n79, CK => clk, RN => n35, Q => Q(14)
                           , QN => net644981);
   Q_reg_13_inst : DFFR_X1 port map( D => n78, CK => clk, RN => n35, Q => Q(13)
                           , QN => net644980);
   Q_reg_12_inst : DFFR_X1 port map( D => n77, CK => clk, RN => n35, Q => Q(12)
                           , QN => net644979);
   Q_reg_11_inst : DFFR_X1 port map( D => n76, CK => clk, RN => n35, Q => Q(11)
                           , QN => net644978);
   Q_reg_10_inst : DFFR_X1 port map( D => n75, CK => clk, RN => n35, Q => Q(10)
                           , QN => net644977);
   Q_reg_9_inst : DFFR_X1 port map( D => n74, CK => clk, RN => n35, Q => Q(9), 
                           QN => net644976);
   Q_reg_8_inst : DFFR_X1 port map( D => n73, CK => clk, RN => n35, Q => Q(8), 
                           QN => net644975);
   Q_reg_7_inst : DFFR_X1 port map( D => n72, CK => clk, RN => n35, Q => Q(7), 
                           QN => net644974);
   Q_reg_6_inst : DFFR_X1 port map( D => n71, CK => clk, RN => n35, Q => Q(6), 
                           QN => net644973);
   Q_reg_5_inst : DFFR_X1 port map( D => n70, CK => clk, RN => n35, Q => Q(5), 
                           QN => net644972);
   Q_reg_4_inst : DFFR_X1 port map( D => n69, CK => clk, RN => n35, Q => Q(4), 
                           QN => net644971);
   Q_reg_3_inst : DFFR_X1 port map( D => n68, CK => clk, RN => n35, Q => Q(3), 
                           QN => net644970);
   Q_reg_2_inst : DFFR_X1 port map( D => n67, CK => clk, RN => n35, Q => Q(2), 
                           QN => net644969);
   Q_reg_1_inst : DFFR_X1 port map( D => n66, CK => clk, RN => n35, Q => Q(1), 
                           QN => net644968);
   Q_reg_0_inst : DFFR_X1 port map( D => n65, CK => clk, RN => n35, Q => Q(0), 
                           QN => net644967);
   Q_reg_31_inst : DFFR_X2 port map( D => n97, CK => clk, RN => n35, Q => Q(31)
                           , QN => net644998);
   U6 : NAND2_X1 port map( A1 => en, A2 => D(30), ZN => n3);
   U5 : OAI21_X1 port map( B1 => en, B2 => net644997, A => n3, ZN => n95);
   U3 : NAND2_X1 port map( A1 => en, A2 => D(31), ZN => n2);
   U2 : OAI21_X1 port map( B1 => en, B2 => net644998, A => n2, ZN => n97);
   U48 : NAND2_X1 port map( A1 => en, A2 => D(9), ZN => n24);
   U47 : OAI21_X1 port map( B1 => en, B2 => net644976, A => n24, ZN => n74);
   U52 : NAND2_X1 port map( A1 => en, A2 => D(7), ZN => n26);
   U51 : OAI21_X1 port map( B1 => en, B2 => net644974, A => n26, ZN => n72);
   U34 : NAND2_X1 port map( A1 => en, A2 => D(16), ZN => n17);
   U33 : OAI21_X1 port map( B1 => en, B2 => net644983, A => n17, ZN => n81);
   U64 : NAND2_X1 port map( A1 => en, A2 => D(1), ZN => n32);
   U63 : OAI21_X1 port map( B1 => n34, B2 => net644968, A => n32, ZN => n66);
   U66 : NAND2_X1 port map( A1 => en, A2 => D(0), ZN => n33);
   U65 : OAI21_X1 port map( B1 => en, B2 => net644967, A => n33, ZN => n65);
   U50 : NAND2_X1 port map( A1 => en, A2 => D(8), ZN => n25);
   U49 : OAI21_X1 port map( B1 => en, B2 => net644975, A => n25, ZN => n73);
   U54 : NAND2_X1 port map( A1 => n34, A2 => D(6), ZN => n27);
   U53 : OAI21_X1 port map( B1 => en, B2 => net644973, A => n27, ZN => n71);
   U62 : NAND2_X1 port map( A1 => n34, A2 => D(2), ZN => n31);
   U61 : OAI21_X1 port map( B1 => en, B2 => net644969, A => n31, ZN => n67);
   U60 : NAND2_X1 port map( A1 => n34, A2 => D(3), ZN => n30);
   U59 : OAI21_X1 port map( B1 => en, B2 => net644970, A => n30, ZN => n68);
   U56 : NAND2_X1 port map( A1 => en, A2 => D(5), ZN => n28);
   U55 : OAI21_X1 port map( B1 => en, B2 => net644972, A => n28, ZN => n70);
   U16 : NAND2_X1 port map( A1 => n34, A2 => D(25), ZN => n8);
   U15 : OAI21_X1 port map( B1 => en, B2 => net644992, A => n8, ZN => n90);
   U24 : NAND2_X1 port map( A1 => n34, A2 => D(21), ZN => n12);
   U23 : OAI21_X1 port map( B1 => en, B2 => net644988, A => n12, ZN => n86);
   U18 : NAND2_X1 port map( A1 => n34, A2 => D(24), ZN => n9);
   U17 : OAI21_X1 port map( B1 => en, B2 => net644991, A => n9, ZN => n89);
   U20 : NAND2_X1 port map( A1 => n34, A2 => D(23), ZN => n10);
   U19 : OAI21_X1 port map( B1 => en, B2 => net644990, A => n10, ZN => n88);
   U8 : NAND2_X1 port map( A1 => n34, A2 => D(29), ZN => n4);
   U7 : OAI21_X1 port map( B1 => en, B2 => net644996, A => n4, ZN => n94);
   U14 : NAND2_X1 port map( A1 => n34, A2 => D(26), ZN => n7);
   U13 : OAI21_X1 port map( B1 => en, B2 => net644993, A => n7, ZN => n91);
   U58 : NAND2_X1 port map( A1 => n34, A2 => D(4), ZN => n29);
   U57 : OAI21_X1 port map( B1 => n34, B2 => net644971, A => n29, ZN => n69);
   U12 : NAND2_X1 port map( A1 => n34, A2 => D(27), ZN => n6);
   U10 : NAND2_X1 port map( A1 => n34, A2 => D(28), ZN => n5);
   U36 : NAND2_X1 port map( A1 => en, A2 => D(15), ZN => n18);
   U35 : OAI21_X1 port map( B1 => n34, B2 => net644982, A => n18, ZN => n80);
   U32 : NAND2_X1 port map( A1 => en, A2 => D(17), ZN => n16);
   U31 : OAI21_X1 port map( B1 => n34, B2 => net644984, A => n16, ZN => n82);
   U30 : NAND2_X1 port map( A1 => en, A2 => D(18), ZN => n15);
   U29 : OAI21_X1 port map( B1 => en, B2 => net644985, A => n15, ZN => n83);
   U26 : NAND2_X1 port map( A1 => en, A2 => D(20), ZN => n13);
   U25 : OAI21_X1 port map( B1 => en, B2 => net644987, A => n13, ZN => n85);
   U40 : NAND2_X1 port map( A1 => en, A2 => D(13), ZN => n20);
   U39 : OAI21_X1 port map( B1 => en, B2 => net644980, A => n20, ZN => n78);
   U38 : NAND2_X1 port map( A1 => en, A2 => D(14), ZN => n19);
   U37 : OAI21_X1 port map( B1 => en, B2 => net644981, A => n19, ZN => n79);
   U42 : NAND2_X1 port map( A1 => en, A2 => D(12), ZN => n21);
   U41 : OAI21_X1 port map( B1 => en, B2 => net644979, A => n21, ZN => n77);
   U22 : NAND2_X1 port map( A1 => en, A2 => D(22), ZN => n11);
   U21 : OAI21_X1 port map( B1 => en, B2 => net644989, A => n11, ZN => n87);
   U46 : NAND2_X1 port map( A1 => en, A2 => D(10), ZN => n23);
   U45 : OAI21_X1 port map( B1 => en, B2 => net644977, A => n23, ZN => n75);
   U28 : NAND2_X1 port map( A1 => en, A2 => D(19), ZN => n14);
   U27 : OAI21_X1 port map( B1 => en, B2 => net644986, A => n14, ZN => n84);
   U44 : NAND2_X1 port map( A1 => en, A2 => D(11), ZN => n22);
   U43 : OAI21_X1 port map( B1 => en, B2 => net644978, A => n22, ZN => n76);
   Q_reg_21_inst : DFFR_X2 port map( D => n86, CK => clk, RN => n35, Q => Q(21)
                           , QN => net644988);
   Q_reg_28_inst : DFFS_X1 port map( D => n93, CK => clk, SN => n35, Q => Q(28)
                           , QN => net644995);
   Q_reg_26_inst : DFFS_X1 port map( D => n91, CK => clk, SN => n35, Q => Q(26)
                           , QN => net644993);
   Q_reg_29_inst : DFFR_X1 port map( D => n94, CK => clk, RN => n35, Q => Q(29)
                           , QN => net644996);
   Q_reg_27_inst : DFFR_X1 port map( D => n92, CK => clk, RN => n35, Q => Q(27)
                           , QN => net644994);
   Q_reg_30_inst : DFFS_X2 port map( D => n95, CK => clk, SN => n35, Q => Q(30)
                           , QN => net644997);
   Q_reg_25_inst : DFFR_X1 port map( D => n90, CK => clk, RN => n35, Q => Q(25)
                           , QN => net644992);
   U4 : INV_X2 port map( A => rst, ZN => n35);
   U9 : BUF_X1 port map( A => en, Z => n34);
   U11 : OAI21_X1 port map( B1 => en, B2 => net644994, A => n6, ZN => n92);
   U67 : OAI21_X1 port map( B1 => en, B2 => net644995, A => n5, ZN => n93);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity ff32_en_1 is

   port( D : in std_logic_vector (31 downto 0);  en, clk, rst : in std_logic;  
         Q : out std_logic_vector (31 downto 0));

end ff32_en_1;

architecture SYN_behavioral of ff32_en_1 is

   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, 
      n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31
      , n32, n33, net645075, net645076, net645077, net645078, net645079, 
      net645080, net645081, net645082, net645083, net645084, net645085, 
      net645086, net645087, net645088, net645089, net645090, net645091, 
      net645092, net645093, net645094, net645095, net645096, net645097, 
      net645098, net645099, net645100, net645101, net645102, net645103, 
      net645104, net645105, net645106, n35, n36, n37, n38, n39, n40, n41, n42, 
      n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57
      , n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68 : std_logic;

begin
   
   Q_reg_31_inst : DFFR_X1 port map( D => n1, CK => clk, RN => n68, Q => Q(31),
                           QN => net645106);
   Q_reg_30_inst : DFFR_X1 port map( D => n3, CK => clk, RN => n68, Q => Q(30),
                           QN => net645105);
   Q_reg_29_inst : DFFR_X1 port map( D => n4, CK => clk, RN => n68, Q => Q(29),
                           QN => net645104);
   Q_reg_28_inst : DFFR_X1 port map( D => n5, CK => clk, RN => n68, Q => Q(28),
                           QN => net645103);
   Q_reg_27_inst : DFFR_X1 port map( D => n6, CK => clk, RN => n68, Q => Q(27),
                           QN => net645102);
   Q_reg_26_inst : DFFR_X1 port map( D => n7, CK => clk, RN => n68, Q => Q(26),
                           QN => net645101);
   Q_reg_25_inst : DFFR_X1 port map( D => n8, CK => clk, RN => n68, Q => Q(25),
                           QN => net645100);
   Q_reg_24_inst : DFFR_X1 port map( D => n9, CK => clk, RN => n68, Q => Q(24),
                           QN => net645099);
   Q_reg_23_inst : DFFR_X1 port map( D => n10, CK => clk, RN => n68, Q => Q(23)
                           , QN => net645098);
   Q_reg_22_inst : DFFR_X1 port map( D => n11, CK => clk, RN => n68, Q => Q(22)
                           , QN => net645097);
   Q_reg_21_inst : DFFR_X1 port map( D => n12, CK => clk, RN => n68, Q => Q(21)
                           , QN => net645096);
   Q_reg_20_inst : DFFR_X1 port map( D => n13, CK => clk, RN => n68, Q => Q(20)
                           , QN => net645095);
   Q_reg_19_inst : DFFR_X1 port map( D => n14, CK => clk, RN => n68, Q => Q(19)
                           , QN => net645094);
   Q_reg_18_inst : DFFR_X1 port map( D => n15, CK => clk, RN => n68, Q => Q(18)
                           , QN => net645093);
   Q_reg_17_inst : DFFR_X1 port map( D => n16, CK => clk, RN => n68, Q => Q(17)
                           , QN => net645092);
   Q_reg_16_inst : DFFR_X1 port map( D => n17, CK => clk, RN => n68, Q => Q(16)
                           , QN => net645091);
   Q_reg_15_inst : DFFR_X1 port map( D => n18, CK => clk, RN => n68, Q => Q(15)
                           , QN => net645090);
   Q_reg_14_inst : DFFR_X1 port map( D => n19, CK => clk, RN => n68, Q => Q(14)
                           , QN => net645089);
   Q_reg_13_inst : DFFR_X1 port map( D => n20, CK => clk, RN => n68, Q => Q(13)
                           , QN => net645088);
   Q_reg_12_inst : DFFR_X1 port map( D => n21, CK => clk, RN => n68, Q => Q(12)
                           , QN => net645087);
   Q_reg_11_inst : DFFR_X1 port map( D => n22, CK => clk, RN => n68, Q => Q(11)
                           , QN => net645086);
   Q_reg_10_inst : DFFR_X1 port map( D => n23, CK => clk, RN => n68, Q => Q(10)
                           , QN => net645085);
   Q_reg_9_inst : DFFR_X1 port map( D => n24, CK => clk, RN => n68, Q => Q(9), 
                           QN => net645084);
   Q_reg_8_inst : DFFR_X1 port map( D => n25, CK => clk, RN => n68, Q => Q(8), 
                           QN => net645083);
   Q_reg_7_inst : DFFR_X1 port map( D => n26, CK => clk, RN => n68, Q => Q(7), 
                           QN => net645082);
   Q_reg_6_inst : DFFR_X1 port map( D => n27, CK => clk, RN => n68, Q => Q(6), 
                           QN => net645081);
   Q_reg_5_inst : DFFR_X1 port map( D => n28, CK => clk, RN => n68, Q => Q(5), 
                           QN => net645080);
   Q_reg_4_inst : DFFR_X1 port map( D => n29, CK => clk, RN => n68, Q => Q(4), 
                           QN => net645079);
   Q_reg_3_inst : DFFR_X1 port map( D => n30, CK => clk, RN => n68, Q => Q(3), 
                           QN => net645078);
   Q_reg_2_inst : DFFR_X1 port map( D => n31, CK => clk, RN => n68, Q => Q(2), 
                           QN => net645077);
   Q_reg_1_inst : DFFR_X1 port map( D => n32, CK => clk, RN => n68, Q => Q(1), 
                           QN => net645076);
   Q_reg_0_inst : DFFR_X1 port map( D => n33, CK => clk, RN => n68, Q => Q(0), 
                           QN => net645075);
   U66 : NAND2_X1 port map( A1 => en, A2 => D(31), ZN => n66);
   U65 : OAI21_X1 port map( B1 => en, B2 => net645106, A => n66, ZN => n1);
   U23 : NAND2_X1 port map( A1 => n67, A2 => D(30), ZN => n45);
   U22 : OAI21_X1 port map( B1 => en, B2 => net645105, A => n45, ZN => n3);
   U13 : NAND2_X1 port map( A1 => en, A2 => D(29), ZN => n40);
   U12 : OAI21_X1 port map( B1 => en, B2 => net645104, A => n40, ZN => n4);
   U11 : NAND2_X1 port map( A1 => en, A2 => D(28), ZN => n39);
   U10 : OAI21_X1 port map( B1 => en, B2 => net645103, A => n39, ZN => n5);
   U9 : NAND2_X1 port map( A1 => n67, A2 => D(27), ZN => n38);
   U8 : OAI21_X1 port map( B1 => en, B2 => net645102, A => n38, ZN => n6);
   U7 : NAND2_X1 port map( A1 => en, A2 => D(26), ZN => n37);
   U6 : OAI21_X1 port map( B1 => en, B2 => net645101, A => n37, ZN => n7);
   U5 : NAND2_X1 port map( A1 => en, A2 => D(25), ZN => n36);
   U4 : OAI21_X1 port map( B1 => en, B2 => net645100, A => n36, ZN => n8);
   U19 : NAND2_X1 port map( A1 => en, A2 => D(2), ZN => n43);
   U18 : OAI21_X1 port map( B1 => en, B2 => net645077, A => n43, ZN => n31);
   U3 : NAND2_X1 port map( A1 => en, A2 => D(24), ZN => n35);
   U2 : OAI21_X1 port map( B1 => en, B2 => net645099, A => n35, ZN => n9);
   U62 : NAND2_X1 port map( A1 => en, A2 => D(22), ZN => n64);
   U61 : OAI21_X1 port map( B1 => n67, B2 => net645097, A => n64, ZN => n11);
   U64 : NAND2_X1 port map( A1 => en, A2 => D(23), ZN => n65);
   U63 : OAI21_X1 port map( B1 => en, B2 => net645098, A => n65, ZN => n10);
   U17 : NAND2_X1 port map( A1 => n67, A2 => D(1), ZN => n42);
   U16 : OAI21_X1 port map( B1 => en, B2 => net645076, A => n42, ZN => n32);
   U52 : NAND2_X1 port map( A1 => n67, A2 => D(17), ZN => n59);
   U51 : OAI21_X1 port map( B1 => en, B2 => net645092, A => n59, ZN => n16);
   U39 : NAND2_X1 port map( A1 => n67, A2 => D(11), ZN => n53);
   U38 : OAI21_X1 port map( B1 => en, B2 => net645086, A => n53, ZN => n22);
   U41 : NAND2_X1 port map( A1 => n67, A2 => D(12), ZN => n54);
   U40 : OAI21_X1 port map( B1 => en, B2 => net645087, A => n54, ZN => n21);
   U35 : NAND2_X1 port map( A1 => n67, A2 => D(9), ZN => n51);
   U34 : OAI21_X1 port map( B1 => en, B2 => net645084, A => n51, ZN => n24);
   U31 : NAND2_X1 port map( A1 => n67, A2 => D(7), ZN => n49);
   U30 : OAI21_X1 port map( B1 => en, B2 => net645082, A => n49, ZN => n26);
   U33 : NAND2_X1 port map( A1 => n67, A2 => D(8), ZN => n50);
   U32 : OAI21_X1 port map( B1 => en, B2 => net645083, A => n50, ZN => n25);
   U48 : NAND2_X1 port map( A1 => n67, A2 => D(15), ZN => n57);
   U47 : OAI21_X1 port map( B1 => en, B2 => net645090, A => n57, ZN => n18);
   U25 : NAND2_X1 port map( A1 => n67, A2 => D(4), ZN => n46);
   U24 : OAI21_X1 port map( B1 => en, B2 => net645079, A => n46, ZN => n29);
   U43 : NAND2_X1 port map( A1 => n67, A2 => D(13), ZN => n55);
   U42 : OAI21_X1 port map( B1 => en, B2 => net645088, A => n55, ZN => n20);
   U29 : NAND2_X1 port map( A1 => n67, A2 => D(6), ZN => n48);
   U28 : OAI21_X1 port map( B1 => en, B2 => net645081, A => n48, ZN => n27);
   U37 : NAND2_X1 port map( A1 => n67, A2 => D(10), ZN => n52);
   U36 : OAI21_X1 port map( B1 => en, B2 => net645085, A => n52, ZN => n23);
   U21 : NAND2_X1 port map( A1 => n67, A2 => D(3), ZN => n44);
   U20 : OAI21_X1 port map( B1 => en, B2 => net645078, A => n44, ZN => n30);
   U46 : NAND2_X1 port map( A1 => n67, A2 => D(14), ZN => n56);
   U45 : OAI21_X1 port map( B1 => en, B2 => net645089, A => n56, ZN => n19);
   U27 : NAND2_X1 port map( A1 => n67, A2 => D(5), ZN => n47);
   U26 : OAI21_X1 port map( B1 => en, B2 => net645080, A => n47, ZN => n28);
   U50 : NAND2_X1 port map( A1 => n67, A2 => D(16), ZN => n58);
   U49 : OAI21_X1 port map( B1 => n67, B2 => net645091, A => n58, ZN => n17);
   U58 : NAND2_X1 port map( A1 => n67, A2 => D(20), ZN => n62);
   U57 : OAI21_X1 port map( B1 => n67, B2 => net645095, A => n62, ZN => n13);
   U54 : NAND2_X1 port map( A1 => n67, A2 => D(18), ZN => n60);
   U53 : OAI21_X1 port map( B1 => n67, B2 => net645093, A => n60, ZN => n15);
   U60 : NAND2_X1 port map( A1 => n67, A2 => D(21), ZN => n63);
   U59 : OAI21_X1 port map( B1 => n67, B2 => net645096, A => n63, ZN => n12);
   U56 : NAND2_X1 port map( A1 => n67, A2 => D(19), ZN => n61);
   U55 : OAI21_X1 port map( B1 => en, B2 => net645094, A => n61, ZN => n14);
   U15 : NAND2_X1 port map( A1 => en, A2 => D(0), ZN => n41);
   U14 : OAI21_X1 port map( B1 => en, B2 => net645075, A => n41, ZN => n33);
   U44 : INV_X2 port map( A => rst, ZN => n68);
   U67 : BUF_X2 port map( A => en, Z => n67);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity predictor_2_15 is

   port( clock, reset, enable, taken_i : in std_logic;  prediction_o : out 
         std_logic);

end predictor_2_15;

architecture SYN_bhe of predictor_2_15 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal prediction_o_port, next_STATE_1_port, next_STATE_0_port, N11, N12, n5
      , n6, n8, n9, n11_port, n10, n12_port, net684298 : std_logic;

begin
   prediction_o <= prediction_o_port;
   
   next_STATE_reg_0_inst : DLH_X1 port map( G => enable, D => N11, Q => 
                           next_STATE_0_port);
   STATE_reg_0_inst : DFFR_X1 port map( D => n6, CK => clock, RN => n12_port, Q
                           => n5, QN => n10);
   next_STATE_reg_1_inst : DLH_X1 port map( G => enable, D => N12, Q => 
                           next_STATE_1_port);
   STATE_reg_1_inst : DFFR_X1 port map( D => n8, CK => clock, RN => n12_port, Q
                           => prediction_o_port, QN => net684298);
   U8 : MUX2_X1 port map( A => prediction_o_port, B => next_STATE_1_port, S => 
                           enable, Z => n8);
   U9 : MUX2_X1 port map( A => n5, B => next_STATE_0_port, S => enable, Z => n6
                           );
   U7 : NOR2_X1 port map( A1 => prediction_o_port, A2 => taken_i, ZN => n9);
   U6 : NAND2_X1 port map( A1 => prediction_o_port, A2 => taken_i, ZN => 
                           n11_port);
   U3 : OAI21_X1 port map( B1 => n9, B2 => n10, A => n11_port, ZN => N12);
   U5 : OAI21_X1 port map( B1 => n5, B2 => n9, A => n11_port, ZN => N11);
   U2 : INV_X1 port map( A => reset, ZN => n12_port);

end SYN_bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity predictor_2_0 is

   port( clock, reset, enable, taken_i : in std_logic;  prediction_o : out 
         std_logic);

end predictor_2_0;

architecture SYN_bhe of predictor_2_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal prediction_o_port, next_STATE_1_port, next_STATE_0_port, N11, N12, n9
      , n11_port, n5, n6, n8, n7, n10, net684297 : std_logic;

begin
   prediction_o <= prediction_o_port;
   
   next_STATE_reg_0_inst : DLH_X1 port map( G => enable, D => N11, Q => 
                           next_STATE_0_port);
   STATE_reg_0_inst : DFFR_X1 port map( D => n11_port, CK => clock, RN => n10, 
                           Q => n5, QN => n7);
   next_STATE_reg_1_inst : DLH_X1 port map( G => enable, D => N12, Q => 
                           next_STATE_1_port);
   STATE_reg_1_inst : DFFR_X1 port map( D => n9, CK => clock, RN => n10, Q => 
                           prediction_o_port, QN => net684297);
   U8 : MUX2_X1 port map( A => prediction_o_port, B => next_STATE_1_port, S => 
                           enable, Z => n9);
   U9 : MUX2_X1 port map( A => n5, B => next_STATE_0_port, S => enable, Z => 
                           n11_port);
   U7 : NOR2_X1 port map( A1 => prediction_o_port, A2 => taken_i, ZN => n6);
   U6 : NAND2_X1 port map( A1 => prediction_o_port, A2 => taken_i, ZN => n8);
   U3 : OAI21_X1 port map( B1 => n6, B2 => n7, A => n8, ZN => N12);
   U5 : OAI21_X1 port map( B1 => n5, B2 => n6, A => n8, ZN => N11);
   U2 : INV_X1 port map( A => reset, ZN => n10);

end SYN_bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity mux41_0 is

   port( IN0, IN1, IN2, IN3 : in std_logic_vector (31 downto 0);  CTRL : in 
         std_logic_vector (1 downto 0);  OUT1 : out std_logic_vector (31 downto
         0));

end mux41_0;

architecture SYN_bhe of mux41_0 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X4
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n194, n4, n5, n6, n7, n10, n11, n18, n19, n60, n61, n62, n63, n68, 
      n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83
      , n84, n85, n86, n87, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, 
      n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, 
      n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, 
      n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, 
      n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, 
      n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, 
      n159, n160, n161, n162, n163, n164, n165, n166, n167, n169, n170, n171, 
      n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, 
      n184, n185, n186, n187, n188, n189, n190, n191, n192, n193 : std_logic;

begin
   
   U87 : AOI22_X1 port map( A1 => n6, A2 => IN1(12), B1 => n193, B2 => IN0(12),
                           ZN => n62);
   U86 : AOI22_X1 port map( A1 => n89, A2 => IN3(12), B1 => n90, B2 => IN2(12),
                           ZN => n63);
   U84 : AOI22_X1 port map( A1 => n6, A2 => IN1(13), B1 => n193, B2 => IN0(13),
                           ZN => n60);
   U83 : AOI22_X1 port map( A1 => n89, A2 => IN3(13), B1 => n90, B2 => IN2(13),
                           ZN => n61);
   U9 : AOI22_X1 port map( A1 => n6, A2 => IN1(7), B1 => n193, B2 => IN0(7), ZN
                           => n10);
   U8 : AOI22_X1 port map( A1 => IN3(7), A2 => n89, B1 => n90, B2 => IN2(7), ZN
                           => n11);
   U98 : AOI22_X1 port map( A1 => n6, A2 => IN1(0), B1 => n193, B2 => IN0(0), 
                           ZN => n68);
   U95 : AOI22_X1 port map( A1 => n89, A2 => IN3(0), B1 => n90, B2 => IN2(0), 
                           ZN => n69);
   U21 : AOI22_X1 port map( A1 => n6, A2 => IN1(3), B1 => n193, B2 => IN0(3), 
                           ZN => n18);
   U20 : AOI22_X1 port map( A1 => n89, A2 => IN3(3), B1 => n90, B2 => IN2(3), 
                           ZN => n19);
   U96 : NOR2_X1 port map( A1 => CTRL(0), A2 => n70, ZN => n5);
   U99 : NOR2_X1 port map( A1 => CTRL(0), A2 => CTRL(1), ZN => n7);
   U101 : INV_X1 port map( A => CTRL(1), ZN => n70);
   U100 : AND2_X2 port map( A1 => n70, A2 => CTRL(0), ZN => n6);
   U1 : NAND3_X1 port map( A1 => n169, A2 => n170, A3 => n171, ZN => OUT1(1));
   U2 : BUF_X2 port map( A => n194, Z => OUT1(7));
   U3 : OR2_X2 port map( A1 => n134, A2 => n135, ZN => OUT1(5));
   U4 : NAND2_X1 port map( A1 => n89, A2 => IN3(10), ZN => n71);
   U5 : NAND2_X1 port map( A1 => n90, A2 => IN2(10), ZN => n72);
   U6 : NAND2_X1 port map( A1 => n6, A2 => IN1(10), ZN => n73);
   U7 : NAND4_X1 port map( A1 => n181, A2 => n71, A3 => n72, A4 => n73, ZN => 
                           OUT1(10));
   U10 : AOI222_X1 port map( A1 => n90, A2 => IN2(8), B1 => IN0(8), B2 => n193,
                           C1 => n6, C2 => IN1(8), ZN => n74);
   U11 : NAND2_X1 port map( A1 => n89, A2 => IN3(8), ZN => n75);
   U12 : NAND2_X1 port map( A1 => n74, A2 => n75, ZN => OUT1(8));
   U13 : NAND2_X1 port map( A1 => n89, A2 => IN3(14), ZN => n76);
   U14 : NAND2_X1 port map( A1 => n90, A2 => IN2(14), ZN => n77);
   U15 : NAND2_X1 port map( A1 => n6, A2 => IN1(14), ZN => n78);
   U16 : NAND4_X1 port map( A1 => n121, A2 => n76, A3 => n77, A4 => n78, ZN => 
                           OUT1(14));
   U17 : AOI222_X1 port map( A1 => n7, A2 => IN0(4), B1 => n6, B2 => IN1(4), C1
                           => n5, C2 => IN2(4), ZN => n187);
   U18 : AOI222_X1 port map( A1 => n90, A2 => IN2(25), B1 => IN0(25), B2 => 
                           n193, C1 => n6, C2 => IN1(25), ZN => n79);
   U19 : NAND2_X1 port map( A1 => n89, A2 => IN3(25), ZN => n80);
   U22 : NAND2_X1 port map( A1 => n79, A2 => n80, ZN => OUT1(25));
   U23 : AOI22_X1 port map( A1 => IN0(29), A2 => n193, B1 => n6, B2 => IN1(29),
                           ZN => n81);
   U24 : INV_X1 port map( A => n81, ZN => n162);
   U25 : AOI22_X1 port map( A1 => IN0(18), A2 => n193, B1 => n6, B2 => IN1(18),
                           ZN => n82);
   U26 : INV_X1 port map( A => n82, ZN => n153);
   U27 : AOI22_X1 port map( A1 => IN0(5), A2 => n7, B1 => IN2(5), B2 => n5, ZN 
                           => n83);
   U28 : INV_X1 port map( A => n83, ZN => n133);
   U29 : NAND2_X1 port map( A1 => n89, A2 => IN3(22), ZN => n84);
   U30 : NAND2_X1 port map( A1 => n90, A2 => IN2(22), ZN => n85);
   U31 : NAND2_X1 port map( A1 => n6, A2 => IN1(22), ZN => n86);
   U32 : NAND4_X1 port map( A1 => n154, A2 => n84, A3 => n85, A4 => n86, ZN => 
                           OUT1(22));
   U33 : NAND2_X1 port map( A1 => n89, A2 => IN3(4), ZN => n87);
   U34 : NAND2_X1 port map( A1 => n187, A2 => n87, ZN => OUT1(4));
   U35 : NAND2_X4 port map( A1 => n151, A2 => n152, ZN => OUT1(18));
   U36 : NAND2_X1 port map( A1 => n11, A2 => n10, ZN => n194);
   U37 : NAND2_X2 port map( A1 => n122, A2 => n123, ZN => OUT1(15));
   U38 : OR3_X2 port map( A1 => n174, A2 => n175, A3 => n173, ZN => OUT1(2));
   U39 : BUF_X2 port map( A => n4, Z => n89);
   U40 : NAND2_X1 port map( A1 => n91, A2 => n92, ZN => OUT1(24));
   U41 : AND2_X1 port map( A1 => IN3(5), A2 => n89, ZN => n134);
   U42 : AND2_X1 port map( A1 => IN3(2), A2 => n89, ZN => n174);
   U43 : INV_X1 port map( A => n132, ZN => n135);
   U44 : INV_X1 port map( A => n172, ZN => n175);
   U45 : BUF_X2 port map( A => n7, Z => n193);
   U46 : BUF_X2 port map( A => n5, Z => n90);
   U47 : AND2_X1 port map( A1 => CTRL(0), A2 => CTRL(1), ZN => n4);
   U48 : NAND2_X1 port map( A1 => n127, A2 => n128, ZN => OUT1(17));
   U49 : NAND2_X1 port map( A1 => n160, A2 => n161, ZN => OUT1(29));
   U50 : NAND2_X1 port map( A1 => n182, A2 => n183, ZN => OUT1(16));
   U51 : NAND2_X1 port map( A1 => n136, A2 => n137, ZN => OUT1(20));
   U52 : AND2_X1 port map( A1 => IN1(2), A2 => n6, ZN => n173);
   U53 : NAND2_X1 port map( A1 => n111, A2 => n112, ZN => OUT1(21));
   U54 : NAND2_X1 port map( A1 => n106, A2 => n107, ZN => OUT1(23));
   U55 : NAND2_X1 port map( A1 => n146, A2 => n147, ZN => OUT1(11));
   U56 : NAND2_X1 port map( A1 => n141, A2 => n142, ZN => OUT1(19));
   U57 : NAND2_X1 port map( A1 => n62, A2 => n63, ZN => OUT1(12));
   U58 : NAND2_X1 port map( A1 => n101, A2 => n102, ZN => OUT1(31));
   U59 : NAND2_X1 port map( A1 => n68, A2 => n69, ZN => OUT1(0));
   U60 : NAND2_X1 port map( A1 => n116, A2 => n117, ZN => OUT1(26));
   U61 : NAND2_X1 port map( A1 => n60, A2 => n61, ZN => OUT1(13));
   U62 : NAND2_X1 port map( A1 => n18, A2 => n19, ZN => OUT1(3));
   U63 : NAND2_X1 port map( A1 => n155, A2 => n156, ZN => OUT1(27));
   U64 : NAND2_X1 port map( A1 => n163, A2 => n164, ZN => OUT1(30));
   U65 : NAND2_X1 port map( A1 => n177, A2 => n176, ZN => OUT1(28));
   U66 : NAND2_X1 port map( A1 => IN3(28), A2 => n89, ZN => n176);
   U67 : NAND2_X2 port map( A1 => n188, A2 => n189, ZN => OUT1(6));
   U68 : NAND2_X2 port map( A1 => n96, A2 => n97, ZN => OUT1(9));
   U69 : AOI21_X1 port map( B1 => IN2(17), B2 => n90, A => n129, ZN => n128);
   U70 : NAND2_X1 port map( A1 => n130, A2 => n131, ZN => n129);
   U71 : NAND2_X1 port map( A1 => n193, A2 => IN0(17), ZN => n131);
   U72 : NAND2_X1 port map( A1 => IN1(17), A2 => n6, ZN => n130);
   U73 : AOI21_X1 port map( B1 => IN2(16), B2 => n90, A => n184, ZN => n183);
   U74 : NAND2_X1 port map( A1 => n185, A2 => n186, ZN => n184);
   U75 : NAND2_X1 port map( A1 => n193, A2 => IN0(16), ZN => n186);
   U76 : NAND2_X1 port map( A1 => IN1(16), A2 => n6, ZN => n185);
   U77 : AOI21_X1 port map( B1 => IN2(19), B2 => n90, A => n143, ZN => n142);
   U78 : NAND2_X1 port map( A1 => n144, A2 => n145, ZN => n143);
   U79 : NAND2_X1 port map( A1 => n193, A2 => IN0(19), ZN => n145);
   U80 : NAND2_X1 port map( A1 => IN1(19), A2 => n6, ZN => n144);
   U81 : AOI21_X1 port map( B1 => IN2(18), B2 => n90, A => n153, ZN => n152);
   U82 : NAND2_X1 port map( A1 => n179, A2 => n180, ZN => n178);
   U85 : NAND2_X1 port map( A1 => n193, A2 => IN0(28), ZN => n180);
   U88 : NAND2_X1 port map( A1 => IN1(28), A2 => n6, ZN => n179);
   U89 : AOI21_X1 port map( B1 => IN2(27), B2 => n90, A => n157, ZN => n156);
   U90 : NAND2_X1 port map( A1 => n158, A2 => n159, ZN => n157);
   U91 : NAND2_X1 port map( A1 => n193, A2 => IN0(27), ZN => n159);
   U92 : NAND2_X1 port map( A1 => IN1(27), A2 => n6, ZN => n158);
   U93 : AOI21_X1 port map( B1 => IN2(30), B2 => n90, A => n165, ZN => n164);
   U94 : NAND2_X1 port map( A1 => n166, A2 => n167, ZN => n165);
   U97 : NAND2_X1 port map( A1 => n193, A2 => IN0(30), ZN => n167);
   U102 : NAND2_X1 port map( A1 => IN1(30), A2 => n6, ZN => n166);
   U103 : AOI21_X1 port map( B1 => IN2(23), B2 => n90, A => n108, ZN => n107);
   U104 : NAND2_X1 port map( A1 => n109, A2 => n110, ZN => n108);
   U105 : NAND2_X1 port map( A1 => n193, A2 => IN0(23), ZN => n110);
   U106 : NAND2_X1 port map( A1 => IN1(23), A2 => n6, ZN => n109);
   U107 : NAND2_X1 port map( A1 => n193, A2 => IN0(22), ZN => n154);
   U108 : AOI21_X1 port map( B1 => IN2(21), B2 => n90, A => n113, ZN => n112);
   U109 : NAND2_X1 port map( A1 => n114, A2 => n115, ZN => n113);
   U110 : NAND2_X1 port map( A1 => n193, A2 => IN0(21), ZN => n115);
   U111 : NAND2_X1 port map( A1 => IN1(21), A2 => n6, ZN => n114);
   U112 : AOI21_X1 port map( B1 => IN2(20), B2 => n90, A => n138, ZN => n137);
   U113 : NAND2_X1 port map( A1 => n139, A2 => n140, ZN => n138);
   U114 : NAND2_X1 port map( A1 => n193, A2 => IN0(20), ZN => n140);
   U115 : NAND2_X1 port map( A1 => IN1(20), A2 => n6, ZN => n139);
   U116 : AOI21_X1 port map( B1 => IN2(26), B2 => n90, A => n118, ZN => n117);
   U117 : NAND2_X1 port map( A1 => n119, A2 => n120, ZN => n118);
   U118 : NAND2_X1 port map( A1 => n193, A2 => IN0(26), ZN => n120);
   U119 : NAND2_X1 port map( A1 => IN1(26), A2 => n6, ZN => n119);
   U120 : AOI21_X1 port map( B1 => IN2(24), B2 => n90, A => n93, ZN => n92);
   U121 : NAND2_X1 port map( A1 => n94, A2 => n95, ZN => n93);
   U122 : NAND2_X1 port map( A1 => n193, A2 => IN0(24), ZN => n95);
   U123 : NAND2_X1 port map( A1 => IN1(24), A2 => n6, ZN => n94);
   U124 : AOI21_X1 port map( B1 => IN2(31), B2 => n90, A => n103, ZN => n102);
   U125 : NAND2_X1 port map( A1 => n104, A2 => n105, ZN => n103);
   U126 : NAND2_X1 port map( A1 => n193, A2 => IN0(31), ZN => n105);
   U127 : NAND2_X1 port map( A1 => IN1(31), A2 => n6, ZN => n104);
   U128 : AOI22_X1 port map( A1 => n90, A2 => IN2(2), B1 => n7, B2 => IN0(2), 
                           ZN => n172);
   U129 : NAND2_X1 port map( A1 => IN1(1), A2 => n6, ZN => n171);
   U130 : AOI22_X1 port map( A1 => n90, A2 => IN2(1), B1 => n193, B2 => IN0(1),
                           ZN => n170);
   U131 : AOI21_X1 port map( B1 => IN1(6), B2 => n6, A => n190, ZN => n189);
   U132 : NAND2_X1 port map( A1 => n191, A2 => n192, ZN => n190);
   U133 : NAND2_X1 port map( A1 => n193, A2 => IN0(6), ZN => n192);
   U134 : NAND2_X1 port map( A1 => n90, A2 => IN2(6), ZN => n191);
   U135 : AOI21_X1 port map( B1 => IN1(5), B2 => n6, A => n133, ZN => n132);
   U136 : AOI21_X1 port map( B1 => IN2(11), B2 => n90, A => n148, ZN => n147);
   U137 : NAND2_X1 port map( A1 => n149, A2 => n150, ZN => n148);
   U138 : NAND2_X1 port map( A1 => n193, A2 => IN0(11), ZN => n150);
   U139 : NAND2_X1 port map( A1 => IN1(11), A2 => n6, ZN => n149);
   U140 : NAND2_X1 port map( A1 => n193, A2 => IN0(10), ZN => n181);
   U141 : AOI21_X1 port map( B1 => IN2(9), B2 => n90, A => n98, ZN => n97);
   U142 : NAND2_X1 port map( A1 => n99, A2 => n100, ZN => n98);
   U143 : NAND2_X1 port map( A1 => n193, A2 => IN0(9), ZN => n100);
   U144 : NAND2_X1 port map( A1 => IN1(9), A2 => n6, ZN => n99);
   U145 : AOI21_X1 port map( B1 => IN2(15), B2 => n90, A => n124, ZN => n123);
   U146 : NAND2_X1 port map( A1 => n125, A2 => n126, ZN => n124);
   U147 : NAND2_X1 port map( A1 => n193, A2 => IN0(15), ZN => n126);
   U148 : NAND2_X1 port map( A1 => IN1(15), A2 => n6, ZN => n125);
   U149 : NAND2_X1 port map( A1 => n193, A2 => IN0(14), ZN => n121);
   U150 : NAND2_X1 port map( A1 => IN3(24), A2 => n4, ZN => n91);
   U151 : NAND2_X1 port map( A1 => IN3(9), A2 => n89, ZN => n96);
   U152 : NAND2_X1 port map( A1 => IN3(31), A2 => n89, ZN => n101);
   U153 : NAND2_X1 port map( A1 => IN3(23), A2 => n89, ZN => n106);
   U154 : NAND2_X1 port map( A1 => IN3(21), A2 => n89, ZN => n111);
   U155 : NAND2_X1 port map( A1 => IN3(26), A2 => n89, ZN => n116);
   U156 : NAND2_X1 port map( A1 => IN3(15), A2 => n89, ZN => n122);
   U157 : NAND2_X1 port map( A1 => IN3(17), A2 => n89, ZN => n127);
   U158 : NAND2_X1 port map( A1 => IN3(20), A2 => n89, ZN => n136);
   U159 : NAND2_X1 port map( A1 => IN3(19), A2 => n89, ZN => n141);
   U160 : NAND2_X1 port map( A1 => IN3(11), A2 => n89, ZN => n146);
   U161 : NAND2_X1 port map( A1 => IN3(18), A2 => n89, ZN => n151);
   U162 : NAND2_X1 port map( A1 => IN3(27), A2 => n89, ZN => n155);
   U163 : NAND2_X1 port map( A1 => IN3(29), A2 => n4, ZN => n160);
   U164 : AOI21_X1 port map( B1 => IN2(29), B2 => n90, A => n162, ZN => n161);
   U165 : NAND2_X1 port map( A1 => IN3(30), A2 => n4, ZN => n163);
   U166 : NAND2_X1 port map( A1 => IN3(1), A2 => n89, ZN => n169);
   U167 : AOI21_X1 port map( B1 => IN2(28), B2 => n90, A => n178, ZN => n177);
   U168 : NAND2_X1 port map( A1 => IN3(16), A2 => n89, ZN => n182);
   U169 : NAND2_X1 port map( A1 => IN3(6), A2 => n89, ZN => n188);

end SYN_bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity add4 is

   port( IN1 : in std_logic_vector (31 downto 0);  OUT1 : out std_logic_vector 
         (31 downto 0));

end add4;

architecture SYN_bhe of add4 is

   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal OUT1_31_port, OUT1_30_port, OUT1_29_port, OUT1_28_port, OUT1_27_port,
      OUT1_26_port, OUT1_25_port, OUT1_24_port, OUT1_23_port, OUT1_22_port, 
      OUT1_21_port, OUT1_20_port, OUT1_19_port, OUT1_18_port, OUT1_17_port, 
      OUT1_16_port, OUT1_15_port, OUT1_14_port, OUT1_13_port, OUT1_12_port, 
      OUT1_11_port, OUT1_10_port, OUT1_9_port, OUT1_8_port, OUT1_7_port, 
      OUT1_6_port, OUT1_5_port, OUT1_4_port, OUT1_3_port, OUT1_2_port, 
      add_27_carry_4_port, add_27_carry_5_port, add_27_carry_6_port, 
      add_27_carry_7_port, add_27_carry_8_port, add_27_carry_9_port, 
      add_27_carry_10_port, add_27_carry_11_port, add_27_carry_12_port, 
      add_27_carry_13_port, add_27_carry_14_port, add_27_carry_15_port, 
      add_27_carry_16_port, add_27_carry_17_port, add_27_carry_18_port, 
      add_27_carry_19_port, add_27_carry_20_port, add_27_carry_21_port, 
      add_27_carry_22_port, add_27_carry_23_port, add_27_carry_24_port, 
      add_27_carry_25_port, add_27_carry_26_port, add_27_carry_27_port, 
      add_27_carry_28_port, add_27_carry_29_port, add_27_carry_30_port, n1 : 
      std_logic;

begin
   OUT1 <= ( OUT1_31_port, OUT1_30_port, OUT1_29_port, OUT1_28_port, 
      OUT1_27_port, OUT1_26_port, OUT1_25_port, OUT1_24_port, OUT1_23_port, 
      OUT1_22_port, OUT1_21_port, OUT1_20_port, OUT1_19_port, OUT1_18_port, 
      OUT1_17_port, OUT1_16_port, OUT1_15_port, OUT1_14_port, OUT1_13_port, 
      OUT1_12_port, OUT1_11_port, OUT1_10_port, OUT1_9_port, OUT1_8_port, 
      OUT1_7_port, OUT1_6_port, OUT1_5_port, OUT1_4_port, OUT1_3_port, 
      OUT1_2_port, IN1(1), IN1(0) );
   
   add_27_U57 : XOR2_X1 port map( A => IN1(3), B => IN1(2), Z => OUT1_3_port);
   add_27_U55 : XOR2_X1 port map( A => IN1(4), B => add_27_carry_4_port, Z => 
                           OUT1_4_port);
   add_27_U53 : XOR2_X1 port map( A => IN1(5), B => add_27_carry_5_port, Z => 
                           OUT1_5_port);
   add_27_U51 : XOR2_X1 port map( A => IN1(6), B => add_27_carry_6_port, Z => 
                           OUT1_6_port);
   add_27_U49 : XOR2_X1 port map( A => IN1(7), B => add_27_carry_7_port, Z => 
                           OUT1_7_port);
   add_27_U47 : XOR2_X1 port map( A => IN1(8), B => add_27_carry_8_port, Z => 
                           OUT1_8_port);
   add_27_U45 : XOR2_X1 port map( A => IN1(9), B => add_27_carry_9_port, Z => 
                           OUT1_9_port);
   add_27_U43 : XOR2_X1 port map( A => IN1(10), B => add_27_carry_10_port, Z =>
                           OUT1_10_port);
   add_27_U41 : XOR2_X1 port map( A => IN1(11), B => add_27_carry_11_port, Z =>
                           OUT1_11_port);
   add_27_U39 : XOR2_X1 port map( A => IN1(12), B => add_27_carry_12_port, Z =>
                           OUT1_12_port);
   add_27_U37 : XOR2_X1 port map( A => IN1(13), B => add_27_carry_13_port, Z =>
                           OUT1_13_port);
   add_27_U35 : XOR2_X1 port map( A => IN1(14), B => add_27_carry_14_port, Z =>
                           OUT1_14_port);
   add_27_U33 : XOR2_X1 port map( A => IN1(15), B => add_27_carry_15_port, Z =>
                           OUT1_15_port);
   add_27_U31 : XOR2_X1 port map( A => IN1(16), B => add_27_carry_16_port, Z =>
                           OUT1_16_port);
   add_27_U29 : XOR2_X1 port map( A => IN1(17), B => add_27_carry_17_port, Z =>
                           OUT1_17_port);
   add_27_U27 : XOR2_X1 port map( A => IN1(18), B => add_27_carry_18_port, Z =>
                           OUT1_18_port);
   add_27_U25 : XOR2_X1 port map( A => IN1(19), B => add_27_carry_19_port, Z =>
                           OUT1_19_port);
   add_27_U23 : XOR2_X1 port map( A => IN1(20), B => add_27_carry_20_port, Z =>
                           OUT1_20_port);
   add_27_U21 : XOR2_X1 port map( A => IN1(21), B => add_27_carry_21_port, Z =>
                           OUT1_21_port);
   add_27_U19 : XOR2_X1 port map( A => IN1(22), B => add_27_carry_22_port, Z =>
                           OUT1_22_port);
   add_27_U17 : XOR2_X1 port map( A => IN1(23), B => add_27_carry_23_port, Z =>
                           OUT1_23_port);
   add_27_U15 : XOR2_X1 port map( A => IN1(24), B => add_27_carry_24_port, Z =>
                           OUT1_24_port);
   add_27_U13 : XOR2_X1 port map( A => IN1(25), B => add_27_carry_25_port, Z =>
                           OUT1_25_port);
   add_27_U11 : XOR2_X1 port map( A => IN1(26), B => add_27_carry_26_port, Z =>
                           OUT1_26_port);
   add_27_U9 : XOR2_X1 port map( A => IN1(27), B => add_27_carry_27_port, Z => 
                           OUT1_27_port);
   add_27_U7 : XOR2_X1 port map( A => IN1(28), B => add_27_carry_28_port, Z => 
                           OUT1_28_port);
   add_27_U5 : XOR2_X1 port map( A => IN1(29), B => add_27_carry_29_port, Z => 
                           OUT1_29_port);
   add_27_U3 : XOR2_X1 port map( A => IN1(30), B => add_27_carry_30_port, Z => 
                           OUT1_30_port);
   add_27_U58 : INV_X1 port map( A => IN1(2), ZN => OUT1_2_port);
   add_27_U36 : AND2_X1 port map( A1 => add_27_carry_13_port, A2 => IN1(13), ZN
                           => add_27_carry_14_port);
   add_27_U34 : AND2_X1 port map( A1 => add_27_carry_14_port, A2 => IN1(14), ZN
                           => add_27_carry_15_port);
   add_27_U32 : AND2_X1 port map( A1 => add_27_carry_15_port, A2 => IN1(15), ZN
                           => add_27_carry_16_port);
   add_27_U30 : AND2_X1 port map( A1 => add_27_carry_16_port, A2 => IN1(16), ZN
                           => add_27_carry_17_port);
   add_27_U28 : AND2_X1 port map( A1 => add_27_carry_17_port, A2 => IN1(17), ZN
                           => add_27_carry_18_port);
   add_27_U26 : AND2_X1 port map( A1 => add_27_carry_18_port, A2 => IN1(18), ZN
                           => add_27_carry_19_port);
   add_27_U12 : AND2_X1 port map( A1 => add_27_carry_25_port, A2 => IN1(25), ZN
                           => add_27_carry_26_port);
   add_27_U10 : AND2_X1 port map( A1 => add_27_carry_26_port, A2 => IN1(26), ZN
                           => add_27_carry_27_port);
   add_27_U8 : AND2_X1 port map( A1 => add_27_carry_27_port, A2 => IN1(27), ZN 
                           => add_27_carry_28_port);
   add_27_U6 : AND2_X1 port map( A1 => add_27_carry_28_port, A2 => IN1(28), ZN 
                           => add_27_carry_29_port);
   add_27_U4 : AND2_X1 port map( A1 => add_27_carry_29_port, A2 => IN1(29), ZN 
                           => add_27_carry_30_port);
   U3 : AND2_X1 port map( A1 => IN1(2), A2 => IN1(3), ZN => add_27_carry_4_port
                           );
   U4 : AND2_X1 port map( A1 => add_27_carry_4_port, A2 => IN1(4), ZN => 
                           add_27_carry_5_port);
   U5 : AND2_X1 port map( A1 => add_27_carry_19_port, A2 => IN1(19), ZN => 
                           add_27_carry_20_port);
   U6 : AND2_X1 port map( A1 => add_27_carry_24_port, A2 => IN1(24), ZN => 
                           add_27_carry_25_port);
   U7 : NAND2_X1 port map( A1 => add_27_carry_30_port, A2 => IN1(30), ZN => n1)
                           ;
   U8 : XNOR2_X1 port map( A => n1, B => IN1(31), ZN => OUT1_31_port);
   U9 : AND2_X2 port map( A1 => add_27_carry_23_port, A2 => IN1(23), ZN => 
                           add_27_carry_24_port);
   U10 : AND2_X2 port map( A1 => add_27_carry_22_port, A2 => IN1(22), ZN => 
                           add_27_carry_23_port);
   U11 : AND2_X2 port map( A1 => add_27_carry_20_port, A2 => IN1(20), ZN => 
                           add_27_carry_21_port);
   U12 : AND2_X2 port map( A1 => add_27_carry_21_port, A2 => IN1(21), ZN => 
                           add_27_carry_22_port);
   U13 : AND2_X2 port map( A1 => add_27_carry_6_port, A2 => IN1(6), ZN => 
                           add_27_carry_7_port);
   U14 : AND2_X2 port map( A1 => add_27_carry_5_port, A2 => IN1(5), ZN => 
                           add_27_carry_6_port);
   U15 : AND2_X2 port map( A1 => add_27_carry_8_port, A2 => IN1(8), ZN => 
                           add_27_carry_9_port);
   U16 : AND2_X2 port map( A1 => add_27_carry_7_port, A2 => IN1(7), ZN => 
                           add_27_carry_8_port);
   U17 : AND2_X2 port map( A1 => add_27_carry_10_port, A2 => IN1(10), ZN => 
                           add_27_carry_11_port);
   U18 : AND2_X2 port map( A1 => add_27_carry_9_port, A2 => IN1(9), ZN => 
                           add_27_carry_10_port);
   U19 : AND2_X2 port map( A1 => add_27_carry_12_port, A2 => IN1(12), ZN => 
                           add_27_carry_13_port);
   U20 : AND2_X2 port map( A1 => add_27_carry_11_port, A2 => IN1(11), ZN => 
                           add_27_carry_12_port);

end SYN_bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity ff32_en_0 is

   port( D : in std_logic_vector (31 downto 0);  en, clk, rst : in std_logic;  
         Q : out std_logic_vector (31 downto 0));

end ff32_en_0;

architecture SYN_behavioral of ff32_en_0 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_31_port, Q_30_port, Q_29_port, Q_28_port, Q_27_port, Q_26_port, 
      Q_25_port, Q_24_port, Q_23_port, Q_22_port, Q_21_port, Q_20_port, 
      Q_19_port, Q_18_port, Q_17_port, Q_16_port, Q_15_port, Q_14_port, 
      Q_13_port, Q_12_port, Q_11_port, Q_10_port, Q_9_port, Q_8_port, Q_7_port,
      Q_6_port, Q_5_port, Q_4_port, Q_3_port, Q_2_port, Q_1_port, Q_0_port, n65
      , n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, 
      n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94
      , n95, n97, net644934, net644935, net644936, net644937, net644938, 
      net644939, net644940, net644941, net644942, net644943, net644944, 
      net644945, net644946, net644947, net644948, net644949, net644950, 
      net644951, net644952, net644953, net644954, net644955, net644956, 
      net644957, net644958, net644959, net644960, net644961, net644962, 
      net644963, net644964, net644965, n3, n5, n8, n9, n12, n13, n20, n25, n27,
      n32, n33, n29, n11, n14, n16, n28, n17, n31, n30, n10, n15, n23, n4, n6, 
      n19, n26, n7, n24, n2, n18, n1, n21, n22, n34, n36, n37, n38, n39 : 
      std_logic;

begin
   Q <= ( Q_31_port, Q_30_port, Q_29_port, Q_28_port, Q_27_port, Q_26_port, 
      Q_25_port, Q_24_port, Q_23_port, Q_22_port, Q_21_port, Q_20_port, 
      Q_19_port, Q_18_port, Q_17_port, Q_16_port, Q_15_port, Q_14_port, 
      Q_13_port, Q_12_port, Q_11_port, Q_10_port, Q_9_port, Q_8_port, Q_7_port,
      Q_6_port, Q_5_port, Q_4_port, Q_3_port, Q_2_port, Q_1_port, Q_0_port );
   
   Q_reg_30_inst : DFFR_X1 port map( D => n95, CK => clk, RN => n39, Q => 
                           Q_30_port, QN => net644964);
   Q_reg_29_inst : DFFR_X1 port map( D => n94, CK => clk, RN => n39, Q => 
                           Q_29_port, QN => net644963);
   Q_reg_28_inst : DFFR_X1 port map( D => n93, CK => clk, RN => n39, Q => 
                           Q_28_port, QN => net644962);
   Q_reg_27_inst : DFFR_X1 port map( D => n92, CK => clk, RN => n39, Q => 
                           Q_27_port, QN => net644961);
   Q_reg_26_inst : DFFR_X1 port map( D => n91, CK => clk, RN => n39, Q => 
                           Q_26_port, QN => net644960);
   Q_reg_25_inst : DFFR_X1 port map( D => n90, CK => clk, RN => n39, Q => 
                           Q_25_port, QN => net644959);
   Q_reg_24_inst : DFFR_X1 port map( D => n89, CK => clk, RN => n39, Q => 
                           Q_24_port, QN => net644958);
   Q_reg_23_inst : DFFR_X1 port map( D => n88, CK => clk, RN => n39, Q => 
                           Q_23_port, QN => net644957);
   Q_reg_22_inst : DFFR_X1 port map( D => n87, CK => clk, RN => n39, Q => 
                           Q_22_port, QN => net644956);
   Q_reg_21_inst : DFFR_X1 port map( D => n86, CK => clk, RN => n39, Q => 
                           Q_21_port, QN => net644955);
   Q_reg_20_inst : DFFR_X1 port map( D => n85, CK => clk, RN => n39, Q => 
                           Q_20_port, QN => net644954);
   Q_reg_19_inst : DFFR_X1 port map( D => n84, CK => clk, RN => n39, Q => 
                           Q_19_port, QN => net644953);
   Q_reg_18_inst : DFFR_X1 port map( D => n83, CK => clk, RN => n39, Q => 
                           Q_18_port, QN => net644952);
   Q_reg_17_inst : DFFR_X1 port map( D => n82, CK => clk, RN => n39, Q => 
                           Q_17_port, QN => net644951);
   Q_reg_16_inst : DFFR_X1 port map( D => n81, CK => clk, RN => n39, Q => 
                           Q_16_port, QN => net644950);
   Q_reg_15_inst : DFFR_X1 port map( D => n80, CK => clk, RN => n39, Q => 
                           Q_15_port, QN => net644949);
   Q_reg_14_inst : DFFR_X1 port map( D => n79, CK => clk, RN => n39, Q => 
                           Q_14_port, QN => net644948);
   Q_reg_12_inst : DFFR_X1 port map( D => n77, CK => clk, RN => n39, Q => 
                           Q_12_port, QN => net644946);
   Q_reg_10_inst : DFFR_X1 port map( D => n75, CK => clk, RN => n39, Q => 
                           Q_10_port, QN => net644944);
   Q_reg_9_inst : DFFR_X1 port map( D => n74, CK => clk, RN => n39, Q => 
                           Q_9_port, QN => net644943);
   Q_reg_8_inst : DFFR_X1 port map( D => n73, CK => clk, RN => n39, Q => 
                           Q_8_port, QN => net644942);
   Q_reg_7_inst : DFFR_X1 port map( D => n72, CK => clk, RN => n39, Q => 
                           Q_7_port, QN => net644941);
   Q_reg_6_inst : DFFR_X1 port map( D => n71, CK => clk, RN => n39, Q => 
                           Q_6_port, QN => net644940);
   Q_reg_5_inst : DFFR_X1 port map( D => n70, CK => clk, RN => n39, Q => 
                           Q_5_port, QN => net644939);
   Q_reg_4_inst : DFFR_X1 port map( D => n69, CK => clk, RN => n39, Q => 
                           Q_4_port, QN => net644938);
   Q_reg_3_inst : DFFR_X1 port map( D => n68, CK => clk, RN => n39, Q => 
                           Q_3_port, QN => net644937);
   Q_reg_2_inst : DFFR_X1 port map( D => n67, CK => clk, RN => n39, Q => 
                           Q_2_port, QN => net644936);
   Q_reg_1_inst : DFFR_X1 port map( D => n66, CK => clk, RN => n39, Q => 
                           Q_1_port, QN => net644935);
   Q_reg_0_inst : DFFR_X1 port map( D => n65, CK => clk, RN => n39, Q => 
                           Q_0_port, QN => net644934);
   Q_reg_13_inst : DFFR_X1 port map( D => n78, CK => clk, RN => n39, Q => 
                           Q_13_port, QN => net644947);
   Q_reg_31_inst : DFFR_X1 port map( D => n97, CK => clk, RN => n39, Q => 
                           Q_31_port, QN => net644965);
   Q_reg_11_inst : DFFR_X1 port map( D => n76, CK => clk, RN => n39, Q => 
                           Q_11_port, QN => net644945);
   U2 : NAND2_X1 port map( A1 => n37, A2 => D(11), ZN => n1);
   U3 : OAI21_X1 port map( B1 => en, B2 => net644945, A => n1, ZN => n76);
   U4 : INV_X1 port map( A => Q_12_port, ZN => n21);
   U5 : NAND2_X1 port map( A1 => D(12), A2 => n36, ZN => n22);
   U6 : OAI21_X1 port map( B1 => n21, B2 => en, A => n22, ZN => n77);
   U7 : OR2_X1 port map( A1 => en, A2 => net644965, ZN => n34);
   U8 : NAND2_X1 port map( A1 => n34, A2 => n2, ZN => n97);
   U9 : INV_X2 port map( A => rst, ZN => n39);
   U10 : BUF_X1 port map( A => en, Z => n36);
   U11 : BUF_X1 port map( A => en, Z => n37);
   U12 : BUF_X1 port map( A => en, Z => n38);
   U13 : OAI21_X1 port map( B1 => en, B2 => net644949, A => n18, ZN => n80);
   U14 : OAI21_X1 port map( B1 => en, B2 => net644944, A => n23, ZN => n75);
   U15 : OAI21_X1 port map( B1 => en, B2 => net644952, A => n15, ZN => n83);
   U16 : OAI21_X1 port map( B1 => en, B2 => net644948, A => n19, ZN => n79);
   U17 : OAI21_X1 port map( B1 => en, B2 => net644950, A => n17, ZN => n81);
   U18 : OAI21_X1 port map( B1 => en, B2 => net644951, A => n16, ZN => n82);
   U19 : NAND2_X1 port map( A1 => D(15), A2 => en, ZN => n18);
   U20 : NAND2_X1 port map( A1 => en, A2 => D(31), ZN => n2);
   U21 : NAND2_X1 port map( A1 => D(9), A2 => en, ZN => n24);
   U22 : OAI21_X1 port map( B1 => en, B2 => net644943, A => n24, ZN => n74);
   U23 : NAND2_X1 port map( A1 => n38, A2 => D(26), ZN => n7);
   U24 : OAI21_X1 port map( B1 => n36, B2 => net644960, A => n7, ZN => n91);
   U25 : NAND2_X1 port map( A1 => D(7), A2 => en, ZN => n26);
   U26 : OAI21_X1 port map( B1 => en, B2 => net644941, A => n26, ZN => n72);
   U27 : NAND2_X1 port map( A1 => D(14), A2 => n37, ZN => n19);
   U28 : NAND2_X1 port map( A1 => n38, A2 => D(27), ZN => n6);
   U29 : OAI21_X1 port map( B1 => n36, B2 => net644961, A => n6, ZN => n92);
   U30 : NAND2_X1 port map( A1 => D(29), A2 => n38, ZN => n4);
   U31 : OAI21_X1 port map( B1 => n36, B2 => net644963, A => n4, ZN => n94);
   U32 : NAND2_X1 port map( A1 => D(10), A2 => n37, ZN => n23);
   U33 : NAND2_X1 port map( A1 => D(18), A2 => en, ZN => n15);
   U34 : NAND2_X1 port map( A1 => n38, A2 => D(23), ZN => n10);
   U35 : OAI21_X1 port map( B1 => n36, B2 => net644957, A => n10, ZN => n88);
   U36 : NAND2_X1 port map( A1 => D(3), A2 => n38, ZN => n30);
   U37 : OAI21_X1 port map( B1 => n37, B2 => net644937, A => n30, ZN => n68);
   U38 : NAND2_X1 port map( A1 => n38, A2 => D(2), ZN => n31);
   U39 : OAI21_X1 port map( B1 => n37, B2 => net644936, A => n31, ZN => n67);
   U40 : NAND2_X1 port map( A1 => D(16), A2 => en, ZN => n17);
   U41 : NAND2_X1 port map( A1 => D(5), A2 => n38, ZN => n28);
   U42 : OAI21_X1 port map( B1 => n37, B2 => net644939, A => n28, ZN => n70);
   U43 : NAND2_X1 port map( A1 => D(17), A2 => en, ZN => n16);
   U44 : NAND2_X1 port map( A1 => D(19), A2 => n38, ZN => n14);
   U45 : OAI21_X1 port map( B1 => n36, B2 => net644953, A => n14, ZN => n84);
   U46 : NAND2_X1 port map( A1 => D(22), A2 => en, ZN => n11);
   U47 : OAI21_X1 port map( B1 => n36, B2 => net644956, A => n11, ZN => n87);
   U48 : NAND2_X1 port map( A1 => n38, A2 => D(4), ZN => n29);
   U49 : OAI21_X1 port map( B1 => n37, B2 => net644938, A => n29, ZN => n69);
   U50 : OAI21_X1 port map( B1 => n37, B2 => net644934, A => n33, ZN => n65);
   U51 : OAI21_X1 port map( B1 => n36, B2 => net644955, A => n12, ZN => n86);
   U52 : OAI21_X1 port map( B1 => n36, B2 => net644962, A => n5, ZN => n93);
   U53 : NAND2_X1 port map( A1 => n38, A2 => D(28), ZN => n5);
   U54 : OAI21_X1 port map( B1 => n36, B2 => net644964, A => n3, ZN => n95);
   U55 : NAND2_X1 port map( A1 => en, A2 => D(30), ZN => n3);
   U56 : OAI21_X1 port map( B1 => n36, B2 => net644958, A => n9, ZN => n89);
   U57 : NAND2_X1 port map( A1 => D(24), A2 => n38, ZN => n9);
   U58 : OAI21_X1 port map( B1 => n36, B2 => net644959, A => n8, ZN => n90);
   U59 : NAND2_X1 port map( A1 => n38, A2 => D(25), ZN => n8);
   U60 : OAI21_X1 port map( B1 => n36, B2 => net644954, A => n13, ZN => n85);
   U61 : NAND2_X1 port map( A1 => D(20), A2 => n36, ZN => n13);
   U62 : OAI21_X1 port map( B1 => n37, B2 => net644942, A => n25, ZN => n73);
   U63 : NAND2_X1 port map( A1 => D(8), A2 => n37, ZN => n25);
   U64 : NAND2_X1 port map( A1 => en, A2 => D(0), ZN => n33);
   U65 : OAI21_X1 port map( B1 => n37, B2 => net644940, A => n27, ZN => n71);
   U66 : NAND2_X1 port map( A1 => D(6), A2 => n38, ZN => n27);
   U67 : OAI21_X1 port map( B1 => n37, B2 => net644935, A => n32, ZN => n66);
   U68 : NAND2_X1 port map( A1 => en, A2 => D(1), ZN => n32);
   U69 : NAND2_X1 port map( A1 => n38, A2 => D(21), ZN => n12);
   U70 : OAI21_X1 port map( B1 => en, B2 => net644947, A => n20, ZN => n78);
   U71 : NAND2_X1 port map( A1 => D(13), A2 => n37, ZN => n20);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity fw_logic is

   port( D1_i, rAdec_i, D2_i, D3_i, rA_i, rB_i : in std_logic_vector (4 downto 
         0);  S_mem_W, S_wb_W, S_exe_W : in std_logic;  S_FWAdec, S_FWA, S_FWB 
         : out std_logic_vector (1 downto 0);  S_mem_LOAD_BAR : in std_logic);

end fw_logic;

architecture SYN_beh of fw_logic is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X2
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n102, n103, n22, n24, n25, n28, n29, n30, n31, n32, n34, n35, n36, 
      n37, n38, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57
      , n58, n59, n60, n61, n62, n63, n64, n44, n43, n42, n41, n40, n39, n101, 
      n65, n66, n67, n69, n70, n71, n73, n74, n75, n76, n77, n78, n79, n80, n81
      , n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, 
      n96, n97, n99, n100 : std_logic;

begin
   
   U53 : XOR2_X1 port map( A => D2_i(2), B => rB_i(2), Z => n29);
   U54 : XOR2_X1 port map( A => D2_i(2), B => rAdec_i(2), Z => n45);
   U55 : XOR2_X1 port map( A => D2_i(2), B => rA_i(2), Z => n60);
   U39 : OAI221_X1 port map( B1 => rA_i(3), B2 => n28, C1 => n59, C2 => n67, A 
                           => S_wb_W, ZN => n50);
   U24 : INV_X1 port map( A => rAdec_i(3), ZN => n44);
   U40 : INV_X1 port map( A => rA_i(3), ZN => n59);
   U37 : INV_X1 port map( A => rA_i(2), ZN => n57);
   U38 : INV_X1 port map( A => rA_i(1), ZN => n56);
   U33 : INV_X1 port map( A => rA_i(0), ZN => n54);
   U34 : INV_X1 port map( A => rA_i(4), ZN => n53);
   U2 : OR2_X1 port map( A1 => n94, A2 => rB_i(1), ZN => n99);
   U3 : CLKBUF_X1 port map( A => n66, Z => n73);
   U4 : INV_X1 port map( A => D2_i(1), ZN => n97);
   U5 : OR2_X1 port map( A1 => n34, A2 => rB_i(3), ZN => n100);
   U6 : INV_X1 port map( A => n90, ZN => n76);
   U7 : CLKBUF_X1 port map( A => D3_i(1), Z => n65);
   U8 : INV_X1 port map( A => D3_i(2), ZN => n25);
   U9 : CLKBUF_X1 port map( A => D3_i(0), Z => n91);
   U10 : OR2_X1 port map( A1 => n96, A2 => rAdec_i(4), ZN => n92);
   U11 : INV_X1 port map( A => D3_i(4), ZN => n66);
   U12 : INV_X1 port map( A => n28, ZN => n67);
   U13 : INV_X1 port map( A => D3_i(3), ZN => n28);
   U14 : NOR4_X1 port map( A1 => n60, A2 => n62, A3 => n61, A4 => n30, ZN => 
                           S_FWA(0));
   U15 : NOR4_X1 port map( A1 => n60, A2 => n62, A3 => n61, A4 => n30, ZN => 
                           n102);
   U16 : INV_X1 port map( A => n91, ZN => n69);
   U17 : OR2_X1 port map( A1 => n37, A2 => rAdec_i(0), ZN => n93);
   U18 : AOI22_X1 port map( A1 => n36, A2 => rAdec_i(4), B1 => rAdec_i(0), B2 
                           => n37, ZN => n49);
   U19 : CLKBUF_X1 port map( A => D3_i(4), Z => n70);
   U20 : INV_X1 port map( A => D2_i(1), ZN => n94);
   U21 : OAI221_X1 port map( B1 => n97, B2 => rAdec_i(1), C1 => n34, C2 => 
                           rAdec_i(3), A => n48, ZN => n47);
   U22 : NAND3_X1 port map( A1 => n92, A2 => n93, A3 => n49, ZN => n46);
   U23 : CLKBUF_X1 port map( A => n30, Z => n71);
   U25 : INV_X1 port map( A => D3_i(0), ZN => n22);
   U26 : NOR3_X1 port map( A1 => n31, A2 => n32, A3 => n95, ZN => S_FWB(0));
   U27 : NAND2_X1 port map( A1 => S_mem_W, A2 => S_mem_LOAD_BAR, ZN => n30);
   U28 : NOR4_X1 port map( A1 => n47, A2 => n46, A3 => n30, A4 => n45, ZN => 
                           n101);
   U29 : NOR4_X1 port map( A1 => n102, A2 => n50, A3 => n51, A4 => n52, ZN => 
                           S_FWA(1));
   U30 : INV_X1 port map( A => D3_i(1), ZN => n88);
   U31 : INV_X1 port map( A => D3_i(1), ZN => n24);
   U32 : OR2_X1 port map( A1 => n41, A2 => n39, ZN => n74);
   U35 : INV_X1 port map( A => S_wb_W, ZN => n83);
   U36 : INV_X1 port map( A => D3_i(3), ZN => n82);
   U41 : NOR3_X1 port map( A1 => n101, A2 => n40, A3 => n74, ZN => S_FWAdec(1))
                           ;
   U42 : INV_X1 port map( A => n79, ZN => n78);
   U43 : NOR3_X1 port map( A1 => n31, A2 => n32, A3 => n95, ZN => n103);
   U44 : OR2_X1 port map( A1 => n29, A2 => n30, ZN => n95);
   U45 : INV_X1 port map( A => D2_i(4), ZN => n36);
   U46 : NOR4_X2 port map( A1 => n45, A2 => n71, A3 => n46, A4 => n47, ZN => 
                           S_FWAdec(0));
   U47 : OAI221_X1 port map( B1 => n24, B2 => rAdec_i(1), C1 => n25, C2 => 
                           rAdec_i(2), A => n43, ZN => n40);
   U48 : OAI22_X1 port map( A1 => rB_i(3), A2 => n28, B1 => n69, B2 => rB_i(0),
                           ZN => n90);
   U49 : NOR2_X1 port map( A1 => n75, A2 => n103, ZN => S_FWB(1));
   U50 : NAND3_X1 port map( A1 => n77, A2 => n76, A3 => n78, ZN => n75);
   U51 : NAND2_X1 port map( A1 => n88, A2 => rB_i(1), ZN => n87);
   U52 : AOI21_X1 port map( B1 => n82, B2 => rB_i(3), A => n83, ZN => n80);
   U56 : OAI211_X1 port map( C1 => n24, C2 => rB_i(1), A => n81, B => n80, ZN 
                           => n79);
   U57 : NAND2_X1 port map( A1 => n66, A2 => rB_i(4), ZN => n89);
   U58 : OAI21_X1 port map( B1 => n73, B2 => rB_i(4), A => n89, ZN => n84);
   U59 : NAND2_X1 port map( A1 => n22, A2 => rB_i(0), ZN => n86);
   U60 : OAI211_X1 port map( C1 => rB_i(2), C2 => n25, A => n86, B => n87, ZN 
                           => n85);
   U61 : NAND2_X1 port map( A1 => n25, A2 => rB_i(2), ZN => n81);
   U62 : NOR2_X1 port map( A1 => n84, A2 => n85, ZN => n77);
   U63 : AOI22_X1 port map( A1 => n66, A2 => rAdec_i(4), B1 => n22, B2 => 
                           rAdec_i(0), ZN => n42);
   U64 : OAI221_X1 port map( B1 => D3_i(3), B2 => n44, C1 => n28, C2 => 
                           rAdec_i(3), A => S_wb_W, ZN => n39);
   U65 : OAI221_X1 port map( B1 => n73, B2 => rAdec_i(4), C1 => n69, C2 => 
                           rAdec_i(0), A => n42, ZN => n41);
   U66 : AOI22_X1 port map( A1 => n24, A2 => rAdec_i(1), B1 => rAdec_i(2), B2 
                           => n25, ZN => n43);
   U67 : INV_X1 port map( A => D2_i(4), ZN => n96);
   U68 : OAI221_X1 port map( B1 => n96, B2 => rA_i(4), C1 => n37, C2 => rA_i(0)
                           , A => n64, ZN => n61);
   U69 : OAI221_X1 port map( B1 => n94, B2 => rA_i(1), C1 => n34, C2 => rA_i(3)
                           , A => n63, ZN => n62);
   U70 : OAI221_X1 port map( B1 => n36, B2 => rB_i(4), C1 => n37, C2 => rB_i(0)
                           , A => n38, ZN => n31);
   U71 : AOI22_X1 port map( A1 => n56, A2 => n65, B1 => D3_i(2), B2 => n57, ZN 
                           => n58);
   U72 : OAI221_X1 port map( B1 => n56, B2 => n65, C1 => n57, C2 => D3_i(2), A 
                           => n58, ZN => n51);
   U73 : OAI221_X1 port map( B1 => n53, B2 => n70, C1 => n54, C2 => n91, A => 
                           n55, ZN => n52);
   U74 : AOI22_X1 port map( A1 => n53, A2 => n70, B1 => n91, B2 => n54, ZN => 
                           n55);
   U75 : NAND3_X1 port map( A1 => n99, A2 => n100, A3 => n35, ZN => n32);
   U76 : AOI22_X1 port map( A1 => n97, A2 => rAdec_i(1), B1 => rAdec_i(3), B2 
                           => n34, ZN => n48);
   U77 : AOI22_X1 port map( A1 => n97, A2 => rA_i(1), B1 => rA_i(3), B2 => n34,
                           ZN => n63);
   U78 : AOI22_X1 port map( A1 => n96, A2 => rA_i(4), B1 => rA_i(0), B2 => n37,
                           ZN => n64);
   U79 : AOI22_X1 port map( A1 => n36, A2 => rB_i(4), B1 => rB_i(0), B2 => n37,
                           ZN => n38);
   U80 : AOI22_X1 port map( A1 => n94, A2 => rB_i(1), B1 => rB_i(3), B2 => n34,
                           ZN => n35);
   U81 : INV_X1 port map( A => D2_i(0), ZN => n37);
   U82 : INV_X1 port map( A => D2_i(3), ZN => n34);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity mem_block is

   port( X_i, LOAD_i : in std_logic_vector (31 downto 0);  W_o : out 
         std_logic_vector (31 downto 0);  S_MUX_MEM_i_BAR : in std_logic);

end mem_block;

architecture SYN_struct of mem_block is

   component mux21_3
      port( IN0, IN1 : in std_logic_vector (31 downto 0);  OUT1 : out 
            std_logic_vector (31 downto 0);  CTRL_BAR : in std_logic);
   end component;

begin
   
   MUXMEM : mux21_3 port map( IN0(31) => X_i(31), IN0(30) => X_i(30), IN0(29) 
                           => X_i(29), IN0(28) => X_i(28), IN0(27) => X_i(27), 
                           IN0(26) => X_i(26), IN0(25) => X_i(25), IN0(24) => 
                           X_i(24), IN0(23) => X_i(23), IN0(22) => X_i(22), 
                           IN0(21) => X_i(21), IN0(20) => X_i(20), IN0(19) => 
                           X_i(19), IN0(18) => X_i(18), IN0(17) => X_i(17), 
                           IN0(16) => X_i(16), IN0(15) => X_i(15), IN0(14) => 
                           X_i(14), IN0(13) => X_i(13), IN0(12) => X_i(12), 
                           IN0(11) => X_i(11), IN0(10) => X_i(10), IN0(9) => 
                           X_i(9), IN0(8) => X_i(8), IN0(7) => X_i(7), IN0(6) 
                           => X_i(6), IN0(5) => X_i(5), IN0(4) => X_i(4), 
                           IN0(3) => X_i(3), IN0(2) => X_i(2), IN0(1) => X_i(1)
                           , IN0(0) => X_i(0), IN1(31) => LOAD_i(31), IN1(30) 
                           => LOAD_i(30), IN1(29) => LOAD_i(29), IN1(28) => 
                           LOAD_i(28), IN1(27) => LOAD_i(27), IN1(26) => 
                           LOAD_i(26), IN1(25) => LOAD_i(25), IN1(24) => 
                           LOAD_i(24), IN1(23) => LOAD_i(23), IN1(22) => 
                           LOAD_i(22), IN1(21) => LOAD_i(21), IN1(20) => 
                           LOAD_i(20), IN1(19) => LOAD_i(19), IN1(18) => 
                           LOAD_i(18), IN1(17) => LOAD_i(17), IN1(16) => 
                           LOAD_i(16), IN1(15) => LOAD_i(15), IN1(14) => 
                           LOAD_i(14), IN1(13) => LOAD_i(13), IN1(12) => 
                           LOAD_i(12), IN1(11) => LOAD_i(11), IN1(10) => 
                           LOAD_i(10), IN1(9) => LOAD_i(9), IN1(8) => LOAD_i(8)
                           , IN1(7) => LOAD_i(7), IN1(6) => LOAD_i(6), IN1(5) 
                           => LOAD_i(5), IN1(4) => LOAD_i(4), IN1(3) => 
                           LOAD_i(3), IN1(2) => LOAD_i(2), IN1(1) => LOAD_i(1),
                           IN1(0) => LOAD_i(0), OUT1(31) => W_o(31), OUT1(30) 
                           => W_o(30), OUT1(29) => W_o(29), OUT1(28) => W_o(28)
                           , OUT1(27) => W_o(27), OUT1(26) => W_o(26), OUT1(25)
                           => W_o(25), OUT1(24) => W_o(24), OUT1(23) => W_o(23)
                           , OUT1(22) => W_o(22), OUT1(21) => W_o(21), OUT1(20)
                           => W_o(20), OUT1(19) => W_o(19), OUT1(18) => W_o(18)
                           , OUT1(17) => W_o(17), OUT1(16) => W_o(16), OUT1(15)
                           => W_o(15), OUT1(14) => W_o(14), OUT1(13) => W_o(13)
                           , OUT1(12) => W_o(12), OUT1(11) => W_o(11), OUT1(10)
                           => W_o(10), OUT1(9) => W_o(9), OUT1(8) => W_o(8), 
                           OUT1(7) => W_o(7), OUT1(6) => W_o(6), OUT1(5) => 
                           W_o(5), OUT1(4) => W_o(4), OUT1(3) => W_o(3), 
                           OUT1(2) => W_o(2), OUT1(1) => W_o(1), OUT1(0) => 
                           W_o(0), CTRL_BAR => S_MUX_MEM_i_BAR);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity mem_regs is

   port( W_i : in std_logic_vector (31 downto 0);  D3_i : in std_logic_vector 
         (4 downto 0);  W_o : out std_logic_vector (31 downto 0);  D3_o : out 
         std_logic_vector (4 downto 0);  clk, rst : in std_logic);

end mem_regs;

architecture SYN_Struct of mem_regs is

   component ff32_SIZE5
      port( D : in std_logic_vector (4 downto 0);  clk, rst : in std_logic;  Q 
            : out std_logic_vector (4 downto 0));
   end component;
   
   component ff32_SIZE32
      port( D : in std_logic_vector (31 downto 0);  clk, rst : in std_logic;  Q
            : out std_logic_vector (31 downto 0));
   end component;

begin
   
   W : ff32_SIZE32 port map( D(31) => W_i(31), D(30) => W_i(30), D(29) => 
                           W_i(29), D(28) => W_i(28), D(27) => W_i(27), D(26) 
                           => W_i(26), D(25) => W_i(25), D(24) => W_i(24), 
                           D(23) => W_i(23), D(22) => W_i(22), D(21) => W_i(21)
                           , D(20) => W_i(20), D(19) => W_i(19), D(18) => 
                           W_i(18), D(17) => W_i(17), D(16) => W_i(16), D(15) 
                           => W_i(15), D(14) => W_i(14), D(13) => W_i(13), 
                           D(12) => W_i(12), D(11) => W_i(11), D(10) => W_i(10)
                           , D(9) => W_i(9), D(8) => W_i(8), D(7) => W_i(7), 
                           D(6) => W_i(6), D(5) => W_i(5), D(4) => W_i(4), D(3)
                           => W_i(3), D(2) => W_i(2), D(1) => W_i(1), D(0) => 
                           W_i(0), clk => clk, rst => rst, Q(31) => W_o(31), 
                           Q(30) => W_o(30), Q(29) => W_o(29), Q(28) => W_o(28)
                           , Q(27) => W_o(27), Q(26) => W_o(26), Q(25) => 
                           W_o(25), Q(24) => W_o(24), Q(23) => W_o(23), Q(22) 
                           => W_o(22), Q(21) => W_o(21), Q(20) => W_o(20), 
                           Q(19) => W_o(19), Q(18) => W_o(18), Q(17) => W_o(17)
                           , Q(16) => W_o(16), Q(15) => W_o(15), Q(14) => 
                           W_o(14), Q(13) => W_o(13), Q(12) => W_o(12), Q(11) 
                           => W_o(11), Q(10) => W_o(10), Q(9) => W_o(9), Q(8) 
                           => W_o(8), Q(7) => W_o(7), Q(6) => W_o(6), Q(5) => 
                           W_o(5), Q(4) => W_o(4), Q(3) => W_o(3), Q(2) => 
                           W_o(2), Q(1) => W_o(1), Q(0) => W_o(0));
   D3 : ff32_SIZE5 port map( D(4) => D3_i(4), D(3) => D3_i(3), D(2) => D3_i(2),
                           D(1) => D3_i(1), D(0) => D3_i(0), clk => clk, rst =>
                           rst, Q(4) => D3_o(4), Q(3) => D3_o(3), Q(2) => 
                           D3_o(2), Q(1) => D3_o(1), Q(0) => D3_o(0));

end SYN_Struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity execute_block is

   port( IMM_i, A_i : in std_logic_vector (31 downto 0);  rB_i, rC_i : in 
         std_logic_vector (4 downto 0);  MUXED_B_i : in std_logic_vector (31 
         downto 0);  S_MUX_ALUIN_i : in std_logic;  FW_X_i, FW_W_i : in 
         std_logic_vector (31 downto 0);  S_FW_A_i, S_FW_B_i : in 
         std_logic_vector (1 downto 0);  muxed_dest : out std_logic_vector (4 
         downto 0);  muxed_B : out std_logic_vector (31 downto 0);  
         S_MUX_DEST_i : in std_logic_vector (1 downto 0);  OP : in 
         std_logic_vector (0 to 4);  ALUW_i : in std_logic_vector (12 downto 0)
         ;  DOUT : out std_logic_vector (31 downto 0);  stall_o : out std_logic
         ;  Clock, Reset : in std_logic);

end execute_block;

architecture SYN_struct of execute_block is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component mux41_MUX_SIZE32_1
      port( IN0, IN1, IN2, IN3 : in std_logic_vector (31 downto 0);  CTRL : in 
            std_logic_vector (1 downto 0);  OUT1 : out std_logic_vector (31 
            downto 0));
   end component;
   
   component mux41_MUX_SIZE32_0
      port( IN0, IN1, IN2, IN3 : in std_logic_vector (31 downto 0);  CTRL : in 
            std_logic_vector (1 downto 0);  OUT1 : out std_logic_vector (31 
            downto 0));
   end component;
   
   component mux41_MUX_SIZE5
      port( IN0, IN1, IN2, IN3 : in std_logic_vector (4 downto 0);  CTRL : in 
            std_logic_vector (1 downto 0);  OUT1 : out std_logic_vector (4 
            downto 0));
   end component;
   
   component real_alu_DATA_SIZE32
      port( IN1, IN2 : in std_logic_vector (31 downto 0);  ALUW_i : in 
            std_logic_vector (12 downto 0);  DOUT : out std_logic_vector (31 
            downto 0);  stall_o : out std_logic;  Clock, Reset : in std_logic);
   end component;
   
   component mux21_0
      port( IN0, IN1 : in std_logic_vector (31 downto 0);  CTRL : in std_logic;
            OUT1 : out std_logic_vector (31 downto 0));
   end component;
   
   signal X_Logic1_port, X_Logic0_port, muxed_B_31_port, muxed_B_30_port, 
      muxed_B_29_port, muxed_B_28_port, muxed_B_27_port, muxed_B_25_port, 
      muxed_B_24_port, muxed_B_23_port, muxed_B_22_port, muxed_B_21_port, 
      muxed_B_20_port, muxed_B_19_port, muxed_B_18_port, muxed_B_16_port, 
      muxed_B_14_port, muxed_B_13_port, muxed_B_12_port, muxed_B_11_port, 
      muxed_B_10_port, n6, muxed_B_8_port, muxed_B_7_port, muxed_B_6_port, 
      muxed_B_5_port, muxed_B_4_port, muxed_B_2_port, muxed_B_1_port, 
      FWB2alu_31_port, FWB2alu_30_port, FWB2alu_29_port, FWB2alu_28_port, 
      FWB2alu_27_port, FWB2alu_26_port, FWB2alu_25_port, FWB2alu_24_port, 
      FWB2alu_23_port, FWB2alu_22_port, FWB2alu_21_port, FWB2alu_20_port, 
      FWB2alu_19_port, FWB2alu_18_port, FWB2alu_17_port, FWB2alu_16_port, 
      FWB2alu_15_port, FWB2alu_14_port, FWB2alu_13_port, FWB2alu_12_port, 
      FWB2alu_11_port, FWB2alu_10_port, FWB2alu_9_port, FWB2alu_8_port, 
      FWB2alu_7_port, FWB2alu_6_port, FWB2alu_5_port, FWB2alu_4_port, 
      FWB2alu_3_port, FWB2alu_2_port, FWB2alu_1_port, FWB2alu_0_port, 
      FWA2alu_31_port, FWA2alu_30_port, FWA2alu_29_port, FWA2alu_28_port, 
      FWA2alu_27_port, FWA2alu_26_port, FWA2alu_25_port, FWA2alu_24_port, 
      FWA2alu_23_port, FWA2alu_22_port, FWA2alu_21_port, FWA2alu_20_port, 
      FWA2alu_19_port, FWA2alu_18_port, FWA2alu_17_port, FWA2alu_16_port, 
      FWA2alu_15_port, FWA2alu_14_port, FWA2alu_13_port, FWA2alu_12_port, 
      FWA2alu_11_port, FWA2alu_10_port, FWA2alu_9_port, FWA2alu_8_port, 
      FWA2alu_7_port, FWA2alu_6_port, FWA2alu_5_port, FWA2alu_4_port, 
      FWA2alu_3_port, FWA2alu_2_port, FWA2alu_1_port, FWA2alu_0_port, n1, 
      muxed_B_15_port, muxed_B_17_port, muxed_B_26_port, muxed_B_0_port, 
      muxed_B_3_port, muxed_B_9_port : std_logic;

begin
   muxed_B <= ( muxed_B_31_port, muxed_B_30_port, muxed_B_29_port, 
      muxed_B_28_port, muxed_B_27_port, muxed_B_26_port, muxed_B_25_port, 
      muxed_B_24_port, muxed_B_23_port, muxed_B_22_port, muxed_B_21_port, 
      muxed_B_20_port, muxed_B_19_port, muxed_B_18_port, muxed_B_17_port, 
      muxed_B_16_port, muxed_B_15_port, muxed_B_14_port, muxed_B_13_port, 
      muxed_B_12_port, muxed_B_11_port, muxed_B_10_port, muxed_B_9_port, 
      muxed_B_8_port, muxed_B_7_port, muxed_B_6_port, muxed_B_5_port, 
      muxed_B_4_port, muxed_B_3_port, muxed_B_2_port, muxed_B_1_port, 
      muxed_B_0_port );
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   n1 <= '0';
   ALUIN_MUX : mux21_0 port map( IN0(31) => muxed_B_31_port, IN0(30) => 
                           muxed_B_30_port, IN0(29) => muxed_B_29_port, IN0(28)
                           => muxed_B_28_port, IN0(27) => muxed_B_27_port, 
                           IN0(26) => muxed_B_26_port, IN0(25) => 
                           muxed_B_25_port, IN0(24) => muxed_B_24_port, IN0(23)
                           => muxed_B_23_port, IN0(22) => muxed_B_22_port, 
                           IN0(21) => muxed_B_21_port, IN0(20) => 
                           muxed_B_20_port, IN0(19) => muxed_B_19_port, IN0(18)
                           => muxed_B_18_port, IN0(17) => muxed_B_17_port, 
                           IN0(16) => muxed_B_16_port, IN0(15) => 
                           muxed_B_15_port, IN0(14) => muxed_B_14_port, IN0(13)
                           => muxed_B_13_port, IN0(12) => muxed_B_12_port, 
                           IN0(11) => muxed_B_11_port, IN0(10) => 
                           muxed_B_10_port, IN0(9) => n6, IN0(8) => 
                           muxed_B_8_port, IN0(7) => muxed_B_7_port, IN0(6) => 
                           muxed_B_6_port, IN0(5) => muxed_B_5_port, IN0(4) => 
                           muxed_B_4_port, IN0(3) => muxed_B_3_port, IN0(2) => 
                           muxed_B_2_port, IN0(1) => muxed_B_1_port, IN0(0) => 
                           muxed_B_0_port, IN1(31) => IMM_i(31), IN1(30) => 
                           IMM_i(30), IN1(29) => IMM_i(29), IN1(28) => 
                           IMM_i(28), IN1(27) => IMM_i(27), IN1(26) => 
                           IMM_i(26), IN1(25) => IMM_i(25), IN1(24) => 
                           IMM_i(24), IN1(23) => IMM_i(23), IN1(22) => 
                           IMM_i(22), IN1(21) => IMM_i(21), IN1(20) => 
                           IMM_i(20), IN1(19) => IMM_i(19), IN1(18) => 
                           IMM_i(18), IN1(17) => IMM_i(17), IN1(16) => 
                           IMM_i(16), IN1(15) => IMM_i(15), IN1(14) => 
                           IMM_i(14), IN1(13) => IMM_i(13), IN1(12) => 
                           IMM_i(12), IN1(11) => IMM_i(11), IN1(10) => 
                           IMM_i(10), IN1(9) => IMM_i(9), IN1(8) => IMM_i(8), 
                           IN1(7) => IMM_i(7), IN1(6) => IMM_i(6), IN1(5) => 
                           IMM_i(5), IN1(4) => IMM_i(4), IN1(3) => IMM_i(3), 
                           IN1(2) => IMM_i(2), IN1(1) => IMM_i(1), IN1(0) => 
                           IMM_i(0), CTRL => S_MUX_ALUIN_i, OUT1(31) => 
                           FWB2alu_31_port, OUT1(30) => FWB2alu_30_port, 
                           OUT1(29) => FWB2alu_29_port, OUT1(28) => 
                           FWB2alu_28_port, OUT1(27) => FWB2alu_27_port, 
                           OUT1(26) => FWB2alu_26_port, OUT1(25) => 
                           FWB2alu_25_port, OUT1(24) => FWB2alu_24_port, 
                           OUT1(23) => FWB2alu_23_port, OUT1(22) => 
                           FWB2alu_22_port, OUT1(21) => FWB2alu_21_port, 
                           OUT1(20) => FWB2alu_20_port, OUT1(19) => 
                           FWB2alu_19_port, OUT1(18) => FWB2alu_18_port, 
                           OUT1(17) => FWB2alu_17_port, OUT1(16) => 
                           FWB2alu_16_port, OUT1(15) => FWB2alu_15_port, 
                           OUT1(14) => FWB2alu_14_port, OUT1(13) => 
                           FWB2alu_13_port, OUT1(12) => FWB2alu_12_port, 
                           OUT1(11) => FWB2alu_11_port, OUT1(10) => 
                           FWB2alu_10_port, OUT1(9) => FWB2alu_9_port, OUT1(8) 
                           => FWB2alu_8_port, OUT1(7) => FWB2alu_7_port, 
                           OUT1(6) => FWB2alu_6_port, OUT1(5) => FWB2alu_5_port
                           , OUT1(4) => FWB2alu_4_port, OUT1(3) => 
                           FWB2alu_3_port, OUT1(2) => FWB2alu_2_port, OUT1(1) 
                           => FWB2alu_1_port, OUT1(0) => FWB2alu_0_port);
   ALU : real_alu_DATA_SIZE32 port map( IN1(31) => FWA2alu_31_port, IN1(30) => 
                           FWA2alu_30_port, IN1(29) => FWA2alu_29_port, IN1(28)
                           => FWA2alu_28_port, IN1(27) => FWA2alu_27_port, 
                           IN1(26) => FWA2alu_26_port, IN1(25) => 
                           FWA2alu_25_port, IN1(24) => FWA2alu_24_port, IN1(23)
                           => FWA2alu_23_port, IN1(22) => FWA2alu_22_port, 
                           IN1(21) => FWA2alu_21_port, IN1(20) => 
                           FWA2alu_20_port, IN1(19) => FWA2alu_19_port, IN1(18)
                           => FWA2alu_18_port, IN1(17) => FWA2alu_17_port, 
                           IN1(16) => FWA2alu_16_port, IN1(15) => 
                           FWA2alu_15_port, IN1(14) => FWA2alu_14_port, IN1(13)
                           => FWA2alu_13_port, IN1(12) => FWA2alu_12_port, 
                           IN1(11) => FWA2alu_11_port, IN1(10) => 
                           FWA2alu_10_port, IN1(9) => FWA2alu_9_port, IN1(8) =>
                           FWA2alu_8_port, IN1(7) => FWA2alu_7_port, IN1(6) => 
                           FWA2alu_6_port, IN1(5) => FWA2alu_5_port, IN1(4) => 
                           FWA2alu_4_port, IN1(3) => FWA2alu_3_port, IN1(2) => 
                           FWA2alu_2_port, IN1(1) => FWA2alu_1_port, IN1(0) => 
                           FWA2alu_0_port, IN2(31) => FWB2alu_31_port, IN2(30) 
                           => FWB2alu_30_port, IN2(29) => FWB2alu_29_port, 
                           IN2(28) => FWB2alu_28_port, IN2(27) => 
                           FWB2alu_27_port, IN2(26) => FWB2alu_26_port, IN2(25)
                           => FWB2alu_25_port, IN2(24) => FWB2alu_24_port, 
                           IN2(23) => FWB2alu_23_port, IN2(22) => 
                           FWB2alu_22_port, IN2(21) => FWB2alu_21_port, IN2(20)
                           => FWB2alu_20_port, IN2(19) => FWB2alu_19_port, 
                           IN2(18) => FWB2alu_18_port, IN2(17) => 
                           FWB2alu_17_port, IN2(16) => FWB2alu_16_port, IN2(15)
                           => FWB2alu_15_port, IN2(14) => FWB2alu_14_port, 
                           IN2(13) => FWB2alu_13_port, IN2(12) => 
                           FWB2alu_12_port, IN2(11) => FWB2alu_11_port, IN2(10)
                           => FWB2alu_10_port, IN2(9) => FWB2alu_9_port, IN2(8)
                           => FWB2alu_8_port, IN2(7) => FWB2alu_7_port, IN2(6) 
                           => FWB2alu_6_port, IN2(5) => FWB2alu_5_port, IN2(4) 
                           => FWB2alu_4_port, IN2(3) => FWB2alu_3_port, IN2(2) 
                           => FWB2alu_2_port, IN2(1) => FWB2alu_1_port, IN2(0) 
                           => FWB2alu_0_port, ALUW_i(12) => ALUW_i(12), 
                           ALUW_i(11) => ALUW_i(11), ALUW_i(10) => ALUW_i(10), 
                           ALUW_i(9) => ALUW_i(9), ALUW_i(8) => ALUW_i(8), 
                           ALUW_i(7) => ALUW_i(7), ALUW_i(6) => ALUW_i(6), 
                           ALUW_i(5) => ALUW_i(5), ALUW_i(4) => ALUW_i(4), 
                           ALUW_i(3) => ALUW_i(3), ALUW_i(2) => ALUW_i(2), 
                           ALUW_i(1) => ALUW_i(1), ALUW_i(0) => ALUW_i(0), 
                           DOUT(31) => DOUT(31), DOUT(30) => DOUT(30), DOUT(29)
                           => DOUT(29), DOUT(28) => DOUT(28), DOUT(27) => 
                           DOUT(27), DOUT(26) => DOUT(26), DOUT(25) => DOUT(25)
                           , DOUT(24) => DOUT(24), DOUT(23) => DOUT(23), 
                           DOUT(22) => DOUT(22), DOUT(21) => DOUT(21), DOUT(20)
                           => DOUT(20), DOUT(19) => DOUT(19), DOUT(18) => 
                           DOUT(18), DOUT(17) => DOUT(17), DOUT(16) => DOUT(16)
                           , DOUT(15) => DOUT(15), DOUT(14) => DOUT(14), 
                           DOUT(13) => DOUT(13), DOUT(12) => DOUT(12), DOUT(11)
                           => DOUT(11), DOUT(10) => DOUT(10), DOUT(9) => 
                           DOUT(9), DOUT(8) => DOUT(8), DOUT(7) => DOUT(7), 
                           DOUT(6) => DOUT(6), DOUT(5) => DOUT(5), DOUT(4) => 
                           DOUT(4), DOUT(3) => DOUT(3), DOUT(2) => DOUT(2), 
                           DOUT(1) => DOUT(1), DOUT(0) => DOUT(0), stall_o => 
                           stall_o, Clock => Clock, Reset => Reset);
   MUXDEST : mux41_MUX_SIZE5 port map( IN0(4) => X_Logic0_port, IN0(3) => 
                           X_Logic0_port, IN0(2) => X_Logic0_port, IN0(1) => 
                           X_Logic0_port, IN0(0) => X_Logic0_port, IN1(4) => 
                           rC_i(4), IN1(3) => rC_i(3), IN1(2) => rC_i(2), 
                           IN1(1) => rC_i(1), IN1(0) => rC_i(0), IN2(4) => 
                           rB_i(4), IN2(3) => rB_i(3), IN2(2) => rB_i(2), 
                           IN2(1) => rB_i(1), IN2(0) => rB_i(0), IN3(4) => 
                           X_Logic1_port, IN3(3) => X_Logic1_port, IN3(2) => 
                           X_Logic1_port, IN3(1) => X_Logic1_port, IN3(0) => 
                           X_Logic1_port, CTRL(1) => S_MUX_DEST_i(1), CTRL(0) 
                           => S_MUX_DEST_i(0), OUT1(4) => muxed_dest(4), 
                           OUT1(3) => muxed_dest(3), OUT1(2) => muxed_dest(2), 
                           OUT1(1) => muxed_dest(1), OUT1(0) => muxed_dest(0));
   MUX_FWA : mux41_MUX_SIZE32_0 port map( IN0(31) => A_i(31), IN0(30) => 
                           A_i(30), IN0(29) => A_i(29), IN0(28) => A_i(28), 
                           IN0(27) => A_i(27), IN0(26) => A_i(26), IN0(25) => 
                           A_i(25), IN0(24) => A_i(24), IN0(23) => A_i(23), 
                           IN0(22) => A_i(22), IN0(21) => A_i(21), IN0(20) => 
                           A_i(20), IN0(19) => A_i(19), IN0(18) => A_i(18), 
                           IN0(17) => A_i(17), IN0(16) => A_i(16), IN0(15) => 
                           A_i(15), IN0(14) => A_i(14), IN0(13) => A_i(13), 
                           IN0(12) => A_i(12), IN0(11) => A_i(11), IN0(10) => 
                           A_i(10), IN0(9) => A_i(9), IN0(8) => A_i(8), IN0(7) 
                           => A_i(7), IN0(6) => A_i(6), IN0(5) => A_i(5), 
                           IN0(4) => A_i(4), IN0(3) => A_i(3), IN0(2) => A_i(2)
                           , IN0(1) => A_i(1), IN0(0) => A_i(0), IN1(31) => 
                           FW_X_i(31), IN1(30) => FW_X_i(30), IN1(29) => 
                           FW_X_i(29), IN1(28) => FW_X_i(28), IN1(27) => 
                           FW_X_i(27), IN1(26) => FW_X_i(26), IN1(25) => 
                           FW_X_i(25), IN1(24) => FW_X_i(24), IN1(23) => 
                           FW_X_i(23), IN1(22) => FW_X_i(22), IN1(21) => 
                           FW_X_i(21), IN1(20) => FW_X_i(20), IN1(19) => 
                           FW_X_i(19), IN1(18) => FW_X_i(18), IN1(17) => 
                           FW_X_i(17), IN1(16) => FW_X_i(16), IN1(15) => 
                           FW_X_i(15), IN1(14) => FW_X_i(14), IN1(13) => 
                           FW_X_i(13), IN1(12) => FW_X_i(12), IN1(11) => 
                           FW_X_i(11), IN1(10) => FW_X_i(10), IN1(9) => 
                           FW_X_i(9), IN1(8) => FW_X_i(8), IN1(7) => FW_X_i(7),
                           IN1(6) => FW_X_i(6), IN1(5) => FW_X_i(5), IN1(4) => 
                           FW_X_i(4), IN1(3) => FW_X_i(3), IN1(2) => FW_X_i(2),
                           IN1(1) => FW_X_i(1), IN1(0) => FW_X_i(0), IN2(31) =>
                           FW_W_i(31), IN2(30) => FW_W_i(30), IN2(29) => 
                           FW_W_i(29), IN2(28) => FW_W_i(28), IN2(27) => 
                           FW_W_i(27), IN2(26) => FW_W_i(26), IN2(25) => 
                           FW_W_i(25), IN2(24) => FW_W_i(24), IN2(23) => 
                           FW_W_i(23), IN2(22) => FW_W_i(22), IN2(21) => 
                           FW_W_i(21), IN2(20) => FW_W_i(20), IN2(19) => 
                           FW_W_i(19), IN2(18) => FW_W_i(18), IN2(17) => 
                           FW_W_i(17), IN2(16) => FW_W_i(16), IN2(15) => 
                           FW_W_i(15), IN2(14) => FW_W_i(14), IN2(13) => 
                           FW_W_i(13), IN2(12) => FW_W_i(12), IN2(11) => 
                           FW_W_i(11), IN2(10) => FW_W_i(10), IN2(9) => 
                           FW_W_i(9), IN2(8) => FW_W_i(8), IN2(7) => FW_W_i(7),
                           IN2(6) => FW_W_i(6), IN2(5) => FW_W_i(5), IN2(4) => 
                           FW_W_i(4), IN2(3) => FW_W_i(3), IN2(2) => FW_W_i(2),
                           IN2(1) => FW_W_i(1), IN2(0) => FW_W_i(0), IN3(31) =>
                           n1, IN3(30) => n1, IN3(29) => n1, IN3(28) => n1, 
                           IN3(27) => n1, IN3(26) => n1, IN3(25) => n1, IN3(24)
                           => n1, IN3(23) => n1, IN3(22) => n1, IN3(21) => n1, 
                           IN3(20) => n1, IN3(19) => n1, IN3(18) => n1, IN3(17)
                           => n1, IN3(16) => n1, IN3(15) => n1, IN3(14) => n1, 
                           IN3(13) => n1, IN3(12) => n1, IN3(11) => n1, IN3(10)
                           => n1, IN3(9) => n1, IN3(8) => n1, IN3(7) => n1, 
                           IN3(6) => n1, IN3(5) => n1, IN3(4) => n1, IN3(3) => 
                           n1, IN3(2) => n1, IN3(1) => n1, IN3(0) => n1, 
                           CTRL(1) => S_FW_A_i(1), CTRL(0) => S_FW_A_i(0), 
                           OUT1(31) => FWA2alu_31_port, OUT1(30) => 
                           FWA2alu_30_port, OUT1(29) => FWA2alu_29_port, 
                           OUT1(28) => FWA2alu_28_port, OUT1(27) => 
                           FWA2alu_27_port, OUT1(26) => FWA2alu_26_port, 
                           OUT1(25) => FWA2alu_25_port, OUT1(24) => 
                           FWA2alu_24_port, OUT1(23) => FWA2alu_23_port, 
                           OUT1(22) => FWA2alu_22_port, OUT1(21) => 
                           FWA2alu_21_port, OUT1(20) => FWA2alu_20_port, 
                           OUT1(19) => FWA2alu_19_port, OUT1(18) => 
                           FWA2alu_18_port, OUT1(17) => FWA2alu_17_port, 
                           OUT1(16) => FWA2alu_16_port, OUT1(15) => 
                           FWA2alu_15_port, OUT1(14) => FWA2alu_14_port, 
                           OUT1(13) => FWA2alu_13_port, OUT1(12) => 
                           FWA2alu_12_port, OUT1(11) => FWA2alu_11_port, 
                           OUT1(10) => FWA2alu_10_port, OUT1(9) => 
                           FWA2alu_9_port, OUT1(8) => FWA2alu_8_port, OUT1(7) 
                           => FWA2alu_7_port, OUT1(6) => FWA2alu_6_port, 
                           OUT1(5) => FWA2alu_5_port, OUT1(4) => FWA2alu_4_port
                           , OUT1(3) => FWA2alu_3_port, OUT1(2) => 
                           FWA2alu_2_port, OUT1(1) => FWA2alu_1_port, OUT1(0) 
                           => FWA2alu_0_port);
   MUX_FWB : mux41_MUX_SIZE32_1 port map( IN0(31) => MUXED_B_i(31), IN0(30) => 
                           MUXED_B_i(30), IN0(29) => MUXED_B_i(29), IN0(28) => 
                           MUXED_B_i(28), IN0(27) => MUXED_B_i(27), IN0(26) => 
                           MUXED_B_i(26), IN0(25) => MUXED_B_i(25), IN0(24) => 
                           MUXED_B_i(24), IN0(23) => MUXED_B_i(23), IN0(22) => 
                           MUXED_B_i(22), IN0(21) => MUXED_B_i(21), IN0(20) => 
                           MUXED_B_i(20), IN0(19) => MUXED_B_i(19), IN0(18) => 
                           MUXED_B_i(18), IN0(17) => MUXED_B_i(17), IN0(16) => 
                           MUXED_B_i(16), IN0(15) => MUXED_B_i(15), IN0(14) => 
                           MUXED_B_i(14), IN0(13) => MUXED_B_i(13), IN0(12) => 
                           MUXED_B_i(12), IN0(11) => MUXED_B_i(11), IN0(10) => 
                           MUXED_B_i(10), IN0(9) => MUXED_B_i(9), IN0(8) => 
                           MUXED_B_i(8), IN0(7) => MUXED_B_i(7), IN0(6) => 
                           MUXED_B_i(6), IN0(5) => MUXED_B_i(5), IN0(4) => 
                           MUXED_B_i(4), IN0(3) => MUXED_B_i(3), IN0(2) => 
                           MUXED_B_i(2), IN0(1) => MUXED_B_i(1), IN0(0) => 
                           MUXED_B_i(0), IN1(31) => FW_X_i(31), IN1(30) => 
                           FW_X_i(30), IN1(29) => FW_X_i(29), IN1(28) => 
                           FW_X_i(28), IN1(27) => FW_X_i(27), IN1(26) => 
                           FW_X_i(26), IN1(25) => FW_X_i(25), IN1(24) => 
                           FW_X_i(24), IN1(23) => FW_X_i(23), IN1(22) => 
                           FW_X_i(22), IN1(21) => FW_X_i(21), IN1(20) => 
                           FW_X_i(20), IN1(19) => FW_X_i(19), IN1(18) => 
                           FW_X_i(18), IN1(17) => FW_X_i(17), IN1(16) => 
                           FW_X_i(16), IN1(15) => FW_X_i(15), IN1(14) => 
                           FW_X_i(14), IN1(13) => FW_X_i(13), IN1(12) => 
                           FW_X_i(12), IN1(11) => FW_X_i(11), IN1(10) => 
                           FW_X_i(10), IN1(9) => FW_X_i(9), IN1(8) => FW_X_i(8)
                           , IN1(7) => FW_X_i(7), IN1(6) => FW_X_i(6), IN1(5) 
                           => FW_X_i(5), IN1(4) => FW_X_i(4), IN1(3) => 
                           FW_X_i(3), IN1(2) => FW_X_i(2), IN1(1) => FW_X_i(1),
                           IN1(0) => FW_X_i(0), IN2(31) => FW_W_i(31), IN2(30) 
                           => FW_W_i(30), IN2(29) => FW_W_i(29), IN2(28) => 
                           FW_W_i(28), IN2(27) => FW_W_i(27), IN2(26) => 
                           FW_W_i(26), IN2(25) => FW_W_i(25), IN2(24) => 
                           FW_W_i(24), IN2(23) => FW_W_i(23), IN2(22) => 
                           FW_W_i(22), IN2(21) => FW_W_i(21), IN2(20) => 
                           FW_W_i(20), IN2(19) => FW_W_i(19), IN2(18) => 
                           FW_W_i(18), IN2(17) => FW_W_i(17), IN2(16) => 
                           FW_W_i(16), IN2(15) => FW_W_i(15), IN2(14) => 
                           FW_W_i(14), IN2(13) => FW_W_i(13), IN2(12) => 
                           FW_W_i(12), IN2(11) => FW_W_i(11), IN2(10) => 
                           FW_W_i(10), IN2(9) => FW_W_i(9), IN2(8) => FW_W_i(8)
                           , IN2(7) => FW_W_i(7), IN2(6) => FW_W_i(6), IN2(5) 
                           => FW_W_i(5), IN2(4) => FW_W_i(4), IN2(3) => 
                           FW_W_i(3), IN2(2) => FW_W_i(2), IN2(1) => FW_W_i(1),
                           IN2(0) => FW_W_i(0), IN3(31) => n1, IN3(30) => n1, 
                           IN3(29) => n1, IN3(28) => n1, IN3(27) => n1, IN3(26)
                           => n1, IN3(25) => n1, IN3(24) => n1, IN3(23) => n1, 
                           IN3(22) => n1, IN3(21) => n1, IN3(20) => n1, IN3(19)
                           => n1, IN3(18) => n1, IN3(17) => n1, IN3(16) => n1, 
                           IN3(15) => n1, IN3(14) => n1, IN3(13) => n1, IN3(12)
                           => n1, IN3(11) => n1, IN3(10) => n1, IN3(9) => n1, 
                           IN3(8) => n1, IN3(7) => n1, IN3(6) => n1, IN3(5) => 
                           n1, IN3(4) => n1, IN3(3) => n1, IN3(2) => n1, IN3(1)
                           => n1, IN3(0) => n1, CTRL(1) => S_FW_B_i(1), CTRL(0)
                           => S_FW_B_i(0), OUT1(31) => muxed_B_31_port, 
                           OUT1(30) => muxed_B_30_port, OUT1(29) => 
                           muxed_B_29_port, OUT1(28) => muxed_B_28_port, 
                           OUT1(27) => muxed_B_27_port, OUT1(26) => 
                           muxed_B_26_port, OUT1(25) => muxed_B_25_port, 
                           OUT1(24) => muxed_B_24_port, OUT1(23) => 
                           muxed_B_23_port, OUT1(22) => muxed_B_22_port, 
                           OUT1(21) => muxed_B_21_port, OUT1(20) => 
                           muxed_B_20_port, OUT1(19) => muxed_B_19_port, 
                           OUT1(18) => muxed_B_18_port, OUT1(17) => 
                           muxed_B_17_port, OUT1(16) => muxed_B_16_port, 
                           OUT1(15) => muxed_B_15_port, OUT1(14) => 
                           muxed_B_14_port, OUT1(13) => muxed_B_13_port, 
                           OUT1(12) => muxed_B_12_port, OUT1(11) => 
                           muxed_B_11_port, OUT1(10) => muxed_B_10_port, 
                           OUT1(9) => n6, OUT1(8) => muxed_B_8_port, OUT1(7) =>
                           muxed_B_7_port, OUT1(6) => muxed_B_6_port, OUT1(5) 
                           => muxed_B_5_port, OUT1(4) => muxed_B_4_port, 
                           OUT1(3) => muxed_B_3_port, OUT1(2) => muxed_B_2_port
                           , OUT1(1) => muxed_B_1_port, OUT1(0) => 
                           muxed_B_0_port);
   U5 : CLKBUF_X1 port map( A => n6, Z => muxed_B_9_port);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity execute_regs is

   port( X_i, S_i : in std_logic_vector (31 downto 0);  D2_i : in 
         std_logic_vector (4 downto 0);  X_o, S_o : out std_logic_vector (31 
         downto 0);  D2_o : out std_logic_vector (4 downto 0);  stall_i, clk, 
         rst : in std_logic);

end execute_regs;

architecture SYN_struct of execute_regs is

   component ff32_en_SIZE5_1
      port( D : in std_logic_vector (4 downto 0);  en, clk, rst : in std_logic;
            Q : out std_logic_vector (4 downto 0));
   end component;
   
   component ff32_en_SIZE32_2
      port( D : in std_logic_vector (31 downto 0);  en, clk, rst : in std_logic
            ;  Q : out std_logic_vector (31 downto 0));
   end component;
   
   component ff32_en_SIZE32_3
      port( D : in std_logic_vector (31 downto 0);  en, clk, rst : in std_logic
            ;  Q : out std_logic_vector (31 downto 0));
   end component;
   
   signal n3 : std_logic;

begin
   
   X : ff32_en_SIZE32_3 port map( D(31) => X_i(31), D(30) => X_i(30), D(29) => 
                           X_i(29), D(28) => X_i(28), D(27) => X_i(27), D(26) 
                           => X_i(26), D(25) => X_i(25), D(24) => X_i(24), 
                           D(23) => X_i(23), D(22) => X_i(22), D(21) => X_i(21)
                           , D(20) => X_i(20), D(19) => X_i(19), D(18) => 
                           X_i(18), D(17) => X_i(17), D(16) => X_i(16), D(15) 
                           => X_i(15), D(14) => X_i(14), D(13) => X_i(13), 
                           D(12) => X_i(12), D(11) => X_i(11), D(10) => X_i(10)
                           , D(9) => X_i(9), D(8) => X_i(8), D(7) => X_i(7), 
                           D(6) => X_i(6), D(5) => X_i(5), D(4) => X_i(4), D(3)
                           => X_i(3), D(2) => X_i(2), D(1) => X_i(1), D(0) => 
                           X_i(0), en => n3, clk => clk, rst => rst, Q(31) => 
                           X_o(31), Q(30) => X_o(30), Q(29) => X_o(29), Q(28) 
                           => X_o(28), Q(27) => X_o(27), Q(26) => X_o(26), 
                           Q(25) => X_o(25), Q(24) => X_o(24), Q(23) => X_o(23)
                           , Q(22) => X_o(22), Q(21) => X_o(21), Q(20) => 
                           X_o(20), Q(19) => X_o(19), Q(18) => X_o(18), Q(17) 
                           => X_o(17), Q(16) => X_o(16), Q(15) => X_o(15), 
                           Q(14) => X_o(14), Q(13) => X_o(13), Q(12) => X_o(12)
                           , Q(11) => X_o(11), Q(10) => X_o(10), Q(9) => X_o(9)
                           , Q(8) => X_o(8), Q(7) => X_o(7), Q(6) => X_o(6), 
                           Q(5) => X_o(5), Q(4) => X_o(4), Q(3) => X_o(3), Q(2)
                           => X_o(2), Q(1) => X_o(1), Q(0) => X_o(0));
   S : ff32_en_SIZE32_2 port map( D(31) => S_i(31), D(30) => S_i(30), D(29) => 
                           S_i(29), D(28) => S_i(28), D(27) => S_i(27), D(26) 
                           => S_i(26), D(25) => S_i(25), D(24) => S_i(24), 
                           D(23) => S_i(23), D(22) => S_i(22), D(21) => S_i(21)
                           , D(20) => S_i(20), D(19) => S_i(19), D(18) => 
                           S_i(18), D(17) => S_i(17), D(16) => S_i(16), D(15) 
                           => S_i(15), D(14) => S_i(14), D(13) => S_i(13), 
                           D(12) => S_i(12), D(11) => S_i(11), D(10) => S_i(10)
                           , D(9) => S_i(9), D(8) => S_i(8), D(7) => S_i(7), 
                           D(6) => S_i(6), D(5) => S_i(5), D(4) => S_i(4), D(3)
                           => S_i(3), D(2) => S_i(2), D(1) => S_i(1), D(0) => 
                           S_i(0), en => n3, clk => clk, rst => rst, Q(31) => 
                           S_o(31), Q(30) => S_o(30), Q(29) => S_o(29), Q(28) 
                           => S_o(28), Q(27) => S_o(27), Q(26) => S_o(26), 
                           Q(25) => S_o(25), Q(24) => S_o(24), Q(23) => S_o(23)
                           , Q(22) => S_o(22), Q(21) => S_o(21), Q(20) => 
                           S_o(20), Q(19) => S_o(19), Q(18) => S_o(18), Q(17) 
                           => S_o(17), Q(16) => S_o(16), Q(15) => S_o(15), 
                           Q(14) => S_o(14), Q(13) => S_o(13), Q(12) => S_o(12)
                           , Q(11) => S_o(11), Q(10) => S_o(10), Q(9) => S_o(9)
                           , Q(8) => S_o(8), Q(7) => S_o(7), Q(6) => S_o(6), 
                           Q(5) => S_o(5), Q(4) => S_o(4), Q(3) => S_o(3), Q(2)
                           => S_o(2), Q(1) => S_o(1), Q(0) => S_o(0));
   D2 : ff32_en_SIZE5_1 port map( D(4) => D2_i(4), D(3) => D2_i(3), D(2) => 
                           D2_i(2), D(1) => D2_i(1), D(0) => D2_i(0), en => n3,
                           clk => clk, rst => rst, Q(4) => D2_o(4), Q(3) => 
                           D2_o(3), Q(2) => D2_o(2), Q(1) => D2_o(1), Q(0) => 
                           D2_o(0));
   n3 <= '1';

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity decode_regs is

   port( A_i, B_i : in std_logic_vector (31 downto 0);  rA_i, rB_i, rC_i : in 
         std_logic_vector (4 downto 0);  IMM_i : in std_logic_vector (31 downto
         0);  ALUW_i : in std_logic_vector (12 downto 0);  A_o, B_o : out 
         std_logic_vector (31 downto 0);  rA_o, rB_o, rC_o : out 
         std_logic_vector (4 downto 0);  IMM_o : out std_logic_vector (31 
         downto 0);  ALUW_o : out std_logic_vector (12 downto 0);  stall_i, clk
         , rst : in std_logic);

end decode_regs;

architecture SYN_struct of decode_regs is

   component INV_X8
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component ff32_en_SIZE13
      port( D : in std_logic_vector (12 downto 0);  en, clk, rst : in std_logic
            ;  Q : out std_logic_vector (12 downto 0));
   end component;
   
   component ff32_en_SIZE32_4
      port( D : in std_logic_vector (31 downto 0);  en, clk, rst : in std_logic
            ;  Q : out std_logic_vector (31 downto 0));
   end component;
   
   component ff32_en_SIZE5_2
      port( D : in std_logic_vector (4 downto 0);  en, clk, rst : in std_logic;
            Q : out std_logic_vector (4 downto 0));
   end component;
   
   component ff32_en_SIZE5_3
      port( D : in std_logic_vector (4 downto 0);  en, clk, rst : in std_logic;
            Q : out std_logic_vector (4 downto 0));
   end component;
   
   component ff32_en_SIZE5_0
      port( D : in std_logic_vector (4 downto 0);  en, clk, rst : in std_logic;
            Q : out std_logic_vector (4 downto 0));
   end component;
   
   component ff32_en_SIZE32_5
      port( D : in std_logic_vector (31 downto 0);  en, clk, rst : in std_logic
            ;  Q : out std_logic_vector (31 downto 0));
   end component;
   
   component ff32_en_SIZE32_0
      port( D : in std_logic_vector (31 downto 0);  en, clk, rst : in std_logic
            ;  Q : out std_logic_vector (31 downto 0));
   end component;
   
   signal enable : std_logic;

begin
   
   A : ff32_en_SIZE32_0 port map( D(31) => A_i(31), D(30) => A_i(30), D(29) => 
                           A_i(29), D(28) => A_i(28), D(27) => A_i(27), D(26) 
                           => A_i(26), D(25) => A_i(25), D(24) => A_i(24), 
                           D(23) => A_i(23), D(22) => A_i(22), D(21) => A_i(21)
                           , D(20) => A_i(20), D(19) => A_i(19), D(18) => 
                           A_i(18), D(17) => A_i(17), D(16) => A_i(16), D(15) 
                           => A_i(15), D(14) => A_i(14), D(13) => A_i(13), 
                           D(12) => A_i(12), D(11) => A_i(11), D(10) => A_i(10)
                           , D(9) => A_i(9), D(8) => A_i(8), D(7) => A_i(7), 
                           D(6) => A_i(6), D(5) => A_i(5), D(4) => A_i(4), D(3)
                           => A_i(3), D(2) => A_i(2), D(1) => A_i(1), D(0) => 
                           A_i(0), en => enable, clk => clk, rst => rst, Q(31) 
                           => A_o(31), Q(30) => A_o(30), Q(29) => A_o(29), 
                           Q(28) => A_o(28), Q(27) => A_o(27), Q(26) => A_o(26)
                           , Q(25) => A_o(25), Q(24) => A_o(24), Q(23) => 
                           A_o(23), Q(22) => A_o(22), Q(21) => A_o(21), Q(20) 
                           => A_o(20), Q(19) => A_o(19), Q(18) => A_o(18), 
                           Q(17) => A_o(17), Q(16) => A_o(16), Q(15) => A_o(15)
                           , Q(14) => A_o(14), Q(13) => A_o(13), Q(12) => 
                           A_o(12), Q(11) => A_o(11), Q(10) => A_o(10), Q(9) =>
                           A_o(9), Q(8) => A_o(8), Q(7) => A_o(7), Q(6) => 
                           A_o(6), Q(5) => A_o(5), Q(4) => A_o(4), Q(3) => 
                           A_o(3), Q(2) => A_o(2), Q(1) => A_o(1), Q(0) => 
                           A_o(0));
   B : ff32_en_SIZE32_5 port map( D(31) => B_i(31), D(30) => B_i(30), D(29) => 
                           B_i(29), D(28) => B_i(28), D(27) => B_i(27), D(26) 
                           => B_i(26), D(25) => B_i(25), D(24) => B_i(24), 
                           D(23) => B_i(23), D(22) => B_i(22), D(21) => B_i(21)
                           , D(20) => B_i(20), D(19) => B_i(19), D(18) => 
                           B_i(18), D(17) => B_i(17), D(16) => B_i(16), D(15) 
                           => B_i(15), D(14) => B_i(14), D(13) => B_i(13), 
                           D(12) => B_i(12), D(11) => B_i(11), D(10) => B_i(10)
                           , D(9) => B_i(9), D(8) => B_i(8), D(7) => B_i(7), 
                           D(6) => B_i(6), D(5) => B_i(5), D(4) => B_i(4), D(3)
                           => B_i(3), D(2) => B_i(2), D(1) => B_i(1), D(0) => 
                           B_i(0), en => enable, clk => clk, rst => rst, Q(31) 
                           => B_o(31), Q(30) => B_o(30), Q(29) => B_o(29), 
                           Q(28) => B_o(28), Q(27) => B_o(27), Q(26) => B_o(26)
                           , Q(25) => B_o(25), Q(24) => B_o(24), Q(23) => 
                           B_o(23), Q(22) => B_o(22), Q(21) => B_o(21), Q(20) 
                           => B_o(20), Q(19) => B_o(19), Q(18) => B_o(18), 
                           Q(17) => B_o(17), Q(16) => B_o(16), Q(15) => B_o(15)
                           , Q(14) => B_o(14), Q(13) => B_o(13), Q(12) => 
                           B_o(12), Q(11) => B_o(11), Q(10) => B_o(10), Q(9) =>
                           B_o(9), Q(8) => B_o(8), Q(7) => B_o(7), Q(6) => 
                           B_o(6), Q(5) => B_o(5), Q(4) => B_o(4), Q(3) => 
                           B_o(3), Q(2) => B_o(2), Q(1) => B_o(1), Q(0) => 
                           B_o(0));
   rA : ff32_en_SIZE5_0 port map( D(4) => rA_i(4), D(3) => rA_i(3), D(2) => 
                           rA_i(2), D(1) => rA_i(1), D(0) => rA_i(0), en => 
                           enable, clk => clk, rst => rst, Q(4) => rA_o(4), 
                           Q(3) => rA_o(3), Q(2) => rA_o(2), Q(1) => rA_o(1), 
                           Q(0) => rA_o(0));
   rB : ff32_en_SIZE5_3 port map( D(4) => rB_i(4), D(3) => rB_i(3), D(2) => 
                           rB_i(2), D(1) => rB_i(1), D(0) => rB_i(0), en => 
                           enable, clk => clk, rst => rst, Q(4) => rB_o(4), 
                           Q(3) => rB_o(3), Q(2) => rB_o(2), Q(1) => rB_o(1), 
                           Q(0) => rB_o(0));
   rC : ff32_en_SIZE5_2 port map( D(4) => rC_i(4), D(3) => rC_i(3), D(2) => 
                           rC_i(2), D(1) => rC_i(1), D(0) => rC_i(0), en => 
                           enable, clk => clk, rst => rst, Q(4) => rC_o(4), 
                           Q(3) => rC_o(3), Q(2) => rC_o(2), Q(1) => rC_o(1), 
                           Q(0) => rC_o(0));
   IMM : ff32_en_SIZE32_4 port map( D(31) => IMM_i(31), D(30) => IMM_i(30), 
                           D(29) => IMM_i(29), D(28) => IMM_i(28), D(27) => 
                           IMM_i(27), D(26) => IMM_i(26), D(25) => IMM_i(25), 
                           D(24) => IMM_i(24), D(23) => IMM_i(23), D(22) => 
                           IMM_i(22), D(21) => IMM_i(21), D(20) => IMM_i(20), 
                           D(19) => IMM_i(19), D(18) => IMM_i(18), D(17) => 
                           IMM_i(17), D(16) => IMM_i(16), D(15) => IMM_i(15), 
                           D(14) => IMM_i(14), D(13) => IMM_i(13), D(12) => 
                           IMM_i(12), D(11) => IMM_i(11), D(10) => IMM_i(10), 
                           D(9) => IMM_i(9), D(8) => IMM_i(8), D(7) => IMM_i(7)
                           , D(6) => IMM_i(6), D(5) => IMM_i(5), D(4) => 
                           IMM_i(4), D(3) => IMM_i(3), D(2) => IMM_i(2), D(1) 
                           => IMM_i(1), D(0) => IMM_i(0), en => enable, clk => 
                           clk, rst => rst, Q(31) => IMM_o(31), Q(30) => 
                           IMM_o(30), Q(29) => IMM_o(29), Q(28) => IMM_o(28), 
                           Q(27) => IMM_o(27), Q(26) => IMM_o(26), Q(25) => 
                           IMM_o(25), Q(24) => IMM_o(24), Q(23) => IMM_o(23), 
                           Q(22) => IMM_o(22), Q(21) => IMM_o(21), Q(20) => 
                           IMM_o(20), Q(19) => IMM_o(19), Q(18) => IMM_o(18), 
                           Q(17) => IMM_o(17), Q(16) => IMM_o(16), Q(15) => 
                           IMM_o(15), Q(14) => IMM_o(14), Q(13) => IMM_o(13), 
                           Q(12) => IMM_o(12), Q(11) => IMM_o(11), Q(10) => 
                           IMM_o(10), Q(9) => IMM_o(9), Q(8) => IMM_o(8), Q(7) 
                           => IMM_o(7), Q(6) => IMM_o(6), Q(5) => IMM_o(5), 
                           Q(4) => IMM_o(4), Q(3) => IMM_o(3), Q(2) => IMM_o(2)
                           , Q(1) => IMM_o(1), Q(0) => IMM_o(0));
   ALUW : ff32_en_SIZE13 port map( D(12) => ALUW_i(12), D(11) => ALUW_i(11), 
                           D(10) => ALUW_i(10), D(9) => ALUW_i(9), D(8) => 
                           ALUW_i(8), D(7) => ALUW_i(7), D(6) => ALUW_i(6), 
                           D(5) => ALUW_i(5), D(4) => ALUW_i(4), D(3) => 
                           ALUW_i(3), D(2) => ALUW_i(2), D(1) => ALUW_i(1), 
                           D(0) => ALUW_i(0), en => enable, clk => clk, rst => 
                           rst, Q(12) => ALUW_o(12), Q(11) => ALUW_o(11), Q(10)
                           => ALUW_o(10), Q(9) => ALUW_o(9), Q(8) => ALUW_o(8),
                           Q(7) => ALUW_o(7), Q(6) => ALUW_o(6), Q(5) => 
                           ALUW_o(5), Q(4) => ALUW_o(4), Q(3) => ALUW_o(3), 
                           Q(2) => ALUW_o(2), Q(1) => ALUW_o(1), Q(0) => 
                           ALUW_o(0));
   U1 : INV_X8 port map( A => stall_i, ZN => enable);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity dlx_regfile is

   port( Clk, Rst, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, 
         ADD_RD2 : in std_logic_vector (4 downto 0);  DATAIN : in 
         std_logic_vector (31 downto 0);  OUT1, OUT2 : out std_logic_vector (31
         downto 0));

end dlx_regfile;

architecture SYN_A of dlx_regfile is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X4
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n2152, n2184, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703,
      n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, 
      n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, 
      n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, 
      n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, 
      n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, 
      n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, 
      n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, 
      n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, 
      n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, 
      n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, 
      n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, 
      n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, 
      n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, 
      n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, 
      n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, 
      n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, 
      n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, 
      n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, 
      n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, 
      n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, 
      n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, 
      n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, 
      n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, 
      n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, 
      n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, 
      n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, 
      n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, 
      n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, 
      n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, 
      n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, 
      n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, 
      n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, 
      n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, 
      n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, 
      n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, 
      n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, 
      n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, 
      n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, 
      n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, 
      n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, 
      n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, 
      n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, 
      n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, 
      n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, 
      n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, 
      n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, 
      n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, 
      n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, 
      n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, 
      n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, 
      n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, 
      n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, 
      n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, 
      n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, 
      n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, 
      n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, 
      n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, 
      n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, 
      n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, 
      n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, 
      n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, 
      n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, 
      n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, 
      n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, 
      n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, 
      n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, 
      n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, 
      n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, 
      n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, 
      n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, 
      n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, 
      n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, 
      n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, 
      n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, 
      n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, 
      n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, 
      n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, 
      n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, 
      n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, 
      n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, 
      n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, 
      n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, 
      n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, 
      n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, 
      n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, 
      n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, 
      n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, 
      n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, 
      n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, 
      n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, 
      n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, 
      n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, 
      n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, 
      n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, 
      n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, 
      n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, 
      n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, 
      n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, 
      n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, 
      n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, 
      n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, 
      n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, 
      n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, 
      n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, 
      n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n222, n353, n354,
      n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, 
      n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, 
      n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, 
      n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, 
      n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, 
      n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, 
      n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, 
      n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, 
      n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, 
      n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, 
      n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, 
      n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, 
      n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, 
      n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, 
      n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, 
      n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, 
      n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, 
      n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, 
      n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, 
      n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, 
      n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, 
      n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, 
      n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, 
      n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, 
      n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, 
      n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, 
      n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, 
      n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, 
      n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, 
      n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, 
      n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, 
      n727, n728, n729, n730, n731, n732, n733, n734, n2087, n2219, n2220, 
      n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, 
      n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, 
      n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2601, n2634, 
      n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, 
      n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, 
      n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, 
      n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, 
      n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, 
      n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, 
      n3784, net644357, net644358, net644359, net644360, net644361, net644362, 
      net644363, net644364, net644365, net644366, net644367, net644368, 
      net644369, net644370, net644371, net644372, net644373, net644374, 
      net644375, net644376, net644377, net644378, net644379, net644380, 
      net644381, net644382, net644383, net644384, net644385, net644386, 
      net644387, net644388, net644389, net644390, net644391, net644392, 
      net644393, net644394, net644395, net644396, net644397, net644398, 
      net644399, net644400, net644401, net644402, net644403, net644404, 
      net644405, net644406, net644407, net644408, net644409, net644410, 
      net644411, net644412, net644413, net644414, net644415, net644416, 
      net644417, net644418, net644419, net644420, net644421, net644422, 
      net644423, net644424, net644425, net644426, net644427, net644428, 
      net644429, net644430, net644431, net644432, net644433, net644434, 
      net644435, net644436, net644437, net644438, net644439, net644440, 
      net644441, net644442, net644443, net644444, net644445, net644446, 
      net644447, net644448, net644449, net644450, net644451, net644452, 
      net644453, net644454, net644455, net644456, net644457, net644458, 
      net644459, net644460, net644461, net644462, net644463, net644464, 
      net644465, net644466, net644467, net644468, net644469, net644470, 
      net644471, net644472, net644473, net644474, net644475, net644476, 
      net644477, net644478, net644479, net644480, net644481, net644482, 
      net644483, net644484, net644485, net644486, net644487, net644488, 
      net644489, net644490, net644491, net644492, net644493, net644494, 
      net644495, net644496, net644497, net644498, net644499, net644500, 
      net644501, net644502, net644503, net644504, net644505, net644506, 
      net644507, net644508, net644509, net644510, net644511, net644512, 
      net644513, net644514, net644515, net644516, net644517, net644518, 
      net644519, net644520, net644521, net644522, net644523, net644524, 
      net644525, net644526, net644527, net644528, net644529, net644530, 
      net644531, net644532, net644533, net644534, net644535, net644536, 
      net644537, net644538, net644539, net644540, net644541, net644542, 
      net644543, net644544, net644545, net644546, net644547, net644548, 
      net644549, net644550, net644551, net644552, net644553, net644554, 
      net644555, net644556, net644557, net644558, net644559, net644560, 
      net644561, net644562, net644563, net644564, net644565, net644566, 
      net644567, net644568, net644569, net644570, net644571, net644572, 
      net644573, net644574, net644575, net644576, net644577, net644578, 
      net644579, net644580, net644581, net644582, net644583, net644584, 
      net644585, net644586, net644587, net644588, net644589, net644590, 
      net644591, net644592, net644593, net644594, net644595, net644596, 
      net644597, net644598, net644599, net644600, net644601, net644602, 
      net644603, net644604, net644605, net644606, net644607, net644608, 
      net644609, net644610, net644611, net644612, net644613, net644614, 
      net644615, net644616, net644617, net644618, net644619, net644620, 
      net644621, net644622, net644623, net644624, net644625, net644626, 
      net644627, net644628, net644629, net644630, net644631, net644632, 
      net644633, net644634, net644635, net644636, net644637, net644638, 
      net644639, net644640, net644641, net644642, net644643, net644644, 
      net644645, net644646, net644647, net644648, net644649, net644650, 
      net644651, net644652, net644653, net644654, net644655, net644656, 
      net644657, net644658, net644659, net644660, net644661, net644662, 
      net644663, net644664, net644665, net644666, net644667, net644668, 
      net644669, net644670, net644671, net644672, net644673, net644674, 
      net644675, net644676, net644677, net644678, net644679, net644680, 
      net644681, net644682, net644683, net644684, net644685, net644686, 
      net644687, net644688, net644689, net644690, net644691, net644692, 
      net644693, net644694, net644695, net644696, net644697, net644698, 
      net644699, net644700, net644701, net644702, net644703, net644704, 
      net644705, net644706, net644707, net644708, net644709, net644710, 
      net644711, net644712, net644713, net644714, net644715, net644716, 
      net644717, net644718, net644719, net644720, net644721, net644722, 
      net644723, net644724, net644725, net644726, net644727, net644728, 
      net644729, net644730, net644731, net644732, net644733, net644734, 
      net644735, net644736, net644737, net644738, net644739, net644740, 
      net644741, net644742, net644743, net644744, net644745, net644746, 
      net644747, net644748, net644749, net644750, net644751, net644752, 
      net644753, net644754, net644755, net644756, net644757, net644758, 
      net644759, net644760, net644761, net644762, net644763, net644764, 
      net644765, net644766, net644767, net644768, net644769, net644770, 
      net644771, net644772, net644773, net644774, net644775, net644776, 
      net644777, net644778, net644779, net644780, net644781, net644782, 
      net644783, net644784, net644785, net644786, net644787, net644788, 
      net644789, net644790, net644791, net644792, net644793, net644794, 
      net644795, net644796, net644797, net644798, net644799, net644800, 
      net644801, net644802, net644803, net644804, net644805, net644806, 
      net644807, net644808, net644809, net644810, net644811, net644812, 
      net644813, net644814, net644815, net644816, net644817, net644818, 
      net644819, net644820, net644821, net644822, net644823, net644824, 
      net644825, net644826, net644827, net644828, net644829, net644830, 
      net644831, net644832, net644833, net644834, net644835, net644836, 
      net644837, net644838, net644839, net644840, net644841, net644842, 
      net644843, net644844, net644845, net644846, net644847, net644848, 
      net644849, net644850, net644851, net644852, net644853, net644854, 
      net644855, net644856, net644857, net644858, net644859, net644860, 
      net644861, net644862, net644863, net644864, net644865, net644866, 
      net644867, net644868, net644869, net644870, net644871, net644872, 
      net644873, net644874, net644875, net644876, net644877, net644878, 
      net644879, net644880, net644881, net644882, net644883, net644884, 
      net644885, net644886, net644887, net644888, net644889, net644890, 
      net644891, net644892, net644893, net644894, net644895, net644896, 
      net644897, net644898, net644899, net644900, net644901, net644902, 
      net644903, net644904, net644905, net644906, net644907, net644908, 
      net644909, net644910, net644911, net644912, net644913, net644914, 
      net644915, net644916, net644917, net644918, net644919, net644920, 
      net644921, net644922, net644923, net644924, net644925, net644926, 
      net644927, net644928, net644929, net644930, net644931, net644932, 
      net644933, n1662, n1663, n1664, n1666, n1668, n1670, n1672, n1674, n1676,
      n1678, n1680, n1682, n1684, n1686, n1688, n1690, n1692, n1694, n1696, 
      n1698, n1700, n1702, n1704, n1706, n1708, n1710, n1712, n1714, n1716, 
      n1718, n1720, n1722, n1724, n1726, n1728, n1729, n1730, n1731, n1733, 
      n1735, n1736, n1768, n1769, n1770, n1772, n1773, n1805, n1806, n1807, 
      n1808, n1811, n1812, n1843, n1844, n1846, n1847, n1848, n1850, n1852, 
      n1853, n1885, n1886, n1917, n1918, n1919, n1921, n1922, n1954, n1956, 
      n1957, n1990, n1991, n2023, n2024, n2025, n2027, n2028, n2060, n2062, 
      n2063, n3888, n3889, n3892, n3893, n3924, n3926, n3927, n3959, n3961, 
      n3962, n3994, n3995, n3996, n3997, n4000, n4001, n4033, n4035, n4036, 
      n4068, n4069, n4073, n4074, n4106, n4107, n4108, n4110, n4111, n4143, 
      n4145, n4146, n4178, n4180, n4181, n4182, n4183, n4184, n4185, n4186, 
      n4187, n4188, n4189, n4190, n4192, n4194, n4195, n4196, n4197, n4198, 
      n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4207, n4208, n4209, 
      n4210, n4211, n4212, n4214, n4215, n4216, n4217, n4218, n4219, n4220, 
      n4221, n4223, n4224, n4225, n4226, n4228, n4229, n4231, n4232, n4233, 
      n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4243, n4246, 
      n4247, n4248, n4249, n4250, n4251, n4252, n4254, n4255, n4256, n4257, 
      n4258, n4259, n4260, n4261, n4264, n4265, n4266, n4267, n4270, n4271, 
      n4272, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4284, n4285, 
      n4286, n4287, n4288, n4289, n4290, n4291, n4294, n4295, n4296, n4297, 
      n4300, n4301, n4302, n4306, n4307, n4308, n4309, n4310, n4311, n4312, 
      n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4324, n4325, 
      n4326, n4327, n4330, n4331, n4332, n4336, n4337, n4338, n4339, n4340, 
      n4341, n4342, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, 
      n4354, n4355, n4356, n4357, n4360, n4361, n4362, n4366, n4367, n4368, 
      n4369, n4370, n4371, n4372, n4374, n4375, n4376, n4377, n4378, n4379, 
      n4380, n4381, n4384, n4385, n4386, n4387, n4390, n4391, n4392, n4396, 
      n4397, n4398, n4399, n4400, n4401, n4402, n4404, n4405, n4406, n4407, 
      n4408, n4409, n4410, n4411, n4414, n4415, n4416, n4417, n4420, n4421, 
      n4422, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4434, n4435, 
      n4436, n4437, n4438, n4439, n4440, n4441, n4444, n4445, n4446, n4447, 
      n4450, n4451, n4452, n4456, n4457, n4458, n4459, n4460, n4461, n4462, 
      n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4474, n4475, 
      n4476, n4477, n4480, n4481, n4482, n4486, n4487, n4488, n4489, n4490, 
      n4491, n4492, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, 
      n4504, n4505, n4506, n4507, n4510, n4511, n4512, n4516, n4517, n4518, 
      n4519, n4520, n4521, n4522, n4524, n4525, n4526, n4527, n4528, n4529, 
      n4530, n4531, n4534, n4535, n4536, n4537, n4540, n4541, n4542, n4546, 
      n4547, n4548, n4549, n4550, n4551, n4552, n4554, n4555, n4556, n4557, 
      n4558, n4559, n4560, n4561, n4564, n4565, n4566, n4567, n4570, n4571, 
      n4572, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4584, n4585, 
      n4586, n4587, n4588, n4589, n4590, n4591, n4594, n4595, n4596, n4597, 
      n4600, n4601, n4602, n4606, n4607, n4608, n4609, n4610, n4611, n4612, 
      n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4624, n4625, 
      n4626, n4627, n4630, n4631, n4632, n4636, n4637, n4638, n4639, n4640, 
      n4641, n4642, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, 
      n4654, n4655, n4656, n4657, n4660, n4661, n4662, n4666, n4667, n4668, 
      n4669, n4670, n4671, n4672, n4674, n4675, n4676, n4677, n4678, n4679, 
      n4680, n4681, n4684, n4685, n4686, n4687, n4690, n4691, n4692, n4696, 
      n4697, n4698, n4699, n4700, n4701, n4702, n4704, n4705, n4706, n4707, 
      n4708, n4709, n4710, n4711, n4714, n4715, n4716, n4717, n4720, n4721, 
      n4722, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4734, n4735, 
      n4736, n4737, n4738, n4739, n4740, n4741, n4744, n4745, n4746, n4747, 
      n4750, n4751, n4752, n4756, n4757, n4758, n4759, n4760, n4761, n4762, 
      n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4774, n4775, 
      n4776, n4777, n4780, n4781, n4782, n4786, n4787, n4788, n4789, n4790, 
      n4791, n4792, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, 
      n4804, n4805, n4806, n4807, n4810, n4811, n4812, n4816, n4817, n4818, 
      n4819, n4820, n4821, n4822, n4824, n4825, n4826, n4827, n4828, n4829, 
      n4830, n4831, n4834, n4835, n4836, n4837, n4840, n4841, n4842, n4846, 
      n4847, n4848, n4849, n4850, n4851, n4852, n4854, n4855, n4856, n4857, 
      n4858, n4859, n4860, n4861, n4864, n4865, n4866, n4867, n4870, n4871, 
      n4872, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4884, n4885, 
      n4886, n4887, n4888, n4889, n4890, n4891, n4894, n4895, n4896, n4897, 
      n4900, n4901, n4902, n4906, n4907, n4908, n4909, n4910, n4911, n4912, 
      n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4924, n4925, 
      n4926, n4927, n4930, n4931, n4932, n4936, n4937, n4938, n4939, n4940, 
      n4941, n4942, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, 
      n4954, n4955, n4956, n4957, n4960, n4961, n4962, n4966, n4967, n4968, 
      n4969, n4970, n4971, n4972, n4974, n4975, n4976, n4977, n4978, n4979, 
      n4980, n4981, n4984, n4985, n4986, n4987, n4990, n4991, n4992, n4996, 
      n4997, n4998, n4999, n5000, n5001, n5002, n5004, n5005, n5006, n5007, 
      n5008, n5009, n5010, n5011, n5014, n5015, n5016, n5017, n5020, n5021, 
      n5022, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5034, n5035, 
      n5036, n5037, n5038, n5039, n5040, n5041, n5044, n5045, n5046, n5047, 
      n5050, n5051, n5052, n5056, n5057, n5058, n5059, n5060, n5061, n5062, 
      n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5074, n5075, 
      n5076, n5077, n5080, n5081, n5082, n5086, n5087, n5088, n5089, n5090, 
      n5091, n5092, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, 
      n5104, n5105, n5106, n5107, n5110, n5111, n5112, n5116, n5117, n5118, 
      n5119, n5120, n5121, n5122, n5124, n5125, n5126, n5127, n5128, n5129, 
      n5130, n5131, n5132, n5135, n5136, n5137, n5138, n5140, n5141, n5142, 
      n5143, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5154, n5155, 
      n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, 
      n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5175, n5176, 
      n5177, n5178, n5179, n5181, n5182, n5184, n5185, n5186, n5187, n5189, 
      n5190, n5191, n5192, n5194, n5195, n5196, n5197, n5198, n5199, n5200, 
      n5201, n5202, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, 
      n5213, n5214, n5215, n5216, n5217, n5219, n5220, n5221, n5222, n5223, 
      n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, 
      n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, 
      n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5253, n5254, 
      n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, 
      n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, 
      n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, 
      n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, 
      n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, 
      n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, 
      n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, 
      n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, 
      n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, 
      n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, 
      n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, 
      n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, 
      n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, 
      n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, 
      n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, 
      n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, 
      n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, 
      n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, 
      n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, 
      n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, 
      n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, 
      n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, 
      n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, 
      n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, 
      n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, 
      n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, 
      n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, 
      n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, 
      n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, 
      n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, 
      n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, 
      n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, 
      n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, 
      n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, 
      n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, 
      n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, 
      n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, 
      n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, 
      n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, 
      n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, 
      n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, 
      n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, 
      n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, 
      n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, 
      n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, 
      n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, 
      n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, 
      n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, 
      n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, 
      n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, 
      n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, 
      n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, 
      n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, 
      n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, 
      n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, 
      n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, 
      n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, 
      n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, 
      n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, 
      n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, 
      n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, 
      n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, 
      n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, 
      n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, 
      n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, 
      n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, 
      n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, 
      n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5934, n5935, 
      n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, 
      n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, 
      n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5966, 
      n5967, n5968, n5969, n5971, n5972, n5973, n5974, n5975, n5976, n5977, 
      n5978, n5979, n5980, n5981, n5982, n5983, n5984, n3880, n3881, n3882, 
      n3883, n3884, n3885, n3886, n3887, n3890, n3891, n3894, n3895, n3896, 
      n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, 
      n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, 
      n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3925, n3928, n3929, 
      n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, 
      n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, 
      n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3960, 
      n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, 
      n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, 
      n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, 
      n3993, n3998, n3999, n4002, n4003, n4004, n4005, n4006, n4007, n4008, 
      n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, 
      n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, 
      n4029, n4030, n4031, n4032, n4034, n4037, n4038, n4039, n4040, n4041, 
      n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, 
      n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, 
      n4062, n4063, n4064, n4065, n4066, n4067, n4070, n4071, n4072, n4075, 
      n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, 
      n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, 
      n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, 
      n4109, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, 
      n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, 
      n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, 
      n4141, n4142, n4144, n4147, n4148, n4149, n4150, n4151, n4152, n4153, 
      n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, 
      n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, 
      n4174, n4175, n4176, n4177, n4179, n4191, n4193, n4206, n4213, n4222, 
      n4227, n4230, n4242, n4244, n4245, n4253, n4262, n4263, n4268, n4269, 
      n4273, n4274, n4275, n4283, n4292, n4293, n4298, n4299, n4303, n4304, 
      n4305, n4313, n4322, n4323, n4328, n4329, n4333, n4334, n4335, n4343, 
      n4352, n4353, n4358, n4359, n4363, n4364, n4365, n4373, n4382, n4383, 
      n4388, n4389, n4393, n4394, n4395, n4403, n4412, n4413, n4418, n4419, 
      n4423, n4424, n4425, n4433, n4442, n4443, n4448, n4449, n4453, n4454, 
      n4455, n4463, n4472, n4473, n4478, n4479, n4483, n4484, n4485, n4493, 
      n4502, n4503, n4508, n4509, n4513, n4514, n4515, n4523, n4532, n4533, 
      n4538, n4539, n4543, n4544, n4545, n4553, n4562, n4563, n4568, n4569, 
      n4573, n4574, n4575, n4583, n4592, n4593, n4598, n4599, n4603, n4604, 
      n4605, n4613, n4622, n4623, n4628, n4629, n4633, n4634, n4635, n4643, 
      n4652, n4653, n4658, n4659, n4663, n4664, n4665, n4673, n4682, n4683, 
      n4688, n4689, n4693, n4694, n4695, n4703, n4712, n4713, n4718, n4719, 
      n4723, n4724, n4725, n4733, n4742, n4743, n4748, n4749, n4753, n4754, 
      n4755, n4763, n4772, n4773, n4778, n4779, n4783, n4784, n4785, n4793, 
      n4802, n4803, n4808, n4809, n4813, n4814, n4815, n4823, n4832, n4833, 
      n4838, n4839, n4843, n4844, n4845, n4853, n4862, n4863, n4868, n4869, 
      n4873, n4874, n4875, n4883, n4892, n4893, n4898, n4899, n4903, n4904, 
      n4905, n4913, n4922, n4923, n4928, n4929, n4933, n4934, n4935, n4943, 
      n4952, n4953, n4958, n4959, n4963, n4964, n4965, n4973, n4982, n4983, 
      n4988, n4989, n4993, n4994, n4995, n5003, n5012, n5013, n5018, n5019, 
      n5023, n5024, n5025, n5033, n5042, n5043, n5048, n5049, n5053, n5054, 
      n5055, n5063, n5072, n5073, n5078, n5079, n5083, n5084, n5085, n5093, 
      n5102, n5103, n5108, n5109, n5113, n5114, n5115, n5123, n5133, n5134, 
      n5139, n5144, n5145, n5153, n5174, n5180, n5183, n5188, n5193, n5203, 
      n5204, n5218, n5252, n5933, n5965, n5970, n5985, n5986, n5987, n5988, 
      n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, 
      n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, 
      n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, 
      n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, 
      n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, 
      n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, 
      n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, 
      n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, 
      n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, 
      n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, 
      n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, 
      n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, 
      n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, 
      n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, 
      n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, 
      n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, 
      n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, 
      n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, 
      n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, 
      n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, 
      n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, 
      n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, 
      n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, 
      n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, 
      n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, 
      n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, 
      n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, 
      n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, 
      n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, 
      n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, 
      n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, 
      n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, 
      n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, 
      n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, 
      n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, 
      n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, 
      n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, 
      n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, 
      n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, 
      n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, 
      n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, 
      n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, 
      n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, 
      n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, 
      n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, 
      n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, net684169, 
      net684170, net684171, net684172, net684173, net684174, net684175, 
      net684176, net684177, net684178, net684179, net684180, net684181, 
      net684182, net684183, net684184, net684185, net684186, net684187, 
      net684188, net684189, net684190, net684191, net684192, net684193, 
      net684194, net684195, net684196, net684197, net684198, net684199, 
      net684200, net684201, net684202, net684203, net684204, net684205, 
      net684206, net684207, net684208, net684209, net684210, net684211, 
      net684212, net684213, net684214, net684215, net684216, net684217, 
      net684218, net684219, net684220, net684221, net684222, net684223, 
      net684224, net684225, net684226, net684227, net684228, net684229, 
      net684230, net684231, net684232, net684233, net684234, net684235, 
      net684236, net684237, net684238, net684239, net684240, net684241, 
      net684242, net684243, net684244, net684245, net684246, net684247, 
      net684248, net684249, net684250, net684251, net684252, net684253, 
      net684254, net684255, net684256, net684257, net684258, net684259, 
      net684260, net684261, net684262, net684263, net684264, net684265, 
      net684266, net684267, net684268, net684269, net684270, net684271, 
      net684272, net684273, net684274, net684275, net684276, net684277, 
      net684278, net684279, net684280, net684281, net684282, net684283, 
      net684284, net684285, net684286, net684287, net684288, net684289, 
      net684290, net684291, net684292, net684293, net684294, net684295, 
      net684296 : std_logic;

begin
   
   REGISTERS_reg_1_31_inst : DFF_X1 port map( D => n3751, CK => Clk, Q => 
                           net644933, QN => n6055);
   REGISTERS_reg_1_30_inst : DFF_X1 port map( D => n3750, CK => Clk, Q => 
                           net644932, QN => n6054);
   REGISTERS_reg_1_29_inst : DFF_X1 port map( D => n3749, CK => Clk, Q => 
                           net644931, QN => n6053);
   REGISTERS_reg_1_28_inst : DFF_X1 port map( D => n3748, CK => Clk, Q => 
                           net644930, QN => n6052);
   REGISTERS_reg_1_27_inst : DFF_X1 port map( D => n3747, CK => Clk, Q => 
                           net644929, QN => n6051);
   REGISTERS_reg_1_26_inst : DFF_X1 port map( D => n3746, CK => Clk, Q => 
                           net644928, QN => n6050);
   REGISTERS_reg_1_25_inst : DFF_X1 port map( D => n3745, CK => Clk, Q => 
                           net644927, QN => n6049);
   REGISTERS_reg_1_24_inst : DFF_X1 port map( D => n3744, CK => Clk, Q => 
                           net644926, QN => n6048);
   REGISTERS_reg_1_23_inst : DFF_X1 port map( D => n3743, CK => Clk, Q => 
                           net644925, QN => n6047);
   REGISTERS_reg_1_22_inst : DFF_X1 port map( D => n3742, CK => Clk, Q => 
                           net644924, QN => n6046);
   REGISTERS_reg_1_21_inst : DFF_X1 port map( D => n3741, CK => Clk, Q => 
                           net644923, QN => n6045);
   REGISTERS_reg_1_20_inst : DFF_X1 port map( D => n3740, CK => Clk, Q => 
                           net644922, QN => n6044);
   REGISTERS_reg_1_19_inst : DFF_X1 port map( D => n3739, CK => Clk, Q => 
                           net644921, QN => n6043);
   REGISTERS_reg_1_18_inst : DFF_X1 port map( D => n3738, CK => Clk, Q => 
                           net644920, QN => n6042);
   REGISTERS_reg_1_17_inst : DFF_X1 port map( D => n3737, CK => Clk, Q => 
                           net644919, QN => n6041);
   REGISTERS_reg_1_16_inst : DFF_X1 port map( D => n3736, CK => Clk, Q => 
                           net644918, QN => n6040);
   REGISTERS_reg_1_15_inst : DFF_X1 port map( D => n3735, CK => Clk, Q => 
                           net644917, QN => n6039);
   REGISTERS_reg_1_14_inst : DFF_X1 port map( D => n3734, CK => Clk, Q => 
                           net644916, QN => n6038);
   REGISTERS_reg_1_13_inst : DFF_X1 port map( D => n3733, CK => Clk, Q => 
                           net644915, QN => n6037);
   REGISTERS_reg_1_12_inst : DFF_X1 port map( D => n3732, CK => Clk, Q => 
                           net644914, QN => n6036);
   REGISTERS_reg_1_11_inst : DFF_X1 port map( D => n3731, CK => Clk, Q => 
                           net644913, QN => n6035);
   REGISTERS_reg_1_10_inst : DFF_X1 port map( D => n3730, CK => Clk, Q => 
                           net644912, QN => n6034);
   REGISTERS_reg_1_9_inst : DFF_X1 port map( D => n3729, CK => Clk, Q => 
                           net644911, QN => n6033);
   REGISTERS_reg_1_8_inst : DFF_X1 port map( D => n3728, CK => Clk, Q => 
                           net644910, QN => n6032);
   REGISTERS_reg_1_7_inst : DFF_X1 port map( D => n3727, CK => Clk, Q => 
                           net644909, QN => n6031);
   REGISTERS_reg_1_6_inst : DFF_X1 port map( D => n3726, CK => Clk, Q => 
                           net644908, QN => n6030);
   REGISTERS_reg_1_5_inst : DFF_X1 port map( D => n3725, CK => Clk, Q => 
                           net644907, QN => n6029);
   REGISTERS_reg_1_4_inst : DFF_X1 port map( D => n3724, CK => Clk, Q => 
                           net644906, QN => n6028);
   REGISTERS_reg_1_3_inst : DFF_X1 port map( D => n3723, CK => Clk, Q => 
                           net644905, QN => n6027);
   REGISTERS_reg_1_2_inst : DFF_X1 port map( D => n3722, CK => Clk, Q => 
                           net644904, QN => n6026);
   REGISTERS_reg_1_1_inst : DFF_X1 port map( D => n3721, CK => Clk, Q => 
                           net644903, QN => n6025);
   REGISTERS_reg_1_0_inst : DFF_X1 port map( D => n3720, CK => Clk, Q => 
                           net644902, QN => n6346);
   REGISTERS_reg_2_31_inst : DFF_X1 port map( D => n3719, CK => Clk, Q => n3949
                           , QN => n577);
   REGISTERS_reg_2_30_inst : DFF_X1 port map( D => n3718, CK => Clk, Q => n3948
                           , QN => n578);
   REGISTERS_reg_2_29_inst : DFF_X1 port map( D => n3717, CK => Clk, Q => n3947
                           , QN => n579);
   REGISTERS_reg_2_28_inst : DFF_X1 port map( D => n3716, CK => Clk, Q => n3946
                           , QN => n580);
   REGISTERS_reg_2_27_inst : DFF_X1 port map( D => n3715, CK => Clk, Q => n3945
                           , QN => n581);
   REGISTERS_reg_2_26_inst : DFF_X1 port map( D => n3714, CK => Clk, Q => n3944
                           , QN => n582);
   REGISTERS_reg_2_25_inst : DFF_X1 port map( D => n3713, CK => Clk, Q => n3943
                           , QN => n583);
   REGISTERS_reg_2_24_inst : DFF_X1 port map( D => n3712, CK => Clk, Q => n3942
                           , QN => n584);
   REGISTERS_reg_2_23_inst : DFF_X1 port map( D => n3711, CK => Clk, Q => n3941
                           , QN => n585);
   REGISTERS_reg_2_22_inst : DFF_X1 port map( D => n3710, CK => Clk, Q => n3940
                           , QN => n586);
   REGISTERS_reg_2_21_inst : DFF_X1 port map( D => n3709, CK => Clk, Q => n3939
                           , QN => n587);
   REGISTERS_reg_2_20_inst : DFF_X1 port map( D => n3708, CK => Clk, Q => n3938
                           , QN => n588);
   REGISTERS_reg_2_19_inst : DFF_X1 port map( D => n3707, CK => Clk, Q => n3937
                           , QN => n589);
   REGISTERS_reg_2_18_inst : DFF_X1 port map( D => n3706, CK => Clk, Q => n3936
                           , QN => n590);
   REGISTERS_reg_2_17_inst : DFF_X1 port map( D => n3705, CK => Clk, Q => n3935
                           , QN => n591);
   REGISTERS_reg_2_16_inst : DFF_X1 port map( D => n3704, CK => Clk, Q => n3934
                           , QN => n592);
   REGISTERS_reg_2_15_inst : DFF_X1 port map( D => n3703, CK => Clk, Q => n3933
                           , QN => n593);
   REGISTERS_reg_2_14_inst : DFF_X1 port map( D => n3702, CK => Clk, Q => n3932
                           , QN => n594);
   REGISTERS_reg_2_13_inst : DFF_X1 port map( D => n3701, CK => Clk, Q => n3931
                           , QN => n595);
   REGISTERS_reg_2_12_inst : DFF_X1 port map( D => n3700, CK => Clk, Q => n3930
                           , QN => n596);
   REGISTERS_reg_2_11_inst : DFF_X1 port map( D => n3699, CK => Clk, Q => n3929
                           , QN => n597);
   REGISTERS_reg_2_10_inst : DFF_X1 port map( D => n3698, CK => Clk, Q => n3928
                           , QN => n598);
   REGISTERS_reg_2_9_inst : DFF_X1 port map( D => n3697, CK => Clk, Q => n3925,
                           QN => n599);
   REGISTERS_reg_2_8_inst : DFF_X1 port map( D => n3696, CK => Clk, Q => n3923,
                           QN => n600);
   REGISTERS_reg_2_7_inst : DFF_X1 port map( D => n3695, CK => Clk, Q => n3922,
                           QN => n601);
   REGISTERS_reg_2_6_inst : DFF_X1 port map( D => n3694, CK => Clk, Q => n3921,
                           QN => n602);
   REGISTERS_reg_2_5_inst : DFF_X1 port map( D => n3693, CK => Clk, Q => n3920,
                           QN => n603);
   REGISTERS_reg_2_4_inst : DFF_X1 port map( D => n3692, CK => Clk, Q => n3919,
                           QN => n604);
   REGISTERS_reg_2_3_inst : DFF_X1 port map( D => n3691, CK => Clk, Q => n3918,
                           QN => n605);
   REGISTERS_reg_2_2_inst : DFF_X1 port map( D => n3690, CK => Clk, Q => n3917,
                           QN => n606);
   REGISTERS_reg_2_1_inst : DFF_X1 port map( D => n3689, CK => Clk, Q => n3916,
                           QN => n607);
   REGISTERS_reg_2_0_inst : DFF_X1 port map( D => n3688, CK => Clk, Q => 
                           net644901, QN => n6345);
   REGISTERS_reg_3_31_inst : DFF_X1 port map( D => n3687, CK => Clk, Q => 
                           net644900, QN => n6024);
   REGISTERS_reg_3_30_inst : DFF_X1 port map( D => n3686, CK => Clk, Q => 
                           net644899, QN => n6023);
   REGISTERS_reg_3_29_inst : DFF_X1 port map( D => n3685, CK => Clk, Q => 
                           net644898, QN => n6022);
   REGISTERS_reg_3_28_inst : DFF_X1 port map( D => n3684, CK => Clk, Q => 
                           net644897, QN => n6021);
   REGISTERS_reg_3_27_inst : DFF_X1 port map( D => n3683, CK => Clk, Q => 
                           net644896, QN => n6020);
   REGISTERS_reg_3_26_inst : DFF_X1 port map( D => n3682, CK => Clk, Q => 
                           net644895, QN => n6019);
   REGISTERS_reg_3_25_inst : DFF_X1 port map( D => n3681, CK => Clk, Q => 
                           net644894, QN => n6018);
   REGISTERS_reg_3_24_inst : DFF_X1 port map( D => n3680, CK => Clk, Q => 
                           net644893, QN => n6017);
   REGISTERS_reg_3_23_inst : DFF_X1 port map( D => n3679, CK => Clk, Q => 
                           net644892, QN => n6016);
   REGISTERS_reg_3_22_inst : DFF_X1 port map( D => n3678, CK => Clk, Q => 
                           net644891, QN => n6015);
   REGISTERS_reg_3_21_inst : DFF_X1 port map( D => n3677, CK => Clk, Q => 
                           net644890, QN => n6014);
   REGISTERS_reg_3_20_inst : DFF_X1 port map( D => n3676, CK => Clk, Q => 
                           net644889, QN => n6013);
   REGISTERS_reg_3_19_inst : DFF_X1 port map( D => n3675, CK => Clk, Q => 
                           net644888, QN => n6012);
   REGISTERS_reg_3_18_inst : DFF_X1 port map( D => n3674, CK => Clk, Q => 
                           net644887, QN => n6011);
   REGISTERS_reg_3_17_inst : DFF_X1 port map( D => n3673, CK => Clk, Q => 
                           net644886, QN => n6010);
   REGISTERS_reg_3_16_inst : DFF_X1 port map( D => n3672, CK => Clk, Q => 
                           net644885, QN => n6009);
   REGISTERS_reg_3_15_inst : DFF_X1 port map( D => n3671, CK => Clk, Q => 
                           net644884, QN => n6008);
   REGISTERS_reg_3_14_inst : DFF_X1 port map( D => n3670, CK => Clk, Q => 
                           net644883, QN => n6007);
   REGISTERS_reg_3_13_inst : DFF_X1 port map( D => n3669, CK => Clk, Q => 
                           net644882, QN => n6006);
   REGISTERS_reg_3_12_inst : DFF_X1 port map( D => n3668, CK => Clk, Q => 
                           net644881, QN => n6005);
   REGISTERS_reg_3_11_inst : DFF_X1 port map( D => n3667, CK => Clk, Q => 
                           net644880, QN => n6004);
   REGISTERS_reg_3_10_inst : DFF_X1 port map( D => n3666, CK => Clk, Q => 
                           net644879, QN => n6003);
   REGISTERS_reg_3_9_inst : DFF_X1 port map( D => n3665, CK => Clk, Q => 
                           net644878, QN => n6002);
   REGISTERS_reg_3_8_inst : DFF_X1 port map( D => n3664, CK => Clk, Q => 
                           net644877, QN => n6001);
   REGISTERS_reg_3_7_inst : DFF_X1 port map( D => n3663, CK => Clk, Q => 
                           net644876, QN => n6000);
   REGISTERS_reg_3_6_inst : DFF_X1 port map( D => n3662, CK => Clk, Q => 
                           net644875, QN => n5999);
   REGISTERS_reg_3_5_inst : DFF_X1 port map( D => n3661, CK => Clk, Q => 
                           net644874, QN => n5998);
   REGISTERS_reg_3_4_inst : DFF_X1 port map( D => n3660, CK => Clk, Q => 
                           net644873, QN => n5997);
   REGISTERS_reg_3_3_inst : DFF_X1 port map( D => n3659, CK => Clk, Q => 
                           net644872, QN => n5996);
   REGISTERS_reg_3_2_inst : DFF_X1 port map( D => n3658, CK => Clk, Q => 
                           net644871, QN => n5995);
   REGISTERS_reg_3_1_inst : DFF_X1 port map( D => n3657, CK => Clk, Q => 
                           net644870, QN => n5994);
   REGISTERS_reg_3_0_inst : DFF_X1 port map( D => n3656, CK => Clk, Q => 
                           net644869, QN => n6354);
   REGISTERS_reg_4_31_inst : DFF_X1 port map( D => n3655, CK => Clk, Q => n388,
                           QN => n4413);
   REGISTERS_reg_4_30_inst : DFF_X1 port map( D => n3654, CK => Clk, Q => n391,
                           QN => n4412);
   REGISTERS_reg_4_29_inst : DFF_X1 port map( D => n3653, CK => Clk, Q => n394,
                           QN => n4403);
   REGISTERS_reg_4_28_inst : DFF_X1 port map( D => n3652, CK => Clk, Q => n397,
                           QN => n4395);
   REGISTERS_reg_4_27_inst : DFF_X1 port map( D => n3651, CK => Clk, Q => n400,
                           QN => n4394);
   REGISTERS_reg_4_26_inst : DFF_X1 port map( D => n3650, CK => Clk, Q => n403,
                           QN => n4393);
   REGISTERS_reg_4_25_inst : DFF_X1 port map( D => n3649, CK => Clk, Q => n406,
                           QN => n4389);
   REGISTERS_reg_4_24_inst : DFF_X1 port map( D => n3648, CK => Clk, Q => n409,
                           QN => n4388);
   REGISTERS_reg_4_23_inst : DFF_X1 port map( D => n3647, CK => Clk, Q => n412,
                           QN => n4383);
   REGISTERS_reg_4_22_inst : DFF_X1 port map( D => n3646, CK => Clk, Q => n415,
                           QN => n4382);
   REGISTERS_reg_4_21_inst : DFF_X1 port map( D => n3645, CK => Clk, Q => n418,
                           QN => n4373);
   REGISTERS_reg_4_20_inst : DFF_X1 port map( D => n3644, CK => Clk, Q => n421,
                           QN => n4365);
   REGISTERS_reg_4_19_inst : DFF_X1 port map( D => n3643, CK => Clk, Q => n424,
                           QN => n4364);
   REGISTERS_reg_4_18_inst : DFF_X1 port map( D => n3642, CK => Clk, Q => n427,
                           QN => n4363);
   REGISTERS_reg_4_17_inst : DFF_X1 port map( D => n3641, CK => Clk, Q => n430,
                           QN => n4359);
   REGISTERS_reg_4_16_inst : DFF_X1 port map( D => n3640, CK => Clk, Q => n433,
                           QN => n4358);
   REGISTERS_reg_4_15_inst : DFF_X1 port map( D => n3639, CK => Clk, Q => n436,
                           QN => n4353);
   REGISTERS_reg_4_14_inst : DFF_X1 port map( D => n3638, CK => Clk, Q => n439,
                           QN => n4352);
   REGISTERS_reg_4_13_inst : DFF_X1 port map( D => n3637, CK => Clk, Q => n442,
                           QN => n4343);
   REGISTERS_reg_4_12_inst : DFF_X1 port map( D => n3636, CK => Clk, Q => n445,
                           QN => n4335);
   REGISTERS_reg_4_11_inst : DFF_X1 port map( D => n3635, CK => Clk, Q => n448,
                           QN => n4334);
   REGISTERS_reg_4_10_inst : DFF_X1 port map( D => n3634, CK => Clk, Q => n451,
                           QN => n4333);
   REGISTERS_reg_4_9_inst : DFF_X1 port map( D => n3633, CK => Clk, Q => n454, 
                           QN => n4329);
   REGISTERS_reg_4_8_inst : DFF_X1 port map( D => n3632, CK => Clk, Q => n457, 
                           QN => n4328);
   REGISTERS_reg_4_7_inst : DFF_X1 port map( D => n3631, CK => Clk, Q => n460, 
                           QN => n4323);
   REGISTERS_reg_4_6_inst : DFF_X1 port map( D => n3630, CK => Clk, Q => n463, 
                           QN => n4322);
   REGISTERS_reg_4_5_inst : DFF_X1 port map( D => n3629, CK => Clk, Q => n466, 
                           QN => n4313);
   REGISTERS_reg_4_4_inst : DFF_X1 port map( D => n3628, CK => Clk, Q => n469, 
                           QN => n4305);
   REGISTERS_reg_4_3_inst : DFF_X1 port map( D => n3627, CK => Clk, Q => n472, 
                           QN => n4304);
   REGISTERS_reg_4_2_inst : DFF_X1 port map( D => n3626, CK => Clk, Q => n475, 
                           QN => n4303);
   REGISTERS_reg_4_1_inst : DFF_X1 port map( D => n3625, CK => Clk, Q => n478, 
                           QN => n4299);
   REGISTERS_reg_4_0_inst : DFF_X1 port map( D => n3624, CK => Clk, Q => 
                           net644868, QN => n6353);
   REGISTERS_reg_5_31_inst : DFF_X1 port map( D => n3623, CK => Clk, Q => n4058
                           , QN => n3784);
   REGISTERS_reg_5_30_inst : DFF_X1 port map( D => n3622, CK => Clk, Q => n4055
                           , QN => n3783);
   REGISTERS_reg_5_29_inst : DFF_X1 port map( D => n3621, CK => Clk, Q => n4052
                           , QN => n3782);
   REGISTERS_reg_5_28_inst : DFF_X1 port map( D => n3620, CK => Clk, Q => n4049
                           , QN => n3781);
   REGISTERS_reg_5_27_inst : DFF_X1 port map( D => n3619, CK => Clk, Q => n4046
                           , QN => n3780);
   REGISTERS_reg_5_26_inst : DFF_X1 port map( D => n3618, CK => Clk, Q => n4043
                           , QN => n3779);
   REGISTERS_reg_5_25_inst : DFF_X1 port map( D => n3617, CK => Clk, Q => n4040
                           , QN => n3778);
   REGISTERS_reg_5_24_inst : DFF_X1 port map( D => n3616, CK => Clk, Q => n4037
                           , QN => n3777);
   REGISTERS_reg_5_23_inst : DFF_X1 port map( D => n3615, CK => Clk, Q => n4031
                           , QN => n3776);
   REGISTERS_reg_5_22_inst : DFF_X1 port map( D => n3614, CK => Clk, Q => n4028
                           , QN => n3775);
   REGISTERS_reg_5_21_inst : DFF_X1 port map( D => n3613, CK => Clk, Q => n4025
                           , QN => n3774);
   REGISTERS_reg_5_20_inst : DFF_X1 port map( D => n3612, CK => Clk, Q => n4022
                           , QN => n3773);
   REGISTERS_reg_5_19_inst : DFF_X1 port map( D => n3611, CK => Clk, Q => n4019
                           , QN => n3772);
   REGISTERS_reg_5_18_inst : DFF_X1 port map( D => n3610, CK => Clk, Q => n4016
                           , QN => n3771);
   REGISTERS_reg_5_17_inst : DFF_X1 port map( D => n3609, CK => Clk, Q => n4013
                           , QN => n3770);
   REGISTERS_reg_5_16_inst : DFF_X1 port map( D => n3608, CK => Clk, Q => n4010
                           , QN => n3769);
   REGISTERS_reg_5_15_inst : DFF_X1 port map( D => n3607, CK => Clk, Q => n4007
                           , QN => n3768);
   REGISTERS_reg_5_14_inst : DFF_X1 port map( D => n3606, CK => Clk, Q => n4004
                           , QN => n3767);
   REGISTERS_reg_5_13_inst : DFF_X1 port map( D => n3605, CK => Clk, Q => n3999
                           , QN => n3766);
   REGISTERS_reg_5_12_inst : DFF_X1 port map( D => n3604, CK => Clk, Q => n3992
                           , QN => n3765);
   REGISTERS_reg_5_11_inst : DFF_X1 port map( D => n3603, CK => Clk, Q => n3989
                           , QN => n3764);
   REGISTERS_reg_5_10_inst : DFF_X1 port map( D => n3602, CK => Clk, Q => n3986
                           , QN => n3763);
   REGISTERS_reg_5_9_inst : DFF_X1 port map( D => n3601, CK => Clk, Q => n3983,
                           QN => n3762);
   REGISTERS_reg_5_8_inst : DFF_X1 port map( D => n3600, CK => Clk, Q => n3980,
                           QN => n3761);
   REGISTERS_reg_5_7_inst : DFF_X1 port map( D => n3599, CK => Clk, Q => n3977,
                           QN => n3760);
   REGISTERS_reg_5_6_inst : DFF_X1 port map( D => n3598, CK => Clk, Q => n3974,
                           QN => n3759);
   REGISTERS_reg_5_5_inst : DFF_X1 port map( D => n3597, CK => Clk, Q => n3971,
                           QN => n3758);
   REGISTERS_reg_5_4_inst : DFF_X1 port map( D => n3596, CK => Clk, Q => n3968,
                           QN => n3757);
   REGISTERS_reg_5_3_inst : DFF_X1 port map( D => n3595, CK => Clk, Q => n3965,
                           QN => n3756);
   REGISTERS_reg_5_2_inst : DFF_X1 port map( D => n3594, CK => Clk, Q => n3960,
                           QN => n3755);
   REGISTERS_reg_5_1_inst : DFF_X1 port map( D => n3593, CK => Clk, Q => n3956,
                           QN => n3754);
   REGISTERS_reg_5_0_inst : DFF_X1 port map( D => n3592, CK => Clk, Q => 
                           net644867, QN => n6344);
   REGISTERS_reg_6_31_inst : DFF_X1 port map( D => n3591, CK => Clk, Q => 
                           net644866, QN => n6336);
   REGISTERS_reg_6_30_inst : DFF_X1 port map( D => n3590, CK => Clk, Q => 
                           net644865, QN => n6335);
   REGISTERS_reg_6_29_inst : DFF_X1 port map( D => n3589, CK => Clk, Q => 
                           net644864, QN => n6334);
   REGISTERS_reg_6_28_inst : DFF_X1 port map( D => n3588, CK => Clk, Q => 
                           net644863, QN => n6333);
   REGISTERS_reg_6_27_inst : DFF_X1 port map( D => n3587, CK => Clk, Q => 
                           net644862, QN => n6332);
   REGISTERS_reg_6_26_inst : DFF_X1 port map( D => n3586, CK => Clk, Q => 
                           net644861, QN => n6331);
   REGISTERS_reg_6_25_inst : DFF_X1 port map( D => n3585, CK => Clk, Q => 
                           net644860, QN => n6330);
   REGISTERS_reg_6_24_inst : DFF_X1 port map( D => n3584, CK => Clk, Q => 
                           net644859, QN => n6329);
   REGISTERS_reg_6_23_inst : DFF_X1 port map( D => n3583, CK => Clk, Q => 
                           net644858, QN => n6328);
   REGISTERS_reg_6_22_inst : DFF_X1 port map( D => n3582, CK => Clk, Q => 
                           net644857, QN => n6327);
   REGISTERS_reg_6_21_inst : DFF_X1 port map( D => n3581, CK => Clk, Q => 
                           net644856, QN => n6326);
   REGISTERS_reg_6_20_inst : DFF_X1 port map( D => n3580, CK => Clk, Q => 
                           net644855, QN => n6325);
   REGISTERS_reg_6_19_inst : DFF_X1 port map( D => n3579, CK => Clk, Q => 
                           net644854, QN => n6324);
   REGISTERS_reg_6_18_inst : DFF_X1 port map( D => n3578, CK => Clk, Q => 
                           net644853, QN => n6323);
   REGISTERS_reg_6_17_inst : DFF_X1 port map( D => n3577, CK => Clk, Q => 
                           net644852, QN => n6322);
   REGISTERS_reg_6_16_inst : DFF_X1 port map( D => n3576, CK => Clk, Q => 
                           net644851, QN => n6321);
   REGISTERS_reg_6_15_inst : DFF_X1 port map( D => n3575, CK => Clk, Q => 
                           net644850, QN => n6320);
   REGISTERS_reg_6_14_inst : DFF_X1 port map( D => n3574, CK => Clk, Q => 
                           net644849, QN => n6319);
   REGISTERS_reg_6_13_inst : DFF_X1 port map( D => n3573, CK => Clk, Q => 
                           net644848, QN => n6318);
   REGISTERS_reg_6_12_inst : DFF_X1 port map( D => n3572, CK => Clk, Q => 
                           net644847, QN => n6317);
   REGISTERS_reg_6_11_inst : DFF_X1 port map( D => n3571, CK => Clk, Q => 
                           net644846, QN => n6316);
   REGISTERS_reg_6_10_inst : DFF_X1 port map( D => n3570, CK => Clk, Q => 
                           net644845, QN => n6315);
   REGISTERS_reg_6_9_inst : DFF_X1 port map( D => n3569, CK => Clk, Q => 
                           net644844, QN => n6314);
   REGISTERS_reg_6_8_inst : DFF_X1 port map( D => n3568, CK => Clk, Q => 
                           net644843, QN => n6313);
   REGISTERS_reg_6_7_inst : DFF_X1 port map( D => n3567, CK => Clk, Q => 
                           net644842, QN => n6312);
   REGISTERS_reg_6_6_inst : DFF_X1 port map( D => n3566, CK => Clk, Q => 
                           net644841, QN => n6311);
   REGISTERS_reg_6_5_inst : DFF_X1 port map( D => n3565, CK => Clk, Q => 
                           net644840, QN => n6310);
   REGISTERS_reg_6_4_inst : DFF_X1 port map( D => n3564, CK => Clk, Q => 
                           net644839, QN => n6309);
   REGISTERS_reg_6_3_inst : DFF_X1 port map( D => n3563, CK => Clk, Q => 
                           net644838, QN => n6308);
   REGISTERS_reg_6_2_inst : DFF_X1 port map( D => n3562, CK => Clk, Q => 
                           net644837, QN => n6307);
   REGISTERS_reg_6_1_inst : DFF_X1 port map( D => n3561, CK => Clk, Q => 
                           net644836, QN => n6306);
   REGISTERS_reg_6_0_inst : DFF_X1 port map( D => n3560, CK => Clk, Q => n4059,
                           QN => n480);
   REGISTERS_reg_7_31_inst : DFF_X1 port map( D => n3559, CK => Clk, Q => 
                           net684296, QN => n608);
   REGISTERS_reg_7_30_inst : DFF_X1 port map( D => n3558, CK => Clk, Q => 
                           net684295, QN => n609);
   REGISTERS_reg_7_29_inst : DFF_X1 port map( D => n3557, CK => Clk, Q => 
                           net684294, QN => n610);
   REGISTERS_reg_7_28_inst : DFF_X1 port map( D => n3556, CK => Clk, Q => 
                           net684293, QN => n611);
   REGISTERS_reg_7_27_inst : DFF_X1 port map( D => n3555, CK => Clk, Q => 
                           net684292, QN => n612);
   REGISTERS_reg_7_26_inst : DFF_X1 port map( D => n3554, CK => Clk, Q => 
                           net684291, QN => n613);
   REGISTERS_reg_7_25_inst : DFF_X1 port map( D => n3553, CK => Clk, Q => 
                           net684290, QN => n614);
   REGISTERS_reg_7_24_inst : DFF_X1 port map( D => n3552, CK => Clk, Q => 
                           net684289, QN => n615);
   REGISTERS_reg_7_23_inst : DFF_X1 port map( D => n3551, CK => Clk, Q => 
                           net684288, QN => n616);
   REGISTERS_reg_7_22_inst : DFF_X1 port map( D => n3550, CK => Clk, Q => 
                           net684287, QN => n617);
   REGISTERS_reg_7_21_inst : DFF_X1 port map( D => n3549, CK => Clk, Q => 
                           net684286, QN => n618);
   REGISTERS_reg_7_20_inst : DFF_X1 port map( D => n3548, CK => Clk, Q => 
                           net684285, QN => n619);
   REGISTERS_reg_7_19_inst : DFF_X1 port map( D => n3547, CK => Clk, Q => 
                           net684284, QN => n620);
   REGISTERS_reg_7_18_inst : DFF_X1 port map( D => n3546, CK => Clk, Q => 
                           net684283, QN => n621);
   REGISTERS_reg_7_17_inst : DFF_X1 port map( D => n3545, CK => Clk, Q => 
                           net684282, QN => n622);
   REGISTERS_reg_7_16_inst : DFF_X1 port map( D => n3544, CK => Clk, Q => 
                           net684281, QN => n623);
   REGISTERS_reg_7_15_inst : DFF_X1 port map( D => n3543, CK => Clk, Q => 
                           net684280, QN => n624);
   REGISTERS_reg_7_14_inst : DFF_X1 port map( D => n3542, CK => Clk, Q => 
                           net684279, QN => n625);
   REGISTERS_reg_7_13_inst : DFF_X1 port map( D => n3541, CK => Clk, Q => 
                           net684278, QN => n626);
   REGISTERS_reg_7_12_inst : DFF_X1 port map( D => n3540, CK => Clk, Q => 
                           net684277, QN => n627);
   REGISTERS_reg_7_11_inst : DFF_X1 port map( D => n3539, CK => Clk, Q => 
                           net684276, QN => n628);
   REGISTERS_reg_7_10_inst : DFF_X1 port map( D => n3538, CK => Clk, Q => 
                           net684275, QN => n629);
   REGISTERS_reg_7_9_inst : DFF_X1 port map( D => n3537, CK => Clk, Q => 
                           net684274, QN => n630);
   REGISTERS_reg_7_8_inst : DFF_X1 port map( D => n3536, CK => Clk, Q => 
                           net684273, QN => n631);
   REGISTERS_reg_7_7_inst : DFF_X1 port map( D => n3535, CK => Clk, Q => 
                           net684272, QN => n632);
   REGISTERS_reg_7_6_inst : DFF_X1 port map( D => n3534, CK => Clk, Q => 
                           net684271, QN => n633);
   REGISTERS_reg_7_5_inst : DFF_X1 port map( D => n3533, CK => Clk, Q => 
                           net684270, QN => n634);
   REGISTERS_reg_7_4_inst : DFF_X1 port map( D => n3532, CK => Clk, Q => 
                           net684269, QN => n635);
   REGISTERS_reg_7_3_inst : DFF_X1 port map( D => n3531, CK => Clk, Q => 
                           net684268, QN => n636);
   REGISTERS_reg_7_2_inst : DFF_X1 port map( D => n3530, CK => Clk, Q => 
                           net684267, QN => n637);
   REGISTERS_reg_7_1_inst : DFF_X1 port map( D => n3529, CK => Clk, Q => 
                           net684266, QN => n638);
   REGISTERS_reg_7_0_inst : DFF_X1 port map( D => n3528, CK => Clk, Q => 
                           net644835, QN => n6343);
   REGISTERS_reg_8_31_inst : DFF_X1 port map( D => n3527, CK => Clk, Q => n4165
                           , QN => n2664);
   REGISTERS_reg_8_30_inst : DFF_X1 port map( D => n3526, CK => Clk, Q => n4162
                           , QN => n2663);
   REGISTERS_reg_8_29_inst : DFF_X1 port map( D => n3525, CK => Clk, Q => n4159
                           , QN => n2662);
   REGISTERS_reg_8_28_inst : DFF_X1 port map( D => n3524, CK => Clk, Q => n4156
                           , QN => n2661);
   REGISTERS_reg_8_27_inst : DFF_X1 port map( D => n3523, CK => Clk, Q => n4153
                           , QN => n2660);
   REGISTERS_reg_8_26_inst : DFF_X1 port map( D => n3522, CK => Clk, Q => n4150
                           , QN => n2659);
   REGISTERS_reg_8_25_inst : DFF_X1 port map( D => n3521, CK => Clk, Q => n4147
                           , QN => n2658);
   REGISTERS_reg_8_24_inst : DFF_X1 port map( D => n3520, CK => Clk, Q => n4141
                           , QN => n2657);
   REGISTERS_reg_8_23_inst : DFF_X1 port map( D => n3519, CK => Clk, Q => n4138
                           , QN => n2656);
   REGISTERS_reg_8_22_inst : DFF_X1 port map( D => n3518, CK => Clk, Q => n4135
                           , QN => n2655);
   REGISTERS_reg_8_21_inst : DFF_X1 port map( D => n3517, CK => Clk, Q => n4132
                           , QN => n2654);
   REGISTERS_reg_8_20_inst : DFF_X1 port map( D => n3516, CK => Clk, Q => n4129
                           , QN => n2653);
   REGISTERS_reg_8_19_inst : DFF_X1 port map( D => n3515, CK => Clk, Q => n4126
                           , QN => n2652);
   REGISTERS_reg_8_18_inst : DFF_X1 port map( D => n3514, CK => Clk, Q => n4123
                           , QN => n2651);
   REGISTERS_reg_8_17_inst : DFF_X1 port map( D => n3513, CK => Clk, Q => n4120
                           , QN => n2650);
   REGISTERS_reg_8_16_inst : DFF_X1 port map( D => n3512, CK => Clk, Q => n4117
                           , QN => n2649);
   REGISTERS_reg_8_15_inst : DFF_X1 port map( D => n3511, CK => Clk, Q => n4114
                           , QN => n2648);
   REGISTERS_reg_8_14_inst : DFF_X1 port map( D => n3510, CK => Clk, Q => n4109
                           , QN => n2647);
   REGISTERS_reg_8_13_inst : DFF_X1 port map( D => n3509, CK => Clk, Q => n4103
                           , QN => n2646);
   REGISTERS_reg_8_12_inst : DFF_X1 port map( D => n3508, CK => Clk, Q => n4100
                           , QN => n2645);
   REGISTERS_reg_8_11_inst : DFF_X1 port map( D => n3507, CK => Clk, Q => n4097
                           , QN => n2644);
   REGISTERS_reg_8_10_inst : DFF_X1 port map( D => n3506, CK => Clk, Q => n4094
                           , QN => n2643);
   REGISTERS_reg_8_9_inst : DFF_X1 port map( D => n3505, CK => Clk, Q => n4091,
                           QN => n2642);
   REGISTERS_reg_8_8_inst : DFF_X1 port map( D => n3504, CK => Clk, Q => n4088,
                           QN => n2641);
   REGISTERS_reg_8_7_inst : DFF_X1 port map( D => n3503, CK => Clk, Q => n4085,
                           QN => n2640);
   REGISTERS_reg_8_6_inst : DFF_X1 port map( D => n3502, CK => Clk, Q => n4082,
                           QN => n2639);
   REGISTERS_reg_8_5_inst : DFF_X1 port map( D => n3501, CK => Clk, Q => n4079,
                           QN => n2638);
   REGISTERS_reg_8_4_inst : DFF_X1 port map( D => n3500, CK => Clk, Q => n4076,
                           QN => n2637);
   REGISTERS_reg_8_3_inst : DFF_X1 port map( D => n3499, CK => Clk, Q => n4071,
                           QN => n2636);
   REGISTERS_reg_8_2_inst : DFF_X1 port map( D => n3498, CK => Clk, Q => n4066,
                           QN => n2635);
   REGISTERS_reg_8_1_inst : DFF_X1 port map( D => n3497, CK => Clk, Q => n4063,
                           QN => n2634);
   REGISTERS_reg_8_0_inst : DFF_X1 port map( D => n3496, CK => Clk, Q => n384, 
                           QN => n4169);
   REGISTERS_reg_9_31_inst : DFF_X1 port map( D => n3495, CK => Clk, Q => n389,
                           QN => n5993);
   REGISTERS_reg_9_30_inst : DFF_X1 port map( D => n3494, CK => Clk, Q => n392,
                           QN => n5992);
   REGISTERS_reg_9_29_inst : DFF_X1 port map( D => n3493, CK => Clk, Q => n395,
                           QN => n5991);
   REGISTERS_reg_9_28_inst : DFF_X1 port map( D => n3492, CK => Clk, Q => n398,
                           QN => n5990);
   REGISTERS_reg_9_27_inst : DFF_X1 port map( D => n3491, CK => Clk, Q => n401,
                           QN => n5989);
   REGISTERS_reg_9_26_inst : DFF_X1 port map( D => n3490, CK => Clk, Q => n404,
                           QN => n5988);
   REGISTERS_reg_9_25_inst : DFF_X1 port map( D => n3489, CK => Clk, Q => n407,
                           QN => n5987);
   REGISTERS_reg_9_24_inst : DFF_X1 port map( D => n3488, CK => Clk, Q => n410,
                           QN => n5986);
   REGISTERS_reg_9_23_inst : DFF_X1 port map( D => n3487, CK => Clk, Q => n413,
                           QN => n5985);
   REGISTERS_reg_9_22_inst : DFF_X1 port map( D => n3486, CK => Clk, Q => n416,
                           QN => n5970);
   REGISTERS_reg_9_21_inst : DFF_X1 port map( D => n3485, CK => Clk, Q => n419,
                           QN => n5965);
   REGISTERS_reg_9_20_inst : DFF_X1 port map( D => n3484, CK => Clk, Q => n422,
                           QN => n5933);
   REGISTERS_reg_9_19_inst : DFF_X1 port map( D => n3483, CK => Clk, Q => n425,
                           QN => n5252);
   REGISTERS_reg_9_18_inst : DFF_X1 port map( D => n3482, CK => Clk, Q => n428,
                           QN => n5218);
   REGISTERS_reg_9_17_inst : DFF_X1 port map( D => n3481, CK => Clk, Q => n431,
                           QN => n5204);
   REGISTERS_reg_9_16_inst : DFF_X1 port map( D => n3480, CK => Clk, Q => n434,
                           QN => n5203);
   REGISTERS_reg_9_15_inst : DFF_X1 port map( D => n3479, CK => Clk, Q => n437,
                           QN => n5193);
   REGISTERS_reg_9_14_inst : DFF_X1 port map( D => n3478, CK => Clk, Q => n440,
                           QN => n5188);
   REGISTERS_reg_9_13_inst : DFF_X1 port map( D => n3477, CK => Clk, Q => n443,
                           QN => n5183);
   REGISTERS_reg_9_12_inst : DFF_X1 port map( D => n3476, CK => Clk, Q => n446,
                           QN => n5180);
   REGISTERS_reg_9_11_inst : DFF_X1 port map( D => n3475, CK => Clk, Q => n449,
                           QN => n5174);
   REGISTERS_reg_9_10_inst : DFF_X1 port map( D => n3474, CK => Clk, Q => n452,
                           QN => n5153);
   REGISTERS_reg_9_9_inst : DFF_X1 port map( D => n3473, CK => Clk, Q => n455, 
                           QN => n5145);
   REGISTERS_reg_9_8_inst : DFF_X1 port map( D => n3472, CK => Clk, Q => n458, 
                           QN => n5144);
   REGISTERS_reg_9_7_inst : DFF_X1 port map( D => n3471, CK => Clk, Q => n461, 
                           QN => n5139);
   REGISTERS_reg_9_6_inst : DFF_X1 port map( D => n3470, CK => Clk, Q => n464, 
                           QN => n5134);
   REGISTERS_reg_9_5_inst : DFF_X1 port map( D => n3469, CK => Clk, Q => n467, 
                           QN => n5133);
   REGISTERS_reg_9_4_inst : DFF_X1 port map( D => n3468, CK => Clk, Q => n470, 
                           QN => n5123);
   REGISTERS_reg_9_3_inst : DFF_X1 port map( D => n3467, CK => Clk, Q => n473, 
                           QN => n5115);
   REGISTERS_reg_9_2_inst : DFF_X1 port map( D => n3466, CK => Clk, Q => n476, 
                           QN => n5114);
   REGISTERS_reg_9_1_inst : DFF_X1 port map( D => n3465, CK => Clk, Q => n479, 
                           QN => n5113);
   REGISTERS_reg_9_0_inst : DFF_X1 port map( D => n3464, CK => Clk, Q => n4062,
                           QN => n2601);
   REGISTERS_reg_10_31_inst : DFF_X1 port map( D => n3463, CK => Clk, Q => 
                           net644834, QN => n5109);
   REGISTERS_reg_10_30_inst : DFF_X1 port map( D => n3462, CK => Clk, Q => 
                           net644833, QN => n5108);
   REGISTERS_reg_10_29_inst : DFF_X1 port map( D => n3461, CK => Clk, Q => 
                           net644832, QN => n5103);
   REGISTERS_reg_10_28_inst : DFF_X1 port map( D => n3460, CK => Clk, Q => 
                           net644831, QN => n5102);
   REGISTERS_reg_10_27_inst : DFF_X1 port map( D => n3459, CK => Clk, Q => 
                           net644830, QN => n5093);
   REGISTERS_reg_10_26_inst : DFF_X1 port map( D => n3458, CK => Clk, Q => 
                           net644829, QN => n5085);
   REGISTERS_reg_10_25_inst : DFF_X1 port map( D => n3457, CK => Clk, Q => 
                           net644828, QN => n5084);
   REGISTERS_reg_10_24_inst : DFF_X1 port map( D => n3456, CK => Clk, Q => 
                           net644827, QN => n5083);
   REGISTERS_reg_10_23_inst : DFF_X1 port map( D => n3455, CK => Clk, Q => 
                           net644826, QN => n5079);
   REGISTERS_reg_10_22_inst : DFF_X1 port map( D => n3454, CK => Clk, Q => 
                           net644825, QN => n5078);
   REGISTERS_reg_10_21_inst : DFF_X1 port map( D => n3453, CK => Clk, Q => 
                           net644824, QN => n5073);
   REGISTERS_reg_10_20_inst : DFF_X1 port map( D => n3452, CK => Clk, Q => 
                           net644823, QN => n5072);
   REGISTERS_reg_10_19_inst : DFF_X1 port map( D => n3451, CK => Clk, Q => 
                           net644822, QN => n5063);
   REGISTERS_reg_10_18_inst : DFF_X1 port map( D => n3450, CK => Clk, Q => 
                           net644821, QN => n5055);
   REGISTERS_reg_10_17_inst : DFF_X1 port map( D => n3449, CK => Clk, Q => 
                           net644820, QN => n5054);
   REGISTERS_reg_10_16_inst : DFF_X1 port map( D => n3448, CK => Clk, Q => 
                           net644819, QN => n5053);
   REGISTERS_reg_10_15_inst : DFF_X1 port map( D => n3447, CK => Clk, Q => 
                           net644818, QN => n5049);
   REGISTERS_reg_10_14_inst : DFF_X1 port map( D => n3446, CK => Clk, Q => 
                           net644817, QN => n5048);
   REGISTERS_reg_10_13_inst : DFF_X1 port map( D => n3445, CK => Clk, Q => 
                           net644816, QN => n5043);
   REGISTERS_reg_10_12_inst : DFF_X1 port map( D => n3444, CK => Clk, Q => 
                           net644815, QN => n5042);
   REGISTERS_reg_10_11_inst : DFF_X1 port map( D => n3443, CK => Clk, Q => 
                           net644814, QN => n5033);
   REGISTERS_reg_10_10_inst : DFF_X1 port map( D => n3442, CK => Clk, Q => 
                           net644813, QN => n5025);
   REGISTERS_reg_10_9_inst : DFF_X1 port map( D => n3441, CK => Clk, Q => 
                           net644812, QN => n5024);
   REGISTERS_reg_10_8_inst : DFF_X1 port map( D => n3440, CK => Clk, Q => 
                           net644811, QN => n5023);
   REGISTERS_reg_10_7_inst : DFF_X1 port map( D => n3439, CK => Clk, Q => 
                           net644810, QN => n5019);
   REGISTERS_reg_10_6_inst : DFF_X1 port map( D => n3438, CK => Clk, Q => 
                           net644809, QN => n5018);
   REGISTERS_reg_10_5_inst : DFF_X1 port map( D => n3437, CK => Clk, Q => 
                           net644808, QN => n5013);
   REGISTERS_reg_10_4_inst : DFF_X1 port map( D => n3436, CK => Clk, Q => 
                           net644807, QN => n5012);
   REGISTERS_reg_10_3_inst : DFF_X1 port map( D => n3435, CK => Clk, Q => 
                           net644806, QN => n5003);
   REGISTERS_reg_10_2_inst : DFF_X1 port map( D => n3434, CK => Clk, Q => 
                           net644805, QN => n4995);
   REGISTERS_reg_10_1_inst : DFF_X1 port map( D => n3433, CK => Clk, Q => 
                           net644804, QN => n4994);
   REGISTERS_reg_10_0_inst : DFF_X1 port map( D => n3432, CK => Clk, Q => 
                           net684265, QN => n481);
   REGISTERS_reg_11_31_inst : DFF_X1 port map( D => n3431, CK => Clk, Q => 
                           n4056, QN => n482);
   REGISTERS_reg_11_30_inst : DFF_X1 port map( D => n3430, CK => Clk, Q => 
                           n4053, QN => n483);
   REGISTERS_reg_11_29_inst : DFF_X1 port map( D => n3429, CK => Clk, Q => 
                           n4050, QN => n484);
   REGISTERS_reg_11_28_inst : DFF_X1 port map( D => n3428, CK => Clk, Q => 
                           n4047, QN => n485);
   REGISTERS_reg_11_27_inst : DFF_X1 port map( D => n3427, CK => Clk, Q => 
                           n4044, QN => n486);
   REGISTERS_reg_11_26_inst : DFF_X1 port map( D => n3426, CK => Clk, Q => 
                           n4041, QN => n487);
   REGISTERS_reg_11_25_inst : DFF_X1 port map( D => n3425, CK => Clk, Q => 
                           n4038, QN => n488);
   REGISTERS_reg_11_24_inst : DFF_X1 port map( D => n3424, CK => Clk, Q => 
                           n4032, QN => n489);
   REGISTERS_reg_11_23_inst : DFF_X1 port map( D => n3423, CK => Clk, Q => 
                           n4029, QN => n490);
   REGISTERS_reg_11_22_inst : DFF_X1 port map( D => n3422, CK => Clk, Q => 
                           n4026, QN => n491);
   REGISTERS_reg_11_21_inst : DFF_X1 port map( D => n3421, CK => Clk, Q => 
                           n4023, QN => n492);
   REGISTERS_reg_11_20_inst : DFF_X1 port map( D => n3420, CK => Clk, Q => 
                           n4020, QN => n493);
   REGISTERS_reg_11_19_inst : DFF_X1 port map( D => n3419, CK => Clk, Q => 
                           n4017, QN => n494);
   REGISTERS_reg_11_18_inst : DFF_X1 port map( D => n3418, CK => Clk, Q => 
                           n4014, QN => n495);
   REGISTERS_reg_11_17_inst : DFF_X1 port map( D => n3417, CK => Clk, Q => 
                           n4011, QN => n496);
   REGISTERS_reg_11_16_inst : DFF_X1 port map( D => n3416, CK => Clk, Q => 
                           n4008, QN => n497);
   REGISTERS_reg_11_15_inst : DFF_X1 port map( D => n3415, CK => Clk, Q => 
                           n4005, QN => n498);
   REGISTERS_reg_11_14_inst : DFF_X1 port map( D => n3414, CK => Clk, Q => 
                           n4002, QN => n499);
   REGISTERS_reg_11_13_inst : DFF_X1 port map( D => n3413, CK => Clk, Q => 
                           n3993, QN => n500);
   REGISTERS_reg_11_12_inst : DFF_X1 port map( D => n3412, CK => Clk, Q => 
                           n3990, QN => n501);
   REGISTERS_reg_11_11_inst : DFF_X1 port map( D => n3411, CK => Clk, Q => 
                           n3987, QN => n502);
   REGISTERS_reg_11_10_inst : DFF_X1 port map( D => n3410, CK => Clk, Q => 
                           n3984, QN => n503);
   REGISTERS_reg_11_9_inst : DFF_X1 port map( D => n3409, CK => Clk, Q => n3981
                           , QN => n504);
   REGISTERS_reg_11_8_inst : DFF_X1 port map( D => n3408, CK => Clk, Q => n3978
                           , QN => n505);
   REGISTERS_reg_11_7_inst : DFF_X1 port map( D => n3407, CK => Clk, Q => n3975
                           , QN => n506);
   REGISTERS_reg_11_6_inst : DFF_X1 port map( D => n3406, CK => Clk, Q => n3972
                           , QN => n507);
   REGISTERS_reg_11_5_inst : DFF_X1 port map( D => n3405, CK => Clk, Q => n3969
                           , QN => n508);
   REGISTERS_reg_11_4_inst : DFF_X1 port map( D => n3404, CK => Clk, Q => n3966
                           , QN => n509);
   REGISTERS_reg_11_3_inst : DFF_X1 port map( D => n3403, CK => Clk, Q => n3963
                           , QN => n510);
   REGISTERS_reg_11_2_inst : DFF_X1 port map( D => n3402, CK => Clk, Q => n3957
                           , QN => n511);
   REGISTERS_reg_11_1_inst : DFF_X1 port map( D => n3401, CK => Clk, Q => n3954
                           , QN => n512);
   REGISTERS_reg_11_0_inst : DFF_X1 port map( D => n3400, CK => Clk, Q => n3915
                           , QN => n639);
   REGISTERS_reg_12_31_inst : DFF_X1 port map( D => n3399, CK => Clk, Q => 
                           net644803, QN => n4993);
   REGISTERS_reg_12_30_inst : DFF_X1 port map( D => n3398, CK => Clk, Q => 
                           net644802, QN => n4989);
   REGISTERS_reg_12_29_inst : DFF_X1 port map( D => n3397, CK => Clk, Q => 
                           net644801, QN => n4988);
   REGISTERS_reg_12_28_inst : DFF_X1 port map( D => n3396, CK => Clk, Q => 
                           net644800, QN => n4983);
   REGISTERS_reg_12_27_inst : DFF_X1 port map( D => n3395, CK => Clk, Q => 
                           net644799, QN => n4982);
   REGISTERS_reg_12_26_inst : DFF_X1 port map( D => n3394, CK => Clk, Q => 
                           net644798, QN => n4973);
   REGISTERS_reg_12_25_inst : DFF_X1 port map( D => n3393, CK => Clk, Q => 
                           net644797, QN => n4965);
   REGISTERS_reg_12_24_inst : DFF_X1 port map( D => n3392, CK => Clk, Q => 
                           net644796, QN => n4964);
   REGISTERS_reg_12_23_inst : DFF_X1 port map( D => n3391, CK => Clk, Q => 
                           net644795, QN => n4963);
   REGISTERS_reg_12_22_inst : DFF_X1 port map( D => n3390, CK => Clk, Q => 
                           net644794, QN => n4959);
   REGISTERS_reg_12_21_inst : DFF_X1 port map( D => n3389, CK => Clk, Q => 
                           net644793, QN => n4958);
   REGISTERS_reg_12_20_inst : DFF_X1 port map( D => n3388, CK => Clk, Q => 
                           net644792, QN => n4953);
   REGISTERS_reg_12_19_inst : DFF_X1 port map( D => n3387, CK => Clk, Q => 
                           net644791, QN => n4952);
   REGISTERS_reg_12_18_inst : DFF_X1 port map( D => n3386, CK => Clk, Q => 
                           net644790, QN => n4943);
   REGISTERS_reg_12_17_inst : DFF_X1 port map( D => n3385, CK => Clk, Q => 
                           net644789, QN => n4935);
   REGISTERS_reg_12_16_inst : DFF_X1 port map( D => n3384, CK => Clk, Q => 
                           net644788, QN => n4934);
   REGISTERS_reg_12_15_inst : DFF_X1 port map( D => n3383, CK => Clk, Q => 
                           net644787, QN => n4933);
   REGISTERS_reg_12_14_inst : DFF_X1 port map( D => n3382, CK => Clk, Q => 
                           net644786, QN => n4929);
   REGISTERS_reg_12_13_inst : DFF_X1 port map( D => n3381, CK => Clk, Q => 
                           net644785, QN => n4928);
   REGISTERS_reg_12_12_inst : DFF_X1 port map( D => n3380, CK => Clk, Q => 
                           net644784, QN => n4923);
   REGISTERS_reg_12_11_inst : DFF_X1 port map( D => n3379, CK => Clk, Q => 
                           net644783, QN => n4922);
   REGISTERS_reg_12_10_inst : DFF_X1 port map( D => n3378, CK => Clk, Q => 
                           net644782, QN => n4913);
   REGISTERS_reg_12_9_inst : DFF_X1 port map( D => n3377, CK => Clk, Q => 
                           net644781, QN => n4905);
   REGISTERS_reg_12_8_inst : DFF_X1 port map( D => n3376, CK => Clk, Q => 
                           net644780, QN => n4904);
   REGISTERS_reg_12_7_inst : DFF_X1 port map( D => n3375, CK => Clk, Q => 
                           net644779, QN => n4903);
   REGISTERS_reg_12_6_inst : DFF_X1 port map( D => n3374, CK => Clk, Q => 
                           net644778, QN => n4899);
   REGISTERS_reg_12_5_inst : DFF_X1 port map( D => n3373, CK => Clk, Q => 
                           net644777, QN => n4898);
   REGISTERS_reg_12_4_inst : DFF_X1 port map( D => n3372, CK => Clk, Q => 
                           net644776, QN => n4893);
   REGISTERS_reg_12_3_inst : DFF_X1 port map( D => n3371, CK => Clk, Q => 
                           net644775, QN => n4892);
   REGISTERS_reg_12_2_inst : DFF_X1 port map( D => n3370, CK => Clk, Q => 
                           net644774, QN => n4883);
   REGISTERS_reg_12_1_inst : DFF_X1 port map( D => n3369, CK => Clk, Q => 
                           net644773, QN => n4875);
   REGISTERS_reg_12_0_inst : DFF_X1 port map( D => n3368, CK => Clk, Q => 
                           net644772, QN => n6342);
   REGISTERS_reg_13_31_inst : DFF_X1 port map( D => n3367, CK => Clk, Q => 
                           net644771, QN => n6305);
   REGISTERS_reg_13_30_inst : DFF_X1 port map( D => n3366, CK => Clk, Q => 
                           net644770, QN => n6304);
   REGISTERS_reg_13_29_inst : DFF_X1 port map( D => n3365, CK => Clk, Q => 
                           net644769, QN => n6303);
   REGISTERS_reg_13_28_inst : DFF_X1 port map( D => n3364, CK => Clk, Q => 
                           net644768, QN => n6302);
   REGISTERS_reg_13_27_inst : DFF_X1 port map( D => n3363, CK => Clk, Q => 
                           net644767, QN => n6301);
   REGISTERS_reg_13_26_inst : DFF_X1 port map( D => n3362, CK => Clk, Q => 
                           net644766, QN => n6300);
   REGISTERS_reg_13_25_inst : DFF_X1 port map( D => n3361, CK => Clk, Q => 
                           net644765, QN => n6299);
   REGISTERS_reg_13_24_inst : DFF_X1 port map( D => n3360, CK => Clk, Q => 
                           net644764, QN => n6298);
   REGISTERS_reg_13_23_inst : DFF_X1 port map( D => n3359, CK => Clk, Q => 
                           net644763, QN => n6297);
   REGISTERS_reg_13_22_inst : DFF_X1 port map( D => n3358, CK => Clk, Q => 
                           net644762, QN => n6296);
   REGISTERS_reg_13_21_inst : DFF_X1 port map( D => n3357, CK => Clk, Q => 
                           net644761, QN => n6295);
   REGISTERS_reg_13_20_inst : DFF_X1 port map( D => n3356, CK => Clk, Q => 
                           net644760, QN => n6294);
   REGISTERS_reg_13_19_inst : DFF_X1 port map( D => n3355, CK => Clk, Q => 
                           net644759, QN => n6293);
   REGISTERS_reg_13_18_inst : DFF_X1 port map( D => n3354, CK => Clk, Q => 
                           net644758, QN => n6292);
   REGISTERS_reg_13_17_inst : DFF_X1 port map( D => n3353, CK => Clk, Q => 
                           net644757, QN => n6291);
   REGISTERS_reg_13_16_inst : DFF_X1 port map( D => n3352, CK => Clk, Q => 
                           net644756, QN => n6290);
   REGISTERS_reg_13_15_inst : DFF_X1 port map( D => n3351, CK => Clk, Q => 
                           net644755, QN => n6289);
   REGISTERS_reg_13_14_inst : DFF_X1 port map( D => n3350, CK => Clk, Q => 
                           net644754, QN => n6288);
   REGISTERS_reg_13_13_inst : DFF_X1 port map( D => n3349, CK => Clk, Q => 
                           net644753, QN => n6287);
   REGISTERS_reg_13_12_inst : DFF_X1 port map( D => n3348, CK => Clk, Q => 
                           net644752, QN => n6286);
   REGISTERS_reg_13_11_inst : DFF_X1 port map( D => n3347, CK => Clk, Q => 
                           net644751, QN => n6285);
   REGISTERS_reg_13_10_inst : DFF_X1 port map( D => n3346, CK => Clk, Q => 
                           net644750, QN => n6284);
   REGISTERS_reg_13_9_inst : DFF_X1 port map( D => n3345, CK => Clk, Q => 
                           net644749, QN => n6283);
   REGISTERS_reg_13_8_inst : DFF_X1 port map( D => n3344, CK => Clk, Q => 
                           net644748, QN => n6282);
   REGISTERS_reg_13_7_inst : DFF_X1 port map( D => n3343, CK => Clk, Q => 
                           net644747, QN => n6281);
   REGISTERS_reg_13_6_inst : DFF_X1 port map( D => n3342, CK => Clk, Q => 
                           net644746, QN => n6280);
   REGISTERS_reg_13_5_inst : DFF_X1 port map( D => n3341, CK => Clk, Q => 
                           net644745, QN => n6279);
   REGISTERS_reg_13_4_inst : DFF_X1 port map( D => n3340, CK => Clk, Q => 
                           net644744, QN => n6278);
   REGISTERS_reg_13_3_inst : DFF_X1 port map( D => n3339, CK => Clk, Q => 
                           net644743, QN => n6277);
   REGISTERS_reg_13_2_inst : DFF_X1 port map( D => n3338, CK => Clk, Q => 
                           net644742, QN => n6276);
   REGISTERS_reg_13_1_inst : DFF_X1 port map( D => n3337, CK => Clk, Q => 
                           net644741, QN => n6275);
   REGISTERS_reg_13_0_inst : DFF_X1 port map( D => n3336, CK => Clk, Q => 
                           net644740, QN => n6352);
   REGISTERS_reg_14_31_inst : DFF_X1 port map( D => n3335, CK => Clk, Q => 
                           net644739, QN => n6118);
   REGISTERS_reg_14_30_inst : DFF_X1 port map( D => n3334, CK => Clk, Q => 
                           net644738, QN => n6117);
   REGISTERS_reg_14_29_inst : DFF_X1 port map( D => n3333, CK => Clk, Q => 
                           net644737, QN => n6116);
   REGISTERS_reg_14_28_inst : DFF_X1 port map( D => n3332, CK => Clk, Q => 
                           net644736, QN => n6115);
   REGISTERS_reg_14_27_inst : DFF_X1 port map( D => n3331, CK => Clk, Q => 
                           net644735, QN => n6114);
   REGISTERS_reg_14_26_inst : DFF_X1 port map( D => n3330, CK => Clk, Q => 
                           net644734, QN => n6113);
   REGISTERS_reg_14_25_inst : DFF_X1 port map( D => n3329, CK => Clk, Q => 
                           net644733, QN => n6112);
   REGISTERS_reg_14_24_inst : DFF_X1 port map( D => n3328, CK => Clk, Q => 
                           net644732, QN => n6111);
   REGISTERS_reg_14_23_inst : DFF_X1 port map( D => n3327, CK => Clk, Q => 
                           net644731, QN => n6110);
   REGISTERS_reg_14_22_inst : DFF_X1 port map( D => n3326, CK => Clk, Q => 
                           net644730, QN => n6109);
   REGISTERS_reg_14_21_inst : DFF_X1 port map( D => n3325, CK => Clk, Q => 
                           net644729, QN => n6108);
   REGISTERS_reg_14_20_inst : DFF_X1 port map( D => n3324, CK => Clk, Q => 
                           net644728, QN => n6107);
   REGISTERS_reg_14_19_inst : DFF_X1 port map( D => n3323, CK => Clk, Q => 
                           net644727, QN => n6106);
   REGISTERS_reg_14_18_inst : DFF_X1 port map( D => n3322, CK => Clk, Q => 
                           net644726, QN => n6105);
   REGISTERS_reg_14_17_inst : DFF_X1 port map( D => n3321, CK => Clk, Q => 
                           net644725, QN => n6104);
   REGISTERS_reg_14_16_inst : DFF_X1 port map( D => n3320, CK => Clk, Q => 
                           net644724, QN => n6103);
   REGISTERS_reg_14_15_inst : DFF_X1 port map( D => n3319, CK => Clk, Q => 
                           net644723, QN => n6102);
   REGISTERS_reg_14_14_inst : DFF_X1 port map( D => n3318, CK => Clk, Q => 
                           net644722, QN => n6101);
   REGISTERS_reg_14_13_inst : DFF_X1 port map( D => n3317, CK => Clk, Q => 
                           net644721, QN => n6100);
   REGISTERS_reg_14_12_inst : DFF_X1 port map( D => n3316, CK => Clk, Q => 
                           net644720, QN => n6099);
   REGISTERS_reg_14_11_inst : DFF_X1 port map( D => n3315, CK => Clk, Q => 
                           net644719, QN => n6098);
   REGISTERS_reg_14_10_inst : DFF_X1 port map( D => n3314, CK => Clk, Q => 
                           net644718, QN => n6097);
   REGISTERS_reg_14_9_inst : DFF_X1 port map( D => n3313, CK => Clk, Q => 
                           net644717, QN => n6096);
   REGISTERS_reg_14_8_inst : DFF_X1 port map( D => n3312, CK => Clk, Q => 
                           net644716, QN => n6095);
   REGISTERS_reg_14_7_inst : DFF_X1 port map( D => n3311, CK => Clk, Q => 
                           net644715, QN => n6094);
   REGISTERS_reg_14_6_inst : DFF_X1 port map( D => n3310, CK => Clk, Q => 
                           net644714, QN => n6093);
   REGISTERS_reg_14_5_inst : DFF_X1 port map( D => n3309, CK => Clk, Q => 
                           net644713, QN => n6092);
   REGISTERS_reg_14_4_inst : DFF_X1 port map( D => n3308, CK => Clk, Q => 
                           net644712, QN => n6091);
   REGISTERS_reg_14_3_inst : DFF_X1 port map( D => n3307, CK => Clk, Q => 
                           net644711, QN => n6090);
   REGISTERS_reg_14_2_inst : DFF_X1 port map( D => n3306, CK => Clk, Q => 
                           net644710, QN => n6089);
   REGISTERS_reg_14_1_inst : DFF_X1 port map( D => n3305, CK => Clk, Q => 
                           net644709, QN => n6088);
   REGISTERS_reg_14_0_inst : DFF_X1 port map( D => n3304, CK => Clk, Q => 
                           net644708, QN => n6087);
   REGISTERS_reg_15_31_inst : DFF_X1 port map( D => n3303, CK => Clk, Q => 
                           n4057, QN => n704);
   REGISTERS_reg_15_30_inst : DFF_X1 port map( D => n3302, CK => Clk, Q => 
                           n4054, QN => n705);
   REGISTERS_reg_15_29_inst : DFF_X1 port map( D => n3301, CK => Clk, Q => 
                           n4051, QN => n706);
   REGISTERS_reg_15_28_inst : DFF_X1 port map( D => n3300, CK => Clk, Q => 
                           n4048, QN => n707);
   REGISTERS_reg_15_27_inst : DFF_X1 port map( D => n3299, CK => Clk, Q => 
                           n4045, QN => n708);
   REGISTERS_reg_15_26_inst : DFF_X1 port map( D => n3298, CK => Clk, Q => 
                           n4042, QN => n709);
   REGISTERS_reg_15_25_inst : DFF_X1 port map( D => n3297, CK => Clk, Q => 
                           n4039, QN => n710);
   REGISTERS_reg_15_24_inst : DFF_X1 port map( D => n3296, CK => Clk, Q => 
                           n4034, QN => n711);
   REGISTERS_reg_15_23_inst : DFF_X1 port map( D => n3295, CK => Clk, Q => 
                           n4030, QN => n712);
   REGISTERS_reg_15_22_inst : DFF_X1 port map( D => n3294, CK => Clk, Q => 
                           n4027, QN => n713);
   REGISTERS_reg_15_21_inst : DFF_X1 port map( D => n3293, CK => Clk, Q => 
                           n4024, QN => n714);
   REGISTERS_reg_15_20_inst : DFF_X1 port map( D => n3292, CK => Clk, Q => 
                           n4021, QN => n715);
   REGISTERS_reg_15_19_inst : DFF_X1 port map( D => n3291, CK => Clk, Q => 
                           n4018, QN => n716);
   REGISTERS_reg_15_18_inst : DFF_X1 port map( D => n3290, CK => Clk, Q => 
                           n4015, QN => n717);
   REGISTERS_reg_15_17_inst : DFF_X1 port map( D => n3289, CK => Clk, Q => 
                           n4012, QN => n718);
   REGISTERS_reg_15_16_inst : DFF_X1 port map( D => n3288, CK => Clk, Q => 
                           n4009, QN => n719);
   REGISTERS_reg_15_15_inst : DFF_X1 port map( D => n3287, CK => Clk, Q => 
                           n4006, QN => n720);
   REGISTERS_reg_15_14_inst : DFF_X1 port map( D => n3286, CK => Clk, Q => 
                           n4003, QN => n721);
   REGISTERS_reg_15_13_inst : DFF_X1 port map( D => n3285, CK => Clk, Q => 
                           n3998, QN => n722);
   REGISTERS_reg_15_12_inst : DFF_X1 port map( D => n3284, CK => Clk, Q => 
                           n3991, QN => n723);
   REGISTERS_reg_15_11_inst : DFF_X1 port map( D => n3283, CK => Clk, Q => 
                           n3988, QN => n724);
   REGISTERS_reg_15_10_inst : DFF_X1 port map( D => n3282, CK => Clk, Q => 
                           n3985, QN => n725);
   REGISTERS_reg_15_9_inst : DFF_X1 port map( D => n3281, CK => Clk, Q => n3982
                           , QN => n726);
   REGISTERS_reg_15_8_inst : DFF_X1 port map( D => n3280, CK => Clk, Q => n3979
                           , QN => n727);
   REGISTERS_reg_15_7_inst : DFF_X1 port map( D => n3279, CK => Clk, Q => n3976
                           , QN => n728);
   REGISTERS_reg_15_6_inst : DFF_X1 port map( D => n3278, CK => Clk, Q => n3973
                           , QN => n729);
   REGISTERS_reg_15_5_inst : DFF_X1 port map( D => n3277, CK => Clk, Q => n3970
                           , QN => n730);
   REGISTERS_reg_15_4_inst : DFF_X1 port map( D => n3276, CK => Clk, Q => n3967
                           , QN => n731);
   REGISTERS_reg_15_3_inst : DFF_X1 port map( D => n3275, CK => Clk, Q => n3964
                           , QN => n732);
   REGISTERS_reg_15_2_inst : DFF_X1 port map( D => n3274, CK => Clk, Q => n3958
                           , QN => n733);
   REGISTERS_reg_15_1_inst : DFF_X1 port map( D => n3273, CK => Clk, Q => n3955
                           , QN => n734);
   REGISTERS_reg_15_0_inst : DFF_X1 port map( D => n3272, CK => Clk, Q => n4061
                           , QN => n513);
   REGISTERS_reg_16_31_inst : DFF_X1 port map( D => n3271, CK => Clk, Q => 
                           net644707, QN => n6274);
   REGISTERS_reg_16_30_inst : DFF_X1 port map( D => n3270, CK => Clk, Q => 
                           net644706, QN => n6273);
   REGISTERS_reg_16_29_inst : DFF_X1 port map( D => n3269, CK => Clk, Q => 
                           net644705, QN => n6272);
   REGISTERS_reg_16_28_inst : DFF_X1 port map( D => n3268, CK => Clk, Q => 
                           net644704, QN => n6271);
   REGISTERS_reg_16_27_inst : DFF_X1 port map( D => n3267, CK => Clk, Q => 
                           net644703, QN => n6270);
   REGISTERS_reg_16_26_inst : DFF_X1 port map( D => n3266, CK => Clk, Q => 
                           net644702, QN => n6269);
   REGISTERS_reg_16_25_inst : DFF_X1 port map( D => n3265, CK => Clk, Q => 
                           net644701, QN => n6268);
   REGISTERS_reg_16_24_inst : DFF_X1 port map( D => n3264, CK => Clk, Q => 
                           net644700, QN => n6267);
   REGISTERS_reg_16_23_inst : DFF_X1 port map( D => n3263, CK => Clk, Q => 
                           net644699, QN => n6266);
   REGISTERS_reg_16_22_inst : DFF_X1 port map( D => n3262, CK => Clk, Q => 
                           net644698, QN => n6265);
   REGISTERS_reg_16_21_inst : DFF_X1 port map( D => n3261, CK => Clk, Q => 
                           net644697, QN => n6264);
   REGISTERS_reg_16_20_inst : DFF_X1 port map( D => n3260, CK => Clk, Q => 
                           net644696, QN => n6263);
   REGISTERS_reg_16_19_inst : DFF_X1 port map( D => n3259, CK => Clk, Q => 
                           net644695, QN => n6262);
   REGISTERS_reg_16_18_inst : DFF_X1 port map( D => n3258, CK => Clk, Q => 
                           net644694, QN => n6261);
   REGISTERS_reg_16_17_inst : DFF_X1 port map( D => n3257, CK => Clk, Q => 
                           net644693, QN => n6260);
   REGISTERS_reg_16_16_inst : DFF_X1 port map( D => n3256, CK => Clk, Q => 
                           net644692, QN => n6259);
   REGISTERS_reg_16_15_inst : DFF_X1 port map( D => n3255, CK => Clk, Q => 
                           net644691, QN => n6258);
   REGISTERS_reg_16_14_inst : DFF_X1 port map( D => n3254, CK => Clk, Q => 
                           net644690, QN => n6257);
   REGISTERS_reg_16_13_inst : DFF_X1 port map( D => n3253, CK => Clk, Q => 
                           net644689, QN => n6256);
   REGISTERS_reg_16_12_inst : DFF_X1 port map( D => n3252, CK => Clk, Q => 
                           net644688, QN => n6255);
   REGISTERS_reg_16_11_inst : DFF_X1 port map( D => n3251, CK => Clk, Q => 
                           net644687, QN => n6254);
   REGISTERS_reg_16_10_inst : DFF_X1 port map( D => n3250, CK => Clk, Q => 
                           net644686, QN => n6253);
   REGISTERS_reg_16_9_inst : DFF_X1 port map( D => n3249, CK => Clk, Q => 
                           net644685, QN => n6252);
   REGISTERS_reg_16_8_inst : DFF_X1 port map( D => n3248, CK => Clk, Q => 
                           net644684, QN => n6251);
   REGISTERS_reg_16_7_inst : DFF_X1 port map( D => n3247, CK => Clk, Q => 
                           net644683, QN => n6250);
   REGISTERS_reg_16_6_inst : DFF_X1 port map( D => n3246, CK => Clk, Q => 
                           net644682, QN => n6249);
   REGISTERS_reg_16_5_inst : DFF_X1 port map( D => n3245, CK => Clk, Q => 
                           net644681, QN => n6248);
   REGISTERS_reg_16_4_inst : DFF_X1 port map( D => n3244, CK => Clk, Q => 
                           net644680, QN => n6247);
   REGISTERS_reg_16_3_inst : DFF_X1 port map( D => n3243, CK => Clk, Q => 
                           net644679, QN => n6246);
   REGISTERS_reg_16_2_inst : DFF_X1 port map( D => n3242, CK => Clk, Q => 
                           net644678, QN => n6245);
   REGISTERS_reg_16_1_inst : DFF_X1 port map( D => n3241, CK => Clk, Q => 
                           net644677, QN => n6244);
   REGISTERS_reg_16_0_inst : DFF_X1 port map( D => n3240, CK => Clk, Q => 
                           net644676, QN => n6351);
   REGISTERS_reg_17_31_inst : DFF_X1 port map( D => n3239, CK => Clk, Q => n353
                           , QN => n4298);
   REGISTERS_reg_17_30_inst : DFF_X1 port map( D => n3238, CK => Clk, Q => n354
                           , QN => n4293);
   REGISTERS_reg_17_29_inst : DFF_X1 port map( D => n3237, CK => Clk, Q => n355
                           , QN => n4292);
   REGISTERS_reg_17_28_inst : DFF_X1 port map( D => n3236, CK => Clk, Q => n356
                           , QN => n4283);
   REGISTERS_reg_17_27_inst : DFF_X1 port map( D => n3235, CK => Clk, Q => n357
                           , QN => n4275);
   REGISTERS_reg_17_26_inst : DFF_X1 port map( D => n3234, CK => Clk, Q => n358
                           , QN => n4274);
   REGISTERS_reg_17_25_inst : DFF_X1 port map( D => n3233, CK => Clk, Q => n359
                           , QN => n4273);
   REGISTERS_reg_17_24_inst : DFF_X1 port map( D => n3232, CK => Clk, Q => n360
                           , QN => n4269);
   REGISTERS_reg_17_23_inst : DFF_X1 port map( D => n3231, CK => Clk, Q => n361
                           , QN => n4268);
   REGISTERS_reg_17_22_inst : DFF_X1 port map( D => n3230, CK => Clk, Q => n362
                           , QN => n4263);
   REGISTERS_reg_17_21_inst : DFF_X1 port map( D => n3229, CK => Clk, Q => n363
                           , QN => n4262);
   REGISTERS_reg_17_20_inst : DFF_X1 port map( D => n3228, CK => Clk, Q => n364
                           , QN => n4253);
   REGISTERS_reg_17_19_inst : DFF_X1 port map( D => n3227, CK => Clk, Q => n365
                           , QN => n4245);
   REGISTERS_reg_17_18_inst : DFF_X1 port map( D => n3226, CK => Clk, Q => n366
                           , QN => n4244);
   REGISTERS_reg_17_17_inst : DFF_X1 port map( D => n3225, CK => Clk, Q => n367
                           , QN => n4242);
   REGISTERS_reg_17_16_inst : DFF_X1 port map( D => n3224, CK => Clk, Q => n368
                           , QN => n4230);
   REGISTERS_reg_17_15_inst : DFF_X1 port map( D => n3223, CK => Clk, Q => n369
                           , QN => n4227);
   REGISTERS_reg_17_14_inst : DFF_X1 port map( D => n3222, CK => Clk, Q => n370
                           , QN => n4222);
   REGISTERS_reg_17_13_inst : DFF_X1 port map( D => n3221, CK => Clk, Q => n371
                           , QN => n4213);
   REGISTERS_reg_17_12_inst : DFF_X1 port map( D => n3220, CK => Clk, Q => n372
                           , QN => n4206);
   REGISTERS_reg_17_11_inst : DFF_X1 port map( D => n3219, CK => Clk, Q => n373
                           , QN => n4193);
   REGISTERS_reg_17_10_inst : DFF_X1 port map( D => n3218, CK => Clk, Q => n374
                           , QN => n4191);
   REGISTERS_reg_17_9_inst : DFF_X1 port map( D => n3217, CK => Clk, Q => n375,
                           QN => n4179);
   REGISTERS_reg_17_8_inst : DFF_X1 port map( D => n3216, CK => Clk, Q => n376,
                           QN => n4177);
   REGISTERS_reg_17_7_inst : DFF_X1 port map( D => n3215, CK => Clk, Q => n377,
                           QN => n4176);
   REGISTERS_reg_17_6_inst : DFF_X1 port map( D => n3214, CK => Clk, Q => n378,
                           QN => n4175);
   REGISTERS_reg_17_5_inst : DFF_X1 port map( D => n3213, CK => Clk, Q => n379,
                           QN => n4174);
   REGISTERS_reg_17_4_inst : DFF_X1 port map( D => n3212, CK => Clk, Q => n380,
                           QN => n4173);
   REGISTERS_reg_17_3_inst : DFF_X1 port map( D => n3211, CK => Clk, Q => n381,
                           QN => n4172);
   REGISTERS_reg_17_2_inst : DFF_X1 port map( D => n3210, CK => Clk, Q => n382,
                           QN => n4171);
   REGISTERS_reg_17_1_inst : DFF_X1 port map( D => n3209, CK => Clk, Q => n383,
                           QN => n4170);
   REGISTERS_reg_17_0_inst : DFF_X1 port map( D => n3208, CK => Clk, Q => n386,
                           QN => n4168);
   REGISTERS_reg_18_31_inst : DFF_X1 port map( D => n3207, CK => Clk, Q => 
                           net684264, QN => n640);
   REGISTERS_reg_18_30_inst : DFF_X1 port map( D => n3206, CK => Clk, Q => 
                           net684263, QN => n641);
   REGISTERS_reg_18_29_inst : DFF_X1 port map( D => n3205, CK => Clk, Q => 
                           net684262, QN => n642);
   REGISTERS_reg_18_28_inst : DFF_X1 port map( D => n3204, CK => Clk, Q => 
                           net684261, QN => n643);
   REGISTERS_reg_18_27_inst : DFF_X1 port map( D => n3203, CK => Clk, Q => 
                           net684260, QN => n644);
   REGISTERS_reg_18_26_inst : DFF_X1 port map( D => n3202, CK => Clk, Q => 
                           net684259, QN => n645);
   REGISTERS_reg_18_25_inst : DFF_X1 port map( D => n3201, CK => Clk, Q => 
                           net684258, QN => n646);
   REGISTERS_reg_18_24_inst : DFF_X1 port map( D => n3200, CK => Clk, Q => 
                           net684257, QN => n647);
   REGISTERS_reg_18_23_inst : DFF_X1 port map( D => n3199, CK => Clk, Q => 
                           net684256, QN => n648);
   REGISTERS_reg_18_22_inst : DFF_X1 port map( D => n3198, CK => Clk, Q => 
                           net684255, QN => n649);
   REGISTERS_reg_18_21_inst : DFF_X1 port map( D => n3197, CK => Clk, Q => 
                           net684254, QN => n650);
   REGISTERS_reg_18_20_inst : DFF_X1 port map( D => n3196, CK => Clk, Q => 
                           net684253, QN => n651);
   REGISTERS_reg_18_19_inst : DFF_X1 port map( D => n3195, CK => Clk, Q => 
                           net684252, QN => n652);
   REGISTERS_reg_18_18_inst : DFF_X1 port map( D => n3194, CK => Clk, Q => 
                           net684251, QN => n653);
   REGISTERS_reg_18_17_inst : DFF_X1 port map( D => n3193, CK => Clk, Q => 
                           net684250, QN => n654);
   REGISTERS_reg_18_16_inst : DFF_X1 port map( D => n3192, CK => Clk, Q => 
                           net684249, QN => n655);
   REGISTERS_reg_18_15_inst : DFF_X1 port map( D => n3191, CK => Clk, Q => 
                           net684248, QN => n656);
   REGISTERS_reg_18_14_inst : DFF_X1 port map( D => n3190, CK => Clk, Q => 
                           net684247, QN => n657);
   REGISTERS_reg_18_13_inst : DFF_X1 port map( D => n3189, CK => Clk, Q => 
                           net684246, QN => n658);
   REGISTERS_reg_18_12_inst : DFF_X1 port map( D => n3188, CK => Clk, Q => 
                           net684245, QN => n659);
   REGISTERS_reg_18_11_inst : DFF_X1 port map( D => n3187, CK => Clk, Q => 
                           net684244, QN => n660);
   REGISTERS_reg_18_10_inst : DFF_X1 port map( D => n3186, CK => Clk, Q => 
                           net684243, QN => n661);
   REGISTERS_reg_18_9_inst : DFF_X1 port map( D => n3185, CK => Clk, Q => 
                           net684242, QN => n662);
   REGISTERS_reg_18_8_inst : DFF_X1 port map( D => n3184, CK => Clk, Q => 
                           net684241, QN => n663);
   REGISTERS_reg_18_7_inst : DFF_X1 port map( D => n3183, CK => Clk, Q => 
                           net684240, QN => n664);
   REGISTERS_reg_18_6_inst : DFF_X1 port map( D => n3182, CK => Clk, Q => 
                           net684239, QN => n665);
   REGISTERS_reg_18_5_inst : DFF_X1 port map( D => n3181, CK => Clk, Q => 
                           net684238, QN => n666);
   REGISTERS_reg_18_4_inst : DFF_X1 port map( D => n3180, CK => Clk, Q => 
                           net684237, QN => n667);
   REGISTERS_reg_18_3_inst : DFF_X1 port map( D => n3179, CK => Clk, Q => 
                           net684236, QN => n668);
   REGISTERS_reg_18_2_inst : DFF_X1 port map( D => n3178, CK => Clk, Q => 
                           net684235, QN => n669);
   REGISTERS_reg_18_1_inst : DFF_X1 port map( D => n3177, CK => Clk, Q => 
                           net684234, QN => n670);
   REGISTERS_reg_18_0_inst : DFF_X1 port map( D => n3176, CK => Clk, Q => 
                           net644675, QN => n6337);
   REGISTERS_reg_19_31_inst : DFF_X1 port map( D => n3175, CK => Clk, Q => 
                           net644674, QN => n6086);
   REGISTERS_reg_19_30_inst : DFF_X1 port map( D => n3174, CK => Clk, Q => 
                           net644673, QN => n6085);
   REGISTERS_reg_19_29_inst : DFF_X1 port map( D => n3173, CK => Clk, Q => 
                           net644672, QN => n6084);
   REGISTERS_reg_19_28_inst : DFF_X1 port map( D => n3172, CK => Clk, Q => 
                           net644671, QN => n6083);
   REGISTERS_reg_19_27_inst : DFF_X1 port map( D => n3171, CK => Clk, Q => 
                           net644670, QN => n6082);
   REGISTERS_reg_19_26_inst : DFF_X1 port map( D => n3170, CK => Clk, Q => 
                           net644669, QN => n6081);
   REGISTERS_reg_19_25_inst : DFF_X1 port map( D => n3169, CK => Clk, Q => 
                           net644668, QN => n6080);
   REGISTERS_reg_19_24_inst : DFF_X1 port map( D => n3168, CK => Clk, Q => 
                           net644667, QN => n6079);
   REGISTERS_reg_19_23_inst : DFF_X1 port map( D => n3167, CK => Clk, Q => 
                           net644666, QN => n6078);
   REGISTERS_reg_19_22_inst : DFF_X1 port map( D => n3166, CK => Clk, Q => 
                           net644665, QN => n6077);
   REGISTERS_reg_19_21_inst : DFF_X1 port map( D => n3165, CK => Clk, Q => 
                           net644664, QN => n6076);
   REGISTERS_reg_19_20_inst : DFF_X1 port map( D => n3164, CK => Clk, Q => 
                           net644663, QN => n6075);
   REGISTERS_reg_19_19_inst : DFF_X1 port map( D => n3163, CK => Clk, Q => 
                           net644662, QN => n6074);
   REGISTERS_reg_19_18_inst : DFF_X1 port map( D => n3162, CK => Clk, Q => 
                           net644661, QN => n6073);
   REGISTERS_reg_19_17_inst : DFF_X1 port map( D => n3161, CK => Clk, Q => 
                           net644660, QN => n6072);
   REGISTERS_reg_19_16_inst : DFF_X1 port map( D => n3160, CK => Clk, Q => 
                           net644659, QN => n6071);
   REGISTERS_reg_19_15_inst : DFF_X1 port map( D => n3159, CK => Clk, Q => 
                           net644658, QN => n6070);
   REGISTERS_reg_19_14_inst : DFF_X1 port map( D => n3158, CK => Clk, Q => 
                           net644657, QN => n6069);
   REGISTERS_reg_19_13_inst : DFF_X1 port map( D => n3157, CK => Clk, Q => 
                           net644656, QN => n6068);
   REGISTERS_reg_19_12_inst : DFF_X1 port map( D => n3156, CK => Clk, Q => 
                           net644655, QN => n6067);
   REGISTERS_reg_19_11_inst : DFF_X1 port map( D => n3155, CK => Clk, Q => 
                           net644654, QN => n6066);
   REGISTERS_reg_19_10_inst : DFF_X1 port map( D => n3154, CK => Clk, Q => 
                           net644653, QN => n6065);
   REGISTERS_reg_19_9_inst : DFF_X1 port map( D => n3153, CK => Clk, Q => 
                           net644652, QN => n6064);
   REGISTERS_reg_19_8_inst : DFF_X1 port map( D => n3152, CK => Clk, Q => 
                           net644651, QN => n6063);
   REGISTERS_reg_19_7_inst : DFF_X1 port map( D => n3151, CK => Clk, Q => 
                           net644650, QN => n6062);
   REGISTERS_reg_19_6_inst : DFF_X1 port map( D => n3150, CK => Clk, Q => 
                           net644649, QN => n6061);
   REGISTERS_reg_19_5_inst : DFF_X1 port map( D => n3149, CK => Clk, Q => 
                           net644648, QN => n6060);
   REGISTERS_reg_19_4_inst : DFF_X1 port map( D => n3148, CK => Clk, Q => 
                           net644647, QN => n6059);
   REGISTERS_reg_19_3_inst : DFF_X1 port map( D => n3147, CK => Clk, Q => 
                           net644646, QN => n6058);
   REGISTERS_reg_19_2_inst : DFF_X1 port map( D => n3146, CK => Clk, Q => 
                           net644645, QN => n6057);
   REGISTERS_reg_19_1_inst : DFF_X1 port map( D => n3145, CK => Clk, Q => 
                           net644644, QN => n6056);
   REGISTERS_reg_19_0_inst : DFF_X1 port map( D => n3144, CK => Clk, Q => 
                           net684233, QN => n514);
   REGISTERS_reg_20_31_inst : DFF_X1 port map( D => n3143, CK => Clk, Q => 
                           net644643, QN => n4874);
   REGISTERS_reg_20_30_inst : DFF_X1 port map( D => n3142, CK => Clk, Q => 
                           net644642, QN => n4873);
   REGISTERS_reg_20_29_inst : DFF_X1 port map( D => n3141, CK => Clk, Q => 
                           net644641, QN => n4869);
   REGISTERS_reg_20_28_inst : DFF_X1 port map( D => n3140, CK => Clk, Q => 
                           net644640, QN => n4868);
   REGISTERS_reg_20_27_inst : DFF_X1 port map( D => n3139, CK => Clk, Q => 
                           net644639, QN => n4863);
   REGISTERS_reg_20_26_inst : DFF_X1 port map( D => n3138, CK => Clk, Q => 
                           net644638, QN => n4862);
   REGISTERS_reg_20_25_inst : DFF_X1 port map( D => n3137, CK => Clk, Q => 
                           net644637, QN => n4853);
   REGISTERS_reg_20_24_inst : DFF_X1 port map( D => n3136, CK => Clk, Q => 
                           net644636, QN => n4845);
   REGISTERS_reg_20_23_inst : DFF_X1 port map( D => n3135, CK => Clk, Q => 
                           net644635, QN => n4844);
   REGISTERS_reg_20_22_inst : DFF_X1 port map( D => n3134, CK => Clk, Q => 
                           net644634, QN => n4843);
   REGISTERS_reg_20_21_inst : DFF_X1 port map( D => n3133, CK => Clk, Q => 
                           net644633, QN => n4839);
   REGISTERS_reg_20_20_inst : DFF_X1 port map( D => n3132, CK => Clk, Q => 
                           net644632, QN => n4838);
   REGISTERS_reg_20_19_inst : DFF_X1 port map( D => n3131, CK => Clk, Q => 
                           net644631, QN => n4833);
   REGISTERS_reg_20_18_inst : DFF_X1 port map( D => n3130, CK => Clk, Q => 
                           net644630, QN => n4832);
   REGISTERS_reg_20_17_inst : DFF_X1 port map( D => n3129, CK => Clk, Q => 
                           net644629, QN => n4823);
   REGISTERS_reg_20_16_inst : DFF_X1 port map( D => n3128, CK => Clk, Q => 
                           net644628, QN => n4815);
   REGISTERS_reg_20_15_inst : DFF_X1 port map( D => n3127, CK => Clk, Q => 
                           net644627, QN => n4814);
   REGISTERS_reg_20_14_inst : DFF_X1 port map( D => n3126, CK => Clk, Q => 
                           net644626, QN => n4813);
   REGISTERS_reg_20_13_inst : DFF_X1 port map( D => n3125, CK => Clk, Q => 
                           net644625, QN => n4809);
   REGISTERS_reg_20_12_inst : DFF_X1 port map( D => n3124, CK => Clk, Q => 
                           net644624, QN => n4808);
   REGISTERS_reg_20_11_inst : DFF_X1 port map( D => n3123, CK => Clk, Q => 
                           net644623, QN => n4803);
   REGISTERS_reg_20_10_inst : DFF_X1 port map( D => n3122, CK => Clk, Q => 
                           net644622, QN => n4802);
   REGISTERS_reg_20_9_inst : DFF_X1 port map( D => n3121, CK => Clk, Q => 
                           net644621, QN => n4793);
   REGISTERS_reg_20_8_inst : DFF_X1 port map( D => n3120, CK => Clk, Q => 
                           net644620, QN => n4785);
   REGISTERS_reg_20_7_inst : DFF_X1 port map( D => n3119, CK => Clk, Q => 
                           net644619, QN => n4784);
   REGISTERS_reg_20_6_inst : DFF_X1 port map( D => n3118, CK => Clk, Q => 
                           net644618, QN => n4783);
   REGISTERS_reg_20_5_inst : DFF_X1 port map( D => n3117, CK => Clk, Q => 
                           net644617, QN => n4779);
   REGISTERS_reg_20_4_inst : DFF_X1 port map( D => n3116, CK => Clk, Q => 
                           net644616, QN => n4778);
   REGISTERS_reg_20_3_inst : DFF_X1 port map( D => n3115, CK => Clk, Q => 
                           net644615, QN => n4773);
   REGISTERS_reg_20_2_inst : DFF_X1 port map( D => n3114, CK => Clk, Q => 
                           net644614, QN => n4772);
   REGISTERS_reg_20_1_inst : DFF_X1 port map( D => n3113, CK => Clk, Q => 
                           net644613, QN => n4763);
   REGISTERS_reg_20_0_inst : DFF_X1 port map( D => n3112, CK => Clk, Q => 
                           net644612, QN => n6341);
   REGISTERS_reg_21_31_inst : DFF_X1 port map( D => n3111, CK => Clk, Q => 
                           net644611, QN => n4755);
   REGISTERS_reg_21_30_inst : DFF_X1 port map( D => n3110, CK => Clk, Q => 
                           net644610, QN => n4754);
   REGISTERS_reg_21_29_inst : DFF_X1 port map( D => n3109, CK => Clk, Q => 
                           net644609, QN => n4753);
   REGISTERS_reg_21_28_inst : DFF_X1 port map( D => n3108, CK => Clk, Q => 
                           net644608, QN => n4749);
   REGISTERS_reg_21_27_inst : DFF_X1 port map( D => n3107, CK => Clk, Q => 
                           net644607, QN => n4748);
   REGISTERS_reg_21_26_inst : DFF_X1 port map( D => n3106, CK => Clk, Q => 
                           net644606, QN => n4743);
   REGISTERS_reg_21_25_inst : DFF_X1 port map( D => n3105, CK => Clk, Q => 
                           net644605, QN => n4742);
   REGISTERS_reg_21_24_inst : DFF_X1 port map( D => n3104, CK => Clk, Q => 
                           net644604, QN => n4733);
   REGISTERS_reg_21_23_inst : DFF_X1 port map( D => n3103, CK => Clk, Q => 
                           net644603, QN => n4725);
   REGISTERS_reg_21_22_inst : DFF_X1 port map( D => n3102, CK => Clk, Q => 
                           net644602, QN => n4724);
   REGISTERS_reg_21_21_inst : DFF_X1 port map( D => n3101, CK => Clk, Q => 
                           net644601, QN => n4723);
   REGISTERS_reg_21_20_inst : DFF_X1 port map( D => n3100, CK => Clk, Q => 
                           net644600, QN => n4719);
   REGISTERS_reg_21_19_inst : DFF_X1 port map( D => n3099, CK => Clk, Q => 
                           net644599, QN => n4718);
   REGISTERS_reg_21_18_inst : DFF_X1 port map( D => n3098, CK => Clk, Q => 
                           net644598, QN => n4713);
   REGISTERS_reg_21_17_inst : DFF_X1 port map( D => n3097, CK => Clk, Q => 
                           net644597, QN => n4712);
   REGISTERS_reg_21_16_inst : DFF_X1 port map( D => n3096, CK => Clk, Q => 
                           net644596, QN => n4703);
   REGISTERS_reg_21_15_inst : DFF_X1 port map( D => n3095, CK => Clk, Q => 
                           net644595, QN => n4695);
   REGISTERS_reg_21_14_inst : DFF_X1 port map( D => n3094, CK => Clk, Q => 
                           net644594, QN => n4694);
   REGISTERS_reg_21_13_inst : DFF_X1 port map( D => n3093, CK => Clk, Q => 
                           net644593, QN => n4693);
   REGISTERS_reg_21_12_inst : DFF_X1 port map( D => n3092, CK => Clk, Q => 
                           net644592, QN => n4689);
   REGISTERS_reg_21_11_inst : DFF_X1 port map( D => n3091, CK => Clk, Q => 
                           net644591, QN => n4688);
   REGISTERS_reg_21_10_inst : DFF_X1 port map( D => n3090, CK => Clk, Q => 
                           net644590, QN => n4683);
   REGISTERS_reg_21_9_inst : DFF_X1 port map( D => n3089, CK => Clk, Q => 
                           net644589, QN => n4682);
   REGISTERS_reg_21_8_inst : DFF_X1 port map( D => n3088, CK => Clk, Q => 
                           net644588, QN => n4673);
   REGISTERS_reg_21_7_inst : DFF_X1 port map( D => n3087, CK => Clk, Q => 
                           net644587, QN => n4665);
   REGISTERS_reg_21_6_inst : DFF_X1 port map( D => n3086, CK => Clk, Q => 
                           net644586, QN => n4664);
   REGISTERS_reg_21_5_inst : DFF_X1 port map( D => n3085, CK => Clk, Q => 
                           net644585, QN => n4663);
   REGISTERS_reg_21_4_inst : DFF_X1 port map( D => n3084, CK => Clk, Q => 
                           net644584, QN => n4659);
   REGISTERS_reg_21_3_inst : DFF_X1 port map( D => n3083, CK => Clk, Q => 
                           net644583, QN => n4658);
   REGISTERS_reg_21_2_inst : DFF_X1 port map( D => n3082, CK => Clk, Q => 
                           net644582, QN => n4653);
   REGISTERS_reg_21_1_inst : DFF_X1 port map( D => n3081, CK => Clk, Q => 
                           net644581, QN => n4652);
   REGISTERS_reg_21_0_inst : DFF_X1 port map( D => n3080, CK => Clk, Q => 
                           net644580, QN => n6340);
   REGISTERS_reg_22_31_inst : DFF_X1 port map( D => n3079, CK => Clk, Q => 
                           net684232, QN => n515);
   REGISTERS_reg_22_30_inst : DFF_X1 port map( D => n3078, CK => Clk, Q => 
                           net684231, QN => n516);
   REGISTERS_reg_22_29_inst : DFF_X1 port map( D => n3077, CK => Clk, Q => 
                           net684230, QN => n517);
   REGISTERS_reg_22_28_inst : DFF_X1 port map( D => n3076, CK => Clk, Q => 
                           net684229, QN => n518);
   REGISTERS_reg_22_27_inst : DFF_X1 port map( D => n3075, CK => Clk, Q => 
                           net684228, QN => n519);
   REGISTERS_reg_22_26_inst : DFF_X1 port map( D => n3074, CK => Clk, Q => 
                           net684227, QN => n520);
   REGISTERS_reg_22_25_inst : DFF_X1 port map( D => n3073, CK => Clk, Q => 
                           net684226, QN => n521);
   REGISTERS_reg_22_24_inst : DFF_X1 port map( D => n3072, CK => Clk, Q => 
                           net684225, QN => n522);
   REGISTERS_reg_22_23_inst : DFF_X1 port map( D => n3071, CK => Clk, Q => 
                           net684224, QN => n523);
   REGISTERS_reg_22_22_inst : DFF_X1 port map( D => n3070, CK => Clk, Q => 
                           net684223, QN => n524);
   REGISTERS_reg_22_21_inst : DFF_X1 port map( D => n3069, CK => Clk, Q => 
                           net684222, QN => n525);
   REGISTERS_reg_22_20_inst : DFF_X1 port map( D => n3068, CK => Clk, Q => 
                           net684221, QN => n526);
   REGISTERS_reg_22_19_inst : DFF_X1 port map( D => n3067, CK => Clk, Q => 
                           net684220, QN => n527);
   REGISTERS_reg_22_18_inst : DFF_X1 port map( D => n3066, CK => Clk, Q => 
                           net684219, QN => n528);
   REGISTERS_reg_22_17_inst : DFF_X1 port map( D => n3065, CK => Clk, Q => 
                           net684218, QN => n529);
   REGISTERS_reg_22_16_inst : DFF_X1 port map( D => n3064, CK => Clk, Q => 
                           net684217, QN => n530);
   REGISTERS_reg_22_15_inst : DFF_X1 port map( D => n3063, CK => Clk, Q => 
                           net684216, QN => n531);
   REGISTERS_reg_22_14_inst : DFF_X1 port map( D => n3062, CK => Clk, Q => 
                           net684215, QN => n532);
   REGISTERS_reg_22_13_inst : DFF_X1 port map( D => n3061, CK => Clk, Q => 
                           net684214, QN => n533);
   REGISTERS_reg_22_12_inst : DFF_X1 port map( D => n3060, CK => Clk, Q => 
                           net684213, QN => n534);
   REGISTERS_reg_22_11_inst : DFF_X1 port map( D => n3059, CK => Clk, Q => 
                           net684212, QN => n535);
   REGISTERS_reg_22_10_inst : DFF_X1 port map( D => n3058, CK => Clk, Q => 
                           net684211, QN => n536);
   REGISTERS_reg_22_9_inst : DFF_X1 port map( D => n3057, CK => Clk, Q => 
                           net684210, QN => n537);
   REGISTERS_reg_22_8_inst : DFF_X1 port map( D => n3056, CK => Clk, Q => 
                           net684209, QN => n538);
   REGISTERS_reg_22_7_inst : DFF_X1 port map( D => n3055, CK => Clk, Q => 
                           net684208, QN => n539);
   REGISTERS_reg_22_6_inst : DFF_X1 port map( D => n3054, CK => Clk, Q => 
                           net684207, QN => n540);
   REGISTERS_reg_22_5_inst : DFF_X1 port map( D => n3053, CK => Clk, Q => 
                           net684206, QN => n541);
   REGISTERS_reg_22_4_inst : DFF_X1 port map( D => n3052, CK => Clk, Q => 
                           net684205, QN => n542);
   REGISTERS_reg_22_3_inst : DFF_X1 port map( D => n3051, CK => Clk, Q => 
                           net684204, QN => n543);
   REGISTERS_reg_22_2_inst : DFF_X1 port map( D => n3050, CK => Clk, Q => 
                           net684203, QN => n544);
   REGISTERS_reg_22_1_inst : DFF_X1 port map( D => n3049, CK => Clk, Q => 
                           net684202, QN => n545);
   REGISTERS_reg_22_0_inst : DFF_X1 port map( D => n3048, CK => Clk, Q => 
                           net684201, QN => n671);
   REGISTERS_reg_23_31_inst : DFF_X1 port map( D => n3047, CK => Clk, Q => 
                           n4166, QN => n672);
   REGISTERS_reg_23_30_inst : DFF_X1 port map( D => n3046, CK => Clk, Q => 
                           n4163, QN => n673);
   REGISTERS_reg_23_29_inst : DFF_X1 port map( D => n3045, CK => Clk, Q => 
                           n4160, QN => n674);
   REGISTERS_reg_23_28_inst : DFF_X1 port map( D => n3044, CK => Clk, Q => 
                           n4157, QN => n675);
   REGISTERS_reg_23_27_inst : DFF_X1 port map( D => n3043, CK => Clk, Q => 
                           n4154, QN => n676);
   REGISTERS_reg_23_26_inst : DFF_X1 port map( D => n3042, CK => Clk, Q => 
                           n4151, QN => n677);
   REGISTERS_reg_23_25_inst : DFF_X1 port map( D => n3041, CK => Clk, Q => 
                           n4148, QN => n678);
   REGISTERS_reg_23_24_inst : DFF_X1 port map( D => n3040, CK => Clk, Q => 
                           n4142, QN => n679);
   REGISTERS_reg_23_23_inst : DFF_X1 port map( D => n3039, CK => Clk, Q => 
                           n4139, QN => n680);
   REGISTERS_reg_23_22_inst : DFF_X1 port map( D => n3038, CK => Clk, Q => 
                           n4136, QN => n681);
   REGISTERS_reg_23_21_inst : DFF_X1 port map( D => n3037, CK => Clk, Q => 
                           n4133, QN => n682);
   REGISTERS_reg_23_20_inst : DFF_X1 port map( D => n3036, CK => Clk, Q => 
                           n4130, QN => n683);
   REGISTERS_reg_23_19_inst : DFF_X1 port map( D => n3035, CK => Clk, Q => 
                           n4127, QN => n684);
   REGISTERS_reg_23_18_inst : DFF_X1 port map( D => n3034, CK => Clk, Q => 
                           n4124, QN => n685);
   REGISTERS_reg_23_17_inst : DFF_X1 port map( D => n3033, CK => Clk, Q => 
                           n4121, QN => n686);
   REGISTERS_reg_23_16_inst : DFF_X1 port map( D => n3032, CK => Clk, Q => 
                           n4118, QN => n687);
   REGISTERS_reg_23_15_inst : DFF_X1 port map( D => n3031, CK => Clk, Q => 
                           n4115, QN => n688);
   REGISTERS_reg_23_14_inst : DFF_X1 port map( D => n3030, CK => Clk, Q => 
                           n4112, QN => n689);
   REGISTERS_reg_23_13_inst : DFF_X1 port map( D => n3029, CK => Clk, Q => 
                           n4104, QN => n690);
   REGISTERS_reg_23_12_inst : DFF_X1 port map( D => n3028, CK => Clk, Q => 
                           n4101, QN => n691);
   REGISTERS_reg_23_11_inst : DFF_X1 port map( D => n3027, CK => Clk, Q => 
                           n4098, QN => n692);
   REGISTERS_reg_23_10_inst : DFF_X1 port map( D => n3026, CK => Clk, Q => 
                           n4095, QN => n693);
   REGISTERS_reg_23_9_inst : DFF_X1 port map( D => n3025, CK => Clk, Q => n4092
                           , QN => n694);
   REGISTERS_reg_23_8_inst : DFF_X1 port map( D => n3024, CK => Clk, Q => n4089
                           , QN => n695);
   REGISTERS_reg_23_7_inst : DFF_X1 port map( D => n3023, CK => Clk, Q => n4086
                           , QN => n696);
   REGISTERS_reg_23_6_inst : DFF_X1 port map( D => n3022, CK => Clk, Q => n4083
                           , QN => n697);
   REGISTERS_reg_23_5_inst : DFF_X1 port map( D => n3021, CK => Clk, Q => n4080
                           , QN => n698);
   REGISTERS_reg_23_4_inst : DFF_X1 port map( D => n3020, CK => Clk, Q => n4077
                           , QN => n699);
   REGISTERS_reg_23_3_inst : DFF_X1 port map( D => n3019, CK => Clk, Q => n4072
                           , QN => n700);
   REGISTERS_reg_23_2_inst : DFF_X1 port map( D => n3018, CK => Clk, Q => n4067
                           , QN => n701);
   REGISTERS_reg_23_1_inst : DFF_X1 port map( D => n3017, CK => Clk, Q => n4064
                           , QN => n702);
   REGISTERS_reg_23_0_inst : DFF_X1 port map( D => n3016, CK => Clk, Q => 
                           net644579, QN => n6350);
   REGISTERS_reg_24_31_inst : DFF_X1 port map( D => n3015, CK => Clk, Q => 
                           net644578, QN => n6149);
   REGISTERS_reg_24_30_inst : DFF_X1 port map( D => n3014, CK => Clk, Q => 
                           net644577, QN => n6148);
   REGISTERS_reg_24_29_inst : DFF_X1 port map( D => n3013, CK => Clk, Q => 
                           net644576, QN => n6147);
   REGISTERS_reg_24_28_inst : DFF_X1 port map( D => n3012, CK => Clk, Q => 
                           net644575, QN => n6146);
   REGISTERS_reg_24_27_inst : DFF_X1 port map( D => n3011, CK => Clk, Q => 
                           net644574, QN => n6145);
   REGISTERS_reg_24_26_inst : DFF_X1 port map( D => n3010, CK => Clk, Q => 
                           net644573, QN => n6144);
   REGISTERS_reg_24_25_inst : DFF_X1 port map( D => n3009, CK => Clk, Q => 
                           net644572, QN => n6143);
   REGISTERS_reg_24_24_inst : DFF_X1 port map( D => n3008, CK => Clk, Q => 
                           net644571, QN => n6142);
   REGISTERS_reg_24_23_inst : DFF_X1 port map( D => n3007, CK => Clk, Q => 
                           net644570, QN => n6141);
   REGISTERS_reg_24_22_inst : DFF_X1 port map( D => n3006, CK => Clk, Q => 
                           net644569, QN => n6140);
   REGISTERS_reg_24_21_inst : DFF_X1 port map( D => n3005, CK => Clk, Q => 
                           net644568, QN => n6139);
   REGISTERS_reg_24_20_inst : DFF_X1 port map( D => n3004, CK => Clk, Q => 
                           net644567, QN => n6138);
   REGISTERS_reg_24_19_inst : DFF_X1 port map( D => n3003, CK => Clk, Q => 
                           net644566, QN => n6137);
   REGISTERS_reg_24_18_inst : DFF_X1 port map( D => n3002, CK => Clk, Q => 
                           net644565, QN => n6136);
   REGISTERS_reg_24_17_inst : DFF_X1 port map( D => n3001, CK => Clk, Q => 
                           net644564, QN => n6135);
   REGISTERS_reg_24_16_inst : DFF_X1 port map( D => n3000, CK => Clk, Q => 
                           net644563, QN => n6134);
   REGISTERS_reg_24_15_inst : DFF_X1 port map( D => n2999, CK => Clk, Q => 
                           net644562, QN => n6133);
   REGISTERS_reg_24_14_inst : DFF_X1 port map( D => n2998, CK => Clk, Q => 
                           net644561, QN => n6132);
   REGISTERS_reg_24_13_inst : DFF_X1 port map( D => n2997, CK => Clk, Q => 
                           net644560, QN => n6131);
   REGISTERS_reg_24_12_inst : DFF_X1 port map( D => n2996, CK => Clk, Q => 
                           net644559, QN => n6130);
   REGISTERS_reg_24_11_inst : DFF_X1 port map( D => n2995, CK => Clk, Q => 
                           net644558, QN => n6129);
   REGISTERS_reg_24_10_inst : DFF_X1 port map( D => n2994, CK => Clk, Q => 
                           net644557, QN => n6128);
   REGISTERS_reg_24_9_inst : DFF_X1 port map( D => n2993, CK => Clk, Q => 
                           net644556, QN => n6127);
   REGISTERS_reg_24_8_inst : DFF_X1 port map( D => n2992, CK => Clk, Q => 
                           net644555, QN => n6126);
   REGISTERS_reg_24_7_inst : DFF_X1 port map( D => n2991, CK => Clk, Q => 
                           net644554, QN => n6125);
   REGISTERS_reg_24_6_inst : DFF_X1 port map( D => n2990, CK => Clk, Q => 
                           net644553, QN => n6124);
   REGISTERS_reg_24_5_inst : DFF_X1 port map( D => n2989, CK => Clk, Q => 
                           net644552, QN => n6123);
   REGISTERS_reg_24_4_inst : DFF_X1 port map( D => n2988, CK => Clk, Q => 
                           net644551, QN => n6122);
   REGISTERS_reg_24_3_inst : DFF_X1 port map( D => n2987, CK => Clk, Q => 
                           net644550, QN => n6121);
   REGISTERS_reg_24_2_inst : DFF_X1 port map( D => n2986, CK => Clk, Q => 
                           net644549, QN => n6120);
   REGISTERS_reg_24_1_inst : DFF_X1 port map( D => n2985, CK => Clk, Q => 
                           net644548, QN => n6119);
   REGISTERS_reg_24_0_inst : DFF_X1 port map( D => n2984, CK => Clk, Q => 
                           net644547, QN => n6349);
   REGISTERS_reg_25_31_inst : DFF_X1 port map( D => n2983, CK => Clk, Q => 
                           net644546, QN => n6180);
   REGISTERS_reg_25_30_inst : DFF_X1 port map( D => n2982, CK => Clk, Q => 
                           net644545, QN => n6179);
   REGISTERS_reg_25_29_inst : DFF_X1 port map( D => n2981, CK => Clk, Q => 
                           net644544, QN => n6178);
   REGISTERS_reg_25_28_inst : DFF_X1 port map( D => n2980, CK => Clk, Q => 
                           net644543, QN => n6177);
   REGISTERS_reg_25_27_inst : DFF_X1 port map( D => n2979, CK => Clk, Q => 
                           net644542, QN => n6176);
   REGISTERS_reg_25_26_inst : DFF_X1 port map( D => n2978, CK => Clk, Q => 
                           net644541, QN => n6175);
   REGISTERS_reg_25_25_inst : DFF_X1 port map( D => n2977, CK => Clk, Q => 
                           net644540, QN => n6174);
   REGISTERS_reg_25_24_inst : DFF_X1 port map( D => n2976, CK => Clk, Q => 
                           net644539, QN => n6173);
   REGISTERS_reg_25_23_inst : DFF_X1 port map( D => n2975, CK => Clk, Q => 
                           net644538, QN => n6172);
   REGISTERS_reg_25_22_inst : DFF_X1 port map( D => n2974, CK => Clk, Q => 
                           net644537, QN => n6171);
   REGISTERS_reg_25_21_inst : DFF_X1 port map( D => n2973, CK => Clk, Q => 
                           net644536, QN => n6170);
   REGISTERS_reg_25_20_inst : DFF_X1 port map( D => n2972, CK => Clk, Q => 
                           net644535, QN => n6169);
   REGISTERS_reg_25_19_inst : DFF_X1 port map( D => n2971, CK => Clk, Q => 
                           net644534, QN => n6168);
   REGISTERS_reg_25_18_inst : DFF_X1 port map( D => n2970, CK => Clk, Q => 
                           net644533, QN => n6167);
   REGISTERS_reg_25_17_inst : DFF_X1 port map( D => n2969, CK => Clk, Q => 
                           net644532, QN => n6166);
   REGISTERS_reg_25_16_inst : DFF_X1 port map( D => n2968, CK => Clk, Q => 
                           net644531, QN => n6165);
   REGISTERS_reg_25_15_inst : DFF_X1 port map( D => n2967, CK => Clk, Q => 
                           net644530, QN => n6164);
   REGISTERS_reg_25_14_inst : DFF_X1 port map( D => n2966, CK => Clk, Q => 
                           net644529, QN => n6163);
   REGISTERS_reg_25_13_inst : DFF_X1 port map( D => n2965, CK => Clk, Q => 
                           net644528, QN => n6162);
   REGISTERS_reg_25_12_inst : DFF_X1 port map( D => n2964, CK => Clk, Q => 
                           net644527, QN => n6161);
   REGISTERS_reg_25_11_inst : DFF_X1 port map( D => n2963, CK => Clk, Q => 
                           net644526, QN => n6160);
   REGISTERS_reg_25_10_inst : DFF_X1 port map( D => n2962, CK => Clk, Q => 
                           net644525, QN => n6159);
   REGISTERS_reg_25_9_inst : DFF_X1 port map( D => n2961, CK => Clk, Q => 
                           net644524, QN => n6158);
   REGISTERS_reg_25_8_inst : DFF_X1 port map( D => n2960, CK => Clk, Q => 
                           net644523, QN => n6157);
   REGISTERS_reg_25_7_inst : DFF_X1 port map( D => n2959, CK => Clk, Q => 
                           net644522, QN => n6156);
   REGISTERS_reg_25_6_inst : DFF_X1 port map( D => n2958, CK => Clk, Q => 
                           net644521, QN => n6155);
   REGISTERS_reg_25_5_inst : DFF_X1 port map( D => n2957, CK => Clk, Q => 
                           net644520, QN => n6154);
   REGISTERS_reg_25_4_inst : DFF_X1 port map( D => n2956, CK => Clk, Q => 
                           net644519, QN => n6153);
   REGISTERS_reg_25_3_inst : DFF_X1 port map( D => n2955, CK => Clk, Q => 
                           net644518, QN => n6152);
   REGISTERS_reg_25_2_inst : DFF_X1 port map( D => n2954, CK => Clk, Q => 
                           net644517, QN => n6151);
   REGISTERS_reg_25_1_inst : DFF_X1 port map( D => n2953, CK => Clk, Q => 
                           net644516, QN => n6150);
   REGISTERS_reg_25_0_inst : DFF_X1 port map( D => n2952, CK => Clk, Q => 
                           net644515, QN => n6339);
   REGISTERS_reg_26_31_inst : DFF_X1 port map( D => n2951, CK => Clk, Q => 
                           n4164, QN => n2248);
   REGISTERS_reg_26_30_inst : DFF_X1 port map( D => n2950, CK => Clk, Q => 
                           n4161, QN => n2247);
   REGISTERS_reg_26_29_inst : DFF_X1 port map( D => n2949, CK => Clk, Q => 
                           n4158, QN => n2246);
   REGISTERS_reg_26_28_inst : DFF_X1 port map( D => n2948, CK => Clk, Q => 
                           n4155, QN => n2245);
   REGISTERS_reg_26_27_inst : DFF_X1 port map( D => n2947, CK => Clk, Q => 
                           n4152, QN => n2244);
   REGISTERS_reg_26_26_inst : DFF_X1 port map( D => n2946, CK => Clk, Q => 
                           n4149, QN => n2243);
   REGISTERS_reg_26_25_inst : DFF_X1 port map( D => n2945, CK => Clk, Q => 
                           n4144, QN => n2242);
   REGISTERS_reg_26_24_inst : DFF_X1 port map( D => n2944, CK => Clk, Q => 
                           n4140, QN => n2241);
   REGISTERS_reg_26_23_inst : DFF_X1 port map( D => n2943, CK => Clk, Q => 
                           n4137, QN => n2240);
   REGISTERS_reg_26_22_inst : DFF_X1 port map( D => n2942, CK => Clk, Q => 
                           n4134, QN => n2239);
   REGISTERS_reg_26_21_inst : DFF_X1 port map( D => n2941, CK => Clk, Q => 
                           n4131, QN => n2238);
   REGISTERS_reg_26_20_inst : DFF_X1 port map( D => n2940, CK => Clk, Q => 
                           n4128, QN => n2237);
   REGISTERS_reg_26_19_inst : DFF_X1 port map( D => n2939, CK => Clk, Q => 
                           n4125, QN => n2236);
   REGISTERS_reg_26_18_inst : DFF_X1 port map( D => n2938, CK => Clk, Q => 
                           n4122, QN => n2235);
   REGISTERS_reg_26_17_inst : DFF_X1 port map( D => n2937, CK => Clk, Q => 
                           n4119, QN => n2234);
   REGISTERS_reg_26_16_inst : DFF_X1 port map( D => n2936, CK => Clk, Q => 
                           n4116, QN => n2233);
   REGISTERS_reg_26_15_inst : DFF_X1 port map( D => n2935, CK => Clk, Q => 
                           n4113, QN => n2232);
   REGISTERS_reg_26_14_inst : DFF_X1 port map( D => n2934, CK => Clk, Q => 
                           n4105, QN => n2231);
   REGISTERS_reg_26_13_inst : DFF_X1 port map( D => n2933, CK => Clk, Q => 
                           n4102, QN => n2230);
   REGISTERS_reg_26_12_inst : DFF_X1 port map( D => n2932, CK => Clk, Q => 
                           n4099, QN => n2229);
   REGISTERS_reg_26_11_inst : DFF_X1 port map( D => n2931, CK => Clk, Q => 
                           n4096, QN => n2228);
   REGISTERS_reg_26_10_inst : DFF_X1 port map( D => n2930, CK => Clk, Q => 
                           n4093, QN => n2227);
   REGISTERS_reg_26_9_inst : DFF_X1 port map( D => n2929, CK => Clk, Q => n4090
                           , QN => n2226);
   REGISTERS_reg_26_8_inst : DFF_X1 port map( D => n2928, CK => Clk, Q => n4087
                           , QN => n2225);
   REGISTERS_reg_26_7_inst : DFF_X1 port map( D => n2927, CK => Clk, Q => n4084
                           , QN => n2224);
   REGISTERS_reg_26_6_inst : DFF_X1 port map( D => n2926, CK => Clk, Q => n4081
                           , QN => n2223);
   REGISTERS_reg_26_5_inst : DFF_X1 port map( D => n2925, CK => Clk, Q => n4078
                           , QN => n2222);
   REGISTERS_reg_26_4_inst : DFF_X1 port map( D => n2924, CK => Clk, Q => n4075
                           , QN => n2221);
   REGISTERS_reg_26_3_inst : DFF_X1 port map( D => n2923, CK => Clk, Q => n4070
                           , QN => n2220);
   REGISTERS_reg_26_2_inst : DFF_X1 port map( D => n2922, CK => Clk, Q => n4065
                           , QN => n2219);
   REGISTERS_reg_26_1_inst : DFF_X1 port map( D => n2921, CK => Clk, Q => n222,
                           QN => n6243);
   REGISTERS_reg_26_0_inst : DFF_X1 port map( D => n2920, CK => Clk, Q => n385,
                           QN => n4167);
   REGISTERS_reg_27_31_inst : DFF_X1 port map( D => n2919, CK => Clk, Q => 
                           net644514, QN => n6242);
   REGISTERS_reg_27_30_inst : DFF_X1 port map( D => n2918, CK => Clk, Q => 
                           net644513, QN => n6241);
   REGISTERS_reg_27_29_inst : DFF_X1 port map( D => n2917, CK => Clk, Q => 
                           net644512, QN => n6240);
   REGISTERS_reg_27_28_inst : DFF_X1 port map( D => n2916, CK => Clk, Q => 
                           net644511, QN => n6239);
   REGISTERS_reg_27_27_inst : DFF_X1 port map( D => n2915, CK => Clk, Q => 
                           net644510, QN => n6238);
   REGISTERS_reg_27_26_inst : DFF_X1 port map( D => n2914, CK => Clk, Q => 
                           net644509, QN => n6237);
   REGISTERS_reg_27_25_inst : DFF_X1 port map( D => n2913, CK => Clk, Q => 
                           net644508, QN => n6236);
   REGISTERS_reg_27_24_inst : DFF_X1 port map( D => n2912, CK => Clk, Q => 
                           net644507, QN => n6235);
   REGISTERS_reg_27_23_inst : DFF_X1 port map( D => n2911, CK => Clk, Q => 
                           net644506, QN => n6234);
   REGISTERS_reg_27_22_inst : DFF_X1 port map( D => n2910, CK => Clk, Q => 
                           net644505, QN => n6233);
   REGISTERS_reg_27_21_inst : DFF_X1 port map( D => n2909, CK => Clk, Q => 
                           net644504, QN => n6232);
   REGISTERS_reg_27_20_inst : DFF_X1 port map( D => n2908, CK => Clk, Q => 
                           net644503, QN => n6231);
   REGISTERS_reg_27_19_inst : DFF_X1 port map( D => n2907, CK => Clk, Q => 
                           net644502, QN => n6230);
   REGISTERS_reg_27_18_inst : DFF_X1 port map( D => n2906, CK => Clk, Q => 
                           net644501, QN => n6229);
   REGISTERS_reg_27_17_inst : DFF_X1 port map( D => n2905, CK => Clk, Q => 
                           net644500, QN => n6228);
   REGISTERS_reg_27_16_inst : DFF_X1 port map( D => n2904, CK => Clk, Q => 
                           net644499, QN => n6227);
   REGISTERS_reg_27_15_inst : DFF_X1 port map( D => n2903, CK => Clk, Q => 
                           net644498, QN => n6226);
   REGISTERS_reg_27_14_inst : DFF_X1 port map( D => n2902, CK => Clk, Q => 
                           net644497, QN => n6225);
   REGISTERS_reg_27_13_inst : DFF_X1 port map( D => n2901, CK => Clk, Q => 
                           net644496, QN => n6224);
   REGISTERS_reg_27_12_inst : DFF_X1 port map( D => n2900, CK => Clk, Q => 
                           net644495, QN => n6223);
   REGISTERS_reg_27_11_inst : DFF_X1 port map( D => n2899, CK => Clk, Q => 
                           net644494, QN => n6222);
   REGISTERS_reg_27_10_inst : DFF_X1 port map( D => n2898, CK => Clk, Q => 
                           net644493, QN => n6221);
   REGISTERS_reg_27_9_inst : DFF_X1 port map( D => n2897, CK => Clk, Q => 
                           net644492, QN => n6220);
   REGISTERS_reg_27_8_inst : DFF_X1 port map( D => n2896, CK => Clk, Q => 
                           net644491, QN => n6219);
   REGISTERS_reg_27_7_inst : DFF_X1 port map( D => n2895, CK => Clk, Q => 
                           net644490, QN => n6218);
   REGISTERS_reg_27_6_inst : DFF_X1 port map( D => n2894, CK => Clk, Q => 
                           net644489, QN => n6217);
   REGISTERS_reg_27_5_inst : DFF_X1 port map( D => n2893, CK => Clk, Q => 
                           net644488, QN => n6216);
   REGISTERS_reg_27_4_inst : DFF_X1 port map( D => n2892, CK => Clk, Q => 
                           net644487, QN => n6215);
   REGISTERS_reg_27_3_inst : DFF_X1 port map( D => n2891, CK => Clk, Q => 
                           net644486, QN => n6214);
   REGISTERS_reg_27_2_inst : DFF_X1 port map( D => n2890, CK => Clk, Q => 
                           net644485, QN => n6213);
   REGISTERS_reg_27_1_inst : DFF_X1 port map( D => n2889, CK => Clk, Q => 
                           net644484, QN => n6212);
   REGISTERS_reg_27_0_inst : DFF_X1 port map( D => n2888, CK => Clk, Q => 
                           net644483, QN => n6348);
   REGISTERS_reg_28_31_inst : DFF_X1 port map( D => n2887, CK => Clk, Q => 
                           net684200, QN => n546);
   REGISTERS_reg_28_30_inst : DFF_X1 port map( D => n2886, CK => Clk, Q => 
                           net684199, QN => n547);
   REGISTERS_reg_28_29_inst : DFF_X1 port map( D => n2885, CK => Clk, Q => 
                           net684198, QN => n548);
   REGISTERS_reg_28_28_inst : DFF_X1 port map( D => n2884, CK => Clk, Q => 
                           net684197, QN => n549);
   REGISTERS_reg_28_27_inst : DFF_X1 port map( D => n2883, CK => Clk, Q => 
                           net684196, QN => n550);
   REGISTERS_reg_28_26_inst : DFF_X1 port map( D => n2882, CK => Clk, Q => 
                           net684195, QN => n551);
   REGISTERS_reg_28_25_inst : DFF_X1 port map( D => n2881, CK => Clk, Q => 
                           net684194, QN => n552);
   REGISTERS_reg_28_24_inst : DFF_X1 port map( D => n2880, CK => Clk, Q => 
                           net684193, QN => n553);
   REGISTERS_reg_28_23_inst : DFF_X1 port map( D => n2879, CK => Clk, Q => 
                           net684192, QN => n554);
   REGISTERS_reg_28_22_inst : DFF_X1 port map( D => n2878, CK => Clk, Q => 
                           net684191, QN => n555);
   REGISTERS_reg_28_21_inst : DFF_X1 port map( D => n2877, CK => Clk, Q => 
                           net684190, QN => n556);
   REGISTERS_reg_28_20_inst : DFF_X1 port map( D => n2876, CK => Clk, Q => 
                           net684189, QN => n557);
   REGISTERS_reg_28_19_inst : DFF_X1 port map( D => n2875, CK => Clk, Q => 
                           net684188, QN => n558);
   REGISTERS_reg_28_18_inst : DFF_X1 port map( D => n2874, CK => Clk, Q => 
                           net684187, QN => n559);
   REGISTERS_reg_28_17_inst : DFF_X1 port map( D => n2873, CK => Clk, Q => 
                           net684186, QN => n560);
   REGISTERS_reg_28_16_inst : DFF_X1 port map( D => n2872, CK => Clk, Q => 
                           net684185, QN => n561);
   REGISTERS_reg_28_15_inst : DFF_X1 port map( D => n2871, CK => Clk, Q => 
                           net684184, QN => n562);
   REGISTERS_reg_28_14_inst : DFF_X1 port map( D => n2870, CK => Clk, Q => 
                           net684183, QN => n563);
   REGISTERS_reg_28_13_inst : DFF_X1 port map( D => n2869, CK => Clk, Q => 
                           net684182, QN => n564);
   REGISTERS_reg_28_12_inst : DFF_X1 port map( D => n2868, CK => Clk, Q => 
                           net684181, QN => n565);
   REGISTERS_reg_28_11_inst : DFF_X1 port map( D => n2867, CK => Clk, Q => 
                           net684180, QN => n566);
   REGISTERS_reg_28_10_inst : DFF_X1 port map( D => n2866, CK => Clk, Q => 
                           net684179, QN => n567);
   REGISTERS_reg_28_9_inst : DFF_X1 port map( D => n2865, CK => Clk, Q => 
                           net684178, QN => n568);
   REGISTERS_reg_28_8_inst : DFF_X1 port map( D => n2864, CK => Clk, Q => 
                           net684177, QN => n569);
   REGISTERS_reg_28_7_inst : DFF_X1 port map( D => n2863, CK => Clk, Q => 
                           net684176, QN => n570);
   REGISTERS_reg_28_6_inst : DFF_X1 port map( D => n2862, CK => Clk, Q => 
                           net684175, QN => n571);
   REGISTERS_reg_28_5_inst : DFF_X1 port map( D => n2861, CK => Clk, Q => 
                           net684174, QN => n572);
   REGISTERS_reg_28_4_inst : DFF_X1 port map( D => n2860, CK => Clk, Q => 
                           net684173, QN => n573);
   REGISTERS_reg_28_3_inst : DFF_X1 port map( D => n2859, CK => Clk, Q => 
                           net684172, QN => n574);
   REGISTERS_reg_28_2_inst : DFF_X1 port map( D => n2858, CK => Clk, Q => 
                           net684171, QN => n575);
   REGISTERS_reg_28_1_inst : DFF_X1 port map( D => n2857, CK => Clk, Q => 
                           net684170, QN => n576);
   REGISTERS_reg_28_0_inst : DFF_X1 port map( D => n2856, CK => Clk, Q => 
                           net684169, QN => n703);
   REGISTERS_reg_29_31_inst : DFF_X1 port map( D => n2855, CK => Clk, Q => 
                           net644482, QN => n4643);
   REGISTERS_reg_29_30_inst : DFF_X1 port map( D => n2854, CK => Clk, Q => 
                           net644481, QN => n4635);
   REGISTERS_reg_29_29_inst : DFF_X1 port map( D => n2853, CK => Clk, Q => 
                           net644480, QN => n4634);
   REGISTERS_reg_29_28_inst : DFF_X1 port map( D => n2852, CK => Clk, Q => 
                           net644479, QN => n4633);
   REGISTERS_reg_29_27_inst : DFF_X1 port map( D => n2851, CK => Clk, Q => 
                           net644478, QN => n4629);
   REGISTERS_reg_29_26_inst : DFF_X1 port map( D => n2850, CK => Clk, Q => 
                           net644477, QN => n4628);
   REGISTERS_reg_29_25_inst : DFF_X1 port map( D => n2849, CK => Clk, Q => 
                           net644476, QN => n4623);
   REGISTERS_reg_29_24_inst : DFF_X1 port map( D => n2848, CK => Clk, Q => 
                           net644475, QN => n4622);
   REGISTERS_reg_29_23_inst : DFF_X1 port map( D => n2847, CK => Clk, Q => 
                           net644474, QN => n4613);
   REGISTERS_reg_29_22_inst : DFF_X1 port map( D => n2846, CK => Clk, Q => 
                           net644473, QN => n4605);
   REGISTERS_reg_29_21_inst : DFF_X1 port map( D => n2845, CK => Clk, Q => 
                           net644472, QN => n4604);
   REGISTERS_reg_29_20_inst : DFF_X1 port map( D => n2844, CK => Clk, Q => 
                           net644471, QN => n4603);
   REGISTERS_reg_29_19_inst : DFF_X1 port map( D => n2843, CK => Clk, Q => 
                           net644470, QN => n4599);
   REGISTERS_reg_29_18_inst : DFF_X1 port map( D => n2842, CK => Clk, Q => 
                           net644469, QN => n4598);
   REGISTERS_reg_29_17_inst : DFF_X1 port map( D => n2841, CK => Clk, Q => 
                           net644468, QN => n4593);
   REGISTERS_reg_29_16_inst : DFF_X1 port map( D => n2840, CK => Clk, Q => 
                           net644467, QN => n4592);
   REGISTERS_reg_29_15_inst : DFF_X1 port map( D => n2839, CK => Clk, Q => 
                           net644466, QN => n4583);
   REGISTERS_reg_29_14_inst : DFF_X1 port map( D => n2838, CK => Clk, Q => 
                           net644465, QN => n4575);
   REGISTERS_reg_29_13_inst : DFF_X1 port map( D => n2837, CK => Clk, Q => 
                           net644464, QN => n4574);
   REGISTERS_reg_29_12_inst : DFF_X1 port map( D => n2836, CK => Clk, Q => 
                           net644463, QN => n4573);
   REGISTERS_reg_29_11_inst : DFF_X1 port map( D => n2835, CK => Clk, Q => 
                           net644462, QN => n4569);
   REGISTERS_reg_29_10_inst : DFF_X1 port map( D => n2834, CK => Clk, Q => 
                           net644461, QN => n4568);
   REGISTERS_reg_29_9_inst : DFF_X1 port map( D => n2833, CK => Clk, Q => 
                           net644460, QN => n4563);
   REGISTERS_reg_29_8_inst : DFF_X1 port map( D => n2832, CK => Clk, Q => 
                           net644459, QN => n4562);
   REGISTERS_reg_29_7_inst : DFF_X1 port map( D => n2831, CK => Clk, Q => 
                           net644458, QN => n4553);
   REGISTERS_reg_29_6_inst : DFF_X1 port map( D => n2830, CK => Clk, Q => 
                           net644457, QN => n4545);
   REGISTERS_reg_29_5_inst : DFF_X1 port map( D => n2829, CK => Clk, Q => 
                           net644456, QN => n4544);
   REGISTERS_reg_29_4_inst : DFF_X1 port map( D => n2828, CK => Clk, Q => 
                           net644455, QN => n4543);
   REGISTERS_reg_29_3_inst : DFF_X1 port map( D => n2827, CK => Clk, Q => 
                           net644454, QN => n4539);
   REGISTERS_reg_29_2_inst : DFF_X1 port map( D => n2826, CK => Clk, Q => 
                           net644453, QN => n4538);
   REGISTERS_reg_29_1_inst : DFF_X1 port map( D => n2825, CK => Clk, Q => 
                           net644452, QN => n4533);
   REGISTERS_reg_29_0_inst : DFF_X1 port map( D => n2824, CK => Clk, Q => 
                           net644451, QN => n6338);
   REGISTERS_reg_30_31_inst : DFF_X1 port map( D => n2823, CK => Clk, Q => 
                           net644450, QN => n6211);
   REGISTERS_reg_30_30_inst : DFF_X1 port map( D => n2822, CK => Clk, Q => 
                           net644449, QN => n6210);
   REGISTERS_reg_30_29_inst : DFF_X1 port map( D => n2821, CK => Clk, Q => 
                           net644448, QN => n6209);
   REGISTERS_reg_30_28_inst : DFF_X1 port map( D => n2820, CK => Clk, Q => 
                           net644447, QN => n6208);
   REGISTERS_reg_30_27_inst : DFF_X1 port map( D => n2819, CK => Clk, Q => 
                           net644446, QN => n6207);
   REGISTERS_reg_30_26_inst : DFF_X1 port map( D => n2818, CK => Clk, Q => 
                           net644445, QN => n6206);
   REGISTERS_reg_30_25_inst : DFF_X1 port map( D => n2817, CK => Clk, Q => 
                           net644444, QN => n6205);
   REGISTERS_reg_30_24_inst : DFF_X1 port map( D => n2816, CK => Clk, Q => 
                           net644443, QN => n6204);
   REGISTERS_reg_30_23_inst : DFF_X1 port map( D => n2815, CK => Clk, Q => 
                           net644442, QN => n6203);
   REGISTERS_reg_30_22_inst : DFF_X1 port map( D => n2814, CK => Clk, Q => 
                           net644441, QN => n6202);
   REGISTERS_reg_30_21_inst : DFF_X1 port map( D => n2813, CK => Clk, Q => 
                           net644440, QN => n6201);
   REGISTERS_reg_30_20_inst : DFF_X1 port map( D => n2812, CK => Clk, Q => 
                           net644439, QN => n6200);
   REGISTERS_reg_30_19_inst : DFF_X1 port map( D => n2811, CK => Clk, Q => 
                           net644438, QN => n6199);
   REGISTERS_reg_30_18_inst : DFF_X1 port map( D => n2810, CK => Clk, Q => 
                           net644437, QN => n6198);
   REGISTERS_reg_30_17_inst : DFF_X1 port map( D => n2809, CK => Clk, Q => 
                           net644436, QN => n6197);
   REGISTERS_reg_30_16_inst : DFF_X1 port map( D => n2808, CK => Clk, Q => 
                           net644435, QN => n6196);
   REGISTERS_reg_30_15_inst : DFF_X1 port map( D => n2807, CK => Clk, Q => 
                           net644434, QN => n6195);
   REGISTERS_reg_30_14_inst : DFF_X1 port map( D => n2806, CK => Clk, Q => 
                           net644433, QN => n6194);
   REGISTERS_reg_30_13_inst : DFF_X1 port map( D => n2805, CK => Clk, Q => 
                           net644432, QN => n6193);
   REGISTERS_reg_30_12_inst : DFF_X1 port map( D => n2804, CK => Clk, Q => 
                           net644431, QN => n6192);
   REGISTERS_reg_30_11_inst : DFF_X1 port map( D => n2803, CK => Clk, Q => 
                           net644430, QN => n6191);
   REGISTERS_reg_30_10_inst : DFF_X1 port map( D => n2802, CK => Clk, Q => 
                           net644429, QN => n6190);
   REGISTERS_reg_30_9_inst : DFF_X1 port map( D => n2801, CK => Clk, Q => 
                           net644428, QN => n6189);
   REGISTERS_reg_30_8_inst : DFF_X1 port map( D => n2800, CK => Clk, Q => 
                           net644427, QN => n6188);
   REGISTERS_reg_30_7_inst : DFF_X1 port map( D => n2799, CK => Clk, Q => 
                           net644426, QN => n6187);
   REGISTERS_reg_30_6_inst : DFF_X1 port map( D => n2798, CK => Clk, Q => 
                           net644425, QN => n6186);
   REGISTERS_reg_30_5_inst : DFF_X1 port map( D => n2797, CK => Clk, Q => 
                           net644424, QN => n6185);
   REGISTERS_reg_30_4_inst : DFF_X1 port map( D => n2796, CK => Clk, Q => 
                           net644423, QN => n6184);
   REGISTERS_reg_30_3_inst : DFF_X1 port map( D => n2795, CK => Clk, Q => 
                           net644422, QN => n6183);
   REGISTERS_reg_30_2_inst : DFF_X1 port map( D => n2794, CK => Clk, Q => 
                           net644421, QN => n6182);
   REGISTERS_reg_30_1_inst : DFF_X1 port map( D => n2793, CK => Clk, Q => 
                           net644420, QN => n6181);
   REGISTERS_reg_30_0_inst : DFF_X1 port map( D => n2792, CK => Clk, Q => 
                           net644419, QN => n6347);
   REGISTERS_reg_31_31_inst : DFF_X1 port map( D => n2791, CK => Clk, Q => n387
                           , QN => n4532);
   OUT2_reg_31_inst : DFF_X1 port map( D => n2790, CK => Clk, Q => OUT2(31), QN
                           => net644418);
   REGISTERS_reg_31_30_inst : DFF_X1 port map( D => n2789, CK => Clk, Q => n390
                           , QN => n4523);
   OUT2_reg_30_inst : DFF_X1 port map( D => n2788, CK => Clk, Q => OUT2(30), QN
                           => net644417);
   REGISTERS_reg_31_29_inst : DFF_X1 port map( D => n2787, CK => Clk, Q => n393
                           , QN => n4515);
   OUT2_reg_29_inst : DFF_X1 port map( D => n2786, CK => Clk, Q => OUT2(29), QN
                           => net644416);
   REGISTERS_reg_31_28_inst : DFF_X1 port map( D => n2785, CK => Clk, Q => n396
                           , QN => n4514);
   OUT2_reg_28_inst : DFF_X1 port map( D => n2784, CK => Clk, Q => OUT2(28), QN
                           => net644415);
   REGISTERS_reg_31_27_inst : DFF_X1 port map( D => n2783, CK => Clk, Q => n399
                           , QN => n4513);
   OUT2_reg_27_inst : DFF_X1 port map( D => n2782, CK => Clk, Q => OUT2(27), QN
                           => net644414);
   REGISTERS_reg_31_26_inst : DFF_X1 port map( D => n2781, CK => Clk, Q => n402
                           , QN => n4509);
   OUT2_reg_26_inst : DFF_X1 port map( D => n2780, CK => Clk, Q => OUT2(26), QN
                           => net644413);
   REGISTERS_reg_31_25_inst : DFF_X1 port map( D => n2779, CK => Clk, Q => n405
                           , QN => n4508);
   OUT2_reg_25_inst : DFF_X1 port map( D => n2778, CK => Clk, Q => OUT2(25), QN
                           => net644412);
   REGISTERS_reg_31_24_inst : DFF_X1 port map( D => n2777, CK => Clk, Q => n408
                           , QN => n4503);
   OUT2_reg_24_inst : DFF_X1 port map( D => n2776, CK => Clk, Q => OUT2(24), QN
                           => net644411);
   REGISTERS_reg_31_23_inst : DFF_X1 port map( D => n2775, CK => Clk, Q => n411
                           , QN => n4502);
   OUT2_reg_23_inst : DFF_X1 port map( D => n2774, CK => Clk, Q => OUT2(23), QN
                           => net644410);
   REGISTERS_reg_31_22_inst : DFF_X1 port map( D => n2773, CK => Clk, Q => n414
                           , QN => n4493);
   OUT2_reg_22_inst : DFF_X1 port map( D => n2772, CK => Clk, Q => OUT2(22), QN
                           => net644409);
   REGISTERS_reg_31_21_inst : DFF_X1 port map( D => n2771, CK => Clk, Q => n417
                           , QN => n4485);
   OUT2_reg_21_inst : DFF_X1 port map( D => n2770, CK => Clk, Q => OUT2(21), QN
                           => net644408);
   REGISTERS_reg_31_20_inst : DFF_X1 port map( D => n2769, CK => Clk, Q => n420
                           , QN => n4484);
   OUT2_reg_20_inst : DFF_X1 port map( D => n2768, CK => Clk, Q => OUT2(20), QN
                           => net644407);
   REGISTERS_reg_31_19_inst : DFF_X1 port map( D => n2767, CK => Clk, Q => n423
                           , QN => n4483);
   OUT2_reg_19_inst : DFF_X1 port map( D => n2766, CK => Clk, Q => OUT2(19), QN
                           => net644406);
   REGISTERS_reg_31_18_inst : DFF_X1 port map( D => n2765, CK => Clk, Q => n426
                           , QN => n4479);
   OUT2_reg_18_inst : DFF_X1 port map( D => n2764, CK => Clk, Q => OUT2(18), QN
                           => net644405);
   REGISTERS_reg_31_17_inst : DFF_X1 port map( D => n2763, CK => Clk, Q => n429
                           , QN => n4478);
   OUT2_reg_17_inst : DFF_X1 port map( D => n2762, CK => Clk, Q => OUT2(17), QN
                           => net644404);
   REGISTERS_reg_31_16_inst : DFF_X1 port map( D => n2761, CK => Clk, Q => n432
                           , QN => n4473);
   OUT2_reg_16_inst : DFF_X1 port map( D => n2760, CK => Clk, Q => OUT2(16), QN
                           => net644403);
   REGISTERS_reg_31_15_inst : DFF_X1 port map( D => n2759, CK => Clk, Q => n435
                           , QN => n4472);
   OUT2_reg_15_inst : DFF_X1 port map( D => n2758, CK => Clk, Q => OUT2(15), QN
                           => net644402);
   REGISTERS_reg_31_14_inst : DFF_X1 port map( D => n2757, CK => Clk, Q => n438
                           , QN => n4463);
   OUT2_reg_14_inst : DFF_X1 port map( D => n2756, CK => Clk, Q => OUT2(14), QN
                           => net644401);
   REGISTERS_reg_31_13_inst : DFF_X1 port map( D => n2755, CK => Clk, Q => n441
                           , QN => n4455);
   OUT2_reg_13_inst : DFF_X1 port map( D => n2754, CK => Clk, Q => OUT2(13), QN
                           => net644400);
   REGISTERS_reg_31_12_inst : DFF_X1 port map( D => n2753, CK => Clk, Q => n444
                           , QN => n4454);
   OUT2_reg_12_inst : DFF_X1 port map( D => n2752, CK => Clk, Q => OUT2(12), QN
                           => net644399);
   REGISTERS_reg_31_11_inst : DFF_X1 port map( D => n2751, CK => Clk, Q => n447
                           , QN => n4453);
   OUT2_reg_11_inst : DFF_X1 port map( D => n2750, CK => Clk, Q => OUT2(11), QN
                           => net644398);
   REGISTERS_reg_31_10_inst : DFF_X1 port map( D => n2749, CK => Clk, Q => n450
                           , QN => n4449);
   OUT2_reg_10_inst : DFF_X1 port map( D => n2748, CK => Clk, Q => OUT2(10), QN
                           => net644397);
   REGISTERS_reg_31_9_inst : DFF_X1 port map( D => n2747, CK => Clk, Q => n453,
                           QN => n4448);
   OUT2_reg_9_inst : DFF_X1 port map( D => n2746, CK => Clk, Q => OUT2(9), QN 
                           => net644396);
   REGISTERS_reg_31_8_inst : DFF_X1 port map( D => n2745, CK => Clk, Q => n456,
                           QN => n4443);
   OUT2_reg_8_inst : DFF_X1 port map( D => n2744, CK => Clk, Q => OUT2(8), QN 
                           => net644395);
   REGISTERS_reg_31_7_inst : DFF_X1 port map( D => n2743, CK => Clk, Q => n459,
                           QN => n4442);
   OUT2_reg_7_inst : DFF_X1 port map( D => n2742, CK => Clk, Q => OUT2(7), QN 
                           => net644394);
   REGISTERS_reg_31_6_inst : DFF_X1 port map( D => n2741, CK => Clk, Q => n462,
                           QN => n4433);
   OUT2_reg_6_inst : DFF_X1 port map( D => n2740, CK => Clk, Q => OUT2(6), QN 
                           => net644393);
   REGISTERS_reg_31_5_inst : DFF_X1 port map( D => n2739, CK => Clk, Q => n465,
                           QN => n4425);
   OUT2_reg_5_inst : DFF_X1 port map( D => n2738, CK => Clk, Q => OUT2(5), QN 
                           => net644392);
   REGISTERS_reg_31_4_inst : DFF_X1 port map( D => n2737, CK => Clk, Q => n468,
                           QN => n4424);
   OUT2_reg_4_inst : DFF_X1 port map( D => n2736, CK => Clk, Q => OUT2(4), QN 
                           => net644391);
   REGISTERS_reg_31_3_inst : DFF_X1 port map( D => n2735, CK => Clk, Q => n471,
                           QN => n4423);
   OUT2_reg_3_inst : DFF_X1 port map( D => n2734, CK => Clk, Q => OUT2(3), QN 
                           => net644390);
   REGISTERS_reg_31_2_inst : DFF_X1 port map( D => n2733, CK => Clk, Q => n474,
                           QN => n4419);
   OUT2_reg_2_inst : DFF_X1 port map( D => n2732, CK => Clk, Q => OUT2(2), QN 
                           => net644389);
   REGISTERS_reg_31_1_inst : DFF_X1 port map( D => n2731, CK => Clk, Q => n477,
                           QN => n4418);
   OUT2_reg_1_inst : DFF_X1 port map( D => n2730, CK => Clk, Q => OUT2(1), QN 
                           => net644388);
   REGISTERS_reg_31_0_inst : DFF_X1 port map( D => n2729, CK => Clk, Q => n4060
                           , QN => n2087);
   OUT2_reg_0_inst : DFF_X1 port map( D => n2728, CK => Clk, Q => OUT2(0), QN 
                           => n2184);
   OUT1_reg_31_inst : DFF_X1 port map( D => n2727, CK => Clk, Q => OUT1(31), QN
                           => net644387);
   OUT1_reg_30_inst : DFF_X1 port map( D => n2726, CK => Clk, Q => OUT1(30), QN
                           => net644386);
   OUT1_reg_29_inst : DFF_X1 port map( D => n2725, CK => Clk, Q => OUT1(29), QN
                           => net644385);
   OUT1_reg_28_inst : DFF_X1 port map( D => n2724, CK => Clk, Q => OUT1(28), QN
                           => net644384);
   OUT1_reg_27_inst : DFF_X1 port map( D => n2723, CK => Clk, Q => OUT1(27), QN
                           => net644383);
   OUT1_reg_26_inst : DFF_X1 port map( D => n2722, CK => Clk, Q => OUT1(26), QN
                           => net644382);
   OUT1_reg_25_inst : DFF_X1 port map( D => n2721, CK => Clk, Q => OUT1(25), QN
                           => net644381);
   OUT1_reg_24_inst : DFF_X1 port map( D => n2720, CK => Clk, Q => OUT1(24), QN
                           => net644380);
   OUT1_reg_23_inst : DFF_X1 port map( D => n2719, CK => Clk, Q => OUT1(23), QN
                           => net644379);
   OUT1_reg_22_inst : DFF_X1 port map( D => n2718, CK => Clk, Q => OUT1(22), QN
                           => net644378);
   OUT1_reg_21_inst : DFF_X1 port map( D => n2717, CK => Clk, Q => OUT1(21), QN
                           => net644377);
   OUT1_reg_20_inst : DFF_X1 port map( D => n2716, CK => Clk, Q => OUT1(20), QN
                           => net644376);
   OUT1_reg_19_inst : DFF_X1 port map( D => n2715, CK => Clk, Q => OUT1(19), QN
                           => net644375);
   OUT1_reg_18_inst : DFF_X1 port map( D => n2714, CK => Clk, Q => OUT1(18), QN
                           => net644374);
   OUT1_reg_17_inst : DFF_X1 port map( D => n2713, CK => Clk, Q => OUT1(17), QN
                           => net644373);
   OUT1_reg_16_inst : DFF_X1 port map( D => n2712, CK => Clk, Q => OUT1(16), QN
                           => net644372);
   OUT1_reg_15_inst : DFF_X1 port map( D => n2711, CK => Clk, Q => OUT1(15), QN
                           => net644371);
   OUT1_reg_14_inst : DFF_X1 port map( D => n2710, CK => Clk, Q => OUT1(14), QN
                           => net644370);
   OUT1_reg_13_inst : DFF_X1 port map( D => n2709, CK => Clk, Q => OUT1(13), QN
                           => net644369);
   OUT1_reg_12_inst : DFF_X1 port map( D => n2708, CK => Clk, Q => OUT1(12), QN
                           => net644368);
   OUT1_reg_11_inst : DFF_X1 port map( D => n2707, CK => Clk, Q => OUT1(11), QN
                           => net644367);
   OUT1_reg_10_inst : DFF_X1 port map( D => n2706, CK => Clk, Q => OUT1(10), QN
                           => net644366);
   OUT1_reg_9_inst : DFF_X1 port map( D => n2705, CK => Clk, Q => OUT1(9), QN 
                           => net644365);
   OUT1_reg_8_inst : DFF_X1 port map( D => n2704, CK => Clk, Q => OUT1(8), QN 
                           => net644364);
   OUT1_reg_7_inst : DFF_X1 port map( D => n2703, CK => Clk, Q => OUT1(7), QN 
                           => net644363);
   OUT1_reg_6_inst : DFF_X1 port map( D => n2702, CK => Clk, Q => OUT1(6), QN 
                           => net644362);
   OUT1_reg_5_inst : DFF_X1 port map( D => n2701, CK => Clk, Q => OUT1(5), QN 
                           => net644361);
   OUT1_reg_4_inst : DFF_X1 port map( D => n2700, CK => Clk, Q => OUT1(4), QN 
                           => net644360);
   OUT1_reg_3_inst : DFF_X1 port map( D => n2699, CK => Clk, Q => OUT1(3), QN 
                           => net644359);
   OUT1_reg_2_inst : DFF_X1 port map( D => n2698, CK => Clk, Q => OUT1(2), QN 
                           => net644358);
   OUT1_reg_1_inst : DFF_X1 port map( D => n2697, CK => Clk, Q => OUT1(1), QN 
                           => net644357);
   OUT1_reg_0_inst : DFF_X1 port map( D => n2696, CK => Clk, Q => OUT1(0), QN 
                           => n2152);
   U3574 : NAND3_X1 port map( A1 => ADD_RD2(4), A2 => ADD_RD2(3), A3 => n5189, 
                           ZN => n5170);
   U3575 : NAND3_X1 port map( A1 => ADD_RD2(3), A2 => n5189, A3 => n5190, ZN =>
                           n5158);
   U3576 : NAND3_X1 port map( A1 => n5194, A2 => ADD_RD2(4), A3 => ADD_RD2(0), 
                           ZN => n5155);
   U3577 : NAND3_X1 port map( A1 => ADD_RD2(0), A2 => ADD_RD2(4), A3 => 
                           ADD_RD2(3), ZN => n5181);
   U3578 : NAND3_X1 port map( A1 => ADD_RD2(4), A2 => n5189, A3 => n5194, ZN =>
                           n5179);
   U3579 : NAND3_X1 port map( A1 => ADD_RD2(0), A2 => n5190, A3 => n5194, ZN =>
                           n5157);
   U3580 : NAND3_X1 port map( A1 => n5189, A2 => n5190, A3 => n5194, ZN => 
                           n5169);
   U3581 : NAND3_X1 port map( A1 => ADD_RD2(0), A2 => ADD_RD2(3), A3 => n5190, 
                           ZN => n5173);
   U3582 : NAND3_X1 port map( A1 => ADD_RD1(3), A2 => ADD_RD1(4), A3 => n5966, 
                           ZN => n5950);
   U3583 : NAND3_X1 port map( A1 => ADD_RD1(3), A2 => n5967, A3 => n5966, ZN =>
                           n5938);
   U3584 : NAND3_X1 port map( A1 => n5971, A2 => ADD_RD1(4), A3 => ADD_RD1(0), 
                           ZN => n5935);
   U3585 : NAND3_X1 port map( A1 => ADD_RD1(4), A2 => ADD_RD1(3), A3 => 
                           ADD_RD1(0), ZN => n5959);
   U3586 : NAND3_X1 port map( A1 => ADD_RD1(4), A2 => n5971, A3 => n5966, ZN =>
                           n5958);
   U3587 : NAND3_X1 port map( A1 => ADD_RD1(0), A2 => n5967, A3 => n5971, ZN =>
                           n5937);
   U3588 : NAND3_X1 port map( A1 => n5967, A2 => n5971, A3 => n5966, ZN => 
                           n5949);
   U3589 : NAND3_X1 port map( A1 => ADD_RD1(3), A2 => ADD_RD1(0), A3 => n5967, 
                           ZN => n5953);
   U3557 : NOR3_X1 port map( A1 => n5979, A2 => n5973, A3 => n5978, ZN => n5980
                           );
   U3553 : NAND2_X1 port map( A1 => n5984, A2 => n1769, ZN => n5983);
   U3549 : AOI22_X1 port map( A1 => n1919, A2 => ADD_RD1(2), B1 => n5146, B2 =>
                           ADD_RD1(4), ZN => n5982);
   U3548 : OAI221_X1 port map( B1 => n1919, B2 => ADD_RD1(2), C1 => n5146, C2 
                           => ADD_RD1(4), A => n5982, ZN => n5981);
   U3534 : AOI22_X1 port map( A1 => n6355, A2 => n3915, B1 => n6357, B2 => 
                           n4059, ZN => n5927);
   U3531 : AOI22_X1 port map( A1 => net644901, A2 => n6356, B1 => net644869, B2
                           => n6358, ZN => n5928);
   U3530 : NOR2_X1 port map( A1 => n5958, A2 => n5939, ZN => n5925);
   U3525 : NOR2_X1 port map( A1 => n5978, A2 => n5979, ZN => n5976);
   U3524 : NAND2_X1 port map( A1 => n5976, A2 => n5977, ZN => n5975);
   U3523 : NOR4_X1 port map( A1 => Rst, A2 => n5973, A3 => n5974, A4 => n5975, 
                           ZN => n5260);
   U3522 : AOI22_X1 port map( A1 => net644451, A2 => n6360, B1 => DATAIN(0), B2
                           => n6359, ZN => n5972);
   U3521 : OAI21_X1 port map( B1 => n5257, B2 => n2152, A => n5972, ZN => n5968
                           );
   U3517 : OAI22_X1 port map( A1 => n671, A2 => n5255, B1 => n514, B2 => n3952,
                           ZN => n5969);
   U3516 : AOI211_X1 port map( C1 => net644675, C2 => n5925, A => n5968, B => 
                           n5969, ZN => n5929);
   U3512 : NAND2_X1 port map( A1 => n5963, A2 => n5964, ZN => n5952);
   U3509 : AOI22_X1 port map( A1 => net644515, A2 => n6363, B1 => net644547, B2
                           => n6362, ZN => n5940);
   U3505 : AOI22_X1 port map( A1 => n6364, A2 => n385, B1 => n5248, B2 => n4060
                           , ZN => n5954);
   U3502 : AOI22_X1 port map( A1 => net644612, A2 => n3911, B1 => net644483, B2
                           => n3912, ZN => n5955);
   U3498 : AOI22_X1 port map( A1 => n6366, A2 => n386, B1 => n5244, B2 => n4061
                           , ZN => n5956);
   U3495 : AOI22_X1 port map( A1 => net644580, A2 => n3913, B1 => net644676, B2
                           => n3914, ZN => n5957);
   U3494 : NAND4_X1 port map( A1 => n5954, A2 => n5955, A3 => n5956, A4 => 
                           n5957, ZN => n5942);
   U3490 : AOI22_X1 port map( A1 => n6368, A2 => n384, B1 => n5236, B2 => n4062
                           , ZN => n5944);
   U3487 : AOI22_X1 port map( A1 => net644772, A2 => n3910, B1 => net644740, B2
                           => n3909, ZN => n5945);
   U3484 : AOI22_X1 port map( A1 => net644902, A2 => n3908, B1 => net644419, B2
                           => n3907, ZN => n5946);
   U3481 : AOI22_X1 port map( A1 => net644867, A2 => n3906, B1 => net644868, B2
                           => n3905, ZN => n5947);
   U3480 : NAND4_X1 port map( A1 => n5944, A2 => n5945, A3 => n5946, A4 => 
                           n5947, ZN => n5943);
   U3479 : OAI21_X1 port map( B1 => n5942, B2 => n5943, A => n6370, ZN => n5941
                           );
   U3478 : OAI211_X1 port map( C1 => n703, C2 => n5220, A => n5940, B => n5941,
                           ZN => n5931);
   U3475 : NOR2_X1 port map( A1 => n5937, A2 => n5936, ZN => n5910);
   U3473 : AOI22_X1 port map( A1 => net644835, A2 => n5910, B1 => net644579, B2
                           => n5219, ZN => n5934);
   U3472 : OAI21_X1 port map( B1 => n481, B2 => n3953, A => n5934, ZN => n5932)
                           ;
   U3471 : AOI211_X1 port map( C1 => n6374, C2 => net644708, A => n5931, B => 
                           n5932, ZN => n5930);
   U3470 : NAND4_X1 port map( A1 => n5927, A2 => n5928, A3 => n5929, A4 => 
                           n5930, ZN => n2696);
   U2534 : AOI22_X1 port map( A1 => ADD_WR(2), A2 => ADD_RD2(2), B1 => n5186, 
                           B2 => n1919, ZN => n5196);
   U2531 : NOR3_X1 port map( A1 => n5202, A2 => n5196, A3 => n5201, ZN => n5205
                           );
   U2530 : AOI22_X1 port map( A1 => n5146, A2 => ADD_RD2(4), B1 => ADD_RD2(3), 
                           B2 => n1846, ZN => n5208);
   U2529 : OAI221_X1 port map( B1 => n5146, B2 => ADD_RD2(4), C1 => n1846, C2 
                           => ADD_RD2(3), A => n5208, ZN => n5207);
   U2528 : NOR2_X1 port map( A1 => n5206, A2 => n5207, ZN => n5200);
   U2517 : AOI22_X1 port map( A1 => n4241, A2 => n3915, B1 => n6377, B2 => 
                           n4059, ZN => n5147);
   U2514 : AOI22_X1 port map( A1 => net644901, A2 => n6375, B1 => net644869, B2
                           => n6378, ZN => n5148);
   U2513 : NOR2_X1 port map( A1 => n5179, A2 => n5159, ZN => n5142);
   U2508 : NOR2_X1 port map( A1 => n5201, A2 => n5202, ZN => n5199);
   U2507 : NAND2_X1 port map( A1 => n5199, A2 => n5200, ZN => n5198);
   U2506 : NOR4_X1 port map( A1 => Rst, A2 => n5196, A3 => n5197, A4 => n5198, 
                           ZN => n4238);
   U2505 : AOI22_X1 port map( A1 => net644451, A2 => n4237, B1 => DATAIN(0), B2
                           => n6379, ZN => n5195);
   U2504 : OAI21_X1 port map( B1 => n4235, B2 => n2184, A => n5195, ZN => n5191
                           );
   U2500 : OAI22_X1 port map( A1 => n671, A2 => n4234, B1 => n514, B2 => n3950,
                           ZN => n5192);
   U2499 : AOI211_X1 port map( C1 => net644675, C2 => n5142, A => n5191, B => 
                           n5192, ZN => n5149);
   U2495 : NAND2_X1 port map( A1 => n5186, A2 => n5187, ZN => n5172);
   U2492 : AOI22_X1 port map( A1 => net644515, A2 => n3880, B1 => net644547, B2
                           => n4228, ZN => n5160);
   U2489 : AOI22_X1 port map( A1 => n3896, A2 => n385, B1 => n4225, B2 => n4060
                           , ZN => n5175);
   U2486 : AOI22_X1 port map( A1 => net644612, A2 => n4223, B1 => net644483, B2
                           => n3894, ZN => n5176);
   U2483 : AOI22_X1 port map( A1 => n6384, A2 => n386, B1 => n3891, B2 => n4061
                           , ZN => n5177);
   U2480 : AOI22_X1 port map( A1 => net644580, A2 => n3890, B1 => net644676, B2
                           => n4219, ZN => n5178);
   U2479 : NAND4_X1 port map( A1 => n5175, A2 => n5176, A3 => n5177, A4 => 
                           n5178, ZN => n5162);
   U2476 : AOI22_X1 port map( A1 => n3903, A2 => n384, B1 => n3904, B2 => n4062
                           , ZN => n5164);
   U2473 : AOI22_X1 port map( A1 => net644772, A2 => n4209, B1 => net644740, B2
                           => n3901, ZN => n5165);
   U2470 : AOI22_X1 port map( A1 => net644902, A2 => n4207, B1 => net644419, B2
                           => n3899, ZN => n5166);
   U2468 : NOR2_X1 port map( A1 => n5168, A2 => n5169, ZN => n4204);
   U2467 : AOI22_X1 port map( A1 => net644867, A2 => n3898, B1 => net644868, B2
                           => n6385, ZN => n5167);
   U2466 : NAND4_X1 port map( A1 => n5164, A2 => n5165, A3 => n5166, A4 => 
                           n5167, ZN => n5163);
   U2465 : OAI21_X1 port map( B1 => n5162, B2 => n5163, A => n6386, ZN => n5161
                           );
   U2464 : OAI211_X1 port map( C1 => n703, C2 => n4194, A => n5160, B => n5161,
                           ZN => n5151);
   U2461 : NOR2_X1 port map( A1 => n5157, A2 => n5156, ZN => n5124);
   U2459 : AOI22_X1 port map( A1 => net644835, A2 => n5124, B1 => net644579, B2
                           => n6388, ZN => n5154);
   U2458 : OAI21_X1 port map( B1 => n481, B2 => n3951, A => n5154, ZN => n5152)
                           ;
   U2457 : AOI211_X1 port map( C1 => net644708, C2 => n4186, A => n5151, B => 
                           n5152, ZN => n5150);
   U2456 : NAND4_X1 port map( A1 => n5147, A2 => n5148, A3 => n5149, A4 => 
                           n5150, ZN => n2728);
   U2596 : AOI22_X1 port map( A1 => n5263, A2 => n3948, B1 => n5264, B2 => 
                           n4053, ZN => n5265);
   U2595 : AOI22_X1 port map( A1 => n5261, A2 => net644899, B1 => n5262, B2 => 
                           net644865, ZN => n5266);
   U2594 : AOI22_X1 port map( A1 => n6360, A2 => net644481, B1 => n6359, B2 => 
                           DATAIN(30), ZN => n5286);
   U2593 : OAI21_X1 port map( B1 => n5257, B2 => net644386, A => n5286, ZN => 
                           n5284);
   U2592 : OAI22_X1 port map( A1 => n516, A2 => n5255, B1 => n641, B2 => n5256,
                           ZN => n5285);
   U2591 : AOI211_X1 port map( C1 => n6361, C2 => net644673, A => n5284, B => 
                           n5285, ZN => n5267);
   U2590 : AOI22_X1 port map( A1 => n6363, A2 => net644545, B1 => n6362, B2 => 
                           net644577, ZN => n5272);
   U2588 : AOI22_X1 port map( A1 => n5248, A2 => n390, B1 => n5249, B2 => n4161
                           , ZN => n5280);
   U2587 : AOI22_X1 port map( A1 => n3911, A2 => net644642, B1 => n3912, B2 => 
                           net644513, ZN => n5281);
   U2585 : AOI22_X1 port map( A1 => n5244, A2 => n4054, B1 => n5245, B2 => n354
                           , ZN => n5282);
   U2584 : AOI22_X1 port map( A1 => n3913, A2 => net644610, B1 => n3914, B2 => 
                           net644706, ZN => n5283);
   U2583 : NAND4_X1 port map( A1 => n5280, A2 => n5281, A3 => n5282, A4 => 
                           n5283, ZN => n5274);
   U2581 : AOI22_X1 port map( A1 => n5236, A2 => n392, B1 => n5237, B2 => n4162
                           , ZN => n5276);
   U2580 : AOI22_X1 port map( A1 => n3910, A2 => net644802, B1 => n3909, B2 => 
                           net644770, ZN => n5277);
   U2579 : AOI22_X1 port map( A1 => n3908, A2 => net644932, B1 => n3907, B2 => 
                           net644449, ZN => n5278);
   U2577 : AOI22_X1 port map( A1 => n3906, A2 => n4055, B1 => n3905, B2 => n391
                           , ZN => n5279);
   U2576 : NAND4_X1 port map( A1 => n5276, A2 => n5277, A3 => n5278, A4 => 
                           n5279, ZN => n5275);
   U2575 : OAI21_X1 port map( B1 => n5274, B2 => n5275, A => n6370, ZN => n5273
                           );
   U2574 : OAI211_X1 port map( C1 => n547, C2 => n5220, A => n5272, B => n5273,
                           ZN => n5269);
   U2572 : AOI22_X1 port map( A1 => n6373, A2 => net644833, B1 => n6372, B2 => 
                           n4163, ZN => n5271);
   U2571 : OAI21_X1 port map( B1 => n609, B2 => n5216, A => n5271, ZN => n5270)
                           ;
   U2570 : AOI211_X1 port map( C1 => n5213, C2 => net644738, A => n5269, B => 
                           n5270, ZN => n5268);
   U2569 : NAND4_X1 port map( A1 => n5265, A2 => n5266, A3 => n5267, A4 => 
                           n5268, ZN => n2726);
   U2626 : AOI22_X1 port map( A1 => n5263, A2 => n3947, B1 => n5264, B2 => 
                           n4050, ZN => n5287);
   U2625 : AOI22_X1 port map( A1 => n5261, A2 => net644898, B1 => n5262, B2 => 
                           net644864, ZN => n5288);
   U2624 : AOI22_X1 port map( A1 => n5259, A2 => net644480, B1 => n5260, B2 => 
                           DATAIN(29), ZN => n5308);
   U2623 : OAI21_X1 port map( B1 => n5257, B2 => net644385, A => n5308, ZN => 
                           n5306);
   U2622 : OAI22_X1 port map( A1 => n517, A2 => n5255, B1 => n642, B2 => n5256,
                           ZN => n5307);
   U2621 : AOI211_X1 port map( C1 => n6361, C2 => net644672, A => n5306, B => 
                           n5307, ZN => n5289);
   U2620 : AOI22_X1 port map( A1 => n5250, A2 => net644544, B1 => n5251, B2 => 
                           net644576, ZN => n5294);
   U2618 : AOI22_X1 port map( A1 => n5248, A2 => n393, B1 => n5249, B2 => n4158
                           , ZN => n5302);
   U2617 : AOI22_X1 port map( A1 => n3911, A2 => net644641, B1 => n3912, B2 => 
                           net644512, ZN => n5303);
   U2615 : AOI22_X1 port map( A1 => n5244, A2 => n4051, B1 => n5245, B2 => n355
                           , ZN => n5304);
   U2614 : AOI22_X1 port map( A1 => n3913, A2 => net644609, B1 => n3914, B2 => 
                           net644705, ZN => n5305);
   U2613 : NAND4_X1 port map( A1 => n5302, A2 => n5303, A3 => n5304, A4 => 
                           n5305, ZN => n5296);
   U2611 : AOI22_X1 port map( A1 => n5236, A2 => n395, B1 => n5237, B2 => n4159
                           , ZN => n5298);
   U2610 : AOI22_X1 port map( A1 => n3910, A2 => net644801, B1 => n3909, B2 => 
                           net644769, ZN => n5299);
   U2609 : AOI22_X1 port map( A1 => n3908, A2 => net644931, B1 => n3907, B2 => 
                           net644448, ZN => n5300);
   U2607 : AOI22_X1 port map( A1 => n3906, A2 => n4052, B1 => n3905, B2 => n394
                           , ZN => n5301);
   U2606 : NAND4_X1 port map( A1 => n5298, A2 => n5299, A3 => n5300, A4 => 
                           n5301, ZN => n5297);
   U2605 : OAI21_X1 port map( B1 => n5296, B2 => n5297, A => n6370, ZN => n5295
                           );
   U2604 : OAI211_X1 port map( C1 => n548, C2 => n5220, A => n5294, B => n5295,
                           ZN => n5291);
   U2602 : AOI22_X1 port map( A1 => n6373, A2 => net644832, B1 => n6372, B2 => 
                           n4160, ZN => n5293);
   U2601 : OAI21_X1 port map( B1 => n610, B2 => n5216, A => n5293, ZN => n5292)
                           ;
   U2600 : AOI211_X1 port map( C1 => n5213, C2 => net644737, A => n5291, B => 
                           n5292, ZN => n5290);
   U2599 : NAND4_X1 port map( A1 => n5287, A2 => n5288, A3 => n5289, A4 => 
                           n5290, ZN => n2725);
   U2656 : AOI22_X1 port map( A1 => n5263, A2 => n3946, B1 => n5264, B2 => 
                           n4047, ZN => n5309);
   U2655 : AOI22_X1 port map( A1 => n5261, A2 => net644897, B1 => n5262, B2 => 
                           net644863, ZN => n5310);
   U2654 : AOI22_X1 port map( A1 => n6360, A2 => net644479, B1 => n5260, B2 => 
                           DATAIN(28), ZN => n5330);
   U2653 : OAI21_X1 port map( B1 => n5257, B2 => net644384, A => n5330, ZN => 
                           n5328);
   U2652 : OAI22_X1 port map( A1 => n518, A2 => n5255, B1 => n643, B2 => n5256,
                           ZN => n5329);
   U2651 : AOI211_X1 port map( C1 => n6361, C2 => net644671, A => n5328, B => 
                           n5329, ZN => n5311);
   U2650 : AOI22_X1 port map( A1 => n6363, A2 => net644543, B1 => n5251, B2 => 
                           net644575, ZN => n5316);
   U2648 : AOI22_X1 port map( A1 => n5248, A2 => n396, B1 => n5249, B2 => n4155
                           , ZN => n5324);
   U2647 : AOI22_X1 port map( A1 => n3911, A2 => net644640, B1 => n3912, B2 => 
                           net644511, ZN => n5325);
   U2645 : AOI22_X1 port map( A1 => n5244, A2 => n4048, B1 => n5245, B2 => n356
                           , ZN => n5326);
   U2644 : AOI22_X1 port map( A1 => n3913, A2 => net644608, B1 => n3914, B2 => 
                           net644704, ZN => n5327);
   U2643 : NAND4_X1 port map( A1 => n5324, A2 => n5325, A3 => n5326, A4 => 
                           n5327, ZN => n5318);
   U2641 : AOI22_X1 port map( A1 => n5236, A2 => n398, B1 => n5237, B2 => n4156
                           , ZN => n5320);
   U2640 : AOI22_X1 port map( A1 => n3910, A2 => net644800, B1 => n3909, B2 => 
                           net644768, ZN => n5321);
   U2639 : AOI22_X1 port map( A1 => n3908, A2 => net644930, B1 => n3907, B2 => 
                           net644447, ZN => n5322);
   U2637 : AOI22_X1 port map( A1 => n3906, A2 => n4049, B1 => n3905, B2 => n397
                           , ZN => n5323);
   U2636 : NAND4_X1 port map( A1 => n5320, A2 => n5321, A3 => n5322, A4 => 
                           n5323, ZN => n5319);
   U2635 : OAI21_X1 port map( B1 => n5318, B2 => n5319, A => n6370, ZN => n5317
                           );
   U2634 : OAI211_X1 port map( C1 => n549, C2 => n5220, A => n5316, B => n5317,
                           ZN => n5313);
   U2632 : AOI22_X1 port map( A1 => n6373, A2 => net644831, B1 => n6372, B2 => 
                           n4157, ZN => n5315);
   U2631 : OAI21_X1 port map( B1 => n611, B2 => n5216, A => n5315, ZN => n5314)
                           ;
   U2630 : AOI211_X1 port map( C1 => n5213, C2 => net644736, A => n5313, B => 
                           n5314, ZN => n5312);
   U2629 : NAND4_X1 port map( A1 => n5309, A2 => n5310, A3 => n5311, A4 => 
                           n5312, ZN => n2724);
   U2566 : AOI22_X1 port map( A1 => n5263, A2 => n3949, B1 => n5264, B2 => 
                           n4056, ZN => n5209);
   U2565 : AOI22_X1 port map( A1 => n6358, A2 => net644900, B1 => n5262, B2 => 
                           net644866, ZN => n5210);
   U2564 : AOI22_X1 port map( A1 => n5259, A2 => net644482, B1 => n6359, B2 => 
                           DATAIN(31), ZN => n5258);
   U2563 : OAI21_X1 port map( B1 => n5257, B2 => net644387, A => n5258, ZN => 
                           n5253);
   U2562 : OAI22_X1 port map( A1 => n515, A2 => n5255, B1 => n640, B2 => n5256,
                           ZN => n5254);
   U2561 : AOI211_X1 port map( C1 => n6361, C2 => net644674, A => n5253, B => 
                           n5254, ZN => n5211);
   U2560 : AOI22_X1 port map( A1 => n5250, A2 => net644546, B1 => n6362, B2 => 
                           net644578, ZN => n5221);
   U2558 : AOI22_X1 port map( A1 => n6365, A2 => n387, B1 => n5249, B2 => n4164
                           , ZN => n5238);
   U2557 : AOI22_X1 port map( A1 => n3911, A2 => net644643, B1 => n3912, B2 => 
                           net644514, ZN => n5239);
   U2555 : AOI22_X1 port map( A1 => n6367, A2 => n4057, B1 => n5245, B2 => n353
                           , ZN => n5240);
   U2554 : AOI22_X1 port map( A1 => n3913, A2 => net644611, B1 => n3914, B2 => 
                           net644707, ZN => n5241);
   U2553 : NAND4_X1 port map( A1 => n5238, A2 => n5239, A3 => n5240, A4 => 
                           n5241, ZN => n5223);
   U2551 : AOI22_X1 port map( A1 => n6369, A2 => n389, B1 => n5237, B2 => n4165
                           , ZN => n5226);
   U2550 : AOI22_X1 port map( A1 => n3910, A2 => net644803, B1 => n3909, B2 => 
                           net644771, ZN => n5227);
   U2549 : AOI22_X1 port map( A1 => n3908, A2 => net644933, B1 => n3907, B2 => 
                           net644450, ZN => n5228);
   U2547 : AOI22_X1 port map( A1 => n3906, A2 => n4058, B1 => n3905, B2 => n388
                           , ZN => n5229);
   U2546 : NAND4_X1 port map( A1 => n5226, A2 => n5227, A3 => n5228, A4 => 
                           n5229, ZN => n5224);
   U2545 : OAI21_X1 port map( B1 => n5223, B2 => n5224, A => n6370, ZN => n5222
                           );
   U2544 : OAI211_X1 port map( C1 => n546, C2 => n5220, A => n5221, B => n5222,
                           ZN => n5214);
   U2542 : AOI22_X1 port map( A1 => n6373, A2 => net644834, B1 => n6372, B2 => 
                           n4166, ZN => n5217);
   U2541 : OAI21_X1 port map( B1 => n608, B2 => n5216, A => n5217, ZN => n5215)
                           ;
   U2540 : AOI211_X1 port map( C1 => n5213, C2 => net644739, A => n5214, B => 
                           n5215, ZN => n5212);
   U2539 : NAND4_X1 port map( A1 => n5209, A2 => n5210, A3 => n5211, A4 => 
                           n5212, ZN => n2727);
   U2746 : AOI22_X1 port map( A1 => n6356, A2 => n3943, B1 => n5264, B2 => 
                           n4038, ZN => n5375);
   U2745 : AOI22_X1 port map( A1 => n6358, A2 => net644894, B1 => n5262, B2 => 
                           net644860, ZN => n5376);
   U2744 : AOI22_X1 port map( A1 => n6360, A2 => net644476, B1 => n6359, B2 => 
                           DATAIN(25), ZN => n5396);
   U2743 : OAI21_X1 port map( B1 => n5257, B2 => net644381, A => n5396, ZN => 
                           n5394);
   U2742 : OAI22_X1 port map( A1 => n521, A2 => n5255, B1 => n646, B2 => n5256,
                           ZN => n5395);
   U2741 : AOI211_X1 port map( C1 => n6361, C2 => net644668, A => n5394, B => 
                           n5395, ZN => n5377);
   U2740 : AOI22_X1 port map( A1 => n6363, A2 => net644540, B1 => n6362, B2 => 
                           net644572, ZN => n5382);
   U2738 : AOI22_X1 port map( A1 => n6365, A2 => n405, B1 => n5249, B2 => n4144
                           , ZN => n5390);
   U2737 : AOI22_X1 port map( A1 => n3911, A2 => net644637, B1 => n3912, B2 => 
                           net644508, ZN => n5391);
   U2735 : AOI22_X1 port map( A1 => n5244, A2 => n4039, B1 => n5245, B2 => n359
                           , ZN => n5392);
   U2734 : AOI22_X1 port map( A1 => n3913, A2 => net644605, B1 => n3914, B2 => 
                           net644701, ZN => n5393);
   U2733 : NAND4_X1 port map( A1 => n5390, A2 => n5391, A3 => n5392, A4 => 
                           n5393, ZN => n5384);
   U2731 : AOI22_X1 port map( A1 => n5236, A2 => n407, B1 => n5237, B2 => n4147
                           , ZN => n5386);
   U2730 : AOI22_X1 port map( A1 => n3910, A2 => net644797, B1 => n3909, B2 => 
                           net644765, ZN => n5387);
   U2729 : AOI22_X1 port map( A1 => n3908, A2 => net644927, B1 => n3907, B2 => 
                           net644444, ZN => n5388);
   U2727 : AOI22_X1 port map( A1 => n3906, A2 => n4040, B1 => n3905, B2 => n406
                           , ZN => n5389);
   U2726 : NAND4_X1 port map( A1 => n5386, A2 => n5387, A3 => n5388, A4 => 
                           n5389, ZN => n5385);
   U2725 : OAI21_X1 port map( B1 => n5384, B2 => n5385, A => n6370, ZN => n5383
                           );
   U2724 : OAI211_X1 port map( C1 => n552, C2 => n5220, A => n5382, B => n5383,
                           ZN => n5379);
   U2722 : AOI22_X1 port map( A1 => n6373, A2 => net644828, B1 => n6372, B2 => 
                           n4148, ZN => n5381);
   U2721 : OAI21_X1 port map( B1 => n614, B2 => n5216, A => n5381, ZN => n5380)
                           ;
   U2720 : AOI211_X1 port map( C1 => n5213, C2 => net644733, A => n5379, B => 
                           n5380, ZN => n5378);
   U2719 : NAND4_X1 port map( A1 => n5375, A2 => n5376, A3 => n5377, A4 => 
                           n5378, ZN => n2721);
   U3046 : AOI22_X1 port map( A1 => n6356, A2 => n3933, B1 => n5264, B2 => 
                           n4005, ZN => n5595);
   U3045 : AOI22_X1 port map( A1 => n6358, A2 => net644884, B1 => n6357, B2 => 
                           net644850, ZN => n5596);
   U3044 : AOI22_X1 port map( A1 => n6360, A2 => net644466, B1 => n6359, B2 => 
                           DATAIN(15), ZN => n5616);
   U3043 : OAI21_X1 port map( B1 => n5257, B2 => net644371, A => n5616, ZN => 
                           n5614);
   U3042 : OAI22_X1 port map( A1 => n531, A2 => n5255, B1 => n656, B2 => n5256,
                           ZN => n5615);
   U3041 : AOI211_X1 port map( C1 => n6361, C2 => net644658, A => n5614, B => 
                           n5615, ZN => n5597);
   U3040 : AOI22_X1 port map( A1 => n6363, A2 => net644530, B1 => n6362, B2 => 
                           net644562, ZN => n5602);
   U3038 : AOI22_X1 port map( A1 => n6365, A2 => n435, B1 => n5249, B2 => n4113
                           , ZN => n5610);
   U3037 : AOI22_X1 port map( A1 => n3911, A2 => net644627, B1 => n3912, B2 => 
                           net644498, ZN => n5611);
   U3035 : AOI22_X1 port map( A1 => n6367, A2 => n4006, B1 => n5245, B2 => n369
                           , ZN => n5612);
   U3034 : AOI22_X1 port map( A1 => n3913, A2 => net644595, B1 => n3914, B2 => 
                           net644691, ZN => n5613);
   U3033 : NAND4_X1 port map( A1 => n5610, A2 => n5611, A3 => n5612, A4 => 
                           n5613, ZN => n5604);
   U3031 : AOI22_X1 port map( A1 => n6369, A2 => n437, B1 => n5237, B2 => n4114
                           , ZN => n5606);
   U3030 : AOI22_X1 port map( A1 => n3910, A2 => net644787, B1 => n3909, B2 => 
                           net644755, ZN => n5607);
   U3029 : AOI22_X1 port map( A1 => n3908, A2 => net644917, B1 => n3907, B2 => 
                           net644434, ZN => n5608);
   U3027 : AOI22_X1 port map( A1 => n3906, A2 => n4007, B1 => n3905, B2 => n436
                           , ZN => n5609);
   U3026 : NAND4_X1 port map( A1 => n5606, A2 => n5607, A3 => n5608, A4 => 
                           n5609, ZN => n5605);
   U3025 : OAI21_X1 port map( B1 => n5604, B2 => n5605, A => n6370, ZN => n5603
                           );
   U3024 : OAI211_X1 port map( C1 => n562, C2 => n5220, A => n5602, B => n5603,
                           ZN => n5599);
   U3022 : AOI22_X1 port map( A1 => n6373, A2 => net644818, B1 => n6372, B2 => 
                           n4115, ZN => n5601);
   U3021 : OAI21_X1 port map( B1 => n624, B2 => n5216, A => n5601, ZN => n5600)
                           ;
   U3020 : AOI211_X1 port map( C1 => n5213, C2 => net644723, A => n5599, B => 
                           n5600, ZN => n5598);
   U3019 : NAND4_X1 port map( A1 => n5595, A2 => n5596, A3 => n5597, A4 => 
                           n5598, ZN => n2711);
   U3076 : AOI22_X1 port map( A1 => n6356, A2 => n3932, B1 => n5264, B2 => 
                           n4002, ZN => n5617);
   U3075 : AOI22_X1 port map( A1 => n6358, A2 => net644883, B1 => n6357, B2 => 
                           net644849, ZN => n5618);
   U3074 : AOI22_X1 port map( A1 => n6360, A2 => net644465, B1 => n6359, B2 => 
                           DATAIN(14), ZN => n5638);
   U3073 : OAI21_X1 port map( B1 => n5257, B2 => net644370, A => n5638, ZN => 
                           n5636);
   U3072 : OAI22_X1 port map( A1 => n532, A2 => n5255, B1 => n657, B2 => n5256,
                           ZN => n5637);
   U3071 : AOI211_X1 port map( C1 => n6361, C2 => net644657, A => n5636, B => 
                           n5637, ZN => n5619);
   U3070 : AOI22_X1 port map( A1 => n6363, A2 => net644529, B1 => n6362, B2 => 
                           net644561, ZN => n5624);
   U3068 : AOI22_X1 port map( A1 => n6365, A2 => n438, B1 => n5249, B2 => n4105
                           , ZN => n5632);
   U3067 : AOI22_X1 port map( A1 => n3911, A2 => net644626, B1 => n3912, B2 => 
                           net644497, ZN => n5633);
   U3065 : AOI22_X1 port map( A1 => n6367, A2 => n4003, B1 => n5245, B2 => n370
                           , ZN => n5634);
   U3064 : AOI22_X1 port map( A1 => n3913, A2 => net644594, B1 => n3914, B2 => 
                           net644690, ZN => n5635);
   U3063 : NAND4_X1 port map( A1 => n5632, A2 => n5633, A3 => n5634, A4 => 
                           n5635, ZN => n5626);
   U3061 : AOI22_X1 port map( A1 => n6369, A2 => n440, B1 => n5237, B2 => n4109
                           , ZN => n5628);
   U3060 : AOI22_X1 port map( A1 => n3910, A2 => net644786, B1 => n3909, B2 => 
                           net644754, ZN => n5629);
   U3059 : AOI22_X1 port map( A1 => n3908, A2 => net644916, B1 => n3907, B2 => 
                           net644433, ZN => n5630);
   U3057 : AOI22_X1 port map( A1 => n3906, A2 => n4004, B1 => n3905, B2 => n439
                           , ZN => n5631);
   U3056 : NAND4_X1 port map( A1 => n5628, A2 => n5629, A3 => n5630, A4 => 
                           n5631, ZN => n5627);
   U3055 : OAI21_X1 port map( B1 => n5626, B2 => n5627, A => n6370, ZN => n5625
                           );
   U3054 : OAI211_X1 port map( C1 => n563, C2 => n5220, A => n5624, B => n5625,
                           ZN => n5621);
   U3052 : AOI22_X1 port map( A1 => n6373, A2 => net644817, B1 => n6372, B2 => 
                           n4112, ZN => n5623);
   U3051 : OAI21_X1 port map( B1 => n625, B2 => n5216, A => n5623, ZN => n5622)
                           ;
   U3050 : AOI211_X1 port map( C1 => n5213, C2 => net644722, A => n5621, B => 
                           n5622, ZN => n5620);
   U3049 : NAND4_X1 port map( A1 => n5617, A2 => n5618, A3 => n5619, A4 => 
                           n5620, ZN => n2710);
   U3226 : AOI22_X1 port map( A1 => n6356, A2 => n3925, B1 => n6355, B2 => 
                           n3981, ZN => n5727);
   U3225 : AOI22_X1 port map( A1 => n6358, A2 => net644878, B1 => n6357, B2 => 
                           net644844, ZN => n5728);
   U3224 : AOI22_X1 port map( A1 => n6360, A2 => net644460, B1 => n6359, B2 => 
                           DATAIN(9), ZN => n5748);
   U3223 : OAI21_X1 port map( B1 => n5257, B2 => net644365, A => n5748, ZN => 
                           n5746);
   U3222 : OAI22_X1 port map( A1 => n537, A2 => n5255, B1 => n662, B2 => n5256,
                           ZN => n5747);
   U3221 : AOI211_X1 port map( C1 => n6361, C2 => net644652, A => n5746, B => 
                           n5747, ZN => n5729);
   U3220 : AOI22_X1 port map( A1 => n6363, A2 => net644524, B1 => n6362, B2 => 
                           net644556, ZN => n5734);
   U3218 : AOI22_X1 port map( A1 => n6365, A2 => n453, B1 => n6364, B2 => n4090
                           , ZN => n5742);
   U3217 : AOI22_X1 port map( A1 => n3911, A2 => net644621, B1 => n3912, B2 => 
                           net644492, ZN => n5743);
   U3215 : AOI22_X1 port map( A1 => n6367, A2 => n3982, B1 => n6366, B2 => n375
                           , ZN => n5744);
   U3214 : AOI22_X1 port map( A1 => n3913, A2 => net644589, B1 => n3914, B2 => 
                           net644685, ZN => n5745);
   U3213 : NAND4_X1 port map( A1 => n5742, A2 => n5743, A3 => n5744, A4 => 
                           n5745, ZN => n5736);
   U3211 : AOI22_X1 port map( A1 => n6369, A2 => n455, B1 => n6368, B2 => n4091
                           , ZN => n5738);
   U3210 : AOI22_X1 port map( A1 => n3910, A2 => net644781, B1 => n3909, B2 => 
                           net644749, ZN => n5739);
   U3209 : AOI22_X1 port map( A1 => n3908, A2 => net644911, B1 => n3907, B2 => 
                           net644428, ZN => n5740);
   U3207 : AOI22_X1 port map( A1 => n3906, A2 => n3983, B1 => n3905, B2 => n454
                           , ZN => n5741);
   U3206 : NAND4_X1 port map( A1 => n5738, A2 => n5739, A3 => n5740, A4 => 
                           n5741, ZN => n5737);
   U3205 : OAI21_X1 port map( B1 => n5736, B2 => n5737, A => n6370, ZN => n5735
                           );
   U3204 : OAI211_X1 port map( C1 => n568, C2 => n5220, A => n5734, B => n5735,
                           ZN => n5731);
   U3202 : AOI22_X1 port map( A1 => n6373, A2 => net644812, B1 => n6372, B2 => 
                           n4092, ZN => n5733);
   U3201 : OAI21_X1 port map( B1 => n630, B2 => n5216, A => n5733, ZN => n5732)
                           ;
   U3200 : AOI211_X1 port map( C1 => n6374, C2 => net644717, A => n5731, B => 
                           n5732, ZN => n5730);
   U3199 : NAND4_X1 port map( A1 => n5727, A2 => n5728, A3 => n5729, A4 => 
                           n5730, ZN => n2705);
   U3106 : AOI22_X1 port map( A1 => n6356, A2 => n3931, B1 => n5264, B2 => 
                           n3993, ZN => n5639);
   U3105 : AOI22_X1 port map( A1 => n6358, A2 => net644882, B1 => n6357, B2 => 
                           net644848, ZN => n5640);
   U3104 : AOI22_X1 port map( A1 => n6360, A2 => net644464, B1 => n6359, B2 => 
                           DATAIN(13), ZN => n5660);
   U3103 : OAI21_X1 port map( B1 => n5257, B2 => net644369, A => n5660, ZN => 
                           n5658);
   U3102 : OAI22_X1 port map( A1 => n533, A2 => n5255, B1 => n658, B2 => n5256,
                           ZN => n5659);
   U3101 : AOI211_X1 port map( C1 => n6361, C2 => net644656, A => n5658, B => 
                           n5659, ZN => n5641);
   U3100 : AOI22_X1 port map( A1 => n6363, A2 => net644528, B1 => n6362, B2 => 
                           net644560, ZN => n5646);
   U3098 : AOI22_X1 port map( A1 => n6365, A2 => n441, B1 => n5249, B2 => n4102
                           , ZN => n5654);
   U3097 : AOI22_X1 port map( A1 => n3911, A2 => net644625, B1 => n3912, B2 => 
                           net644496, ZN => n5655);
   U3095 : AOI22_X1 port map( A1 => n6367, A2 => n3998, B1 => n5245, B2 => n371
                           , ZN => n5656);
   U3094 : AOI22_X1 port map( A1 => n3913, A2 => net644593, B1 => n3914, B2 => 
                           net644689, ZN => n5657);
   U3093 : NAND4_X1 port map( A1 => n5654, A2 => n5655, A3 => n5656, A4 => 
                           n5657, ZN => n5648);
   U3091 : AOI22_X1 port map( A1 => n6369, A2 => n443, B1 => n5237, B2 => n4103
                           , ZN => n5650);
   U3090 : AOI22_X1 port map( A1 => n3910, A2 => net644785, B1 => n3909, B2 => 
                           net644753, ZN => n5651);
   U3089 : AOI22_X1 port map( A1 => n3908, A2 => net644915, B1 => n3907, B2 => 
                           net644432, ZN => n5652);
   U3087 : AOI22_X1 port map( A1 => n3906, A2 => n3999, B1 => n3905, B2 => n442
                           , ZN => n5653);
   U3086 : NAND4_X1 port map( A1 => n5650, A2 => n5651, A3 => n5652, A4 => 
                           n5653, ZN => n5649);
   U3085 : OAI21_X1 port map( B1 => n5648, B2 => n5649, A => n6370, ZN => n5647
                           );
   U3084 : OAI211_X1 port map( C1 => n564, C2 => n5220, A => n5646, B => n5647,
                           ZN => n5643);
   U3082 : AOI22_X1 port map( A1 => n6373, A2 => net644816, B1 => n6372, B2 => 
                           n4104, ZN => n5645);
   U3081 : OAI21_X1 port map( B1 => n626, B2 => n5216, A => n5645, ZN => n5644)
                           ;
   U3080 : AOI211_X1 port map( C1 => n5213, C2 => net644721, A => n5643, B => 
                           n5644, ZN => n5642);
   U3079 : NAND4_X1 port map( A1 => n5639, A2 => n5640, A3 => n5641, A4 => 
                           n5642, ZN => n2709);
   U2986 : AOI22_X1 port map( A1 => n5263, A2 => n3935, B1 => n5264, B2 => 
                           n4011, ZN => n5551);
   U2985 : AOI22_X1 port map( A1 => n6358, A2 => net644886, B1 => n6357, B2 => 
                           net644852, ZN => n5552);
   U2984 : AOI22_X1 port map( A1 => n5259, A2 => net644468, B1 => n6359, B2 => 
                           DATAIN(17), ZN => n5572);
   U2983 : OAI21_X1 port map( B1 => n5257, B2 => net644373, A => n5572, ZN => 
                           n5570);
   U2982 : OAI22_X1 port map( A1 => n529, A2 => n5255, B1 => n654, B2 => n5256,
                           ZN => n5571);
   U2981 : AOI211_X1 port map( C1 => n6361, C2 => net644660, A => n5570, B => 
                           n5571, ZN => n5553);
   U2980 : AOI22_X1 port map( A1 => n5250, A2 => net644532, B1 => n6362, B2 => 
                           net644564, ZN => n5558);
   U2978 : AOI22_X1 port map( A1 => n6365, A2 => n429, B1 => n5249, B2 => n4119
                           , ZN => n5566);
   U2977 : AOI22_X1 port map( A1 => n3911, A2 => net644629, B1 => n3912, B2 => 
                           net644500, ZN => n5567);
   U2975 : AOI22_X1 port map( A1 => n6367, A2 => n4012, B1 => n5245, B2 => n367
                           , ZN => n5568);
   U2974 : AOI22_X1 port map( A1 => n3913, A2 => net644597, B1 => n3914, B2 => 
                           net644693, ZN => n5569);
   U2973 : NAND4_X1 port map( A1 => n5566, A2 => n5567, A3 => n5568, A4 => 
                           n5569, ZN => n5560);
   U2971 : AOI22_X1 port map( A1 => n6369, A2 => n431, B1 => n5237, B2 => n4120
                           , ZN => n5562);
   U2970 : AOI22_X1 port map( A1 => n3910, A2 => net644789, B1 => n3909, B2 => 
                           net644757, ZN => n5563);
   U2969 : AOI22_X1 port map( A1 => n3908, A2 => net644919, B1 => n3907, B2 => 
                           net644436, ZN => n5564);
   U2967 : AOI22_X1 port map( A1 => n3906, A2 => n4013, B1 => n3905, B2 => n430
                           , ZN => n5565);
   U2966 : NAND4_X1 port map( A1 => n5562, A2 => n5563, A3 => n5564, A4 => 
                           n5565, ZN => n5561);
   U2965 : OAI21_X1 port map( B1 => n5560, B2 => n5561, A => n6370, ZN => n5559
                           );
   U2964 : OAI211_X1 port map( C1 => n560, C2 => n5220, A => n5558, B => n5559,
                           ZN => n5555);
   U2962 : AOI22_X1 port map( A1 => n6373, A2 => net644820, B1 => n6372, B2 => 
                           n4121, ZN => n5557);
   U2961 : OAI21_X1 port map( B1 => n622, B2 => n5216, A => n5557, ZN => n5556)
                           ;
   U2960 : AOI211_X1 port map( C1 => n5213, C2 => net644725, A => n5555, B => 
                           n5556, ZN => n5554);
   U2959 : NAND4_X1 port map( A1 => n5551, A2 => n5552, A3 => n5553, A4 => 
                           n5554, ZN => n2713);
   U3436 : AOI22_X1 port map( A1 => n6356, A2 => n3917, B1 => n6355, B2 => 
                           n3957, ZN => n5881);
   U3435 : AOI22_X1 port map( A1 => n6358, A2 => net644871, B1 => n5262, B2 => 
                           net644837, ZN => n5882);
   U3434 : AOI22_X1 port map( A1 => n6360, A2 => net644453, B1 => n6359, B2 => 
                           DATAIN(2), ZN => n5902);
   U3433 : OAI21_X1 port map( B1 => n5257, B2 => net644358, A => n5902, ZN => 
                           n5900);
   U3432 : OAI22_X1 port map( A1 => n544, A2 => n5255, B1 => n669, B2 => n5256,
                           ZN => n5901);
   U3431 : AOI211_X1 port map( C1 => n6361, C2 => net644645, A => n5900, B => 
                           n5901, ZN => n5883);
   U3430 : AOI22_X1 port map( A1 => n6363, A2 => net644517, B1 => n6362, B2 => 
                           net644549, ZN => n5888);
   U3428 : AOI22_X1 port map( A1 => n5248, A2 => n474, B1 => n6364, B2 => n4065
                           , ZN => n5896);
   U3427 : AOI22_X1 port map( A1 => n3911, A2 => net644614, B1 => n3912, B2 => 
                           net644485, ZN => n5897);
   U3425 : AOI22_X1 port map( A1 => n5244, A2 => n3958, B1 => n6366, B2 => n382
                           , ZN => n5898);
   U3424 : AOI22_X1 port map( A1 => n3913, A2 => net644582, B1 => n3914, B2 => 
                           net644678, ZN => n5899);
   U3423 : NAND4_X1 port map( A1 => n5896, A2 => n5897, A3 => n5898, A4 => 
                           n5899, ZN => n5890);
   U3421 : AOI22_X1 port map( A1 => n5236, A2 => n476, B1 => n6368, B2 => n4066
                           , ZN => n5892);
   U3420 : AOI22_X1 port map( A1 => n3910, A2 => net644774, B1 => n3909, B2 => 
                           net644742, ZN => n5893);
   U3419 : AOI22_X1 port map( A1 => n3908, A2 => net644904, B1 => n3907, B2 => 
                           net644421, ZN => n5894);
   U3417 : AOI22_X1 port map( A1 => n3906, A2 => n3960, B1 => n3905, B2 => n475
                           , ZN => n5895);
   U3416 : NAND4_X1 port map( A1 => n5892, A2 => n5893, A3 => n5894, A4 => 
                           n5895, ZN => n5891);
   U3415 : OAI21_X1 port map( B1 => n5890, B2 => n5891, A => n6370, ZN => n5889
                           );
   U3414 : OAI211_X1 port map( C1 => n575, C2 => n5220, A => n5888, B => n5889,
                           ZN => n5885);
   U3412 : AOI22_X1 port map( A1 => n6373, A2 => net644805, B1 => n6372, B2 => 
                           n4067, ZN => n5887);
   U3411 : OAI21_X1 port map( B1 => n637, B2 => n5216, A => n5887, ZN => n5886)
                           ;
   U3410 : AOI211_X1 port map( C1 => n6374, C2 => net644710, A => n5885, B => 
                           n5886, ZN => n5884);
   U3409 : NAND4_X1 port map( A1 => n5881, A2 => n5882, A3 => n5883, A4 => 
                           n5884, ZN => n2698);
   U3136 : AOI22_X1 port map( A1 => n6356, A2 => n3930, B1 => n6355, B2 => 
                           n3990, ZN => n5661);
   U3135 : AOI22_X1 port map( A1 => n6358, A2 => net644881, B1 => n6357, B2 => 
                           net644847, ZN => n5662);
   U3134 : AOI22_X1 port map( A1 => n6360, A2 => net644463, B1 => n6359, B2 => 
                           DATAIN(12), ZN => n5682);
   U3133 : OAI21_X1 port map( B1 => n5257, B2 => net644368, A => n5682, ZN => 
                           n5680);
   U3132 : OAI22_X1 port map( A1 => n534, A2 => n5255, B1 => n659, B2 => n5256,
                           ZN => n5681);
   U3131 : AOI211_X1 port map( C1 => n6361, C2 => net644655, A => n5680, B => 
                           n5681, ZN => n5663);
   U3130 : AOI22_X1 port map( A1 => n6363, A2 => net644527, B1 => n6362, B2 => 
                           net644559, ZN => n5668);
   U3128 : AOI22_X1 port map( A1 => n6365, A2 => n444, B1 => n6364, B2 => n4099
                           , ZN => n5676);
   U3127 : AOI22_X1 port map( A1 => n3911, A2 => net644624, B1 => n3912, B2 => 
                           net644495, ZN => n5677);
   U3125 : AOI22_X1 port map( A1 => n6367, A2 => n3991, B1 => n6366, B2 => n372
                           , ZN => n5678);
   U3124 : AOI22_X1 port map( A1 => n3913, A2 => net644592, B1 => n3914, B2 => 
                           net644688, ZN => n5679);
   U3123 : NAND4_X1 port map( A1 => n5676, A2 => n5677, A3 => n5678, A4 => 
                           n5679, ZN => n5670);
   U3121 : AOI22_X1 port map( A1 => n6369, A2 => n446, B1 => n6368, B2 => n4100
                           , ZN => n5672);
   U3120 : AOI22_X1 port map( A1 => n3910, A2 => net644784, B1 => n3909, B2 => 
                           net644752, ZN => n5673);
   U3119 : AOI22_X1 port map( A1 => n3908, A2 => net644914, B1 => n3907, B2 => 
                           net644431, ZN => n5674);
   U3117 : AOI22_X1 port map( A1 => n3906, A2 => n3992, B1 => n3905, B2 => n445
                           , ZN => n5675);
   U3116 : NAND4_X1 port map( A1 => n5672, A2 => n5673, A3 => n5674, A4 => 
                           n5675, ZN => n5671);
   U3115 : OAI21_X1 port map( B1 => n5670, B2 => n5671, A => n5225, ZN => n5669
                           );
   U3114 : OAI211_X1 port map( C1 => n565, C2 => n5220, A => n5668, B => n5669,
                           ZN => n5665);
   U3112 : AOI22_X1 port map( A1 => n6373, A2 => net644815, B1 => n6372, B2 => 
                           n4101, ZN => n5667);
   U3111 : OAI21_X1 port map( B1 => n627, B2 => n5216, A => n5667, ZN => n5666)
                           ;
   U3110 : AOI211_X1 port map( C1 => n6374, C2 => net644720, A => n5665, B => 
                           n5666, ZN => n5664);
   U3109 : NAND4_X1 port map( A1 => n5661, A2 => n5662, A3 => n5663, A4 => 
                           n5664, ZN => n2708);
   U3196 : AOI22_X1 port map( A1 => n6356, A2 => n3928, B1 => n6355, B2 => 
                           n3984, ZN => n5705);
   U3195 : AOI22_X1 port map( A1 => n6358, A2 => net644879, B1 => n6357, B2 => 
                           net644845, ZN => n5706);
   U3194 : AOI22_X1 port map( A1 => n6360, A2 => net644461, B1 => n6359, B2 => 
                           DATAIN(10), ZN => n5726);
   U3193 : OAI21_X1 port map( B1 => n5257, B2 => net644366, A => n5726, ZN => 
                           n5724);
   U3192 : OAI22_X1 port map( A1 => n536, A2 => n5255, B1 => n661, B2 => n5256,
                           ZN => n5725);
   U3191 : AOI211_X1 port map( C1 => n6361, C2 => net644653, A => n5724, B => 
                           n5725, ZN => n5707);
   U3190 : AOI22_X1 port map( A1 => n6363, A2 => net644525, B1 => n6362, B2 => 
                           net644557, ZN => n5712);
   U3188 : AOI22_X1 port map( A1 => n6365, A2 => n450, B1 => n6364, B2 => n4093
                           , ZN => n5720);
   U3187 : AOI22_X1 port map( A1 => n3911, A2 => net644622, B1 => n3912, B2 => 
                           net644493, ZN => n5721);
   U3185 : AOI22_X1 port map( A1 => n6367, A2 => n3985, B1 => n6366, B2 => n374
                           , ZN => n5722);
   U3184 : AOI22_X1 port map( A1 => n3913, A2 => net644590, B1 => n3914, B2 => 
                           net644686, ZN => n5723);
   U3183 : NAND4_X1 port map( A1 => n5720, A2 => n5721, A3 => n5722, A4 => 
                           n5723, ZN => n5714);
   U3181 : AOI22_X1 port map( A1 => n6369, A2 => n452, B1 => n6368, B2 => n4094
                           , ZN => n5716);
   U3180 : AOI22_X1 port map( A1 => n3910, A2 => net644782, B1 => n3909, B2 => 
                           net644750, ZN => n5717);
   U3179 : AOI22_X1 port map( A1 => n3908, A2 => net644912, B1 => n3907, B2 => 
                           net644429, ZN => n5718);
   U3177 : AOI22_X1 port map( A1 => n3906, A2 => n3986, B1 => n3905, B2 => n451
                           , ZN => n5719);
   U3176 : NAND4_X1 port map( A1 => n5716, A2 => n5717, A3 => n5718, A4 => 
                           n5719, ZN => n5715);
   U3175 : OAI21_X1 port map( B1 => n5714, B2 => n5715, A => n6370, ZN => n5713
                           );
   U3174 : OAI211_X1 port map( C1 => n567, C2 => n5220, A => n5712, B => n5713,
                           ZN => n5709);
   U3172 : AOI22_X1 port map( A1 => n6373, A2 => net644813, B1 => n6372, B2 => 
                           n4095, ZN => n5711);
   U3171 : OAI21_X1 port map( B1 => n629, B2 => n5216, A => n5711, ZN => n5710)
                           ;
   U3170 : AOI211_X1 port map( C1 => n6374, C2 => net644718, A => n5709, B => 
                           n5710, ZN => n5708);
   U3169 : NAND4_X1 port map( A1 => n5705, A2 => n5706, A3 => n5707, A4 => 
                           n5708, ZN => n2706);
   U3166 : AOI22_X1 port map( A1 => n6356, A2 => n3929, B1 => n6355, B2 => 
                           n3987, ZN => n5683);
   U3165 : AOI22_X1 port map( A1 => n6358, A2 => net644880, B1 => n6357, B2 => 
                           net644846, ZN => n5684);
   U3164 : AOI22_X1 port map( A1 => n6360, A2 => net644462, B1 => n6359, B2 => 
                           DATAIN(11), ZN => n5704);
   U3163 : OAI21_X1 port map( B1 => n5257, B2 => net644367, A => n5704, ZN => 
                           n5702);
   U3162 : OAI22_X1 port map( A1 => n535, A2 => n5255, B1 => n660, B2 => n5256,
                           ZN => n5703);
   U3161 : AOI211_X1 port map( C1 => n6361, C2 => net644654, A => n5702, B => 
                           n5703, ZN => n5685);
   U3160 : AOI22_X1 port map( A1 => n6363, A2 => net644526, B1 => n6362, B2 => 
                           net644558, ZN => n5690);
   U3158 : AOI22_X1 port map( A1 => n6365, A2 => n447, B1 => n6364, B2 => n4096
                           , ZN => n5698);
   U3157 : AOI22_X1 port map( A1 => n3911, A2 => net644623, B1 => n3912, B2 => 
                           net644494, ZN => n5699);
   U3155 : AOI22_X1 port map( A1 => n6367, A2 => n3988, B1 => n6366, B2 => n373
                           , ZN => n5700);
   U3154 : AOI22_X1 port map( A1 => n3913, A2 => net644591, B1 => n3914, B2 => 
                           net644687, ZN => n5701);
   U3153 : NAND4_X1 port map( A1 => n5698, A2 => n5699, A3 => n5700, A4 => 
                           n5701, ZN => n5692);
   U3151 : AOI22_X1 port map( A1 => n6369, A2 => n449, B1 => n6368, B2 => n4097
                           , ZN => n5694);
   U3150 : AOI22_X1 port map( A1 => n3910, A2 => net644783, B1 => n3909, B2 => 
                           net644751, ZN => n5695);
   U3149 : AOI22_X1 port map( A1 => n3908, A2 => net644913, B1 => n3907, B2 => 
                           net644430, ZN => n5696);
   U3147 : AOI22_X1 port map( A1 => n3906, A2 => n3989, B1 => n3905, B2 => n448
                           , ZN => n5697);
   U3146 : NAND4_X1 port map( A1 => n5694, A2 => n5695, A3 => n5696, A4 => 
                           n5697, ZN => n5693);
   U3145 : OAI21_X1 port map( B1 => n5692, B2 => n5693, A => n6370, ZN => n5691
                           );
   U3144 : OAI211_X1 port map( C1 => n566, C2 => n5220, A => n5690, B => n5691,
                           ZN => n5687);
   U3142 : AOI22_X1 port map( A1 => n6373, A2 => net644814, B1 => n6372, B2 => 
                           n4098, ZN => n5689);
   U3141 : OAI21_X1 port map( B1 => n628, B2 => n5216, A => n5689, ZN => n5688)
                           ;
   U3140 : AOI211_X1 port map( C1 => n6374, C2 => net644719, A => n5687, B => 
                           n5688, ZN => n5686);
   U3139 : NAND4_X1 port map( A1 => n5683, A2 => n5684, A3 => n5685, A4 => 
                           n5686, ZN => n2707);
   U3406 : AOI22_X1 port map( A1 => n6356, A2 => n3918, B1 => n6355, B2 => 
                           n3963, ZN => n5859);
   U3405 : AOI22_X1 port map( A1 => n6358, A2 => net644872, B1 => n5262, B2 => 
                           net644838, ZN => n5860);
   U3404 : AOI22_X1 port map( A1 => n6360, A2 => net644454, B1 => n6359, B2 => 
                           DATAIN(3), ZN => n5880);
   U3403 : OAI21_X1 port map( B1 => n5257, B2 => net644359, A => n5880, ZN => 
                           n5878);
   U3402 : OAI22_X1 port map( A1 => n543, A2 => n5255, B1 => n668, B2 => n5256,
                           ZN => n5879);
   U3401 : AOI211_X1 port map( C1 => n6361, C2 => net644646, A => n5878, B => 
                           n5879, ZN => n5861);
   U3400 : AOI22_X1 port map( A1 => n6363, A2 => net644518, B1 => n6362, B2 => 
                           net644550, ZN => n5866);
   U3398 : AOI22_X1 port map( A1 => n5248, A2 => n471, B1 => n6364, B2 => n4070
                           , ZN => n5874);
   U3397 : AOI22_X1 port map( A1 => n3911, A2 => net644615, B1 => n3912, B2 => 
                           net644486, ZN => n5875);
   U3395 : AOI22_X1 port map( A1 => n5244, A2 => n3964, B1 => n6366, B2 => n381
                           , ZN => n5876);
   U3394 : AOI22_X1 port map( A1 => n3913, A2 => net644583, B1 => n3914, B2 => 
                           net644679, ZN => n5877);
   U3393 : NAND4_X1 port map( A1 => n5874, A2 => n5875, A3 => n5876, A4 => 
                           n5877, ZN => n5868);
   U3391 : AOI22_X1 port map( A1 => n5236, A2 => n473, B1 => n6368, B2 => n4071
                           , ZN => n5870);
   U3390 : AOI22_X1 port map( A1 => n3910, A2 => net644775, B1 => n3909, B2 => 
                           net644743, ZN => n5871);
   U3389 : AOI22_X1 port map( A1 => n3908, A2 => net644905, B1 => n3907, B2 => 
                           net644422, ZN => n5872);
   U3387 : AOI22_X1 port map( A1 => n3906, A2 => n3965, B1 => n3905, B2 => n472
                           , ZN => n5873);
   U3386 : NAND4_X1 port map( A1 => n5870, A2 => n5871, A3 => n5872, A4 => 
                           n5873, ZN => n5869);
   U3385 : OAI21_X1 port map( B1 => n5868, B2 => n5869, A => n6370, ZN => n5867
                           );
   U3384 : OAI211_X1 port map( C1 => n574, C2 => n5220, A => n5866, B => n5867,
                           ZN => n5863);
   U3382 : AOI22_X1 port map( A1 => n6373, A2 => net644806, B1 => n6372, B2 => 
                           n4072, ZN => n5865);
   U3381 : OAI21_X1 port map( B1 => n636, B2 => n5216, A => n5865, ZN => n5864)
                           ;
   U3380 : AOI211_X1 port map( C1 => n6374, C2 => net644711, A => n5863, B => 
                           n5864, ZN => n5862);
   U3379 : NAND4_X1 port map( A1 => n5859, A2 => n5860, A3 => n5861, A4 => 
                           n5862, ZN => n2699);
   U2926 : AOI22_X1 port map( A1 => n5263, A2 => n3937, B1 => n6355, B2 => 
                           n4017, ZN => n5507);
   U2925 : AOI22_X1 port map( A1 => n5261, A2 => net644888, B1 => n6357, B2 => 
                           net644854, ZN => n5508);
   U2924 : AOI22_X1 port map( A1 => n6360, A2 => net644470, B1 => n6359, B2 => 
                           DATAIN(19), ZN => n5528);
   U2923 : OAI21_X1 port map( B1 => n5257, B2 => net644375, A => n5528, ZN => 
                           n5526);
   U2922 : OAI22_X1 port map( A1 => n527, A2 => n5255, B1 => n652, B2 => n5256,
                           ZN => n5527);
   U2921 : AOI211_X1 port map( C1 => n6361, C2 => net644662, A => n5526, B => 
                           n5527, ZN => n5509);
   U2920 : AOI22_X1 port map( A1 => n6363, A2 => net644534, B1 => n6362, B2 => 
                           net644566, ZN => n5514);
   U2918 : AOI22_X1 port map( A1 => n6365, A2 => n423, B1 => n6364, B2 => n4125
                           , ZN => n5522);
   U2917 : AOI22_X1 port map( A1 => n3911, A2 => net644631, B1 => n3912, B2 => 
                           net644502, ZN => n5523);
   U2915 : AOI22_X1 port map( A1 => n6367, A2 => n4018, B1 => n6366, B2 => n365
                           , ZN => n5524);
   U2914 : AOI22_X1 port map( A1 => n3913, A2 => net644599, B1 => n3914, B2 => 
                           net644695, ZN => n5525);
   U2913 : NAND4_X1 port map( A1 => n5522, A2 => n5523, A3 => n5524, A4 => 
                           n5525, ZN => n5516);
   U2911 : AOI22_X1 port map( A1 => n6369, A2 => n425, B1 => n6368, B2 => n4126
                           , ZN => n5518);
   U2910 : AOI22_X1 port map( A1 => n3910, A2 => net644791, B1 => n3909, B2 => 
                           net644759, ZN => n5519);
   U2909 : AOI22_X1 port map( A1 => n3908, A2 => net644921, B1 => n3907, B2 => 
                           net644438, ZN => n5520);
   U2907 : AOI22_X1 port map( A1 => n3906, A2 => n4019, B1 => n3905, B2 => n424
                           , ZN => n5521);
   U2906 : NAND4_X1 port map( A1 => n5518, A2 => n5519, A3 => n5520, A4 => 
                           n5521, ZN => n5517);
   U2905 : OAI21_X1 port map( B1 => n5516, B2 => n5517, A => n6370, ZN => n5515
                           );
   U2904 : OAI211_X1 port map( C1 => n558, C2 => n5220, A => n5514, B => n5515,
                           ZN => n5511);
   U2902 : AOI22_X1 port map( A1 => n6373, A2 => net644822, B1 => n6372, B2 => 
                           n4127, ZN => n5513);
   U2901 : OAI21_X1 port map( B1 => n620, B2 => n5216, A => n5513, ZN => n5512)
                           ;
   U2900 : AOI211_X1 port map( C1 => n6374, C2 => net644727, A => n5511, B => 
                           n5512, ZN => n5510);
   U2899 : NAND4_X1 port map( A1 => n5507, A2 => n5508, A3 => n5509, A4 => 
                           n5510, ZN => n2715);
   U2896 : AOI22_X1 port map( A1 => n6356, A2 => n3938, B1 => n6355, B2 => 
                           n4020, ZN => n5485);
   U2895 : AOI22_X1 port map( A1 => n6358, A2 => net644889, B1 => n6357, B2 => 
                           net644855, ZN => n5486);
   U2894 : AOI22_X1 port map( A1 => n6360, A2 => net644471, B1 => n6359, B2 => 
                           DATAIN(20), ZN => n5506);
   U2893 : OAI21_X1 port map( B1 => n5257, B2 => net644376, A => n5506, ZN => 
                           n5504);
   U2892 : OAI22_X1 port map( A1 => n526, A2 => n5255, B1 => n651, B2 => n5256,
                           ZN => n5505);
   U2891 : AOI211_X1 port map( C1 => n6361, C2 => net644663, A => n5504, B => 
                           n5505, ZN => n5487);
   U2890 : AOI22_X1 port map( A1 => n6363, A2 => net644535, B1 => n6362, B2 => 
                           net644567, ZN => n5492);
   U2888 : AOI22_X1 port map( A1 => n6365, A2 => n420, B1 => n6364, B2 => n4128
                           , ZN => n5500);
   U2887 : AOI22_X1 port map( A1 => n3911, A2 => net644632, B1 => n3912, B2 => 
                           net644503, ZN => n5501);
   U2885 : AOI22_X1 port map( A1 => n6367, A2 => n4021, B1 => n6366, B2 => n364
                           , ZN => n5502);
   U2884 : AOI22_X1 port map( A1 => n3913, A2 => net644600, B1 => n3914, B2 => 
                           net644696, ZN => n5503);
   U2883 : NAND4_X1 port map( A1 => n5500, A2 => n5501, A3 => n5502, A4 => 
                           n5503, ZN => n5494);
   U2881 : AOI22_X1 port map( A1 => n6369, A2 => n422, B1 => n6368, B2 => n4129
                           , ZN => n5496);
   U2880 : AOI22_X1 port map( A1 => n3910, A2 => net644792, B1 => n3909, B2 => 
                           net644760, ZN => n5497);
   U2879 : AOI22_X1 port map( A1 => n3908, A2 => net644922, B1 => n3907, B2 => 
                           net644439, ZN => n5498);
   U2877 : AOI22_X1 port map( A1 => n3906, A2 => n4022, B1 => n3905, B2 => n421
                           , ZN => n5499);
   U2876 : NAND4_X1 port map( A1 => n5496, A2 => n5497, A3 => n5498, A4 => 
                           n5499, ZN => n5495);
   U2875 : OAI21_X1 port map( B1 => n5494, B2 => n5495, A => n6370, ZN => n5493
                           );
   U2874 : OAI211_X1 port map( C1 => n557, C2 => n5220, A => n5492, B => n5493,
                           ZN => n5489);
   U2872 : AOI22_X1 port map( A1 => n6373, A2 => net644823, B1 => n6372, B2 => 
                           n4130, ZN => n5491);
   U2871 : OAI21_X1 port map( B1 => n619, B2 => n5216, A => n5491, ZN => n5490)
                           ;
   U2870 : AOI211_X1 port map( C1 => n6374, C2 => net644728, A => n5489, B => 
                           n5490, ZN => n5488);
   U2869 : NAND4_X1 port map( A1 => n5485, A2 => n5486, A3 => n5487, A4 => 
                           n5488, ZN => n2716);
   U2956 : AOI22_X1 port map( A1 => n6356, A2 => n3936, B1 => n5264, B2 => 
                           n4014, ZN => n5529);
   U2955 : AOI22_X1 port map( A1 => n5261, A2 => net644887, B1 => n6357, B2 => 
                           net644853, ZN => n5530);
   U2954 : AOI22_X1 port map( A1 => n6360, A2 => net644469, B1 => n6359, B2 => 
                           DATAIN(18), ZN => n5550);
   U2953 : OAI21_X1 port map( B1 => n5257, B2 => net644374, A => n5550, ZN => 
                           n5548);
   U2952 : OAI22_X1 port map( A1 => n528, A2 => n5255, B1 => n653, B2 => n5256,
                           ZN => n5549);
   U2951 : AOI211_X1 port map( C1 => n6361, C2 => net644661, A => n5548, B => 
                           n5549, ZN => n5531);
   U2950 : AOI22_X1 port map( A1 => n6363, A2 => net644533, B1 => n5251, B2 => 
                           net644565, ZN => n5536);
   U2948 : AOI22_X1 port map( A1 => n6365, A2 => n426, B1 => n5249, B2 => n4122
                           , ZN => n5544);
   U2947 : AOI22_X1 port map( A1 => n3911, A2 => net644630, B1 => n3912, B2 => 
                           net644501, ZN => n5545);
   U2945 : AOI22_X1 port map( A1 => n6367, A2 => n4015, B1 => n5245, B2 => n366
                           , ZN => n5546);
   U2944 : AOI22_X1 port map( A1 => n3913, A2 => net644598, B1 => n3914, B2 => 
                           net644694, ZN => n5547);
   U2943 : NAND4_X1 port map( A1 => n5544, A2 => n5545, A3 => n5546, A4 => 
                           n5547, ZN => n5538);
   U2941 : AOI22_X1 port map( A1 => n6369, A2 => n428, B1 => n5237, B2 => n4123
                           , ZN => n5540);
   U2940 : AOI22_X1 port map( A1 => n3910, A2 => net644790, B1 => n3909, B2 => 
                           net644758, ZN => n5541);
   U2939 : AOI22_X1 port map( A1 => n3908, A2 => net644920, B1 => n3907, B2 => 
                           net644437, ZN => n5542);
   U2937 : AOI22_X1 port map( A1 => n3906, A2 => n4016, B1 => n3905, B2 => n427
                           , ZN => n5543);
   U2936 : NAND4_X1 port map( A1 => n5540, A2 => n5541, A3 => n5542, A4 => 
                           n5543, ZN => n5539);
   U2935 : OAI21_X1 port map( B1 => n5538, B2 => n5539, A => n6370, ZN => n5537
                           );
   U2934 : OAI211_X1 port map( C1 => n559, C2 => n5220, A => n5536, B => n5537,
                           ZN => n5533);
   U2932 : AOI22_X1 port map( A1 => n6373, A2 => net644821, B1 => n6372, B2 => 
                           n4124, ZN => n5535);
   U2931 : OAI21_X1 port map( B1 => n621, B2 => n5216, A => n5535, ZN => n5534)
                           ;
   U2930 : AOI211_X1 port map( C1 => n6374, C2 => net644726, A => n5533, B => 
                           n5534, ZN => n5532);
   U2929 : NAND4_X1 port map( A1 => n5529, A2 => n5530, A3 => n5531, A4 => 
                           n5532, ZN => n2714);
   U2776 : AOI22_X1 port map( A1 => n6356, A2 => n3942, B1 => n5264, B2 => 
                           n4032, ZN => n5397);
   U2775 : AOI22_X1 port map( A1 => n6358, A2 => net644893, B1 => n5262, B2 => 
                           net644859, ZN => n5398);
   U2774 : AOI22_X1 port map( A1 => n6360, A2 => net644475, B1 => n6359, B2 => 
                           DATAIN(24), ZN => n5418);
   U2773 : OAI21_X1 port map( B1 => n5257, B2 => net644380, A => n5418, ZN => 
                           n5416);
   U2772 : OAI22_X1 port map( A1 => n522, A2 => n5255, B1 => n647, B2 => n5256,
                           ZN => n5417);
   U2771 : AOI211_X1 port map( C1 => n6361, C2 => net644667, A => n5416, B => 
                           n5417, ZN => n5399);
   U2770 : AOI22_X1 port map( A1 => n6363, A2 => net644539, B1 => n6362, B2 => 
                           net644571, ZN => n5404);
   U2768 : AOI22_X1 port map( A1 => n6365, A2 => n408, B1 => n5249, B2 => n4140
                           , ZN => n5412);
   U2767 : AOI22_X1 port map( A1 => n3911, A2 => net644636, B1 => n3912, B2 => 
                           net644507, ZN => n5413);
   U2765 : AOI22_X1 port map( A1 => n6367, A2 => n4034, B1 => n5245, B2 => n360
                           , ZN => n5414);
   U2764 : AOI22_X1 port map( A1 => n3913, A2 => net644604, B1 => n3914, B2 => 
                           net644700, ZN => n5415);
   U2763 : NAND4_X1 port map( A1 => n5412, A2 => n5413, A3 => n5414, A4 => 
                           n5415, ZN => n5406);
   U2761 : AOI22_X1 port map( A1 => n6369, A2 => n410, B1 => n5237, B2 => n4141
                           , ZN => n5408);
   U2760 : AOI22_X1 port map( A1 => n3910, A2 => net644796, B1 => n3909, B2 => 
                           net644764, ZN => n5409);
   U2759 : AOI22_X1 port map( A1 => n3908, A2 => net644926, B1 => n3907, B2 => 
                           net644443, ZN => n5410);
   U2757 : AOI22_X1 port map( A1 => n3906, A2 => n4037, B1 => n3905, B2 => n409
                           , ZN => n5411);
   U2756 : NAND4_X1 port map( A1 => n5408, A2 => n5409, A3 => n5410, A4 => 
                           n5411, ZN => n5407);
   U2755 : OAI21_X1 port map( B1 => n5406, B2 => n5407, A => n6370, ZN => n5405
                           );
   U2754 : OAI211_X1 port map( C1 => n553, C2 => n5220, A => n5404, B => n5405,
                           ZN => n5401);
   U2752 : AOI22_X1 port map( A1 => n6373, A2 => net644827, B1 => n6372, B2 => 
                           n4142, ZN => n5403);
   U2751 : OAI21_X1 port map( B1 => n615, B2 => n5216, A => n5403, ZN => n5402)
                           ;
   U2750 : AOI211_X1 port map( C1 => n5213, C2 => net644732, A => n5401, B => 
                           n5402, ZN => n5400);
   U2749 : NAND4_X1 port map( A1 => n5397, A2 => n5398, A3 => n5399, A4 => 
                           n5400, ZN => n2720);
   U2866 : AOI22_X1 port map( A1 => n6356, A2 => n3939, B1 => n6355, B2 => 
                           n4023, ZN => n5463);
   U2865 : AOI22_X1 port map( A1 => n6358, A2 => net644890, B1 => n6357, B2 => 
                           net644856, ZN => n5464);
   U2864 : AOI22_X1 port map( A1 => n6360, A2 => net644472, B1 => n6359, B2 => 
                           DATAIN(21), ZN => n5484);
   U2863 : OAI21_X1 port map( B1 => n5257, B2 => net644377, A => n5484, ZN => 
                           n5482);
   U2862 : OAI22_X1 port map( A1 => n525, A2 => n5255, B1 => n650, B2 => n5256,
                           ZN => n5483);
   U2861 : AOI211_X1 port map( C1 => n6361, C2 => net644664, A => n5482, B => 
                           n5483, ZN => n5465);
   U2860 : AOI22_X1 port map( A1 => n6363, A2 => net644536, B1 => n6362, B2 => 
                           net644568, ZN => n5470);
   U2858 : AOI22_X1 port map( A1 => n6365, A2 => n417, B1 => n6364, B2 => n4131
                           , ZN => n5478);
   U2857 : AOI22_X1 port map( A1 => n3911, A2 => net644633, B1 => n3912, B2 => 
                           net644504, ZN => n5479);
   U2855 : AOI22_X1 port map( A1 => n6367, A2 => n4024, B1 => n6366, B2 => n363
                           , ZN => n5480);
   U2854 : AOI22_X1 port map( A1 => n3913, A2 => net644601, B1 => n3914, B2 => 
                           net644697, ZN => n5481);
   U2853 : NAND4_X1 port map( A1 => n5478, A2 => n5479, A3 => n5480, A4 => 
                           n5481, ZN => n5472);
   U2851 : AOI22_X1 port map( A1 => n6369, A2 => n419, B1 => n6368, B2 => n4132
                           , ZN => n5474);
   U2850 : AOI22_X1 port map( A1 => n3910, A2 => net644793, B1 => n3909, B2 => 
                           net644761, ZN => n5475);
   U2849 : AOI22_X1 port map( A1 => n3908, A2 => net644923, B1 => n3907, B2 => 
                           net644440, ZN => n5476);
   U2847 : AOI22_X1 port map( A1 => n3906, A2 => n4025, B1 => n3905, B2 => n418
                           , ZN => n5477);
   U2846 : NAND4_X1 port map( A1 => n5474, A2 => n5475, A3 => n5476, A4 => 
                           n5477, ZN => n5473);
   U2845 : OAI21_X1 port map( B1 => n5472, B2 => n5473, A => n6370, ZN => n5471
                           );
   U2844 : OAI211_X1 port map( C1 => n556, C2 => n5220, A => n5470, B => n5471,
                           ZN => n5467);
   U2842 : AOI22_X1 port map( A1 => n6373, A2 => net644824, B1 => n6372, B2 => 
                           n4133, ZN => n5469);
   U2841 : OAI21_X1 port map( B1 => n618, B2 => n5216, A => n5469, ZN => n5468)
                           ;
   U2840 : AOI211_X1 port map( C1 => n6374, C2 => net644729, A => n5467, B => 
                           n5468, ZN => n5466);
   U2839 : NAND4_X1 port map( A1 => n5463, A2 => n5464, A3 => n5465, A4 => 
                           n5466, ZN => n2717);
   U3016 : AOI22_X1 port map( A1 => n6356, A2 => n3934, B1 => n5264, B2 => 
                           n4008, ZN => n5573);
   U3015 : AOI22_X1 port map( A1 => n6358, A2 => net644885, B1 => n6357, B2 => 
                           net644851, ZN => n5574);
   U3014 : AOI22_X1 port map( A1 => n6360, A2 => net644467, B1 => n6359, B2 => 
                           DATAIN(16), ZN => n5594);
   U3013 : OAI21_X1 port map( B1 => n5257, B2 => net644372, A => n5594, ZN => 
                           n5592);
   U3012 : OAI22_X1 port map( A1 => n530, A2 => n5255, B1 => n655, B2 => n5256,
                           ZN => n5593);
   U3011 : AOI211_X1 port map( C1 => n6361, C2 => net644659, A => n5592, B => 
                           n5593, ZN => n5575);
   U3010 : AOI22_X1 port map( A1 => n6363, A2 => net644531, B1 => n6362, B2 => 
                           net644563, ZN => n5580);
   U3008 : AOI22_X1 port map( A1 => n6365, A2 => n432, B1 => n5249, B2 => n4116
                           , ZN => n5588);
   U3007 : AOI22_X1 port map( A1 => n3911, A2 => net644628, B1 => n3912, B2 => 
                           net644499, ZN => n5589);
   U3005 : AOI22_X1 port map( A1 => n6367, A2 => n4009, B1 => n5245, B2 => n368
                           , ZN => n5590);
   U3004 : AOI22_X1 port map( A1 => n3913, A2 => net644596, B1 => n3914, B2 => 
                           net644692, ZN => n5591);
   U3003 : NAND4_X1 port map( A1 => n5588, A2 => n5589, A3 => n5590, A4 => 
                           n5591, ZN => n5582);
   U3001 : AOI22_X1 port map( A1 => n6369, A2 => n434, B1 => n5237, B2 => n4117
                           , ZN => n5584);
   U3000 : AOI22_X1 port map( A1 => n3910, A2 => net644788, B1 => n3909, B2 => 
                           net644756, ZN => n5585);
   U2999 : AOI22_X1 port map( A1 => n3908, A2 => net644918, B1 => n3907, B2 => 
                           net644435, ZN => n5586);
   U2997 : AOI22_X1 port map( A1 => n3906, A2 => n4010, B1 => n3905, B2 => n433
                           , ZN => n5587);
   U2996 : NAND4_X1 port map( A1 => n5584, A2 => n5585, A3 => n5586, A4 => 
                           n5587, ZN => n5583);
   U2995 : OAI21_X1 port map( B1 => n5582, B2 => n5583, A => n6370, ZN => n5581
                           );
   U2994 : OAI211_X1 port map( C1 => n561, C2 => n5220, A => n5580, B => n5581,
                           ZN => n5577);
   U2992 : AOI22_X1 port map( A1 => n6373, A2 => net644819, B1 => n6372, B2 => 
                           n4118, ZN => n5579);
   U2991 : OAI21_X1 port map( B1 => n623, B2 => n5216, A => n5579, ZN => n5578)
                           ;
   U2990 : AOI211_X1 port map( C1 => n5213, C2 => net644724, A => n5577, B => 
                           n5578, ZN => n5576);
   U2989 : NAND4_X1 port map( A1 => n5573, A2 => n5574, A3 => n5575, A4 => 
                           n5576, ZN => n2712);
   U3256 : AOI22_X1 port map( A1 => n6356, A2 => n3923, B1 => n6355, B2 => 
                           n3978, ZN => n5749);
   U3255 : AOI22_X1 port map( A1 => n6358, A2 => net644877, B1 => n6357, B2 => 
                           net644843, ZN => n5750);
   U3254 : AOI22_X1 port map( A1 => n6360, A2 => net644459, B1 => n6359, B2 => 
                           DATAIN(8), ZN => n5770);
   U3253 : OAI21_X1 port map( B1 => n5257, B2 => net644364, A => n5770, ZN => 
                           n5768);
   U3252 : OAI22_X1 port map( A1 => n538, A2 => n5255, B1 => n663, B2 => n5256,
                           ZN => n5769);
   U3251 : AOI211_X1 port map( C1 => n6361, C2 => net644651, A => n5768, B => 
                           n5769, ZN => n5751);
   U3250 : AOI22_X1 port map( A1 => n6363, A2 => net644523, B1 => n6362, B2 => 
                           net644555, ZN => n5756);
   U3248 : AOI22_X1 port map( A1 => n6365, A2 => n456, B1 => n6364, B2 => n4087
                           , ZN => n5764);
   U3247 : AOI22_X1 port map( A1 => n3911, A2 => net644620, B1 => n3912, B2 => 
                           net644491, ZN => n5765);
   U3245 : AOI22_X1 port map( A1 => n6367, A2 => n3979, B1 => n6366, B2 => n376
                           , ZN => n5766);
   U3244 : AOI22_X1 port map( A1 => n3913, A2 => net644588, B1 => n3914, B2 => 
                           net644684, ZN => n5767);
   U3243 : NAND4_X1 port map( A1 => n5764, A2 => n5765, A3 => n5766, A4 => 
                           n5767, ZN => n5758);
   U3241 : AOI22_X1 port map( A1 => n6369, A2 => n458, B1 => n6368, B2 => n4088
                           , ZN => n5760);
   U3240 : AOI22_X1 port map( A1 => n3910, A2 => net644780, B1 => n3909, B2 => 
                           net644748, ZN => n5761);
   U3239 : AOI22_X1 port map( A1 => n3908, A2 => net644910, B1 => n3907, B2 => 
                           net644427, ZN => n5762);
   U3237 : AOI22_X1 port map( A1 => n3906, A2 => n3980, B1 => n3905, B2 => n457
                           , ZN => n5763);
   U3236 : NAND4_X1 port map( A1 => n5760, A2 => n5761, A3 => n5762, A4 => 
                           n5763, ZN => n5759);
   U3235 : OAI21_X1 port map( B1 => n5758, B2 => n5759, A => n6370, ZN => n5757
                           );
   U3234 : OAI211_X1 port map( C1 => n569, C2 => n5220, A => n5756, B => n5757,
                           ZN => n5753);
   U3232 : AOI22_X1 port map( A1 => n6373, A2 => net644811, B1 => n6372, B2 => 
                           n4089, ZN => n5755);
   U3231 : OAI21_X1 port map( B1 => n631, B2 => n5216, A => n5755, ZN => n5754)
                           ;
   U3230 : AOI211_X1 port map( C1 => n6374, C2 => net644716, A => n5753, B => 
                           n5754, ZN => n5752);
   U3229 : NAND4_X1 port map( A1 => n5749, A2 => n5750, A3 => n5751, A4 => 
                           n5752, ZN => n2704);
   U3316 : AOI22_X1 port map( A1 => n6356, A2 => n3921, B1 => n6355, B2 => 
                           n3972, ZN => n5793);
   U3315 : AOI22_X1 port map( A1 => n6358, A2 => net644875, B1 => n5262, B2 => 
                           net644841, ZN => n5794);
   U3314 : AOI22_X1 port map( A1 => n6360, A2 => net644457, B1 => n6359, B2 => 
                           DATAIN(6), ZN => n5814);
   U3313 : OAI21_X1 port map( B1 => n5257, B2 => net644362, A => n5814, ZN => 
                           n5812);
   U3312 : OAI22_X1 port map( A1 => n540, A2 => n5255, B1 => n665, B2 => n5256,
                           ZN => n5813);
   U3311 : AOI211_X1 port map( C1 => n6361, C2 => net644649, A => n5812, B => 
                           n5813, ZN => n5795);
   U3310 : AOI22_X1 port map( A1 => n6363, A2 => net644521, B1 => n6362, B2 => 
                           net644553, ZN => n5800);
   U3308 : AOI22_X1 port map( A1 => n5248, A2 => n462, B1 => n6364, B2 => n4081
                           , ZN => n5808);
   U3307 : AOI22_X1 port map( A1 => n3911, A2 => net644618, B1 => n3912, B2 => 
                           net644489, ZN => n5809);
   U3305 : AOI22_X1 port map( A1 => n5244, A2 => n3973, B1 => n6366, B2 => n378
                           , ZN => n5810);
   U3304 : AOI22_X1 port map( A1 => n3913, A2 => net644586, B1 => n3914, B2 => 
                           net644682, ZN => n5811);
   U3303 : NAND4_X1 port map( A1 => n5808, A2 => n5809, A3 => n5810, A4 => 
                           n5811, ZN => n5802);
   U3301 : AOI22_X1 port map( A1 => n5236, A2 => n464, B1 => n6368, B2 => n4082
                           , ZN => n5804);
   U3300 : AOI22_X1 port map( A1 => n3910, A2 => net644778, B1 => n3909, B2 => 
                           net644746, ZN => n5805);
   U3299 : AOI22_X1 port map( A1 => n3908, A2 => net644908, B1 => n3907, B2 => 
                           net644425, ZN => n5806);
   U3297 : AOI22_X1 port map( A1 => n3906, A2 => n3974, B1 => n3905, B2 => n463
                           , ZN => n5807);
   U3296 : NAND4_X1 port map( A1 => n5804, A2 => n5805, A3 => n5806, A4 => 
                           n5807, ZN => n5803);
   U3295 : OAI21_X1 port map( B1 => n5802, B2 => n5803, A => n6370, ZN => n5801
                           );
   U3294 : OAI211_X1 port map( C1 => n571, C2 => n5220, A => n5800, B => n5801,
                           ZN => n5797);
   U3292 : AOI22_X1 port map( A1 => n6373, A2 => net644809, B1 => n6372, B2 => 
                           n4083, ZN => n5799);
   U3291 : OAI21_X1 port map( B1 => n633, B2 => n5216, A => n5799, ZN => n5798)
                           ;
   U3290 : AOI211_X1 port map( C1 => n6374, C2 => net644714, A => n5797, B => 
                           n5798, ZN => n5796);
   U3289 : NAND4_X1 port map( A1 => n5793, A2 => n5794, A3 => n5795, A4 => 
                           n5796, ZN => n2702);
   U2836 : AOI22_X1 port map( A1 => n6356, A2 => n3940, B1 => n6355, B2 => 
                           n4026, ZN => n5441);
   U2835 : AOI22_X1 port map( A1 => n6358, A2 => net644891, B1 => n6357, B2 => 
                           net644857, ZN => n5442);
   U2834 : AOI22_X1 port map( A1 => n6360, A2 => net644473, B1 => n6359, B2 => 
                           DATAIN(22), ZN => n5462);
   U2833 : OAI21_X1 port map( B1 => n5257, B2 => net644378, A => n5462, ZN => 
                           n5460);
   U2832 : OAI22_X1 port map( A1 => n524, A2 => n5255, B1 => n649, B2 => n5256,
                           ZN => n5461);
   U2831 : AOI211_X1 port map( C1 => n6361, C2 => net644665, A => n5460, B => 
                           n5461, ZN => n5443);
   U2830 : AOI22_X1 port map( A1 => n6363, A2 => net644537, B1 => n6362, B2 => 
                           net644569, ZN => n5448);
   U2828 : AOI22_X1 port map( A1 => n6365, A2 => n414, B1 => n6364, B2 => n4134
                           , ZN => n5456);
   U2827 : AOI22_X1 port map( A1 => n3911, A2 => net644634, B1 => n3912, B2 => 
                           net644505, ZN => n5457);
   U2825 : AOI22_X1 port map( A1 => n6367, A2 => n4027, B1 => n6366, B2 => n362
                           , ZN => n5458);
   U2824 : AOI22_X1 port map( A1 => n3913, A2 => net644602, B1 => n3914, B2 => 
                           net644698, ZN => n5459);
   U2823 : NAND4_X1 port map( A1 => n5456, A2 => n5457, A3 => n5458, A4 => 
                           n5459, ZN => n5450);
   U2821 : AOI22_X1 port map( A1 => n6369, A2 => n416, B1 => n6368, B2 => n4135
                           , ZN => n5452);
   U2820 : AOI22_X1 port map( A1 => n3910, A2 => net644794, B1 => n3909, B2 => 
                           net644762, ZN => n5453);
   U2819 : AOI22_X1 port map( A1 => n3908, A2 => net644924, B1 => n3907, B2 => 
                           net644441, ZN => n5454);
   U2817 : AOI22_X1 port map( A1 => n3906, A2 => n4028, B1 => n3905, B2 => n415
                           , ZN => n5455);
   U2816 : NAND4_X1 port map( A1 => n5452, A2 => n5453, A3 => n5454, A4 => 
                           n5455, ZN => n5451);
   U2815 : OAI21_X1 port map( B1 => n5450, B2 => n5451, A => n6370, ZN => n5449
                           );
   U2814 : OAI211_X1 port map( C1 => n555, C2 => n5220, A => n5448, B => n5449,
                           ZN => n5445);
   U2812 : AOI22_X1 port map( A1 => n6373, A2 => net644825, B1 => n6372, B2 => 
                           n4136, ZN => n5447);
   U2811 : OAI21_X1 port map( B1 => n617, B2 => n5216, A => n5447, ZN => n5446)
                           ;
   U2810 : AOI211_X1 port map( C1 => n6374, C2 => net644730, A => n5445, B => 
                           n5446, ZN => n5444);
   U2809 : NAND4_X1 port map( A1 => n5441, A2 => n5442, A3 => n5443, A4 => 
                           n5444, ZN => n2718);
   U2686 : AOI22_X1 port map( A1 => n6356, A2 => n3945, B1 => n5264, B2 => 
                           n4044, ZN => n5331);
   U2685 : AOI22_X1 port map( A1 => n5261, A2 => net644896, B1 => n5262, B2 => 
                           net644862, ZN => n5332);
   U2684 : AOI22_X1 port map( A1 => n5259, A2 => net644478, B1 => n5260, B2 => 
                           DATAIN(27), ZN => n5352);
   U2683 : OAI21_X1 port map( B1 => n5257, B2 => net644383, A => n5352, ZN => 
                           n5350);
   U2682 : OAI22_X1 port map( A1 => n519, A2 => n5255, B1 => n644, B2 => n5256,
                           ZN => n5351);
   U2681 : AOI211_X1 port map( C1 => n6361, C2 => net644670, A => n5350, B => 
                           n5351, ZN => n5333);
   U2680 : AOI22_X1 port map( A1 => n5250, A2 => net644542, B1 => n5251, B2 => 
                           net644574, ZN => n5338);
   U2678 : AOI22_X1 port map( A1 => n5248, A2 => n399, B1 => n5249, B2 => n4152
                           , ZN => n5346);
   U2677 : AOI22_X1 port map( A1 => n3911, A2 => net644639, B1 => n3912, B2 => 
                           net644510, ZN => n5347);
   U2675 : AOI22_X1 port map( A1 => n6367, A2 => n4045, B1 => n5245, B2 => n357
                           , ZN => n5348);
   U2674 : AOI22_X1 port map( A1 => n3913, A2 => net644607, B1 => n3914, B2 => 
                           net644703, ZN => n5349);
   U2673 : NAND4_X1 port map( A1 => n5346, A2 => n5347, A3 => n5348, A4 => 
                           n5349, ZN => n5340);
   U2671 : AOI22_X1 port map( A1 => n6369, A2 => n401, B1 => n5237, B2 => n4153
                           , ZN => n5342);
   U2670 : AOI22_X1 port map( A1 => n3910, A2 => net644799, B1 => n3909, B2 => 
                           net644767, ZN => n5343);
   U2669 : AOI22_X1 port map( A1 => n3908, A2 => net644929, B1 => n3907, B2 => 
                           net644446, ZN => n5344);
   U2667 : AOI22_X1 port map( A1 => n3906, A2 => n4046, B1 => n3905, B2 => n400
                           , ZN => n5345);
   U2666 : NAND4_X1 port map( A1 => n5342, A2 => n5343, A3 => n5344, A4 => 
                           n5345, ZN => n5341);
   U2665 : OAI21_X1 port map( B1 => n5340, B2 => n5341, A => n6370, ZN => n5339
                           );
   U2664 : OAI211_X1 port map( C1 => n550, C2 => n5220, A => n5338, B => n5339,
                           ZN => n5335);
   U2662 : AOI22_X1 port map( A1 => n6373, A2 => net644830, B1 => n6372, B2 => 
                           n4154, ZN => n5337);
   U2661 : OAI21_X1 port map( B1 => n612, B2 => n5216, A => n5337, ZN => n5336)
                           ;
   U2660 : AOI211_X1 port map( C1 => n5213, C2 => net644735, A => n5335, B => 
                           n5336, ZN => n5334);
   U2659 : NAND4_X1 port map( A1 => n5331, A2 => n5332, A3 => n5333, A4 => 
                           n5334, ZN => n2723);
   U2806 : AOI22_X1 port map( A1 => n6356, A2 => n3941, B1 => n6355, B2 => 
                           n4029, ZN => n5419);
   U2805 : AOI22_X1 port map( A1 => n6358, A2 => net644892, B1 => n6357, B2 => 
                           net644858, ZN => n5420);
   U2804 : AOI22_X1 port map( A1 => n5259, A2 => net644474, B1 => n6359, B2 => 
                           DATAIN(23), ZN => n5440);
   U2803 : OAI21_X1 port map( B1 => n5257, B2 => net644379, A => n5440, ZN => 
                           n5438);
   U2802 : OAI22_X1 port map( A1 => n523, A2 => n5255, B1 => n648, B2 => n5256,
                           ZN => n5439);
   U2801 : AOI211_X1 port map( C1 => n6361, C2 => net644666, A => n5438, B => 
                           n5439, ZN => n5421);
   U2800 : AOI22_X1 port map( A1 => n5250, A2 => net644538, B1 => n5251, B2 => 
                           net644570, ZN => n5426);
   U2798 : AOI22_X1 port map( A1 => n6365, A2 => n411, B1 => n6364, B2 => n4137
                           , ZN => n5434);
   U2797 : AOI22_X1 port map( A1 => n3911, A2 => net644635, B1 => n3912, B2 => 
                           net644506, ZN => n5435);
   U2795 : AOI22_X1 port map( A1 => n6367, A2 => n4030, B1 => n6366, B2 => n361
                           , ZN => n5436);
   U2794 : AOI22_X1 port map( A1 => n3913, A2 => net644603, B1 => n3914, B2 => 
                           net644699, ZN => n5437);
   U2793 : NAND4_X1 port map( A1 => n5434, A2 => n5435, A3 => n5436, A4 => 
                           n5437, ZN => n5428);
   U2791 : AOI22_X1 port map( A1 => n6369, A2 => n413, B1 => n6368, B2 => n4138
                           , ZN => n5430);
   U2790 : AOI22_X1 port map( A1 => n3910, A2 => net644795, B1 => n3909, B2 => 
                           net644763, ZN => n5431);
   U2789 : AOI22_X1 port map( A1 => n3908, A2 => net644925, B1 => n3907, B2 => 
                           net644442, ZN => n5432);
   U2787 : AOI22_X1 port map( A1 => n3906, A2 => n4031, B1 => n3905, B2 => n412
                           , ZN => n5433);
   U2786 : NAND4_X1 port map( A1 => n5430, A2 => n5431, A3 => n5432, A4 => 
                           n5433, ZN => n5429);
   U2785 : OAI21_X1 port map( B1 => n5428, B2 => n5429, A => n6370, ZN => n5427
                           );
   U2784 : OAI211_X1 port map( C1 => n554, C2 => n5220, A => n5426, B => n5427,
                           ZN => n5423);
   U2782 : AOI22_X1 port map( A1 => n6373, A2 => net644826, B1 => n6372, B2 => 
                           n4139, ZN => n5425);
   U2781 : OAI21_X1 port map( B1 => n616, B2 => n5216, A => n5425, ZN => n5424)
                           ;
   U2780 : AOI211_X1 port map( C1 => n6374, C2 => net644731, A => n5423, B => 
                           n5424, ZN => n5422);
   U2779 : NAND4_X1 port map( A1 => n5419, A2 => n5420, A3 => n5421, A4 => 
                           n5422, ZN => n2719);
   U1691 : AOI22_X1 port map( A1 => n4241, A2 => n4053, B1 => n6375, B2 => 
                           n3948, ZN => n4246);
   U1690 : AOI22_X1 port map( A1 => net644899, A2 => n4239, B1 => net644865, B2
                           => n4240, ZN => n4247);
   U1689 : AOI22_X1 port map( A1 => net644481, A2 => n6380, B1 => DATAIN(30), 
                           B2 => n6379, ZN => n4272);
   U1688 : OAI21_X1 port map( B1 => n4235, B2 => net644417, A => n4272, ZN => 
                           n4270);
   U1687 : OAI22_X1 port map( A1 => n641, A2 => n4233, B1 => n516, B2 => n4234,
                           ZN => n4271);
   U1686 : AOI211_X1 port map( C1 => net644673, C2 => n6381, A => n4270, B => 
                           n4271, ZN => n4248);
   U1685 : AOI22_X1 port map( A1 => net644577, A2 => n6382, B1 => net644545, B2
                           => n3880, ZN => n4254);
   U1684 : AOI22_X1 port map( A1 => n390, A2 => n6383, B1 => n3896, B2 => n4161
                           , ZN => n4264);
   U1683 : AOI22_X1 port map( A1 => net644642, A2 => n3895, B1 => net644513, B2
                           => n3894, ZN => n4265);
   U1682 : AOI22_X1 port map( A1 => n4220, A2 => n354, B1 => n3891, B2 => n4054
                           , ZN => n4266);
   U1681 : AOI22_X1 port map( A1 => net644610, A2 => n3890, B1 => net644706, B2
                           => n3897, ZN => n4267);
   U1680 : NAND4_X1 port map( A1 => n4264, A2 => n4265, A3 => n4266, A4 => 
                           n4267, ZN => n4256);
   U1679 : AOI22_X1 port map( A1 => n392, A2 => n3904, B1 => n3903, B2 => n4162
                           , ZN => n4258);
   U1678 : AOI22_X1 port map( A1 => net644802, A2 => n3902, B1 => net644770, B2
                           => n3901, ZN => n4259);
   U1677 : AOI22_X1 port map( A1 => net644932, A2 => n3900, B1 => net644449, B2
                           => n3899, ZN => n4260);
   U1676 : AOI22_X1 port map( A1 => n4204, A2 => n391, B1 => n3898, B2 => n4055
                           , ZN => n4261);
   U1675 : NAND4_X1 port map( A1 => n4258, A2 => n4259, A3 => n4260, A4 => 
                           n4261, ZN => n4257);
   U1674 : OAI21_X1 port map( B1 => n4256, B2 => n4257, A => n6386, ZN => n4255
                           );
   U1673 : OAI211_X1 port map( C1 => n547, C2 => n4194, A => n4254, B => n4255,
                           ZN => n4250);
   U1672 : AOI22_X1 port map( A1 => net644833, A2 => n6389, B1 => n6388, B2 => 
                           n4163, ZN => n4252);
   U1671 : OAI21_X1 port map( B1 => n609, B2 => n4189, A => n4252, ZN => n4251)
                           ;
   U1670 : AOI211_X1 port map( C1 => net644738, C2 => n6390, A => n4250, B => 
                           n4251, ZN => n4249);
   U1669 : NAND4_X1 port map( A1 => n4246, A2 => n4247, A3 => n4248, A4 => 
                           n4249, ZN => n2788);
   U1743 : AOI22_X1 port map( A1 => n4241, A2 => n4047, B1 => n4243, B2 => 
                           n3946, ZN => n4306);
   U1742 : AOI22_X1 port map( A1 => net644897, A2 => n6378, B1 => net644863, B2
                           => n4240, ZN => n4307);
   U1741 : AOI22_X1 port map( A1 => net644479, A2 => n6380, B1 => DATAIN(28), 
                           B2 => n6379, ZN => n4332);
   U1740 : OAI21_X1 port map( B1 => n4235, B2 => net644415, A => n4332, ZN => 
                           n4330);
   U1739 : OAI22_X1 port map( A1 => n643, A2 => n4233, B1 => n518, B2 => n4234,
                           ZN => n4331);
   U1738 : AOI211_X1 port map( C1 => net644671, C2 => n6381, A => n4330, B => 
                           n4331, ZN => n4308);
   U1737 : AOI22_X1 port map( A1 => net644575, A2 => n6382, B1 => net644543, B2
                           => n3880, ZN => n4314);
   U1736 : AOI22_X1 port map( A1 => n396, A2 => n6383, B1 => n3896, B2 => n4155
                           , ZN => n4324);
   U1735 : AOI22_X1 port map( A1 => net644640, A2 => n3895, B1 => net644511, B2
                           => n3894, ZN => n4325);
   U1734 : AOI22_X1 port map( A1 => n4220, A2 => n356, B1 => n4221, B2 => n4048
                           , ZN => n4326);
   U1733 : AOI22_X1 port map( A1 => net644608, A2 => n3890, B1 => net644704, B2
                           => n3897, ZN => n4327);
   U1732 : NAND4_X1 port map( A1 => n4324, A2 => n4325, A3 => n4326, A4 => 
                           n4327, ZN => n4316);
   U1731 : AOI22_X1 port map( A1 => n398, A2 => n3904, B1 => n4212, B2 => n4156
                           , ZN => n4318);
   U1730 : AOI22_X1 port map( A1 => net644800, A2 => n3902, B1 => net644768, B2
                           => n3901, ZN => n4319);
   U1729 : AOI22_X1 port map( A1 => net644930, A2 => n3900, B1 => net644447, B2
                           => n3899, ZN => n4320);
   U1728 : AOI22_X1 port map( A1 => n4204, A2 => n397, B1 => n3898, B2 => n4049
                           , ZN => n4321);
   U1727 : NAND4_X1 port map( A1 => n4318, A2 => n4319, A3 => n4320, A4 => 
                           n4321, ZN => n4317);
   U1726 : OAI21_X1 port map( B1 => n4316, B2 => n4317, A => n6386, ZN => n4315
                           );
   U1725 : OAI211_X1 port map( C1 => n549, C2 => n4194, A => n4314, B => n4315,
                           ZN => n4310);
   U1724 : AOI22_X1 port map( A1 => net644831, A2 => n6389, B1 => n4192, B2 => 
                           n4157, ZN => n4312);
   U1723 : OAI21_X1 port map( B1 => n611, B2 => n4189, A => n4312, ZN => n4311)
                           ;
   U1722 : AOI211_X1 port map( C1 => net644736, C2 => n6390, A => n4310, B => 
                           n4311, ZN => n4309);
   U1721 : NAND4_X1 port map( A1 => n4306, A2 => n4307, A3 => n4308, A4 => 
                           n4309, ZN => n2784);
   U1665 : AOI22_X1 port map( A1 => n4241, A2 => n4056, B1 => n4243, B2 => 
                           n3949, ZN => n4182);
   U1664 : AOI22_X1 port map( A1 => net644900, A2 => n4239, B1 => net644866, B2
                           => n4240, ZN => n4183);
   U1663 : AOI22_X1 port map( A1 => net644482, A2 => n6380, B1 => DATAIN(31), 
                           B2 => n6379, ZN => n4236);
   U1662 : OAI21_X1 port map( B1 => n4235, B2 => net644418, A => n4236, ZN => 
                           n4231);
   U1661 : OAI22_X1 port map( A1 => n640, A2 => n4233, B1 => n515, B2 => n4234,
                           ZN => n4232);
   U1660 : AOI211_X1 port map( C1 => net644674, C2 => n6381, A => n4231, B => 
                           n4232, ZN => n4184);
   U1659 : AOI22_X1 port map( A1 => net644578, A2 => n4228, B1 => net644546, B2
                           => n3880, ZN => n4195);
   U1658 : AOI22_X1 port map( A1 => n387, A2 => n6383, B1 => n3896, B2 => n4164
                           , ZN => n4214);
   U1657 : AOI22_X1 port map( A1 => net644643, A2 => n3895, B1 => net644514, B2
                           => n3894, ZN => n4215);
   U1656 : AOI22_X1 port map( A1 => n4220, A2 => n353, B1 => n3891, B2 => n4057
                           , ZN => n4216);
   U1655 : AOI22_X1 port map( A1 => net644611, A2 => n3890, B1 => net644707, B2
                           => n3897, ZN => n4217);
   U1654 : NAND4_X1 port map( A1 => n4214, A2 => n4215, A3 => n4216, A4 => 
                           n4217, ZN => n4197);
   U1653 : AOI22_X1 port map( A1 => n389, A2 => n3904, B1 => n3903, B2 => n4165
                           , ZN => n4200);
   U1652 : AOI22_X1 port map( A1 => net644803, A2 => n3902, B1 => net644771, B2
                           => n3901, ZN => n4201);
   U1651 : AOI22_X1 port map( A1 => net644933, A2 => n3900, B1 => net644450, B2
                           => n3899, ZN => n4202);
   U1650 : AOI22_X1 port map( A1 => n6385, A2 => n388, B1 => n3898, B2 => n4058
                           , ZN => n4203);
   U1649 : NAND4_X1 port map( A1 => n4200, A2 => n4201, A3 => n4202, A4 => 
                           n4203, ZN => n4198);
   U1648 : OAI21_X1 port map( B1 => n4197, B2 => n4198, A => n6386, ZN => n4196
                           );
   U1647 : OAI211_X1 port map( C1 => n546, C2 => n4194, A => n4195, B => n4196,
                           ZN => n4187);
   U1646 : AOI22_X1 port map( A1 => net644834, A2 => n6389, B1 => n4192, B2 => 
                           n4166, ZN => n4190);
   U1645 : OAI21_X1 port map( B1 => n608, B2 => n4189, A => n4190, ZN => n4188)
                           ;
   U1644 : AOI211_X1 port map( C1 => net644739, C2 => n6390, A => n4187, B => 
                           n4188, ZN => n4185);
   U1643 : NAND4_X1 port map( A1 => n4182, A2 => n4183, A3 => n4184, A4 => 
                           n4185, ZN => n2790);
   U1717 : AOI22_X1 port map( A1 => n4241, A2 => n4050, B1 => n6375, B2 => 
                           n3947, ZN => n4276);
   U1716 : AOI22_X1 port map( A1 => net644898, A2 => n6378, B1 => net644864, B2
                           => n4240, ZN => n4277);
   U1715 : AOI22_X1 port map( A1 => net644480, A2 => n6380, B1 => DATAIN(29), 
                           B2 => n6379, ZN => n4302);
   U1714 : OAI21_X1 port map( B1 => n4235, B2 => net644416, A => n4302, ZN => 
                           n4300);
   U1713 : OAI22_X1 port map( A1 => n642, A2 => n4233, B1 => n517, B2 => n4234,
                           ZN => n4301);
   U1712 : AOI211_X1 port map( C1 => net644672, C2 => n6381, A => n4300, B => 
                           n4301, ZN => n4278);
   U1711 : AOI22_X1 port map( A1 => net644576, A2 => n6382, B1 => net644544, B2
                           => n3880, ZN => n4284);
   U1710 : AOI22_X1 port map( A1 => n393, A2 => n6383, B1 => n3896, B2 => n4158
                           , ZN => n4294);
   U1709 : AOI22_X1 port map( A1 => net644641, A2 => n3895, B1 => net644512, B2
                           => n3894, ZN => n4295);
   U1708 : AOI22_X1 port map( A1 => n4220, A2 => n355, B1 => n4221, B2 => n4051
                           , ZN => n4296);
   U1707 : AOI22_X1 port map( A1 => net644609, A2 => n3890, B1 => net644705, B2
                           => n3897, ZN => n4297);
   U1706 : NAND4_X1 port map( A1 => n4294, A2 => n4295, A3 => n4296, A4 => 
                           n4297, ZN => n4286);
   U1705 : AOI22_X1 port map( A1 => n395, A2 => n3904, B1 => n4212, B2 => n4159
                           , ZN => n4288);
   U1704 : AOI22_X1 port map( A1 => net644801, A2 => n3902, B1 => net644769, B2
                           => n3901, ZN => n4289);
   U1703 : AOI22_X1 port map( A1 => net644931, A2 => n3900, B1 => net644448, B2
                           => n3899, ZN => n4290);
   U1702 : AOI22_X1 port map( A1 => n6385, A2 => n394, B1 => n3898, B2 => n4052
                           , ZN => n4291);
   U1701 : NAND4_X1 port map( A1 => n4288, A2 => n4289, A3 => n4290, A4 => 
                           n4291, ZN => n4287);
   U1700 : OAI21_X1 port map( B1 => n4286, B2 => n4287, A => n6386, ZN => n4285
                           );
   U1699 : OAI211_X1 port map( C1 => n548, C2 => n4194, A => n4284, B => n4285,
                           ZN => n4280);
   U1698 : AOI22_X1 port map( A1 => net644832, A2 => n6389, B1 => n6388, B2 => 
                           n4160, ZN => n4282);
   U1697 : OAI21_X1 port map( B1 => n610, B2 => n4189, A => n4282, ZN => n4281)
                           ;
   U1696 : AOI211_X1 port map( C1 => net644737, C2 => n6390, A => n4280, B => 
                           n4281, ZN => n4279);
   U1695 : NAND4_X1 port map( A1 => n4276, A2 => n4277, A3 => n4278, A4 => 
                           n4279, ZN => n2786);
   U1821 : AOI22_X1 port map( A1 => n4241, A2 => n4038, B1 => n6375, B2 => 
                           n3943, ZN => n4396);
   U1820 : AOI22_X1 port map( A1 => net644894, A2 => n4239, B1 => net644860, B2
                           => n4240, ZN => n4397);
   U1819 : AOI22_X1 port map( A1 => net644476, A2 => n6380, B1 => DATAIN(25), 
                           B2 => n6379, ZN => n4422);
   U1818 : OAI21_X1 port map( B1 => n4235, B2 => net644412, A => n4422, ZN => 
                           n4420);
   U1817 : OAI22_X1 port map( A1 => n646, A2 => n4233, B1 => n521, B2 => n4234,
                           ZN => n4421);
   U1816 : AOI211_X1 port map( C1 => net644668, C2 => n6381, A => n4420, B => 
                           n4421, ZN => n4398);
   U1815 : AOI22_X1 port map( A1 => net644572, A2 => n6382, B1 => net644540, B2
                           => n3880, ZN => n4404);
   U1814 : AOI22_X1 port map( A1 => n405, A2 => n6383, B1 => n3896, B2 => n4144
                           , ZN => n4414);
   U1813 : AOI22_X1 port map( A1 => net644637, A2 => n3895, B1 => net644508, B2
                           => n3894, ZN => n4415);
   U1812 : AOI22_X1 port map( A1 => n4220, A2 => n359, B1 => n4221, B2 => n4039
                           , ZN => n4416);
   U1811 : AOI22_X1 port map( A1 => net644605, A2 => n3890, B1 => net644701, B2
                           => n3897, ZN => n4417);
   U1810 : NAND4_X1 port map( A1 => n4414, A2 => n4415, A3 => n4416, A4 => 
                           n4417, ZN => n4406);
   U1809 : AOI22_X1 port map( A1 => n407, A2 => n3904, B1 => n4212, B2 => n4147
                           , ZN => n4408);
   U1808 : AOI22_X1 port map( A1 => net644797, A2 => n3902, B1 => net644765, B2
                           => n3901, ZN => n4409);
   U1807 : AOI22_X1 port map( A1 => net644927, A2 => n3900, B1 => net644444, B2
                           => n3899, ZN => n4410);
   U1806 : AOI22_X1 port map( A1 => n6385, A2 => n406, B1 => n3898, B2 => n4040
                           , ZN => n4411);
   U1805 : NAND4_X1 port map( A1 => n4408, A2 => n4409, A3 => n4410, A4 => 
                           n4411, ZN => n4407);
   U1804 : OAI21_X1 port map( B1 => n4406, B2 => n4407, A => n6386, ZN => n4405
                           );
   U1803 : OAI211_X1 port map( C1 => n552, C2 => n4194, A => n4404, B => n4405,
                           ZN => n4400);
   U1802 : AOI22_X1 port map( A1 => net644828, A2 => n6389, B1 => n4192, B2 => 
                           n4148, ZN => n4402);
   U1801 : OAI21_X1 port map( B1 => n614, B2 => n4189, A => n4402, ZN => n4401)
                           ;
   U1800 : AOI211_X1 port map( C1 => net644733, C2 => n6390, A => n4400, B => 
                           n4401, ZN => n4399);
   U1799 : NAND4_X1 port map( A1 => n4396, A2 => n4397, A3 => n4398, A4 => 
                           n4399, ZN => n2778);
   U2341 : AOI22_X1 port map( A1 => n6376, A2 => n3969, B1 => n6375, B2 => 
                           n3920, ZN => n4996);
   U2340 : AOI22_X1 port map( A1 => net644874, A2 => n6378, B1 => net644840, B2
                           => n6377, ZN => n4997);
   U2339 : AOI22_X1 port map( A1 => net644456, A2 => n6380, B1 => DATAIN(5), B2
                           => n6379, ZN => n5022);
   U2338 : OAI21_X1 port map( B1 => n4235, B2 => net644392, A => n5022, ZN => 
                           n5020);
   U2337 : OAI22_X1 port map( A1 => n666, A2 => n4233, B1 => n541, B2 => n4234,
                           ZN => n5021);
   U2336 : AOI211_X1 port map( C1 => net644648, C2 => n6381, A => n5020, B => 
                           n5021, ZN => n4998);
   U2335 : AOI22_X1 port map( A1 => net644552, A2 => n6382, B1 => net644520, B2
                           => n3880, ZN => n5004);
   U2334 : AOI22_X1 port map( A1 => n465, A2 => n4225, B1 => n3896, B2 => n4078
                           , ZN => n5014);
   U2333 : AOI22_X1 port map( A1 => net644617, A2 => n3895, B1 => net644488, B2
                           => n3894, ZN => n5015);
   U2332 : AOI22_X1 port map( A1 => n6384, A2 => n379, B1 => n3891, B2 => n3970
                           , ZN => n5016);
   U2331 : AOI22_X1 port map( A1 => net644585, A2 => n3890, B1 => net644681, B2
                           => n3897, ZN => n5017);
   U2330 : NAND4_X1 port map( A1 => n5014, A2 => n5015, A3 => n5016, A4 => 
                           n5017, ZN => n5006);
   U2329 : AOI22_X1 port map( A1 => n467, A2 => n3904, B1 => n3903, B2 => n4079
                           , ZN => n5008);
   U2328 : AOI22_X1 port map( A1 => net644777, A2 => n3902, B1 => net644745, B2
                           => n3901, ZN => n5009);
   U2327 : AOI22_X1 port map( A1 => net644907, A2 => n3900, B1 => net644424, B2
                           => n3899, ZN => n5010);
   U2326 : AOI22_X1 port map( A1 => n6385, A2 => n466, B1 => n3898, B2 => n3971
                           , ZN => n5011);
   U2325 : NAND4_X1 port map( A1 => n5008, A2 => n5009, A3 => n5010, A4 => 
                           n5011, ZN => n5007);
   U2324 : OAI21_X1 port map( B1 => n5006, B2 => n5007, A => n6386, ZN => n5005
                           );
   U2323 : OAI211_X1 port map( C1 => n572, C2 => n4194, A => n5004, B => n5005,
                           ZN => n5000);
   U2322 : AOI22_X1 port map( A1 => net644808, A2 => n6389, B1 => n6388, B2 => 
                           n4080, ZN => n5002);
   U2321 : OAI21_X1 port map( B1 => n634, B2 => n4189, A => n5002, ZN => n5001)
                           ;
   U2320 : AOI211_X1 port map( C1 => net644713, C2 => n6390, A => n5000, B => 
                           n5001, ZN => n4999);
   U2319 : NAND4_X1 port map( A1 => n4996, A2 => n4997, A3 => n4998, A4 => 
                           n4999, ZN => n2738);
   U2185 : AOI22_X1 port map( A1 => n6376, A2 => n3987, B1 => n6375, B2 => 
                           n3929, ZN => n4816);
   U2184 : AOI22_X1 port map( A1 => net644880, A2 => n6378, B1 => net644846, B2
                           => n6377, ZN => n4817);
   U2183 : AOI22_X1 port map( A1 => net644462, A2 => n4237, B1 => DATAIN(11), 
                           B2 => n4238, ZN => n4842);
   U2182 : OAI21_X1 port map( B1 => n4235, B2 => net644398, A => n4842, ZN => 
                           n4840);
   U2181 : OAI22_X1 port map( A1 => n660, A2 => n4233, B1 => n535, B2 => n4234,
                           ZN => n4841);
   U2180 : AOI211_X1 port map( C1 => net644654, C2 => n6381, A => n4840, B => 
                           n4841, ZN => n4818);
   U2179 : AOI22_X1 port map( A1 => net644558, A2 => n6382, B1 => net644526, B2
                           => n3880, ZN => n4824);
   U2178 : AOI22_X1 port map( A1 => n447, A2 => n6383, B1 => n3896, B2 => n4096
                           , ZN => n4834);
   U2177 : AOI22_X1 port map( A1 => net644623, A2 => n3895, B1 => net644494, B2
                           => n3894, ZN => n4835);
   U2176 : AOI22_X1 port map( A1 => n6384, A2 => n373, B1 => n3891, B2 => n3988
                           , ZN => n4836);
   U2175 : AOI22_X1 port map( A1 => net644591, A2 => n3890, B1 => net644687, B2
                           => n4219, ZN => n4837);
   U2174 : NAND4_X1 port map( A1 => n4834, A2 => n4835, A3 => n4836, A4 => 
                           n4837, ZN => n4826);
   U2173 : AOI22_X1 port map( A1 => n449, A2 => n3904, B1 => n3903, B2 => n4097
                           , ZN => n4828);
   U2172 : AOI22_X1 port map( A1 => net644783, A2 => n3902, B1 => net644751, B2
                           => n3901, ZN => n4829);
   U2171 : AOI22_X1 port map( A1 => net644913, A2 => n3900, B1 => net644430, B2
                           => n3899, ZN => n4830);
   U2170 : AOI22_X1 port map( A1 => n6385, A2 => n448, B1 => n3898, B2 => n3989
                           , ZN => n4831);
   U2169 : NAND4_X1 port map( A1 => n4828, A2 => n4829, A3 => n4830, A4 => 
                           n4831, ZN => n4827);
   U2168 : OAI21_X1 port map( B1 => n4826, B2 => n4827, A => n6386, ZN => n4825
                           );
   U2167 : OAI211_X1 port map( C1 => n566, C2 => n4194, A => n4824, B => n4825,
                           ZN => n4820);
   U2166 : AOI22_X1 port map( A1 => net644814, A2 => n6389, B1 => n6388, B2 => 
                           n4098, ZN => n4822);
   U2165 : OAI21_X1 port map( B1 => n628, B2 => n4189, A => n4822, ZN => n4821)
                           ;
   U2164 : AOI211_X1 port map( C1 => net644719, C2 => n4186, A => n4820, B => 
                           n4821, ZN => n4819);
   U2163 : NAND4_X1 port map( A1 => n4816, A2 => n4817, A3 => n4818, A4 => 
                           n4819, ZN => n2750);
   U2159 : AOI22_X1 port map( A1 => n6376, A2 => n3990, B1 => n6375, B2 => 
                           n3930, ZN => n4786);
   U2158 : AOI22_X1 port map( A1 => net644881, A2 => n6378, B1 => net644847, B2
                           => n6377, ZN => n4787);
   U2157 : AOI22_X1 port map( A1 => net644463, A2 => n6380, B1 => DATAIN(12), 
                           B2 => n6379, ZN => n4812);
   U2156 : OAI21_X1 port map( B1 => n4235, B2 => net644399, A => n4812, ZN => 
                           n4810);
   U2155 : OAI22_X1 port map( A1 => n659, A2 => n4233, B1 => n534, B2 => n4234,
                           ZN => n4811);
   U2154 : AOI211_X1 port map( C1 => net644655, C2 => n6381, A => n4810, B => 
                           n4811, ZN => n4788);
   U2153 : AOI22_X1 port map( A1 => net644559, A2 => n6382, B1 => net644527, B2
                           => n4229, ZN => n4794);
   U2152 : AOI22_X1 port map( A1 => n444, A2 => n4225, B1 => n3896, B2 => n4099
                           , ZN => n4804);
   U2151 : AOI22_X1 port map( A1 => net644624, A2 => n3895, B1 => net644495, B2
                           => n4224, ZN => n4805);
   U2150 : AOI22_X1 port map( A1 => n6384, A2 => n372, B1 => n3891, B2 => n3991
                           , ZN => n4806);
   U2149 : AOI22_X1 port map( A1 => net644592, A2 => n4218, B1 => net644688, B2
                           => n3897, ZN => n4807);
   U2148 : NAND4_X1 port map( A1 => n4804, A2 => n4805, A3 => n4806, A4 => 
                           n4807, ZN => n4796);
   U2147 : AOI22_X1 port map( A1 => n446, A2 => n3904, B1 => n3903, B2 => n4100
                           , ZN => n4798);
   U2146 : AOI22_X1 port map( A1 => net644784, A2 => n3902, B1 => net644752, B2
                           => n4210, ZN => n4799);
   U2145 : AOI22_X1 port map( A1 => net644914, A2 => n3900, B1 => net644431, B2
                           => n4208, ZN => n4800);
   U2144 : AOI22_X1 port map( A1 => n6385, A2 => n445, B1 => n3898, B2 => n3992
                           , ZN => n4801);
   U2143 : NAND4_X1 port map( A1 => n4798, A2 => n4799, A3 => n4800, A4 => 
                           n4801, ZN => n4797);
   U2142 : OAI21_X1 port map( B1 => n4796, B2 => n4797, A => n4199, ZN => n4795
                           );
   U2141 : OAI211_X1 port map( C1 => n565, C2 => n4194, A => n4794, B => n4795,
                           ZN => n4790);
   U2140 : AOI22_X1 port map( A1 => net644815, A2 => n6389, B1 => n6388, B2 => 
                           n4101, ZN => n4792);
   U2139 : OAI21_X1 port map( B1 => n627, B2 => n4189, A => n4792, ZN => n4791)
                           ;
   U2138 : AOI211_X1 port map( C1 => net644720, C2 => n6390, A => n4790, B => 
                           n4791, ZN => n4789);
   U2137 : NAND4_X1 port map( A1 => n4786, A2 => n4787, A3 => n4788, A4 => 
                           n4789, ZN => n2752);
   U2447 : AOI22_X1 port map( A1 => n4241, A2 => n3954, B1 => n6375, B2 => 
                           n3916, ZN => n5116);
   U2446 : AOI22_X1 port map( A1 => net644870, A2 => n6378, B1 => net644836, B2
                           => n6377, ZN => n5117);
   U2445 : AOI22_X1 port map( A1 => net644452, A2 => n4237, B1 => DATAIN(1), B2
                           => n6379, ZN => n5143);
   U2444 : OAI21_X1 port map( B1 => n4235, B2 => net644388, A => n5143, ZN => 
                           n5140);
   U2442 : OAI22_X1 port map( A1 => n670, A2 => n4233, B1 => n545, B2 => n4234,
                           ZN => n5141);
   U2441 : AOI211_X1 port map( C1 => net644644, C2 => n6381, A => n5140, B => 
                           n5141, ZN => n5118);
   U2440 : AOI22_X1 port map( A1 => net644548, A2 => n6382, B1 => net644516, B2
                           => n3880, ZN => n5125);
   U2439 : AOI22_X1 port map( A1 => n477, A2 => n4225, B1 => n222, B2 => n3896,
                           ZN => n5135);
   U2438 : AOI22_X1 port map( A1 => net644613, A2 => n3895, B1 => net644484, B2
                           => n3894, ZN => n5136);
   U2437 : AOI22_X1 port map( A1 => n6384, A2 => n383, B1 => n3891, B2 => n3955
                           , ZN => n5137);
   U2436 : AOI22_X1 port map( A1 => net644581, A2 => n3890, B1 => net644677, B2
                           => n3897, ZN => n5138);
   U2435 : NAND4_X1 port map( A1 => n5135, A2 => n5136, A3 => n5137, A4 => 
                           n5138, ZN => n5127);
   U2434 : AOI22_X1 port map( A1 => n479, A2 => n3904, B1 => n3903, B2 => n4063
                           , ZN => n5129);
   U2433 : AOI22_X1 port map( A1 => net644773, A2 => n3902, B1 => net644741, B2
                           => n3901, ZN => n5130);
   U2432 : AOI22_X1 port map( A1 => net644903, A2 => n3900, B1 => net644420, B2
                           => n3899, ZN => n5131);
   U2431 : AOI22_X1 port map( A1 => n6385, A2 => n478, B1 => n3898, B2 => n3956
                           , ZN => n5132);
   U2430 : NAND4_X1 port map( A1 => n5129, A2 => n5130, A3 => n5131, A4 => 
                           n5132, ZN => n5128);
   U2429 : OAI21_X1 port map( B1 => n5127, B2 => n5128, A => n6386, ZN => n5126
                           );
   U2428 : OAI211_X1 port map( C1 => n576, C2 => n4194, A => n5125, B => n5126,
                           ZN => n5120);
   U2426 : AOI22_X1 port map( A1 => net644804, A2 => n6389, B1 => n6388, B2 => 
                           n4064, ZN => n5122);
   U2425 : OAI21_X1 port map( B1 => n638, B2 => n4189, A => n5122, ZN => n5121)
                           ;
   U2424 : AOI211_X1 port map( C1 => net644709, C2 => n4186, A => n5120, B => 
                           n5121, ZN => n5119);
   U2423 : NAND4_X1 port map( A1 => n5116, A2 => n5117, A3 => n5118, A4 => 
                           n5119, ZN => n2730);
   U2419 : AOI22_X1 port map( A1 => n4241, A2 => n3957, B1 => n6375, B2 => 
                           n3917, ZN => n5086);
   U2418 : AOI22_X1 port map( A1 => net644871, A2 => n6378, B1 => net644837, B2
                           => n6377, ZN => n5087);
   U2417 : AOI22_X1 port map( A1 => net644453, A2 => n4237, B1 => DATAIN(2), B2
                           => n6379, ZN => n5112);
   U2416 : OAI21_X1 port map( B1 => n4235, B2 => net644389, A => n5112, ZN => 
                           n5110);
   U2415 : OAI22_X1 port map( A1 => n669, A2 => n4233, B1 => n544, B2 => n4234,
                           ZN => n5111);
   U2414 : AOI211_X1 port map( C1 => net644645, C2 => n6381, A => n5110, B => 
                           n5111, ZN => n5088);
   U2413 : AOI22_X1 port map( A1 => net644549, A2 => n4228, B1 => net644517, B2
                           => n3880, ZN => n5094);
   U2412 : AOI22_X1 port map( A1 => n474, A2 => n4225, B1 => n3896, B2 => n4065
                           , ZN => n5104);
   U2411 : AOI22_X1 port map( A1 => net644614, A2 => n3895, B1 => net644485, B2
                           => n3894, ZN => n5105);
   U2410 : AOI22_X1 port map( A1 => n6384, A2 => n382, B1 => n3891, B2 => n3958
                           , ZN => n5106);
   U2409 : AOI22_X1 port map( A1 => net644582, A2 => n3890, B1 => net644678, B2
                           => n3897, ZN => n5107);
   U2408 : NAND4_X1 port map( A1 => n5104, A2 => n5105, A3 => n5106, A4 => 
                           n5107, ZN => n5096);
   U2407 : AOI22_X1 port map( A1 => n476, A2 => n3904, B1 => n3903, B2 => n4066
                           , ZN => n5098);
   U2406 : AOI22_X1 port map( A1 => net644774, A2 => n3902, B1 => net644742, B2
                           => n3901, ZN => n5099);
   U2405 : AOI22_X1 port map( A1 => net644904, A2 => n3900, B1 => net644421, B2
                           => n3899, ZN => n5100);
   U2404 : AOI22_X1 port map( A1 => n6385, A2 => n475, B1 => n3898, B2 => n3960
                           , ZN => n5101);
   U2403 : NAND4_X1 port map( A1 => n5098, A2 => n5099, A3 => n5100, A4 => 
                           n5101, ZN => n5097);
   U2402 : OAI21_X1 port map( B1 => n5096, B2 => n5097, A => n6386, ZN => n5095
                           );
   U2401 : OAI211_X1 port map( C1 => n575, C2 => n4194, A => n5094, B => n5095,
                           ZN => n5090);
   U2400 : AOI22_X1 port map( A1 => net644805, A2 => n6389, B1 => n6388, B2 => 
                           n4067, ZN => n5092);
   U2399 : OAI21_X1 port map( B1 => n637, B2 => n4189, A => n5092, ZN => n5091)
                           ;
   U2398 : AOI211_X1 port map( C1 => net644710, C2 => n4186, A => n5090, B => 
                           n5091, ZN => n5089);
   U2397 : NAND4_X1 port map( A1 => n5086, A2 => n5087, A3 => n5088, A4 => 
                           n5089, ZN => n2732);
   U2393 : AOI22_X1 port map( A1 => n6376, A2 => n3963, B1 => n6375, B2 => 
                           n3918, ZN => n5056);
   U2392 : AOI22_X1 port map( A1 => net644872, A2 => n6378, B1 => net644838, B2
                           => n6377, ZN => n5057);
   U2391 : AOI22_X1 port map( A1 => net644454, A2 => n4237, B1 => DATAIN(3), B2
                           => n4238, ZN => n5082);
   U2390 : OAI21_X1 port map( B1 => n4235, B2 => net644390, A => n5082, ZN => 
                           n5080);
   U2389 : OAI22_X1 port map( A1 => n668, A2 => n4233, B1 => n543, B2 => n4234,
                           ZN => n5081);
   U2388 : AOI211_X1 port map( C1 => net644646, C2 => n6381, A => n5080, B => 
                           n5081, ZN => n5058);
   U2387 : AOI22_X1 port map( A1 => net644550, A2 => n6382, B1 => net644518, B2
                           => n3880, ZN => n5064);
   U2386 : AOI22_X1 port map( A1 => n471, A2 => n6383, B1 => n3896, B2 => n4070
                           , ZN => n5074);
   U2385 : AOI22_X1 port map( A1 => net644615, A2 => n3895, B1 => net644486, B2
                           => n3894, ZN => n5075);
   U2384 : AOI22_X1 port map( A1 => n6384, A2 => n381, B1 => n3891, B2 => n3964
                           , ZN => n5076);
   U2383 : AOI22_X1 port map( A1 => net644583, A2 => n3890, B1 => net644679, B2
                           => n3897, ZN => n5077);
   U2382 : NAND4_X1 port map( A1 => n5074, A2 => n5075, A3 => n5076, A4 => 
                           n5077, ZN => n5066);
   U2381 : AOI22_X1 port map( A1 => n473, A2 => n3904, B1 => n3903, B2 => n4071
                           , ZN => n5068);
   U2380 : AOI22_X1 port map( A1 => net644775, A2 => n3902, B1 => net644743, B2
                           => n3901, ZN => n5069);
   U2379 : AOI22_X1 port map( A1 => net644905, A2 => n3900, B1 => net644422, B2
                           => n3899, ZN => n5070);
   U2378 : AOI22_X1 port map( A1 => n6385, A2 => n472, B1 => n3898, B2 => n3965
                           , ZN => n5071);
   U2377 : NAND4_X1 port map( A1 => n5068, A2 => n5069, A3 => n5070, A4 => 
                           n5071, ZN => n5067);
   U2376 : OAI21_X1 port map( B1 => n5066, B2 => n5067, A => n6386, ZN => n5065
                           );
   U2375 : OAI211_X1 port map( C1 => n574, C2 => n4194, A => n5064, B => n5065,
                           ZN => n5060);
   U2374 : AOI22_X1 port map( A1 => net644806, A2 => n6389, B1 => n6388, B2 => 
                           n4072, ZN => n5062);
   U2373 : OAI21_X1 port map( B1 => n636, B2 => n4189, A => n5062, ZN => n5061)
                           ;
   U2372 : AOI211_X1 port map( C1 => net644711, C2 => n6390, A => n5060, B => 
                           n5061, ZN => n5059);
   U2371 : NAND4_X1 port map( A1 => n5056, A2 => n5057, A3 => n5058, A4 => 
                           n5059, ZN => n2734);
   U2055 : AOI22_X1 port map( A1 => n6376, A2 => n4008, B1 => n6375, B2 => 
                           n3934, ZN => n4666);
   U2054 : AOI22_X1 port map( A1 => net644885, A2 => n6378, B1 => net644851, B2
                           => n6377, ZN => n4667);
   U2053 : AOI22_X1 port map( A1 => net644467, A2 => n4237, B1 => DATAIN(16), 
                           B2 => n6379, ZN => n4692);
   U2052 : OAI21_X1 port map( B1 => n4235, B2 => net644403, A => n4692, ZN => 
                           n4690);
   U2051 : OAI22_X1 port map( A1 => n655, A2 => n4233, B1 => n530, B2 => n4234,
                           ZN => n4691);
   U2050 : AOI211_X1 port map( C1 => net644659, C2 => n6381, A => n4690, B => 
                           n4691, ZN => n4668);
   U2049 : AOI22_X1 port map( A1 => net644563, A2 => n6382, B1 => net644531, B2
                           => n3880, ZN => n4674);
   U2048 : AOI22_X1 port map( A1 => n432, A2 => n6383, B1 => n3896, B2 => n4116
                           , ZN => n4684);
   U2047 : AOI22_X1 port map( A1 => net644628, A2 => n3895, B1 => net644499, B2
                           => n3894, ZN => n4685);
   U2046 : AOI22_X1 port map( A1 => n6384, A2 => n368, B1 => n3891, B2 => n4009
                           , ZN => n4686);
   U2045 : AOI22_X1 port map( A1 => net644596, A2 => n3890, B1 => net644692, B2
                           => n3897, ZN => n4687);
   U2044 : NAND4_X1 port map( A1 => n4684, A2 => n4685, A3 => n4686, A4 => 
                           n4687, ZN => n4676);
   U2043 : AOI22_X1 port map( A1 => n434, A2 => n3904, B1 => n3903, B2 => n4117
                           , ZN => n4678);
   U2042 : AOI22_X1 port map( A1 => net644788, A2 => n3902, B1 => net644756, B2
                           => n3901, ZN => n4679);
   U2041 : AOI22_X1 port map( A1 => net644918, A2 => n3900, B1 => net644435, B2
                           => n3899, ZN => n4680);
   U2040 : AOI22_X1 port map( A1 => n6385, A2 => n433, B1 => n3898, B2 => n4010
                           , ZN => n4681);
   U2039 : NAND4_X1 port map( A1 => n4678, A2 => n4679, A3 => n4680, A4 => 
                           n4681, ZN => n4677);
   U2038 : OAI21_X1 port map( B1 => n4676, B2 => n4677, A => n6386, ZN => n4675
                           );
   U2037 : OAI211_X1 port map( C1 => n561, C2 => n4194, A => n4674, B => n4675,
                           ZN => n4670);
   U2036 : AOI22_X1 port map( A1 => net644819, A2 => n6389, B1 => n4192, B2 => 
                           n4118, ZN => n4672);
   U2035 : OAI21_X1 port map( B1 => n623, B2 => n4189, A => n4672, ZN => n4671)
                           ;
   U2034 : AOI211_X1 port map( C1 => net644724, C2 => n4186, A => n4670, B => 
                           n4671, ZN => n4669);
   U2033 : NAND4_X1 port map( A1 => n4666, A2 => n4667, A3 => n4668, A4 => 
                           n4669, ZN => n2760);
   U2367 : AOI22_X1 port map( A1 => n4241, A2 => n3966, B1 => n6375, B2 => 
                           n3919, ZN => n5026);
   U2366 : AOI22_X1 port map( A1 => net644873, A2 => n6378, B1 => net644839, B2
                           => n6377, ZN => n5027);
   U2365 : AOI22_X1 port map( A1 => net644455, A2 => n4237, B1 => DATAIN(4), B2
                           => n6379, ZN => n5052);
   U2364 : OAI21_X1 port map( B1 => n4235, B2 => net644391, A => n5052, ZN => 
                           n5050);
   U2363 : OAI22_X1 port map( A1 => n667, A2 => n4233, B1 => n542, B2 => n4234,
                           ZN => n5051);
   U2362 : AOI211_X1 port map( C1 => net644647, C2 => n6381, A => n5050, B => 
                           n5051, ZN => n5028);
   U2361 : AOI22_X1 port map( A1 => net644551, A2 => n6382, B1 => net644519, B2
                           => n3880, ZN => n5034);
   U2360 : AOI22_X1 port map( A1 => n468, A2 => n4225, B1 => n3896, B2 => n4075
                           , ZN => n5044);
   U2359 : AOI22_X1 port map( A1 => net644616, A2 => n3895, B1 => net644487, B2
                           => n3894, ZN => n5045);
   U2358 : AOI22_X1 port map( A1 => n6384, A2 => n380, B1 => n3891, B2 => n3967
                           , ZN => n5046);
   U2357 : AOI22_X1 port map( A1 => net644584, A2 => n3890, B1 => net644680, B2
                           => n3897, ZN => n5047);
   U2356 : NAND4_X1 port map( A1 => n5044, A2 => n5045, A3 => n5046, A4 => 
                           n5047, ZN => n5036);
   U2355 : AOI22_X1 port map( A1 => n470, A2 => n3904, B1 => n3903, B2 => n4076
                           , ZN => n5038);
   U2354 : AOI22_X1 port map( A1 => net644776, A2 => n3902, B1 => net644744, B2
                           => n3901, ZN => n5039);
   U2353 : AOI22_X1 port map( A1 => net644906, A2 => n3900, B1 => net644423, B2
                           => n3899, ZN => n5040);
   U2352 : AOI22_X1 port map( A1 => n6385, A2 => n469, B1 => n3898, B2 => n3968
                           , ZN => n5041);
   U2351 : NAND4_X1 port map( A1 => n5038, A2 => n5039, A3 => n5040, A4 => 
                           n5041, ZN => n5037);
   U2350 : OAI21_X1 port map( B1 => n5036, B2 => n5037, A => n6386, ZN => n5035
                           );
   U2349 : OAI211_X1 port map( C1 => n573, C2 => n4194, A => n5034, B => n5035,
                           ZN => n5030);
   U2348 : AOI22_X1 port map( A1 => net644807, A2 => n6389, B1 => n6388, B2 => 
                           n4077, ZN => n5032);
   U2347 : OAI21_X1 port map( B1 => n635, B2 => n4189, A => n5032, ZN => n5031)
                           ;
   U2346 : AOI211_X1 port map( C1 => net644712, C2 => n4186, A => n5030, B => 
                           n5031, ZN => n5029);
   U2345 : NAND4_X1 port map( A1 => n5026, A2 => n5027, A3 => n5028, A4 => 
                           n5029, ZN => n2736);
   U2315 : AOI22_X1 port map( A1 => n6376, A2 => n3972, B1 => n6375, B2 => 
                           n3921, ZN => n4966);
   U2314 : AOI22_X1 port map( A1 => net644875, A2 => n6378, B1 => net644841, B2
                           => n6377, ZN => n4967);
   U2313 : AOI22_X1 port map( A1 => net644457, A2 => n6380, B1 => DATAIN(6), B2
                           => n6379, ZN => n4992);
   U2312 : OAI21_X1 port map( B1 => n4235, B2 => net644393, A => n4992, ZN => 
                           n4990);
   U2311 : OAI22_X1 port map( A1 => n665, A2 => n4233, B1 => n540, B2 => n4234,
                           ZN => n4991);
   U2310 : AOI211_X1 port map( C1 => net644649, C2 => n6381, A => n4990, B => 
                           n4991, ZN => n4968);
   U2309 : AOI22_X1 port map( A1 => net644553, A2 => n4228, B1 => net644521, B2
                           => n3880, ZN => n4974);
   U2308 : AOI22_X1 port map( A1 => n462, A2 => n4225, B1 => n3896, B2 => n4081
                           , ZN => n4984);
   U2307 : AOI22_X1 port map( A1 => net644618, A2 => n3895, B1 => net644489, B2
                           => n3894, ZN => n4985);
   U2306 : AOI22_X1 port map( A1 => n6384, A2 => n378, B1 => n3891, B2 => n3973
                           , ZN => n4986);
   U2305 : AOI22_X1 port map( A1 => net644586, A2 => n3890, B1 => net644682, B2
                           => n3897, ZN => n4987);
   U2304 : NAND4_X1 port map( A1 => n4984, A2 => n4985, A3 => n4986, A4 => 
                           n4987, ZN => n4976);
   U2303 : AOI22_X1 port map( A1 => n464, A2 => n3904, B1 => n3903, B2 => n4082
                           , ZN => n4978);
   U2302 : AOI22_X1 port map( A1 => net644778, A2 => n3902, B1 => net644746, B2
                           => n3901, ZN => n4979);
   U2301 : AOI22_X1 port map( A1 => net644908, A2 => n3900, B1 => net644425, B2
                           => n3899, ZN => n4980);
   U2300 : AOI22_X1 port map( A1 => n6385, A2 => n463, B1 => n3898, B2 => n3974
                           , ZN => n4981);
   U2299 : NAND4_X1 port map( A1 => n4978, A2 => n4979, A3 => n4980, A4 => 
                           n4981, ZN => n4977);
   U2298 : OAI21_X1 port map( B1 => n4976, B2 => n4977, A => n6386, ZN => n4975
                           );
   U2297 : OAI211_X1 port map( C1 => n571, C2 => n4194, A => n4974, B => n4975,
                           ZN => n4970);
   U2296 : AOI22_X1 port map( A1 => net644809, A2 => n6389, B1 => n6388, B2 => 
                           n4083, ZN => n4972);
   U2295 : OAI21_X1 port map( B1 => n633, B2 => n4189, A => n4972, ZN => n4971)
                           ;
   U2294 : AOI211_X1 port map( C1 => net644714, C2 => n6390, A => n4970, B => 
                           n4971, ZN => n4969);
   U2293 : NAND4_X1 port map( A1 => n4966, A2 => n4967, A3 => n4968, A4 => 
                           n4969, ZN => n2740);
   U2289 : AOI22_X1 port map( A1 => n6376, A2 => n3975, B1 => n6375, B2 => 
                           n3922, ZN => n4936);
   U2288 : AOI22_X1 port map( A1 => net644876, A2 => n6378, B1 => net644842, B2
                           => n6377, ZN => n4937);
   U2287 : AOI22_X1 port map( A1 => net644458, A2 => n6380, B1 => DATAIN(7), B2
                           => n4238, ZN => n4962);
   U2286 : OAI21_X1 port map( B1 => n4235, B2 => net644394, A => n4962, ZN => 
                           n4960);
   U2285 : OAI22_X1 port map( A1 => n664, A2 => n4233, B1 => n539, B2 => n4234,
                           ZN => n4961);
   U2284 : AOI211_X1 port map( C1 => net644650, C2 => n6381, A => n4960, B => 
                           n4961, ZN => n4938);
   U2283 : AOI22_X1 port map( A1 => net644554, A2 => n4228, B1 => net644522, B2
                           => n3880, ZN => n4944);
   U2282 : AOI22_X1 port map( A1 => n459, A2 => n6383, B1 => n3896, B2 => n4084
                           , ZN => n4954);
   U2281 : AOI22_X1 port map( A1 => net644619, A2 => n3895, B1 => net644490, B2
                           => n3894, ZN => n4955);
   U2280 : AOI22_X1 port map( A1 => n6384, A2 => n377, B1 => n3891, B2 => n3976
                           , ZN => n4956);
   U2279 : AOI22_X1 port map( A1 => net644587, A2 => n3890, B1 => net644683, B2
                           => n3897, ZN => n4957);
   U2278 : NAND4_X1 port map( A1 => n4954, A2 => n4955, A3 => n4956, A4 => 
                           n4957, ZN => n4946);
   U2277 : AOI22_X1 port map( A1 => n461, A2 => n3904, B1 => n3903, B2 => n4085
                           , ZN => n4948);
   U2276 : AOI22_X1 port map( A1 => net644779, A2 => n3902, B1 => net644747, B2
                           => n3901, ZN => n4949);
   U2275 : AOI22_X1 port map( A1 => net644909, A2 => n3900, B1 => net644426, B2
                           => n3899, ZN => n4950);
   U2274 : AOI22_X1 port map( A1 => n6385, A2 => n460, B1 => n3898, B2 => n3977
                           , ZN => n4951);
   U2273 : NAND4_X1 port map( A1 => n4948, A2 => n4949, A3 => n4950, A4 => 
                           n4951, ZN => n4947);
   U2272 : OAI21_X1 port map( B1 => n4946, B2 => n4947, A => n6386, ZN => n4945
                           );
   U2271 : OAI211_X1 port map( C1 => n570, C2 => n4194, A => n4944, B => n4945,
                           ZN => n4940);
   U2270 : AOI22_X1 port map( A1 => net644810, A2 => n6389, B1 => n6388, B2 => 
                           n4086, ZN => n4942);
   U2269 : OAI21_X1 port map( B1 => n632, B2 => n4189, A => n4942, ZN => n4941)
                           ;
   U2268 : AOI211_X1 port map( C1 => net644715, C2 => n4186, A => n4940, B => 
                           n4941, ZN => n4939);
   U2267 : NAND4_X1 port map( A1 => n4936, A2 => n4937, A3 => n4938, A4 => 
                           n4939, ZN => n2742);
   U2263 : AOI22_X1 port map( A1 => n6376, A2 => n3978, B1 => n6375, B2 => 
                           n3923, ZN => n4906);
   U2262 : AOI22_X1 port map( A1 => net644877, A2 => n6378, B1 => net644843, B2
                           => n6377, ZN => n4907);
   U2261 : AOI22_X1 port map( A1 => net644459, A2 => n4237, B1 => DATAIN(8), B2
                           => n4238, ZN => n4932);
   U2260 : OAI21_X1 port map( B1 => n4235, B2 => net644395, A => n4932, ZN => 
                           n4930);
   U2259 : OAI22_X1 port map( A1 => n663, A2 => n4233, B1 => n538, B2 => n4234,
                           ZN => n4931);
   U2258 : AOI211_X1 port map( C1 => net644651, C2 => n6381, A => n4930, B => 
                           n4931, ZN => n4908);
   U2257 : AOI22_X1 port map( A1 => net644555, A2 => n6382, B1 => net644523, B2
                           => n3880, ZN => n4914);
   U2256 : AOI22_X1 port map( A1 => n456, A2 => n6383, B1 => n4226, B2 => n4087
                           , ZN => n4924);
   U2255 : AOI22_X1 port map( A1 => net644620, A2 => n4223, B1 => net644491, B2
                           => n3894, ZN => n4925);
   U2254 : AOI22_X1 port map( A1 => n6384, A2 => n376, B1 => n3891, B2 => n3979
                           , ZN => n4926);
   U2253 : AOI22_X1 port map( A1 => net644588, A2 => n3890, B1 => net644684, B2
                           => n4219, ZN => n4927);
   U2252 : NAND4_X1 port map( A1 => n4924, A2 => n4925, A3 => n4926, A4 => 
                           n4927, ZN => n4916);
   U2251 : AOI22_X1 port map( A1 => n458, A2 => n3904, B1 => n3903, B2 => n4088
                           , ZN => n4918);
   U2250 : AOI22_X1 port map( A1 => net644780, A2 => n4209, B1 => net644748, B2
                           => n3901, ZN => n4919);
   U2249 : AOI22_X1 port map( A1 => net644910, A2 => n4207, B1 => net644427, B2
                           => n3899, ZN => n4920);
   U2248 : AOI22_X1 port map( A1 => n6385, A2 => n457, B1 => n3898, B2 => n3980
                           , ZN => n4921);
   U2247 : NAND4_X1 port map( A1 => n4918, A2 => n4919, A3 => n4920, A4 => 
                           n4921, ZN => n4917);
   U2246 : OAI21_X1 port map( B1 => n4916, B2 => n4917, A => n6386, ZN => n4915
                           );
   U2245 : OAI211_X1 port map( C1 => n569, C2 => n4194, A => n4914, B => n4915,
                           ZN => n4910);
   U2244 : AOI22_X1 port map( A1 => net644811, A2 => n6389, B1 => n6388, B2 => 
                           n4089, ZN => n4912);
   U2243 : OAI21_X1 port map( B1 => n631, B2 => n4189, A => n4912, ZN => n4911)
                           ;
   U2242 : AOI211_X1 port map( C1 => net644716, C2 => n4186, A => n4910, B => 
                           n4911, ZN => n4909);
   U2241 : NAND4_X1 port map( A1 => n4906, A2 => n4907, A3 => n4908, A4 => 
                           n4909, ZN => n2744);
   U2237 : AOI22_X1 port map( A1 => n6376, A2 => n3981, B1 => n6375, B2 => 
                           n3925, ZN => n4876);
   U2236 : AOI22_X1 port map( A1 => net644878, A2 => n6378, B1 => net644844, B2
                           => n4240, ZN => n4877);
   U2235 : AOI22_X1 port map( A1 => net644460, A2 => n4237, B1 => DATAIN(9), B2
                           => n6379, ZN => n4902);
   U2234 : OAI21_X1 port map( B1 => n4235, B2 => net644396, A => n4902, ZN => 
                           n4900);
   U2233 : OAI22_X1 port map( A1 => n662, A2 => n4233, B1 => n537, B2 => n4234,
                           ZN => n4901);
   U2232 : AOI211_X1 port map( C1 => net644652, C2 => n6381, A => n4900, B => 
                           n4901, ZN => n4878);
   U2231 : AOI22_X1 port map( A1 => net644556, A2 => n6382, B1 => net644524, B2
                           => n3880, ZN => n4884);
   U2230 : AOI22_X1 port map( A1 => n453, A2 => n6383, B1 => n3896, B2 => n4090
                           , ZN => n4894);
   U2229 : AOI22_X1 port map( A1 => net644621, A2 => n4223, B1 => net644492, B2
                           => n3894, ZN => n4895);
   U2228 : AOI22_X1 port map( A1 => n6384, A2 => n375, B1 => n3891, B2 => n3982
                           , ZN => n4896);
   U2227 : AOI22_X1 port map( A1 => net644589, A2 => n3890, B1 => net644685, B2
                           => n4219, ZN => n4897);
   U2226 : NAND4_X1 port map( A1 => n4894, A2 => n4895, A3 => n4896, A4 => 
                           n4897, ZN => n4886);
   U2225 : AOI22_X1 port map( A1 => n455, A2 => n3904, B1 => n3903, B2 => n4091
                           , ZN => n4888);
   U2224 : AOI22_X1 port map( A1 => net644781, A2 => n4209, B1 => net644749, B2
                           => n3901, ZN => n4889);
   U2223 : AOI22_X1 port map( A1 => net644911, A2 => n4207, B1 => net644428, B2
                           => n3899, ZN => n4890);
   U2222 : AOI22_X1 port map( A1 => n6385, A2 => n454, B1 => n3898, B2 => n3983
                           , ZN => n4891);
   U2221 : NAND4_X1 port map( A1 => n4888, A2 => n4889, A3 => n4890, A4 => 
                           n4891, ZN => n4887);
   U2220 : OAI21_X1 port map( B1 => n4886, B2 => n4887, A => n6386, ZN => n4885
                           );
   U2219 : OAI211_X1 port map( C1 => n568, C2 => n4194, A => n4884, B => n4885,
                           ZN => n4880);
   U2218 : AOI22_X1 port map( A1 => net644812, A2 => n6389, B1 => n6388, B2 => 
                           n4092, ZN => n4882);
   U2217 : OAI21_X1 port map( B1 => n630, B2 => n4189, A => n4882, ZN => n4881)
                           ;
   U2216 : AOI211_X1 port map( C1 => net644717, C2 => n4186, A => n4880, B => 
                           n4881, ZN => n4879);
   U2215 : NAND4_X1 port map( A1 => n4876, A2 => n4877, A3 => n4878, A4 => 
                           n4879, ZN => n2746);
   U2211 : AOI22_X1 port map( A1 => n4241, A2 => n3984, B1 => n6375, B2 => 
                           n3928, ZN => n4846);
   U2210 : AOI22_X1 port map( A1 => net644879, A2 => n6378, B1 => net644845, B2
                           => n4240, ZN => n4847);
   U2209 : AOI22_X1 port map( A1 => net644461, A2 => n4237, B1 => DATAIN(10), 
                           B2 => n6379, ZN => n4872);
   U2208 : OAI21_X1 port map( B1 => n4235, B2 => net644397, A => n4872, ZN => 
                           n4870);
   U2207 : OAI22_X1 port map( A1 => n661, A2 => n4233, B1 => n536, B2 => n4234,
                           ZN => n4871);
   U2206 : AOI211_X1 port map( C1 => net644653, C2 => n6381, A => n4870, B => 
                           n4871, ZN => n4848);
   U2205 : AOI22_X1 port map( A1 => net644557, A2 => n6382, B1 => net644525, B2
                           => n3880, ZN => n4854);
   U2204 : AOI22_X1 port map( A1 => n450, A2 => n6383, B1 => n3896, B2 => n4093
                           , ZN => n4864);
   U2203 : AOI22_X1 port map( A1 => net644622, A2 => n4223, B1 => net644493, B2
                           => n3894, ZN => n4865);
   U2202 : AOI22_X1 port map( A1 => n6384, A2 => n374, B1 => n3891, B2 => n3985
                           , ZN => n4866);
   U2201 : AOI22_X1 port map( A1 => net644590, A2 => n3890, B1 => net644686, B2
                           => n4219, ZN => n4867);
   U2200 : NAND4_X1 port map( A1 => n4864, A2 => n4865, A3 => n4866, A4 => 
                           n4867, ZN => n4856);
   U2199 : AOI22_X1 port map( A1 => n452, A2 => n3904, B1 => n3903, B2 => n4094
                           , ZN => n4858);
   U2198 : AOI22_X1 port map( A1 => net644782, A2 => n4209, B1 => net644750, B2
                           => n3901, ZN => n4859);
   U2197 : AOI22_X1 port map( A1 => net644912, A2 => n4207, B1 => net644429, B2
                           => n3899, ZN => n4860);
   U2196 : AOI22_X1 port map( A1 => n6385, A2 => n451, B1 => n3898, B2 => n3986
                           , ZN => n4861);
   U2195 : NAND4_X1 port map( A1 => n4858, A2 => n4859, A3 => n4860, A4 => 
                           n4861, ZN => n4857);
   U2194 : OAI21_X1 port map( B1 => n4856, B2 => n4857, A => n6386, ZN => n4855
                           );
   U2193 : OAI211_X1 port map( C1 => n567, C2 => n4194, A => n4854, B => n4855,
                           ZN => n4850);
   U2192 : AOI22_X1 port map( A1 => net644813, A2 => n6389, B1 => n6388, B2 => 
                           n4095, ZN => n4852);
   U2191 : OAI21_X1 port map( B1 => n629, B2 => n4189, A => n4852, ZN => n4851)
                           ;
   U2190 : AOI211_X1 port map( C1 => net644718, C2 => n4186, A => n4850, B => 
                           n4851, ZN => n4849);
   U2189 : NAND4_X1 port map( A1 => n4846, A2 => n4847, A3 => n4848, A4 => 
                           n4849, ZN => n2748);
   U1873 : AOI22_X1 port map( A1 => n6376, A2 => n4029, B1 => n4243, B2 => 
                           n3941, ZN => n4456);
   U1872 : AOI22_X1 port map( A1 => net644892, A2 => n6378, B1 => net644858, B2
                           => n4240, ZN => n4457);
   U1871 : AOI22_X1 port map( A1 => net644474, A2 => n6380, B1 => DATAIN(23), 
                           B2 => n6379, ZN => n4482);
   U1870 : OAI21_X1 port map( B1 => n4235, B2 => net644410, A => n4482, ZN => 
                           n4480);
   U1869 : OAI22_X1 port map( A1 => n648, A2 => n4233, B1 => n523, B2 => n4234,
                           ZN => n4481);
   U1868 : AOI211_X1 port map( C1 => net644666, C2 => n6381, A => n4480, B => 
                           n4481, ZN => n4458);
   U1867 : AOI22_X1 port map( A1 => net644570, A2 => n6382, B1 => net644538, B2
                           => n4229, ZN => n4464);
   U1866 : AOI22_X1 port map( A1 => n411, A2 => n6383, B1 => n3896, B2 => n4137
                           , ZN => n4474);
   U1865 : AOI22_X1 port map( A1 => net644635, A2 => n3895, B1 => net644506, B2
                           => n4224, ZN => n4475);
   U1864 : AOI22_X1 port map( A1 => n4220, A2 => n361, B1 => n3891, B2 => n4030
                           , ZN => n4476);
   U1863 : AOI22_X1 port map( A1 => net644603, A2 => n4218, B1 => net644699, B2
                           => n3897, ZN => n4477);
   U1862 : NAND4_X1 port map( A1 => n4474, A2 => n4475, A3 => n4476, A4 => 
                           n4477, ZN => n4466);
   U1861 : AOI22_X1 port map( A1 => n413, A2 => n4211, B1 => n3903, B2 => n4138
                           , ZN => n4468);
   U1860 : AOI22_X1 port map( A1 => net644795, A2 => n3902, B1 => net644763, B2
                           => n4210, ZN => n4469);
   U1859 : AOI22_X1 port map( A1 => net644925, A2 => n3900, B1 => net644442, B2
                           => n4208, ZN => n4470);
   U1858 : AOI22_X1 port map( A1 => n6385, A2 => n412, B1 => n3898, B2 => n4031
                           , ZN => n4471);
   U1857 : NAND4_X1 port map( A1 => n4468, A2 => n4469, A3 => n4470, A4 => 
                           n4471, ZN => n4467);
   U1856 : OAI21_X1 port map( B1 => n4466, B2 => n4467, A => n6386, ZN => n4465
                           );
   U1855 : OAI211_X1 port map( C1 => n554, C2 => n4194, A => n4464, B => n4465,
                           ZN => n4460);
   U1854 : AOI22_X1 port map( A1 => net644826, A2 => n6389, B1 => n6388, B2 => 
                           n4139, ZN => n4462);
   U1853 : OAI21_X1 port map( B1 => n616, B2 => n4189, A => n4462, ZN => n4461)
                           ;
   U1852 : AOI211_X1 port map( C1 => net644731, C2 => n6390, A => n4460, B => 
                           n4461, ZN => n4459);
   U1851 : NAND4_X1 port map( A1 => n4456, A2 => n4457, A3 => n4458, A4 => 
                           n4459, ZN => n2774);
   U1847 : AOI22_X1 port map( A1 => n4241, A2 => n4032, B1 => n6375, B2 => 
                           n3942, ZN => n4426);
   U1846 : AOI22_X1 port map( A1 => net644893, A2 => n6378, B1 => net644859, B2
                           => n6377, ZN => n4427);
   U1845 : AOI22_X1 port map( A1 => net644475, A2 => n6380, B1 => DATAIN(24), 
                           B2 => n6379, ZN => n4452);
   U1844 : OAI21_X1 port map( B1 => n4235, B2 => net644411, A => n4452, ZN => 
                           n4450);
   U1843 : OAI22_X1 port map( A1 => n647, A2 => n4233, B1 => n522, B2 => n4234,
                           ZN => n4451);
   U1842 : AOI211_X1 port map( C1 => net644667, C2 => n6381, A => n4450, B => 
                           n4451, ZN => n4428);
   U1841 : AOI22_X1 port map( A1 => net644571, A2 => n6382, B1 => net644539, B2
                           => n3880, ZN => n4434);
   U1840 : AOI22_X1 port map( A1 => n408, A2 => n6383, B1 => n3896, B2 => n4140
                           , ZN => n4444);
   U1839 : AOI22_X1 port map( A1 => net644636, A2 => n3895, B1 => net644507, B2
                           => n3894, ZN => n4445);
   U1838 : AOI22_X1 port map( A1 => n4220, A2 => n360, B1 => n4221, B2 => n4034
                           , ZN => n4446);
   U1837 : AOI22_X1 port map( A1 => net644604, A2 => n3890, B1 => net644700, B2
                           => n3897, ZN => n4447);
   U1836 : NAND4_X1 port map( A1 => n4444, A2 => n4445, A3 => n4446, A4 => 
                           n4447, ZN => n4436);
   U1835 : AOI22_X1 port map( A1 => n410, A2 => n4211, B1 => n4212, B2 => n4141
                           , ZN => n4438);
   U1834 : AOI22_X1 port map( A1 => net644796, A2 => n3902, B1 => net644764, B2
                           => n3901, ZN => n4439);
   U1833 : AOI22_X1 port map( A1 => net644926, A2 => n3900, B1 => net644443, B2
                           => n3899, ZN => n4440);
   U1832 : AOI22_X1 port map( A1 => n6385, A2 => n409, B1 => n3898, B2 => n4037
                           , ZN => n4441);
   U1831 : NAND4_X1 port map( A1 => n4438, A2 => n4439, A3 => n4440, A4 => 
                           n4441, ZN => n4437);
   U1830 : OAI21_X1 port map( B1 => n4436, B2 => n4437, A => n6386, ZN => n4435
                           );
   U1829 : OAI211_X1 port map( C1 => n553, C2 => n4194, A => n4434, B => n4435,
                           ZN => n4430);
   U1828 : AOI22_X1 port map( A1 => net644827, A2 => n6389, B1 => n6388, B2 => 
                           n4142, ZN => n4432);
   U1827 : OAI21_X1 port map( B1 => n615, B2 => n4189, A => n4432, ZN => n4431)
                           ;
   U1826 : AOI211_X1 port map( C1 => net644732, C2 => n6390, A => n4430, B => 
                           n4431, ZN => n4429);
   U1825 : NAND4_X1 port map( A1 => n4426, A2 => n4427, A3 => n4428, A4 => 
                           n4429, ZN => n2776);
   U2133 : AOI22_X1 port map( A1 => n6376, A2 => n3993, B1 => n6375, B2 => 
                           n3931, ZN => n4756);
   U2132 : AOI22_X1 port map( A1 => net644882, A2 => n6378, B1 => net644848, B2
                           => n6377, ZN => n4757);
   U2131 : AOI22_X1 port map( A1 => net644464, A2 => n6380, B1 => DATAIN(13), 
                           B2 => n6379, ZN => n4782);
   U2130 : OAI21_X1 port map( B1 => n4235, B2 => net644400, A => n4782, ZN => 
                           n4780);
   U2129 : OAI22_X1 port map( A1 => n658, A2 => n4233, B1 => n533, B2 => n4234,
                           ZN => n4781);
   U2128 : AOI211_X1 port map( C1 => net644656, C2 => n6381, A => n4780, B => 
                           n4781, ZN => n4758);
   U2127 : AOI22_X1 port map( A1 => net644560, A2 => n6382, B1 => net644528, B2
                           => n3880, ZN => n4764);
   U2126 : AOI22_X1 port map( A1 => n441, A2 => n4225, B1 => n3896, B2 => n4102
                           , ZN => n4774);
   U2125 : AOI22_X1 port map( A1 => net644625, A2 => n3895, B1 => net644496, B2
                           => n3894, ZN => n4775);
   U2124 : AOI22_X1 port map( A1 => n6384, A2 => n371, B1 => n3891, B2 => n3998
                           , ZN => n4776);
   U2123 : AOI22_X1 port map( A1 => net644593, A2 => n3890, B1 => net644689, B2
                           => n3897, ZN => n4777);
   U2122 : NAND4_X1 port map( A1 => n4774, A2 => n4775, A3 => n4776, A4 => 
                           n4777, ZN => n4766);
   U2121 : AOI22_X1 port map( A1 => n443, A2 => n3904, B1 => n3903, B2 => n4103
                           , ZN => n4768);
   U2120 : AOI22_X1 port map( A1 => net644785, A2 => n3902, B1 => net644753, B2
                           => n3901, ZN => n4769);
   U2119 : AOI22_X1 port map( A1 => net644915, A2 => n3900, B1 => net644432, B2
                           => n3899, ZN => n4770);
   U2118 : AOI22_X1 port map( A1 => n6385, A2 => n442, B1 => n3898, B2 => n3999
                           , ZN => n4771);
   U2117 : NAND4_X1 port map( A1 => n4768, A2 => n4769, A3 => n4770, A4 => 
                           n4771, ZN => n4767);
   U2116 : OAI21_X1 port map( B1 => n4766, B2 => n4767, A => n6386, ZN => n4765
                           );
   U2115 : OAI211_X1 port map( C1 => n564, C2 => n4194, A => n4764, B => n4765,
                           ZN => n4760);
   U2114 : AOI22_X1 port map( A1 => net644816, A2 => n6389, B1 => n6388, B2 => 
                           n4104, ZN => n4762);
   U2113 : OAI21_X1 port map( B1 => n626, B2 => n4189, A => n4762, ZN => n4761)
                           ;
   U2112 : AOI211_X1 port map( C1 => net644721, C2 => n6390, A => n4760, B => 
                           n4761, ZN => n4759);
   U2111 : NAND4_X1 port map( A1 => n4756, A2 => n4757, A3 => n4758, A4 => 
                           n4759, ZN => n2754);
   U2107 : AOI22_X1 port map( A1 => n6376, A2 => n4002, B1 => n6375, B2 => 
                           n3932, ZN => n4726);
   U2106 : AOI22_X1 port map( A1 => net644883, A2 => n6378, B1 => net644849, B2
                           => n6377, ZN => n4727);
   U2105 : AOI22_X1 port map( A1 => net644465, A2 => n6380, B1 => DATAIN(14), 
                           B2 => n6379, ZN => n4752);
   U2104 : OAI21_X1 port map( B1 => n4235, B2 => net644401, A => n4752, ZN => 
                           n4750);
   U2103 : OAI22_X1 port map( A1 => n657, A2 => n4233, B1 => n532, B2 => n4234,
                           ZN => n4751);
   U2102 : AOI211_X1 port map( C1 => net644657, C2 => n6381, A => n4750, B => 
                           n4751, ZN => n4728);
   U2101 : AOI22_X1 port map( A1 => net644561, A2 => n6382, B1 => net644529, B2
                           => n3880, ZN => n4734);
   U2100 : AOI22_X1 port map( A1 => n438, A2 => n4225, B1 => n3896, B2 => n4105
                           , ZN => n4744);
   U2099 : AOI22_X1 port map( A1 => net644626, A2 => n3895, B1 => net644497, B2
                           => n3894, ZN => n4745);
   U2098 : AOI22_X1 port map( A1 => n6384, A2 => n370, B1 => n3891, B2 => n4003
                           , ZN => n4746);
   U2097 : AOI22_X1 port map( A1 => net644594, A2 => n3890, B1 => net644690, B2
                           => n3897, ZN => n4747);
   U2096 : NAND4_X1 port map( A1 => n4744, A2 => n4745, A3 => n4746, A4 => 
                           n4747, ZN => n4736);
   U2095 : AOI22_X1 port map( A1 => n440, A2 => n3904, B1 => n3903, B2 => n4109
                           , ZN => n4738);
   U2094 : AOI22_X1 port map( A1 => net644786, A2 => n3902, B1 => net644754, B2
                           => n3901, ZN => n4739);
   U2093 : AOI22_X1 port map( A1 => net644916, A2 => n3900, B1 => net644433, B2
                           => n3899, ZN => n4740);
   U2092 : AOI22_X1 port map( A1 => n6385, A2 => n439, B1 => n3898, B2 => n4004
                           , ZN => n4741);
   U2091 : NAND4_X1 port map( A1 => n4738, A2 => n4739, A3 => n4740, A4 => 
                           n4741, ZN => n4737);
   U2090 : OAI21_X1 port map( B1 => n4736, B2 => n4737, A => n6386, ZN => n4735
                           );
   U2089 : OAI211_X1 port map( C1 => n563, C2 => n4194, A => n4734, B => n4735,
                           ZN => n4730);
   U2088 : AOI22_X1 port map( A1 => net644817, A2 => n6389, B1 => n6388, B2 => 
                           n4112, ZN => n4732);
   U2087 : OAI21_X1 port map( B1 => n625, B2 => n4189, A => n4732, ZN => n4731)
                           ;
   U2086 : AOI211_X1 port map( C1 => net644722, C2 => n6390, A => n4730, B => 
                           n4731, ZN => n4729);
   U2085 : NAND4_X1 port map( A1 => n4726, A2 => n4727, A3 => n4728, A4 => 
                           n4729, ZN => n2756);
   U2081 : AOI22_X1 port map( A1 => n6376, A2 => n4005, B1 => n4243, B2 => 
                           n3933, ZN => n4696);
   U2080 : AOI22_X1 port map( A1 => net644884, A2 => n6378, B1 => net644850, B2
                           => n4240, ZN => n4697);
   U2079 : AOI22_X1 port map( A1 => net644466, A2 => n6380, B1 => DATAIN(15), 
                           B2 => n6379, ZN => n4722);
   U2078 : OAI21_X1 port map( B1 => n4235, B2 => net644402, A => n4722, ZN => 
                           n4720);
   U2077 : OAI22_X1 port map( A1 => n656, A2 => n4233, B1 => n531, B2 => n4234,
                           ZN => n4721);
   U2076 : AOI211_X1 port map( C1 => net644658, C2 => n6381, A => n4720, B => 
                           n4721, ZN => n4698);
   U2075 : AOI22_X1 port map( A1 => net644562, A2 => n6382, B1 => net644530, B2
                           => n3880, ZN => n4704);
   U2074 : AOI22_X1 port map( A1 => n435, A2 => n6383, B1 => n3896, B2 => n4113
                           , ZN => n4714);
   U2073 : AOI22_X1 port map( A1 => net644627, A2 => n3895, B1 => net644498, B2
                           => n3894, ZN => n4715);
   U2072 : AOI22_X1 port map( A1 => n4220, A2 => n369, B1 => n3891, B2 => n4006
                           , ZN => n4716);
   U2071 : AOI22_X1 port map( A1 => net644595, A2 => n3890, B1 => net644691, B2
                           => n3897, ZN => n4717);
   U2070 : NAND4_X1 port map( A1 => n4714, A2 => n4715, A3 => n4716, A4 => 
                           n4717, ZN => n4706);
   U2069 : AOI22_X1 port map( A1 => n437, A2 => n3904, B1 => n3903, B2 => n4114
                           , ZN => n4708);
   U2068 : AOI22_X1 port map( A1 => net644787, A2 => n3902, B1 => net644755, B2
                           => n3901, ZN => n4709);
   U2067 : AOI22_X1 port map( A1 => net644917, A2 => n3900, B1 => net644434, B2
                           => n3899, ZN => n4710);
   U2066 : AOI22_X1 port map( A1 => n6385, A2 => n436, B1 => n3898, B2 => n4007
                           , ZN => n4711);
   U2065 : NAND4_X1 port map( A1 => n4708, A2 => n4709, A3 => n4710, A4 => 
                           n4711, ZN => n4707);
   U2064 : OAI21_X1 port map( B1 => n4706, B2 => n4707, A => n6386, ZN => n4705
                           );
   U2063 : OAI211_X1 port map( C1 => n562, C2 => n4194, A => n4704, B => n4705,
                           ZN => n4700);
   U2062 : AOI22_X1 port map( A1 => net644818, A2 => n6389, B1 => n6388, B2 => 
                           n4115, ZN => n4702);
   U2061 : OAI21_X1 port map( B1 => n624, B2 => n4189, A => n4702, ZN => n4701)
                           ;
   U2060 : AOI211_X1 port map( C1 => net644723, C2 => n6390, A => n4700, B => 
                           n4701, ZN => n4699);
   U2059 : NAND4_X1 port map( A1 => n4696, A2 => n4697, A3 => n4698, A4 => 
                           n4699, ZN => n2758);
   U1925 : AOI22_X1 port map( A1 => n6376, A2 => n4023, B1 => n6375, B2 => 
                           n3939, ZN => n4516);
   U1924 : AOI22_X1 port map( A1 => net644890, A2 => n4239, B1 => net644856, B2
                           => n4240, ZN => n4517);
   U1923 : AOI22_X1 port map( A1 => net644472, A2 => n4237, B1 => DATAIN(21), 
                           B2 => n6379, ZN => n4542);
   U1922 : OAI21_X1 port map( B1 => n4235, B2 => net644408, A => n4542, ZN => 
                           n4540);
   U1921 : OAI22_X1 port map( A1 => n650, A2 => n4233, B1 => n525, B2 => n4234,
                           ZN => n4541);
   U1920 : AOI211_X1 port map( C1 => net644664, C2 => n6381, A => n4540, B => 
                           n4541, ZN => n4518);
   U1919 : AOI22_X1 port map( A1 => net644568, A2 => n6382, B1 => net644536, B2
                           => n4229, ZN => n4524);
   U1918 : AOI22_X1 port map( A1 => n417, A2 => n6383, B1 => n3896, B2 => n4131
                           , ZN => n4534);
   U1917 : AOI22_X1 port map( A1 => net644633, A2 => n3895, B1 => net644504, B2
                           => n4224, ZN => n4535);
   U1916 : AOI22_X1 port map( A1 => n4220, A2 => n363, B1 => n3891, B2 => n4024
                           , ZN => n4536);
   U1915 : AOI22_X1 port map( A1 => net644601, A2 => n4218, B1 => net644697, B2
                           => n3897, ZN => n4537);
   U1914 : NAND4_X1 port map( A1 => n4534, A2 => n4535, A3 => n4536, A4 => 
                           n4537, ZN => n4526);
   U1913 : AOI22_X1 port map( A1 => n419, A2 => n3904, B1 => n3903, B2 => n4132
                           , ZN => n4528);
   U1912 : AOI22_X1 port map( A1 => net644793, A2 => n3902, B1 => net644761, B2
                           => n4210, ZN => n4529);
   U1911 : AOI22_X1 port map( A1 => net644923, A2 => n3900, B1 => net644440, B2
                           => n4208, ZN => n4530);
   U1910 : AOI22_X1 port map( A1 => n6385, A2 => n418, B1 => n3898, B2 => n4025
                           , ZN => n4531);
   U1909 : NAND4_X1 port map( A1 => n4528, A2 => n4529, A3 => n4530, A4 => 
                           n4531, ZN => n4527);
   U1908 : OAI21_X1 port map( B1 => n4526, B2 => n4527, A => n6386, ZN => n4525
                           );
   U1907 : OAI211_X1 port map( C1 => n556, C2 => n4194, A => n4524, B => n4525,
                           ZN => n4520);
   U1906 : AOI22_X1 port map( A1 => net644824, A2 => n6389, B1 => n6388, B2 => 
                           n4133, ZN => n4522);
   U1905 : OAI21_X1 port map( B1 => n618, B2 => n4189, A => n4522, ZN => n4521)
                           ;
   U1904 : AOI211_X1 port map( C1 => net644729, C2 => n4186, A => n4520, B => 
                           n4521, ZN => n4519);
   U1903 : NAND4_X1 port map( A1 => n4516, A2 => n4517, A3 => n4518, A4 => 
                           n4519, ZN => n2770);
   U2029 : AOI22_X1 port map( A1 => n6376, A2 => n4011, B1 => n6375, B2 => 
                           n3935, ZN => n4636);
   U2028 : AOI22_X1 port map( A1 => net644886, A2 => n6378, B1 => net644852, B2
                           => n6377, ZN => n4637);
   U2027 : AOI22_X1 port map( A1 => net644468, A2 => n6380, B1 => DATAIN(17), 
                           B2 => n6379, ZN => n4662);
   U2026 : OAI21_X1 port map( B1 => n4235, B2 => net644404, A => n4662, ZN => 
                           n4660);
   U2025 : OAI22_X1 port map( A1 => n654, A2 => n4233, B1 => n529, B2 => n4234,
                           ZN => n4661);
   U2024 : AOI211_X1 port map( C1 => net644660, C2 => n6381, A => n4660, B => 
                           n4661, ZN => n4638);
   U2023 : AOI22_X1 port map( A1 => net644564, A2 => n6382, B1 => net644532, B2
                           => n3880, ZN => n4644);
   U2022 : AOI22_X1 port map( A1 => n429, A2 => n4225, B1 => n3896, B2 => n4119
                           , ZN => n4654);
   U2021 : AOI22_X1 port map( A1 => net644629, A2 => n3895, B1 => net644500, B2
                           => n3894, ZN => n4655);
   U2020 : AOI22_X1 port map( A1 => n6384, A2 => n367, B1 => n3891, B2 => n4012
                           , ZN => n4656);
   U2019 : AOI22_X1 port map( A1 => net644597, A2 => n3890, B1 => net644693, B2
                           => n3897, ZN => n4657);
   U2018 : NAND4_X1 port map( A1 => n4654, A2 => n4655, A3 => n4656, A4 => 
                           n4657, ZN => n4646);
   U2017 : AOI22_X1 port map( A1 => n431, A2 => n3904, B1 => n3903, B2 => n4120
                           , ZN => n4648);
   U2016 : AOI22_X1 port map( A1 => net644789, A2 => n3902, B1 => net644757, B2
                           => n3901, ZN => n4649);
   U2015 : AOI22_X1 port map( A1 => net644919, A2 => n3900, B1 => net644436, B2
                           => n3899, ZN => n4650);
   U2014 : AOI22_X1 port map( A1 => n6385, A2 => n430, B1 => n3898, B2 => n4013
                           , ZN => n4651);
   U2013 : NAND4_X1 port map( A1 => n4648, A2 => n4649, A3 => n4650, A4 => 
                           n4651, ZN => n4647);
   U2012 : OAI21_X1 port map( B1 => n4646, B2 => n4647, A => n6386, ZN => n4645
                           );
   U2011 : OAI211_X1 port map( C1 => n560, C2 => n4194, A => n4644, B => n4645,
                           ZN => n4640);
   U2010 : AOI22_X1 port map( A1 => net644820, A2 => n6389, B1 => n6388, B2 => 
                           n4121, ZN => n4642);
   U2009 : OAI21_X1 port map( B1 => n622, B2 => n4189, A => n4642, ZN => n4641)
                           ;
   U2008 : AOI211_X1 port map( C1 => net644725, C2 => n6390, A => n4640, B => 
                           n4641, ZN => n4639);
   U2007 : NAND4_X1 port map( A1 => n4636, A2 => n4637, A3 => n4638, A4 => 
                           n4639, ZN => n2762);
   U2003 : AOI22_X1 port map( A1 => n6376, A2 => n4014, B1 => n6375, B2 => 
                           n3936, ZN => n4606);
   U2002 : AOI22_X1 port map( A1 => net644887, A2 => n6378, B1 => net644853, B2
                           => n6377, ZN => n4607);
   U2001 : AOI22_X1 port map( A1 => net644469, A2 => n6380, B1 => DATAIN(18), 
                           B2 => n6379, ZN => n4632);
   U2000 : OAI21_X1 port map( B1 => n4235, B2 => net644405, A => n4632, ZN => 
                           n4630);
   U1999 : OAI22_X1 port map( A1 => n653, A2 => n4233, B1 => n528, B2 => n4234,
                           ZN => n4631);
   U1998 : AOI211_X1 port map( C1 => net644661, C2 => n6381, A => n4630, B => 
                           n4631, ZN => n4608);
   U1997 : AOI22_X1 port map( A1 => net644565, A2 => n6382, B1 => net644533, B2
                           => n3880, ZN => n4614);
   U1996 : AOI22_X1 port map( A1 => n426, A2 => n4225, B1 => n3896, B2 => n4122
                           , ZN => n4624);
   U1995 : AOI22_X1 port map( A1 => net644630, A2 => n3895, B1 => net644501, B2
                           => n3894, ZN => n4625);
   U1994 : AOI22_X1 port map( A1 => n6384, A2 => n366, B1 => n3891, B2 => n4015
                           , ZN => n4626);
   U1993 : AOI22_X1 port map( A1 => net644598, A2 => n3890, B1 => net644694, B2
                           => n3897, ZN => n4627);
   U1992 : NAND4_X1 port map( A1 => n4624, A2 => n4625, A3 => n4626, A4 => 
                           n4627, ZN => n4616);
   U1991 : AOI22_X1 port map( A1 => n428, A2 => n3904, B1 => n3903, B2 => n4123
                           , ZN => n4618);
   U1990 : AOI22_X1 port map( A1 => net644790, A2 => n3902, B1 => net644758, B2
                           => n3901, ZN => n4619);
   U1989 : AOI22_X1 port map( A1 => net644920, A2 => n3900, B1 => net644437, B2
                           => n3899, ZN => n4620);
   U1988 : AOI22_X1 port map( A1 => n6385, A2 => n427, B1 => n3898, B2 => n4016
                           , ZN => n4621);
   U1987 : NAND4_X1 port map( A1 => n4618, A2 => n4619, A3 => n4620, A4 => 
                           n4621, ZN => n4617);
   U1986 : OAI21_X1 port map( B1 => n4616, B2 => n4617, A => n6386, ZN => n4615
                           );
   U1985 : OAI211_X1 port map( C1 => n559, C2 => n4194, A => n4614, B => n4615,
                           ZN => n4610);
   U1984 : AOI22_X1 port map( A1 => net644821, A2 => n6389, B1 => n6388, B2 => 
                           n4124, ZN => n4612);
   U1983 : OAI21_X1 port map( B1 => n621, B2 => n4189, A => n4612, ZN => n4611)
                           ;
   U1982 : AOI211_X1 port map( C1 => net644726, C2 => n6390, A => n4610, B => 
                           n4611, ZN => n4609);
   U1981 : NAND4_X1 port map( A1 => n4606, A2 => n4607, A3 => n4608, A4 => 
                           n4609, ZN => n2764);
   U1977 : AOI22_X1 port map( A1 => n6376, A2 => n4017, B1 => n6375, B2 => 
                           n3937, ZN => n4576);
   U1976 : AOI22_X1 port map( A1 => net644888, A2 => n6378, B1 => net644854, B2
                           => n6377, ZN => n4577);
   U1975 : AOI22_X1 port map( A1 => net644470, A2 => n6380, B1 => DATAIN(19), 
                           B2 => n6379, ZN => n4602);
   U1974 : OAI21_X1 port map( B1 => n4235, B2 => net644406, A => n4602, ZN => 
                           n4600);
   U1973 : OAI22_X1 port map( A1 => n652, A2 => n4233, B1 => n527, B2 => n4234,
                           ZN => n4601);
   U1972 : AOI211_X1 port map( C1 => net644662, C2 => n6381, A => n4600, B => 
                           n4601, ZN => n4578);
   U1971 : AOI22_X1 port map( A1 => net644566, A2 => n6382, B1 => net644534, B2
                           => n3880, ZN => n4584);
   U1970 : AOI22_X1 port map( A1 => n423, A2 => n4225, B1 => n3896, B2 => n4125
                           , ZN => n4594);
   U1969 : AOI22_X1 port map( A1 => net644631, A2 => n3895, B1 => net644502, B2
                           => n3894, ZN => n4595);
   U1968 : AOI22_X1 port map( A1 => n6384, A2 => n365, B1 => n3891, B2 => n4018
                           , ZN => n4596);
   U1967 : AOI22_X1 port map( A1 => net644599, A2 => n3890, B1 => net644695, B2
                           => n3897, ZN => n4597);
   U1966 : NAND4_X1 port map( A1 => n4594, A2 => n4595, A3 => n4596, A4 => 
                           n4597, ZN => n4586);
   U1965 : AOI22_X1 port map( A1 => n425, A2 => n3904, B1 => n3903, B2 => n4126
                           , ZN => n4588);
   U1964 : AOI22_X1 port map( A1 => net644791, A2 => n3902, B1 => net644759, B2
                           => n3901, ZN => n4589);
   U1963 : AOI22_X1 port map( A1 => net644921, A2 => n3900, B1 => net644438, B2
                           => n3899, ZN => n4590);
   U1962 : AOI22_X1 port map( A1 => n6385, A2 => n424, B1 => n3898, B2 => n4019
                           , ZN => n4591);
   U1961 : NAND4_X1 port map( A1 => n4588, A2 => n4589, A3 => n4590, A4 => 
                           n4591, ZN => n4587);
   U1960 : OAI21_X1 port map( B1 => n4586, B2 => n4587, A => n6386, ZN => n4585
                           );
   U1959 : OAI211_X1 port map( C1 => n558, C2 => n4194, A => n4584, B => n4585,
                           ZN => n4580);
   U1958 : AOI22_X1 port map( A1 => net644822, A2 => n6389, B1 => n6388, B2 => 
                           n4127, ZN => n4582);
   U1957 : OAI21_X1 port map( B1 => n620, B2 => n4189, A => n4582, ZN => n4581)
                           ;
   U1956 : AOI211_X1 port map( C1 => net644727, C2 => n6390, A => n4580, B => 
                           n4581, ZN => n4579);
   U1955 : NAND4_X1 port map( A1 => n4576, A2 => n4577, A3 => n4578, A4 => 
                           n4579, ZN => n2766);
   U1951 : AOI22_X1 port map( A1 => n6376, A2 => n4020, B1 => n6375, B2 => 
                           n3938, ZN => n4546);
   U1950 : AOI22_X1 port map( A1 => net644889, A2 => n4239, B1 => net644855, B2
                           => n4240, ZN => n4547);
   U1949 : AOI22_X1 port map( A1 => net644471, A2 => n6380, B1 => DATAIN(20), 
                           B2 => n6379, ZN => n4572);
   U1948 : OAI21_X1 port map( B1 => n4235, B2 => net644407, A => n4572, ZN => 
                           n4570);
   U1947 : OAI22_X1 port map( A1 => n651, A2 => n4233, B1 => n526, B2 => n4234,
                           ZN => n4571);
   U1946 : AOI211_X1 port map( C1 => net644663, C2 => n6381, A => n4570, B => 
                           n4571, ZN => n4548);
   U1945 : AOI22_X1 port map( A1 => net644567, A2 => n6382, B1 => net644535, B2
                           => n4229, ZN => n4554);
   U1944 : AOI22_X1 port map( A1 => n420, A2 => n6383, B1 => n3896, B2 => n4128
                           , ZN => n4564);
   U1943 : AOI22_X1 port map( A1 => net644632, A2 => n3895, B1 => net644503, B2
                           => n4224, ZN => n4565);
   U1942 : AOI22_X1 port map( A1 => n4220, A2 => n364, B1 => n3891, B2 => n4021
                           , ZN => n4566);
   U1941 : AOI22_X1 port map( A1 => net644600, A2 => n3890, B1 => net644696, B2
                           => n3897, ZN => n4567);
   U1940 : NAND4_X1 port map( A1 => n4564, A2 => n4565, A3 => n4566, A4 => 
                           n4567, ZN => n4556);
   U1939 : AOI22_X1 port map( A1 => n422, A2 => n3904, B1 => n3903, B2 => n4129
                           , ZN => n4558);
   U1938 : AOI22_X1 port map( A1 => net644792, A2 => n3902, B1 => net644760, B2
                           => n4210, ZN => n4559);
   U1937 : AOI22_X1 port map( A1 => net644922, A2 => n3900, B1 => net644439, B2
                           => n4208, ZN => n4560);
   U1936 : AOI22_X1 port map( A1 => n4204, A2 => n421, B1 => n3898, B2 => n4022
                           , ZN => n4561);
   U1935 : NAND4_X1 port map( A1 => n4558, A2 => n4559, A3 => n4560, A4 => 
                           n4561, ZN => n4557);
   U1934 : OAI21_X1 port map( B1 => n4556, B2 => n4557, A => n6386, ZN => n4555
                           );
   U1933 : OAI211_X1 port map( C1 => n557, C2 => n4194, A => n4554, B => n4555,
                           ZN => n4550);
   U1932 : AOI22_X1 port map( A1 => net644823, A2 => n6389, B1 => n6388, B2 => 
                           n4130, ZN => n4552);
   U1931 : OAI21_X1 port map( B1 => n619, B2 => n4189, A => n4552, ZN => n4551)
                           ;
   U1930 : AOI211_X1 port map( C1 => net644728, C2 => n6390, A => n4550, B => 
                           n4551, ZN => n4549);
   U1929 : NAND4_X1 port map( A1 => n4546, A2 => n4547, A3 => n4548, A4 => 
                           n4549, ZN => n2768);
   U1769 : AOI22_X1 port map( A1 => n4241, A2 => n4044, B1 => n4243, B2 => 
                           n3945, ZN => n4336);
   U1768 : AOI22_X1 port map( A1 => net644896, A2 => n4239, B1 => net644862, B2
                           => n6377, ZN => n4337);
   U1767 : AOI22_X1 port map( A1 => net644478, A2 => n6380, B1 => DATAIN(27), 
                           B2 => n6379, ZN => n4362);
   U1766 : OAI21_X1 port map( B1 => n4235, B2 => net644414, A => n4362, ZN => 
                           n4360);
   U1765 : OAI22_X1 port map( A1 => n644, A2 => n4233, B1 => n519, B2 => n4234,
                           ZN => n4361);
   U1764 : AOI211_X1 port map( C1 => net644670, C2 => n6381, A => n4360, B => 
                           n4361, ZN => n4338);
   U1763 : AOI22_X1 port map( A1 => net644574, A2 => n6382, B1 => net644542, B2
                           => n3880, ZN => n4344);
   U1762 : AOI22_X1 port map( A1 => n399, A2 => n6383, B1 => n3896, B2 => n4152
                           , ZN => n4354);
   U1761 : AOI22_X1 port map( A1 => net644639, A2 => n3895, B1 => net644510, B2
                           => n3894, ZN => n4355);
   U1760 : AOI22_X1 port map( A1 => n4220, A2 => n357, B1 => n4221, B2 => n4045
                           , ZN => n4356);
   U1759 : AOI22_X1 port map( A1 => net644607, A2 => n3890, B1 => net644703, B2
                           => n3897, ZN => n4357);
   U1758 : NAND4_X1 port map( A1 => n4354, A2 => n4355, A3 => n4356, A4 => 
                           n4357, ZN => n4346);
   U1757 : AOI22_X1 port map( A1 => n401, A2 => n4211, B1 => n4212, B2 => n4153
                           , ZN => n4348);
   U1756 : AOI22_X1 port map( A1 => net644799, A2 => n3902, B1 => net644767, B2
                           => n3901, ZN => n4349);
   U1755 : AOI22_X1 port map( A1 => net644929, A2 => n3900, B1 => net644446, B2
                           => n3899, ZN => n4350);
   U1754 : AOI22_X1 port map( A1 => n4204, A2 => n400, B1 => n4205, B2 => n4046
                           , ZN => n4351);
   U1753 : NAND4_X1 port map( A1 => n4348, A2 => n4349, A3 => n4350, A4 => 
                           n4351, ZN => n4347);
   U1752 : OAI21_X1 port map( B1 => n4346, B2 => n4347, A => n6386, ZN => n4345
                           );
   U1751 : OAI211_X1 port map( C1 => n550, C2 => n4194, A => n4344, B => n4345,
                           ZN => n4340);
   U1750 : AOI22_X1 port map( A1 => net644830, A2 => n6389, B1 => n4192, B2 => 
                           n4154, ZN => n4342);
   U1749 : OAI21_X1 port map( B1 => n612, B2 => n4189, A => n4342, ZN => n4341)
                           ;
   U1748 : AOI211_X1 port map( C1 => net644735, C2 => n6390, A => n4340, B => 
                           n4341, ZN => n4339);
   U1747 : NAND4_X1 port map( A1 => n4336, A2 => n4337, A3 => n4338, A4 => 
                           n4339, ZN => n2782);
   U1899 : AOI22_X1 port map( A1 => n6376, A2 => n4026, B1 => n4243, B2 => 
                           n3940, ZN => n4486);
   U1898 : AOI22_X1 port map( A1 => net644891, A2 => n6378, B1 => net644857, B2
                           => n4240, ZN => n4487);
   U1897 : AOI22_X1 port map( A1 => net644473, A2 => n4237, B1 => DATAIN(22), 
                           B2 => n6379, ZN => n4512);
   U1896 : OAI21_X1 port map( B1 => n4235, B2 => net644409, A => n4512, ZN => 
                           n4510);
   U1895 : OAI22_X1 port map( A1 => n649, A2 => n4233, B1 => n524, B2 => n4234,
                           ZN => n4511);
   U1894 : AOI211_X1 port map( C1 => net644665, C2 => n6381, A => n4510, B => 
                           n4511, ZN => n4488);
   U1893 : AOI22_X1 port map( A1 => net644569, A2 => n6382, B1 => net644537, B2
                           => n4229, ZN => n4494);
   U1892 : AOI22_X1 port map( A1 => n414, A2 => n6383, B1 => n3896, B2 => n4134
                           , ZN => n4504);
   U1891 : AOI22_X1 port map( A1 => net644634, A2 => n3895, B1 => net644505, B2
                           => n4224, ZN => n4505);
   U1890 : AOI22_X1 port map( A1 => n4220, A2 => n362, B1 => n3891, B2 => n4027
                           , ZN => n4506);
   U1889 : AOI22_X1 port map( A1 => net644602, A2 => n4218, B1 => net644698, B2
                           => n3897, ZN => n4507);
   U1888 : NAND4_X1 port map( A1 => n4504, A2 => n4505, A3 => n4506, A4 => 
                           n4507, ZN => n4496);
   U1887 : AOI22_X1 port map( A1 => n416, A2 => n4211, B1 => n3903, B2 => n4135
                           , ZN => n4498);
   U1886 : AOI22_X1 port map( A1 => net644794, A2 => n3902, B1 => net644762, B2
                           => n4210, ZN => n4499);
   U1885 : AOI22_X1 port map( A1 => net644924, A2 => n3900, B1 => net644441, B2
                           => n4208, ZN => n4500);
   U1884 : AOI22_X1 port map( A1 => n4204, A2 => n415, B1 => n3898, B2 => n4028
                           , ZN => n4501);
   U1883 : NAND4_X1 port map( A1 => n4498, A2 => n4499, A3 => n4500, A4 => 
                           n4501, ZN => n4497);
   U1882 : OAI21_X1 port map( B1 => n4496, B2 => n4497, A => n6386, ZN => n4495
                           );
   U1881 : OAI211_X1 port map( C1 => n555, C2 => n4194, A => n4494, B => n4495,
                           ZN => n4490);
   U1880 : AOI22_X1 port map( A1 => net644825, A2 => n6389, B1 => n6388, B2 => 
                           n4136, ZN => n4492);
   U1879 : OAI21_X1 port map( B1 => n617, B2 => n4189, A => n4492, ZN => n4491)
                           ;
   U1878 : AOI211_X1 port map( C1 => net644730, C2 => n4186, A => n4490, B => 
                           n4491, ZN => n4489);
   U1877 : NAND4_X1 port map( A1 => n4486, A2 => n4487, A3 => n4488, A4 => 
                           n4489, ZN => n2772);
   U1795 : AOI22_X1 port map( A1 => n4241, A2 => n4041, B1 => n6375, B2 => 
                           n3944, ZN => n4366);
   U1794 : AOI22_X1 port map( A1 => net644895, A2 => n6378, B1 => net644861, B2
                           => n6377, ZN => n4367);
   U1793 : AOI22_X1 port map( A1 => net644477, A2 => n6380, B1 => DATAIN(26), 
                           B2 => n6379, ZN => n4392);
   U1792 : OAI21_X1 port map( B1 => n4235, B2 => net644413, A => n4392, ZN => 
                           n4390);
   U1791 : OAI22_X1 port map( A1 => n645, A2 => n4233, B1 => n520, B2 => n4234,
                           ZN => n4391);
   U1790 : AOI211_X1 port map( C1 => net644669, C2 => n6381, A => n4390, B => 
                           n4391, ZN => n4368);
   U1789 : AOI22_X1 port map( A1 => net644573, A2 => n6382, B1 => net644541, B2
                           => n3880, ZN => n4374);
   U1788 : AOI22_X1 port map( A1 => n402, A2 => n6383, B1 => n3896, B2 => n4149
                           , ZN => n4384);
   U1787 : AOI22_X1 port map( A1 => net644638, A2 => n3895, B1 => net644509, B2
                           => n3894, ZN => n4385);
   U1786 : AOI22_X1 port map( A1 => n4220, A2 => n358, B1 => n4221, B2 => n4042
                           , ZN => n4386);
   U1785 : AOI22_X1 port map( A1 => net644606, A2 => n3890, B1 => net644702, B2
                           => n3897, ZN => n4387);
   U1784 : NAND4_X1 port map( A1 => n4384, A2 => n4385, A3 => n4386, A4 => 
                           n4387, ZN => n4376);
   U1783 : AOI22_X1 port map( A1 => n404, A2 => n4211, B1 => n4212, B2 => n4150
                           , ZN => n4378);
   U1782 : AOI22_X1 port map( A1 => net644798, A2 => n3902, B1 => net644766, B2
                           => n3901, ZN => n4379);
   U1781 : AOI22_X1 port map( A1 => net644928, A2 => n3900, B1 => net644445, B2
                           => n3899, ZN => n4380);
   U1780 : AOI22_X1 port map( A1 => n4204, A2 => n403, B1 => n3898, B2 => n4043
                           , ZN => n4381);
   U1779 : NAND4_X1 port map( A1 => n4378, A2 => n4379, A3 => n4380, A4 => 
                           n4381, ZN => n4377);
   U1778 : OAI21_X1 port map( B1 => n4376, B2 => n4377, A => n6386, ZN => n4375
                           );
   U1777 : OAI211_X1 port map( C1 => n551, C2 => n4194, A => n4374, B => n4375,
                           ZN => n4370);
   U1776 : AOI22_X1 port map( A1 => net644829, A2 => n6389, B1 => n4192, B2 => 
                           n4151, ZN => n4372);
   U1775 : OAI21_X1 port map( B1 => n613, B2 => n4189, A => n4372, ZN => n4371)
                           ;
   U1774 : AOI211_X1 port map( C1 => net644734, C2 => n6390, A => n4370, B => 
                           n4371, ZN => n4369);
   U1773 : NAND4_X1 port map( A1 => n4366, A2 => n4367, A3 => n4368, A4 => 
                           n4369, ZN => n2780);
   U3467 : AOI22_X1 port map( A1 => n6356, A2 => n3916, B1 => n6355, B2 => 
                           n3954, ZN => n5903);
   U3466 : AOI22_X1 port map( A1 => n6358, A2 => net644870, B1 => n5262, B2 => 
                           net644836, ZN => n5904);
   U3465 : AOI22_X1 port map( A1 => n6360, A2 => net644452, B1 => n6359, B2 => 
                           DATAIN(1), ZN => n5926);
   U3464 : OAI21_X1 port map( B1 => n5257, B2 => net644357, A => n5926, ZN => 
                           n5923);
   U3462 : OAI22_X1 port map( A1 => n545, A2 => n5255, B1 => n670, B2 => n5256,
                           ZN => n5924);
   U3461 : AOI211_X1 port map( C1 => n6361, C2 => net644644, A => n5923, B => 
                           n5924, ZN => n5905);
   U3460 : AOI22_X1 port map( A1 => n6363, A2 => net644516, B1 => n6362, B2 => 
                           net644548, ZN => n5911);
   U3459 : AOI22_X1 port map( A1 => n5248, A2 => n477, B1 => n6364, B2 => n222,
                           ZN => n5919);
   U3458 : AOI22_X1 port map( A1 => n3911, A2 => net644613, B1 => n3912, B2 => 
                           net644484, ZN => n5920);
   U3456 : AOI22_X1 port map( A1 => n5244, A2 => n3955, B1 => n6366, B2 => n383
                           , ZN => n5921);
   U3455 : AOI22_X1 port map( A1 => n3913, A2 => net644581, B1 => n3914, B2 => 
                           net644677, ZN => n5922);
   U3454 : NAND4_X1 port map( A1 => n5919, A2 => n5920, A3 => n5921, A4 => 
                           n5922, ZN => n5913);
   U3452 : AOI22_X1 port map( A1 => n5236, A2 => n479, B1 => n6368, B2 => n4063
                           , ZN => n5915);
   U3451 : AOI22_X1 port map( A1 => n3910, A2 => net644773, B1 => n3909, B2 => 
                           net644741, ZN => n5916);
   U3450 : AOI22_X1 port map( A1 => n3908, A2 => net644903, B1 => n3907, B2 => 
                           net644420, ZN => n5917);
   U3448 : AOI22_X1 port map( A1 => n3906, A2 => n3956, B1 => n3905, B2 => n478
                           , ZN => n5918);
   U3447 : NAND4_X1 port map( A1 => n5915, A2 => n5916, A3 => n5917, A4 => 
                           n5918, ZN => n5914);
   U3446 : OAI21_X1 port map( B1 => n5913, B2 => n5914, A => n6370, ZN => n5912
                           );
   U3445 : OAI211_X1 port map( C1 => n576, C2 => n5220, A => n5911, B => n5912,
                           ZN => n5907);
   U3442 : AOI22_X1 port map( A1 => n6373, A2 => net644804, B1 => n5219, B2 => 
                           n4064, ZN => n5909);
   U3441 : OAI21_X1 port map( B1 => n638, B2 => n5216, A => n5909, ZN => n5908)
                           ;
   U3440 : AOI211_X1 port map( C1 => n6374, C2 => net644709, A => n5907, B => 
                           n5908, ZN => n5906);
   U3439 : NAND4_X1 port map( A1 => n5903, A2 => n5904, A3 => n5905, A4 => 
                           n5906, ZN => n2697);
   U3286 : AOI22_X1 port map( A1 => n6356, A2 => n3922, B1 => n6355, B2 => 
                           n3975, ZN => n5771);
   U3285 : AOI22_X1 port map( A1 => n6358, A2 => net644876, B1 => n6357, B2 => 
                           net644842, ZN => n5772);
   U3284 : AOI22_X1 port map( A1 => n6360, A2 => net644458, B1 => n6359, B2 => 
                           DATAIN(7), ZN => n5792);
   U3283 : OAI21_X1 port map( B1 => n5257, B2 => net644363, A => n5792, ZN => 
                           n5790);
   U3282 : OAI22_X1 port map( A1 => n539, A2 => n5255, B1 => n664, B2 => n5256,
                           ZN => n5791);
   U3281 : AOI211_X1 port map( C1 => n6361, C2 => net644650, A => n5790, B => 
                           n5791, ZN => n5773);
   U3280 : AOI22_X1 port map( A1 => n6363, A2 => net644522, B1 => n6362, B2 => 
                           net644554, ZN => n5778);
   U3278 : AOI22_X1 port map( A1 => n5248, A2 => n459, B1 => n6364, B2 => n4084
                           , ZN => n5786);
   U3277 : AOI22_X1 port map( A1 => n3911, A2 => net644619, B1 => n3912, B2 => 
                           net644490, ZN => n5787);
   U3275 : AOI22_X1 port map( A1 => n5244, A2 => n3976, B1 => n6366, B2 => n377
                           , ZN => n5788);
   U3274 : AOI22_X1 port map( A1 => n3913, A2 => net644587, B1 => n3914, B2 => 
                           net644683, ZN => n5789);
   U3273 : NAND4_X1 port map( A1 => n5786, A2 => n5787, A3 => n5788, A4 => 
                           n5789, ZN => n5780);
   U3271 : AOI22_X1 port map( A1 => n5236, A2 => n461, B1 => n6368, B2 => n4085
                           , ZN => n5782);
   U3270 : AOI22_X1 port map( A1 => n3910, A2 => net644779, B1 => n3909, B2 => 
                           net644747, ZN => n5783);
   U3269 : AOI22_X1 port map( A1 => n3908, A2 => net644909, B1 => n3907, B2 => 
                           net644426, ZN => n5784);
   U3267 : AOI22_X1 port map( A1 => n3906, A2 => n3977, B1 => n3905, B2 => n460
                           , ZN => n5785);
   U3266 : NAND4_X1 port map( A1 => n5782, A2 => n5783, A3 => n5784, A4 => 
                           n5785, ZN => n5781);
   U3265 : OAI21_X1 port map( B1 => n5780, B2 => n5781, A => n6370, ZN => n5779
                           );
   U3264 : OAI211_X1 port map( C1 => n570, C2 => n5220, A => n5778, B => n5779,
                           ZN => n5775);
   U3262 : AOI22_X1 port map( A1 => n6373, A2 => net644810, B1 => n5219, B2 => 
                           n4086, ZN => n5777);
   U3261 : OAI21_X1 port map( B1 => n632, B2 => n5216, A => n5777, ZN => n5776)
                           ;
   U3260 : AOI211_X1 port map( C1 => n6374, C2 => net644715, A => n5775, B => 
                           n5776, ZN => n5774);
   U3259 : NAND4_X1 port map( A1 => n5771, A2 => n5772, A3 => n5773, A4 => 
                           n5774, ZN => n2703);
   U3346 : AOI22_X1 port map( A1 => n6356, A2 => n3920, B1 => n6355, B2 => 
                           n3969, ZN => n5815);
   U3345 : AOI22_X1 port map( A1 => n6358, A2 => net644874, B1 => n5262, B2 => 
                           net644840, ZN => n5816);
   U3344 : AOI22_X1 port map( A1 => n6360, A2 => net644456, B1 => n6359, B2 => 
                           DATAIN(5), ZN => n5836);
   U3343 : OAI21_X1 port map( B1 => n5257, B2 => net644361, A => n5836, ZN => 
                           n5834);
   U3342 : OAI22_X1 port map( A1 => n541, A2 => n5255, B1 => n666, B2 => n5256,
                           ZN => n5835);
   U3341 : AOI211_X1 port map( C1 => n6361, C2 => net644648, A => n5834, B => 
                           n5835, ZN => n5817);
   U3340 : AOI22_X1 port map( A1 => n6363, A2 => net644520, B1 => n6362, B2 => 
                           net644552, ZN => n5822);
   U3338 : AOI22_X1 port map( A1 => n5248, A2 => n465, B1 => n6364, B2 => n4078
                           , ZN => n5830);
   U3337 : AOI22_X1 port map( A1 => n3911, A2 => net644617, B1 => n3912, B2 => 
                           net644488, ZN => n5831);
   U3335 : AOI22_X1 port map( A1 => n5244, A2 => n3970, B1 => n6366, B2 => n379
                           , ZN => n5832);
   U3334 : AOI22_X1 port map( A1 => n3913, A2 => net644585, B1 => n3914, B2 => 
                           net644681, ZN => n5833);
   U3333 : NAND4_X1 port map( A1 => n5830, A2 => n5831, A3 => n5832, A4 => 
                           n5833, ZN => n5824);
   U3331 : AOI22_X1 port map( A1 => n5236, A2 => n467, B1 => n6368, B2 => n4079
                           , ZN => n5826);
   U3330 : AOI22_X1 port map( A1 => n3910, A2 => net644777, B1 => n3909, B2 => 
                           net644745, ZN => n5827);
   U3329 : AOI22_X1 port map( A1 => n3908, A2 => net644907, B1 => n3907, B2 => 
                           net644424, ZN => n5828);
   U3327 : AOI22_X1 port map( A1 => n3906, A2 => n3971, B1 => n3905, B2 => n466
                           , ZN => n5829);
   U3326 : NAND4_X1 port map( A1 => n5826, A2 => n5827, A3 => n5828, A4 => 
                           n5829, ZN => n5825);
   U3325 : OAI21_X1 port map( B1 => n5824, B2 => n5825, A => n6370, ZN => n5823
                           );
   U3324 : OAI211_X1 port map( C1 => n572, C2 => n5220, A => n5822, B => n5823,
                           ZN => n5819);
   U3322 : AOI22_X1 port map( A1 => n6373, A2 => net644808, B1 => n5219, B2 => 
                           n4080, ZN => n5821);
   U3321 : OAI21_X1 port map( B1 => n634, B2 => n5216, A => n5821, ZN => n5820)
                           ;
   U3320 : AOI211_X1 port map( C1 => n6374, C2 => net644713, A => n5819, B => 
                           n5820, ZN => n5818);
   U3319 : NAND4_X1 port map( A1 => n5815, A2 => n5816, A3 => n5817, A4 => 
                           n5818, ZN => n2701);
   U3376 : AOI22_X1 port map( A1 => n6356, A2 => n3919, B1 => n6355, B2 => 
                           n3966, ZN => n5837);
   U3375 : AOI22_X1 port map( A1 => n6358, A2 => net644873, B1 => n5262, B2 => 
                           net644839, ZN => n5838);
   U3374 : AOI22_X1 port map( A1 => n6360, A2 => net644455, B1 => n6359, B2 => 
                           DATAIN(4), ZN => n5858);
   U3373 : OAI21_X1 port map( B1 => n5257, B2 => net644360, A => n5858, ZN => 
                           n5856);
   U3372 : OAI22_X1 port map( A1 => n542, A2 => n5255, B1 => n667, B2 => n5256,
                           ZN => n5857);
   U3371 : AOI211_X1 port map( C1 => n6361, C2 => net644647, A => n5856, B => 
                           n5857, ZN => n5839);
   U3370 : AOI22_X1 port map( A1 => n6363, A2 => net644519, B1 => n6362, B2 => 
                           net644551, ZN => n5844);
   U3368 : AOI22_X1 port map( A1 => n5248, A2 => n468, B1 => n6364, B2 => n4075
                           , ZN => n5852);
   U3367 : AOI22_X1 port map( A1 => n3911, A2 => net644616, B1 => n3912, B2 => 
                           net644487, ZN => n5853);
   U3365 : AOI22_X1 port map( A1 => n5244, A2 => n3967, B1 => n6366, B2 => n380
                           , ZN => n5854);
   U3364 : AOI22_X1 port map( A1 => n3913, A2 => net644584, B1 => n3914, B2 => 
                           net644680, ZN => n5855);
   U3363 : NAND4_X1 port map( A1 => n5852, A2 => n5853, A3 => n5854, A4 => 
                           n5855, ZN => n5846);
   U3361 : AOI22_X1 port map( A1 => n5236, A2 => n470, B1 => n6368, B2 => n4076
                           , ZN => n5848);
   U3360 : AOI22_X1 port map( A1 => n3910, A2 => net644776, B1 => n3909, B2 => 
                           net644744, ZN => n5849);
   U3359 : AOI22_X1 port map( A1 => n3908, A2 => net644906, B1 => n3907, B2 => 
                           net644423, ZN => n5850);
   U3357 : AOI22_X1 port map( A1 => n3906, A2 => n3968, B1 => n3905, B2 => n469
                           , ZN => n5851);
   U3356 : NAND4_X1 port map( A1 => n5848, A2 => n5849, A3 => n5850, A4 => 
                           n5851, ZN => n5847);
   U3355 : OAI21_X1 port map( B1 => n5846, B2 => n5847, A => n6370, ZN => n5845
                           );
   U3354 : OAI211_X1 port map( C1 => n573, C2 => n5220, A => n5844, B => n5845,
                           ZN => n5841);
   U3352 : AOI22_X1 port map( A1 => n6373, A2 => net644807, B1 => n5219, B2 => 
                           n4077, ZN => n5843);
   U3351 : OAI21_X1 port map( B1 => n635, B2 => n5216, A => n5843, ZN => n5842)
                           ;
   U3350 : AOI211_X1 port map( C1 => n6374, C2 => net644712, A => n5841, B => 
                           n5842, ZN => n5840);
   U3349 : NAND4_X1 port map( A1 => n5837, A2 => n5838, A3 => n5839, A4 => 
                           n5840, ZN => n2700);
   U2716 : AOI22_X1 port map( A1 => n6356, A2 => n3944, B1 => n5264, B2 => 
                           n4041, ZN => n5353);
   U2715 : AOI22_X1 port map( A1 => n6358, A2 => net644895, B1 => n5262, B2 => 
                           net644861, ZN => n5354);
   U2714 : AOI22_X1 port map( A1 => n5259, A2 => net644477, B1 => n5260, B2 => 
                           DATAIN(26), ZN => n5374);
   U2713 : OAI21_X1 port map( B1 => n5257, B2 => net644382, A => n5374, ZN => 
                           n5372);
   U2712 : OAI22_X1 port map( A1 => n520, A2 => n5255, B1 => n645, B2 => n5256,
                           ZN => n5373);
   U2711 : AOI211_X1 port map( C1 => n6361, C2 => net644669, A => n5372, B => 
                           n5373, ZN => n5355);
   U2710 : AOI22_X1 port map( A1 => n5250, A2 => net644541, B1 => n5251, B2 => 
                           net644573, ZN => n5360);
   U2708 : AOI22_X1 port map( A1 => n5248, A2 => n402, B1 => n5249, B2 => n4149
                           , ZN => n5368);
   U2707 : AOI22_X1 port map( A1 => n5246, A2 => net644638, B1 => n5247, B2 => 
                           net644509, ZN => n5369);
   U2705 : AOI22_X1 port map( A1 => n5244, A2 => n4042, B1 => n5245, B2 => n358
                           , ZN => n5370);
   U2704 : AOI22_X1 port map( A1 => n5242, A2 => net644606, B1 => n5243, B2 => 
                           net644702, ZN => n5371);
   U2703 : NAND4_X1 port map( A1 => n5368, A2 => n5369, A3 => n5370, A4 => 
                           n5371, ZN => n5362);
   U2701 : AOI22_X1 port map( A1 => n5236, A2 => n404, B1 => n5237, B2 => n4150
                           , ZN => n5364);
   U2700 : AOI22_X1 port map( A1 => n5234, A2 => net644798, B1 => n5235, B2 => 
                           net644766, ZN => n5365);
   U2699 : AOI22_X1 port map( A1 => n5232, A2 => net644928, B1 => n5233, B2 => 
                           net644445, ZN => n5366);
   U2697 : AOI22_X1 port map( A1 => n5230, A2 => n4043, B1 => n5231, B2 => n403
                           , ZN => n5367);
   U2696 : NAND4_X1 port map( A1 => n5364, A2 => n5365, A3 => n5366, A4 => 
                           n5367, ZN => n5363);
   U2695 : OAI21_X1 port map( B1 => n5362, B2 => n5363, A => n6370, ZN => n5361
                           );
   U2694 : OAI211_X1 port map( C1 => n551, C2 => n5220, A => n5360, B => n5361,
                           ZN => n5357);
   U2692 : AOI22_X1 port map( A1 => n6373, A2 => net644829, B1 => n5219, B2 => 
                           n4151, ZN => n5359);
   U2691 : OAI21_X1 port map( B1 => n613, B2 => n5216, A => n5359, ZN => n5358)
                           ;
   U2690 : AOI211_X1 port map( C1 => n5213, C2 => net644734, A => n5357, B => 
                           n5358, ZN => n5356);
   U2689 : NAND4_X1 port map( A1 => n5353, A2 => n5354, A3 => n5355, A4 => 
                           n5356, ZN => n2722);
   U496 : OAI22_X1 port map( A1 => n5063, A2 => n6431, B1 => n1688, B2 => n6430
                           , ZN => n3451);
   U484 : OAI22_X1 port map( A1 => n5084, A2 => n1885, B1 => n1676, B2 => n6430
                           , ZN => n3457);
   U431 : OAI22_X1 port map( A1 => n5252, A2 => n6433, B1 => n1688, B2 => n6432
                           , ZN => n3483);
   U518 : OAI22_X1 port map( A1 => n5023, A2 => n6431, B1 => n1710, B2 => n6430
                           , ZN => n3440);
   U478 : OAI22_X1 port map( A1 => n5102, A2 => n1885, B1 => n1670, B2 => n6430
                           , ZN => n3460);
   U453 : OAI22_X1 port map( A1 => n5144, A2 => n6433, B1 => n1710, B2 => n6432
                           , ZN => n3472);
   U498 : OAI22_X1 port map( A1 => n5055, A2 => n6431, B1 => n1690, B2 => n6430
                           , ZN => n3450);
   U502 : OAI22_X1 port map( A1 => n5053, A2 => n6431, B1 => n1694, B2 => n6430
                           , ZN => n3448);
   U486 : OAI22_X1 port map( A1 => n5083, A2 => n1885, B1 => n1678, B2 => n6430
                           , ZN => n3456);
   U506 : OAI22_X1 port map( A1 => n5048, A2 => n6431, B1 => n1698, B2 => n6430
                           , ZN => n3446);
   U445 : OAI22_X1 port map( A1 => n5180, A2 => n6433, B1 => n1702, B2 => n6432
                           , ZN => n3476);
   U516 : OAI22_X1 port map( A1 => n5024, A2 => n6431, B1 => n1708, B2 => n6430
                           , ZN => n3441);
   U441 : OAI22_X1 port map( A1 => n5188, A2 => n6433, B1 => n1698, B2 => n6432
                           , ZN => n3478);
   U451 : OAI22_X1 port map( A1 => n5145, A2 => n6433, B1 => n1708, B2 => n6432
                           , ZN => n3473);
   U439 : OAI22_X1 port map( A1 => n5193, A2 => n6433, B1 => n1696, B2 => n6432
                           , ZN => n3479);
   U500 : OAI22_X1 port map( A1 => n5054, A2 => n6431, B1 => n1692, B2 => n6430
                           , ZN => n3449);
   U512 : OAI22_X1 port map( A1 => n5033, A2 => n6431, B1 => n1704, B2 => n6430
                           , ZN => n3443);
   U474 : OAI22_X1 port map( A1 => n5108, A2 => n6431, B1 => n1666, B2 => n6430
                           , ZN => n3462);
   U443 : OAI22_X1 port map( A1 => n5183, A2 => n6433, B1 => n1700, B2 => n6432
                           , ZN => n3477);
   U476 : OAI22_X1 port map( A1 => n5103, A2 => n1885, B1 => n1668, B2 => n6430
                           , ZN => n3461);
   U504 : OAI22_X1 port map( A1 => n5049, A2 => n6431, B1 => n1696, B2 => n6430
                           , ZN => n3447);
   U435 : OAI22_X1 port map( A1 => n5204, A2 => n6433, B1 => n1692, B2 => n6432
                           , ZN => n3481);
   U514 : OAI22_X1 port map( A1 => n5025, A2 => n6431, B1 => n1706, B2 => n6430
                           , ZN => n3442);
   U411 : OAI22_X1 port map( A1 => n5991, A2 => n1852, B1 => n1668, B2 => n6432
                           , ZN => n3493);
   U510 : OAI22_X1 port map( A1 => n5042, A2 => n6431, B1 => n1702, B2 => n6430
                           , ZN => n3444);
   U508 : OAI22_X1 port map( A1 => n5043, A2 => n6431, B1 => n1700, B2 => n6430
                           , ZN => n3445);
   U413 : OAI22_X1 port map( A1 => n5990, A2 => n1852, B1 => n1670, B2 => n6432
                           , ZN => n3492);
   U421 : OAI22_X1 port map( A1 => n5986, A2 => n1852, B1 => n1678, B2 => n6432
                           , ZN => n3488);
   U449 : OAI22_X1 port map( A1 => n5153, A2 => n6433, B1 => n1706, B2 => n6432
                           , ZN => n3474);
   U447 : OAI22_X1 port map( A1 => n5174, A2 => n6433, B1 => n1704, B2 => n6432
                           , ZN => n3475);
   U437 : OAI22_X1 port map( A1 => n5203, A2 => n6433, B1 => n1694, B2 => n6432
                           , ZN => n3480);
   U433 : OAI22_X1 port map( A1 => n5218, A2 => n6433, B1 => n1690, B2 => n6432
                           , ZN => n3482);
   U409 : OAI22_X1 port map( A1 => n5992, A2 => n6433, B1 => n1666, B2 => n6432
                           , ZN => n3494);
   U419 : OAI22_X1 port map( A1 => n5987, A2 => n1852, B1 => n1676, B2 => n6432
                           , ZN => n3489);
   U469 : OAI22_X1 port map( A1 => n2601, A2 => n6433, B1 => n6432, B2 => n1726
                           , ZN => n3464);
   U534 : OAI22_X1 port map( A1 => n481, A2 => n6431, B1 => n6430, B2 => n1726,
                           ZN => n3432);
   U1444 : OAI22_X1 port map( A1 => n6223, A2 => n6400, B1 => n1702, B2 => 
                           n6399, ZN => n2900);
   U1436 : OAI22_X1 port map( A1 => n6227, A2 => n6400, B1 => n1694, B2 => 
                           n6399, ZN => n2904);
   U1456 : OAI22_X1 port map( A1 => n6217, A2 => n6400, B1 => n1714, B2 => 
                           n6399, ZN => n2894);
   U1438 : OAI22_X1 port map( A1 => n6226, A2 => n6400, B1 => n1696, B2 => 
                           n6399, ZN => n2903);
   U1440 : OAI22_X1 port map( A1 => n6225, A2 => n6400, B1 => n1698, B2 => 
                           n6399, ZN => n2902);
   U1466 : OAI22_X1 port map( A1 => n6212, A2 => n6400, B1 => n1724, B2 => 
                           n6399, ZN => n2889);
   U1452 : OAI22_X1 port map( A1 => n6219, A2 => n6400, B1 => n1710, B2 => 
                           n6399, ZN => n2896);
   U1442 : OAI22_X1 port map( A1 => n6224, A2 => n6400, B1 => n1700, B2 => 
                           n6399, ZN => n2901);
   U1364 : OAI22_X1 port map( A1 => n6150, A2 => n6403, B1 => n1724, B2 => 
                           n6402, ZN => n2953);
   U1362 : OAI22_X1 port map( A1 => n6151, A2 => n6403, B1 => n1722, B2 => 
                           n6402, ZN => n2954);
   U1360 : OAI22_X1 port map( A1 => n6152, A2 => n6403, B1 => n1720, B2 => 
                           n6402, ZN => n2955);
   U1354 : OAI22_X1 port map( A1 => n6155, A2 => n6403, B1 => n1714, B2 => 
                           n6402, ZN => n2958);
   U1352 : OAI22_X1 port map( A1 => n6156, A2 => n6403, B1 => n1712, B2 => 
                           n6402, ZN => n2959);
   U1350 : OAI22_X1 port map( A1 => n6157, A2 => n6403, B1 => n1710, B2 => 
                           n6402, ZN => n2960);
   U1430 : OAI22_X1 port map( A1 => n6230, A2 => n6400, B1 => n1688, B2 => 
                           n6399, ZN => n2907);
   U1454 : OAI22_X1 port map( A1 => n6218, A2 => n6400, B1 => n1712, B2 => 
                           n6399, ZN => n2895);
   U1434 : OAI22_X1 port map( A1 => n6228, A2 => n6400, B1 => n1692, B2 => 
                           n6399, ZN => n2905);
   U1432 : OAI22_X1 port map( A1 => n6229, A2 => n6400, B1 => n1690, B2 => 
                           n6399, ZN => n2906);
   U1462 : OAI22_X1 port map( A1 => n6214, A2 => n6400, B1 => n1720, B2 => 
                           n6399, ZN => n2891);
   U1428 : OAI22_X1 port map( A1 => n6231, A2 => n6400, B1 => n1686, B2 => 
                           n6399, ZN => n2908);
   U1426 : OAI22_X1 port map( A1 => n6232, A2 => n6400, B1 => n1684, B2 => 
                           n6399, ZN => n2909);
   U1424 : OAI22_X1 port map( A1 => n6233, A2 => n6400, B1 => n1682, B2 => 
                           n6399, ZN => n2910);
   U1422 : OAI22_X1 port map( A1 => n6234, A2 => n4073, B1 => n1680, B2 => 
                           n6399, ZN => n2911);
   U1342 : OAI22_X1 port map( A1 => n6161, A2 => n6403, B1 => n1702, B2 => 
                           n6402, ZN => n2964);
   U1464 : OAI22_X1 port map( A1 => n6213, A2 => n6400, B1 => n1722, B2 => 
                           n6399, ZN => n2890);
   U1320 : OAI22_X1 port map( A1 => n6172, A2 => n4035, B1 => n1680, B2 => 
                           n6402, ZN => n2975);
   U1340 : OAI22_X1 port map( A1 => n6162, A2 => n6403, B1 => n1700, B2 => 
                           n6402, ZN => n2965);
   U1322 : OAI22_X1 port map( A1 => n6171, A2 => n6403, B1 => n1682, B2 => 
                           n6402, ZN => n2974);
   U1338 : OAI22_X1 port map( A1 => n6163, A2 => n6403, B1 => n1698, B2 => 
                           n6402, ZN => n2966);
   U1324 : OAI22_X1 port map( A1 => n6170, A2 => n6403, B1 => n1684, B2 => 
                           n6402, ZN => n2973);
   U1326 : OAI22_X1 port map( A1 => n6169, A2 => n6403, B1 => n1686, B2 => 
                           n6402, ZN => n2972);
   U1328 : OAI22_X1 port map( A1 => n6168, A2 => n6403, B1 => n1688, B2 => 
                           n6402, ZN => n2971);
   U1330 : OAI22_X1 port map( A1 => n6167, A2 => n6403, B1 => n1690, B2 => 
                           n6402, ZN => n2970);
   U1332 : OAI22_X1 port map( A1 => n6166, A2 => n6403, B1 => n1692, B2 => 
                           n6402, ZN => n2969);
   U1334 : OAI22_X1 port map( A1 => n6165, A2 => n6403, B1 => n1694, B2 => 
                           n6402, ZN => n2968);
   U1336 : OAI22_X1 port map( A1 => n6164, A2 => n6403, B1 => n1696, B2 => 
                           n6402, ZN => n2967);
   U1256 : OAI22_X1 port map( A1 => n6140, A2 => n6405, B1 => n1682, B2 => 
                           n6404, ZN => n3006);
   U1274 : OAI22_X1 port map( A1 => n6131, A2 => n6405, B1 => n1700, B2 => 
                           n6404, ZN => n2997);
   U1272 : OAI22_X1 port map( A1 => n6132, A2 => n6405, B1 => n1698, B2 => 
                           n6404, ZN => n2998);
   U1270 : OAI22_X1 port map( A1 => n6133, A2 => n6405, B1 => n1696, B2 => 
                           n6404, ZN => n2999);
   U1268 : OAI22_X1 port map( A1 => n6134, A2 => n6405, B1 => n1694, B2 => 
                           n6404, ZN => n3000);
   U1300 : OAI22_X1 port map( A1 => n6349, A2 => n6405, B1 => n1726, B2 => 
                           n6404, ZN => n2984);
   U1266 : OAI22_X1 port map( A1 => n6135, A2 => n6405, B1 => n1692, B2 => 
                           n6404, ZN => n3001);
   U1296 : OAI22_X1 port map( A1 => n6120, A2 => n6405, B1 => n1722, B2 => 
                           n6404, ZN => n2986);
   U1262 : OAI22_X1 port map( A1 => n6137, A2 => n6405, B1 => n1688, B2 => 
                           n6404, ZN => n3003);
   U1294 : OAI22_X1 port map( A1 => n6121, A2 => n6405, B1 => n1720, B2 => 
                           n6404, ZN => n2987);
   U1258 : OAI22_X1 port map( A1 => n6139, A2 => n6405, B1 => n1684, B2 => 
                           n6404, ZN => n3005);
   U1254 : OAI22_X1 port map( A1 => n6141, A2 => n4000, B1 => n1680, B2 => 
                           n6404, ZN => n3007);
   U1260 : OAI22_X1 port map( A1 => n6138, A2 => n6405, B1 => n1686, B2 => 
                           n6404, ZN => n3004);
   U1288 : OAI22_X1 port map( A1 => n6124, A2 => n6405, B1 => n1714, B2 => 
                           n6404, ZN => n2990);
   U1284 : OAI22_X1 port map( A1 => n6126, A2 => n6405, B1 => n1710, B2 => 
                           n6404, ZN => n2992);
   U1286 : OAI22_X1 port map( A1 => n6125, A2 => n6405, B1 => n1712, B2 => 
                           n6404, ZN => n2991);
   U1276 : OAI22_X1 port map( A1 => n6130, A2 => n6405, B1 => n1702, B2 => 
                           n6404, ZN => n2996);
   U1264 : OAI22_X1 port map( A1 => n6136, A2 => n6405, B1 => n1690, B2 => 
                           n6404, ZN => n3002);
   U308 : OAI22_X1 port map( A1 => n6318, A2 => n6437, B1 => n1700, B2 => n6436
                           , ZN => n3573);
   U304 : OAI22_X1 port map( A1 => n6320, A2 => n6437, B1 => n1696, B2 => n6436
                           , ZN => n3575);
   U274 : OAI22_X1 port map( A1 => n6335, A2 => n6437, B1 => n1666, B2 => n6436
                           , ZN => n3590);
   U318 : OAI22_X1 port map( A1 => n6313, A2 => n6437, B1 => n1710, B2 => n6436
                           , ZN => n3568);
   U316 : OAI22_X1 port map( A1 => n6314, A2 => n6437, B1 => n1708, B2 => n6436
                           , ZN => n3569);
   U314 : OAI22_X1 port map( A1 => n6315, A2 => n6437, B1 => n1706, B2 => n6436
                           , ZN => n3570);
   U300 : OAI22_X1 port map( A1 => n6322, A2 => n6437, B1 => n1692, B2 => n6436
                           , ZN => n3577);
   U312 : OAI22_X1 port map( A1 => n6316, A2 => n6437, B1 => n1704, B2 => n6436
                           , ZN => n3571);
   U306 : OAI22_X1 port map( A1 => n6319, A2 => n6437, B1 => n1698, B2 => n6436
                           , ZN => n3574);
   U278 : OAI22_X1 port map( A1 => n6333, A2 => n1811, B1 => n1670, B2 => n6436
                           , ZN => n3588);
   U302 : OAI22_X1 port map( A1 => n6321, A2 => n6437, B1 => n1694, B2 => n6436
                           , ZN => n3576);
   U286 : OAI22_X1 port map( A1 => n6329, A2 => n1811, B1 => n1678, B2 => n6436
                           , ZN => n3584);
   U310 : OAI22_X1 port map( A1 => n6317, A2 => n6437, B1 => n1702, B2 => n6436
                           , ZN => n3572);
   U296 : OAI22_X1 port map( A1 => n6324, A2 => n6437, B1 => n1688, B2 => n6436
                           , ZN => n3579);
   U284 : OAI22_X1 port map( A1 => n6330, A2 => n1811, B1 => n1676, B2 => n6436
                           , ZN => n3585);
   U298 : OAI22_X1 port map( A1 => n6323, A2 => n6437, B1 => n1690, B2 => n6436
                           , ZN => n3578);
   U276 : OAI22_X1 port map( A1 => n6334, A2 => n1811, B1 => n1668, B2 => n6436
                           , ZN => n3589);
   U334 : OAI22_X1 port map( A1 => n480, A2 => n6437, B1 => n6436, B2 => n1726,
                           ZN => n3560);
   U169 : NAND2_X1 port map( A1 => n1769, A2 => n1770, ZN => n1729);
   U31 : OAI22_X1 port map( A1 => n6041, A2 => n6445, B1 => n1692, B2 => n6444,
                           ZN => n3737);
   U37 : OAI22_X1 port map( A1 => n6038, A2 => n6445, B1 => n1698, B2 => n6444,
                           ZN => n3734);
   U33 : OAI22_X1 port map( A1 => n6040, A2 => n6445, B1 => n1694, B2 => n6444,
                           ZN => n3736);
   U63 : OAI22_X1 port map( A1 => n6025, A2 => n6445, B1 => n1724, B2 => n6444,
                           ZN => n3721);
   U25 : OAI22_X1 port map( A1 => n6044, A2 => n6445, B1 => n1686, B2 => n6444,
                           ZN => n3740);
   U61 : OAI22_X1 port map( A1 => n6026, A2 => n6445, B1 => n1722, B2 => n6444,
                           ZN => n3722);
   U21 : OAI22_X1 port map( A1 => n6046, A2 => n6445, B1 => n1682, B2 => n6444,
                           ZN => n3742);
   U35 : OAI22_X1 port map( A1 => n6039, A2 => n6445, B1 => n1696, B2 => n6444,
                           ZN => n3735);
   U23 : OAI22_X1 port map( A1 => n6045, A2 => n6445, B1 => n1684, B2 => n6444,
                           ZN => n3741);
   U27 : OAI22_X1 port map( A1 => n6043, A2 => n6445, B1 => n1688, B2 => n6444,
                           ZN => n3739);
   U49 : OAI22_X1 port map( A1 => n6032, A2 => n6445, B1 => n1710, B2 => n6444,
                           ZN => n3728);
   U41 : OAI22_X1 port map( A1 => n6036, A2 => n6445, B1 => n1702, B2 => n6444,
                           ZN => n3732);
   U29 : OAI22_X1 port map( A1 => n6042, A2 => n6445, B1 => n1690, B2 => n6444,
                           ZN => n3738);
   U39 : OAI22_X1 port map( A1 => n6037, A2 => n6445, B1 => n1700, B2 => n6444,
                           ZN => n3733);
   U53 : OAI22_X1 port map( A1 => n6030, A2 => n6445, B1 => n1714, B2 => n6444,
                           ZN => n3726);
   U59 : OAI22_X1 port map( A1 => n6027, A2 => n6445, B1 => n1720, B2 => n6444,
                           ZN => n3723);
   U19 : OAI22_X1 port map( A1 => n6047, A2 => n1662, B1 => n1680, B2 => n6444,
                           ZN => n3743);
   U51 : OAI22_X1 port map( A1 => n6031, A2 => n6445, B1 => n1712, B2 => n6444,
                           ZN => n3727);
   U565 : OAI22_X1 port map( A1 => n510, A2 => n6429, B1 => n6428, B2 => n1720,
                           ZN => n3403);
   U552 : OAI22_X1 port map( A1 => n497, A2 => n6429, B1 => n6428, B2 => n1694,
                           ZN => n3416);
   U557 : OAI22_X1 port map( A1 => n502, A2 => n6429, B1 => n6428, B2 => n1704,
                           ZN => n3411);
   U547 : OAI22_X1 port map( A1 => n492, A2 => n6429, B1 => n6428, B2 => n1684,
                           ZN => n3421);
   U549 : OAI22_X1 port map( A1 => n494, A2 => n6429, B1 => n6428, B2 => n1688,
                           ZN => n3419);
   U562 : OAI22_X1 port map( A1 => n507, A2 => n6429, B1 => n6428, B2 => n1714,
                           ZN => n3406);
   U554 : OAI22_X1 port map( A1 => n499, A2 => n6429, B1 => n6428, B2 => n1698,
                           ZN => n3414);
   U550 : OAI22_X1 port map( A1 => n495, A2 => n6429, B1 => n6428, B2 => n1690,
                           ZN => n3418);
   U553 : OAI22_X1 port map( A1 => n498, A2 => n6429, B1 => n6428, B2 => n1696,
                           ZN => n3415);
   U548 : OAI22_X1 port map( A1 => n493, A2 => n6429, B1 => n6428, B2 => n1686,
                           ZN => n3420);
   U545 : OAI22_X1 port map( A1 => n490, A2 => n1917, B1 => n6428, B2 => n1680,
                           ZN => n3423);
   U560 : OAI22_X1 port map( A1 => n505, A2 => n6429, B1 => n6428, B2 => n1710,
                           ZN => n3408);
   U561 : OAI22_X1 port map( A1 => n506, A2 => n6429, B1 => n6428, B2 => n1712,
                           ZN => n3407);
   U546 : OAI22_X1 port map( A1 => n491, A2 => n6429, B1 => n6428, B2 => n1682,
                           ZN => n3422);
   U555 : OAI22_X1 port map( A1 => n500, A2 => n6429, B1 => n6428, B2 => n1700,
                           ZN => n3413);
   U556 : OAI22_X1 port map( A1 => n501, A2 => n6429, B1 => n6428, B2 => n1702,
                           ZN => n3412);
   U566 : OAI22_X1 port map( A1 => n511, A2 => n6429, B1 => n6428, B2 => n1722,
                           ZN => n3402);
   U551 : OAI22_X1 port map( A1 => n496, A2 => n6429, B1 => n6428, B2 => n1692,
                           ZN => n3417);
   U195 : OAI22_X1 port map( A1 => n4364, A2 => n6440, B1 => n1688, B2 => n6439
                           , ZN => n3643);
   U199 : OAI22_X1 port map( A1 => n4359, A2 => n6440, B1 => n1692, B2 => n6439
                           , ZN => n3641);
   U227 : OAI22_X1 port map( A1 => n4304, A2 => n6440, B1 => n1720, B2 => n6439
                           , ZN => n3627);
   U191 : OAI22_X1 port map( A1 => n4373, A2 => n6440, B1 => n1684, B2 => n6439
                           , ZN => n3645);
   U193 : OAI22_X1 port map( A1 => n4365, A2 => n6440, B1 => n1686, B2 => n6439
                           , ZN => n3644);
   U201 : OAI22_X1 port map( A1 => n4358, A2 => n6440, B1 => n1694, B2 => n6439
                           , ZN => n3640);
   U221 : OAI22_X1 port map( A1 => n4322, A2 => n6440, B1 => n1714, B2 => n6439
                           , ZN => n3630);
   U203 : OAI22_X1 port map( A1 => n4353, A2 => n6440, B1 => n1696, B2 => n6439
                           , ZN => n3639);
   U197 : OAI22_X1 port map( A1 => n4363, A2 => n6440, B1 => n1690, B2 => n6439
                           , ZN => n3642);
   U205 : OAI22_X1 port map( A1 => n4352, A2 => n6440, B1 => n1698, B2 => n6439
                           , ZN => n3638);
   U219 : OAI22_X1 port map( A1 => n4323, A2 => n6440, B1 => n1712, B2 => n6439
                           , ZN => n3631);
   U217 : OAI22_X1 port map( A1 => n4328, A2 => n6440, B1 => n1710, B2 => n6439
                           , ZN => n3632);
   U189 : OAI22_X1 port map( A1 => n4382, A2 => n6440, B1 => n1682, B2 => n6439
                           , ZN => n3646);
   U233 : OAI22_X1 port map( A1 => n6353, A2 => n6440, B1 => n1726, B2 => n6439
                           , ZN => n3624);
   U209 : OAI22_X1 port map( A1 => n4335, A2 => n6440, B1 => n1702, B2 => n6439
                           , ZN => n3636);
   U187 : OAI22_X1 port map( A1 => n4383, A2 => n1772, B1 => n1680, B2 => n6439
                           , ZN => n3647);
   U207 : OAI22_X1 port map( A1 => n4343, A2 => n6440, B1 => n1700, B2 => n6439
                           , ZN => n3637);
   U229 : OAI22_X1 port map( A1 => n4303, A2 => n6440, B1 => n1722, B2 => n6439
                           , ZN => n3626);
   U1536 : OAI22_X1 port map( A1 => n4592, A2 => n6396, B1 => n1694, B2 => 
                           n6395, ZN => n2840);
   U1542 : OAI22_X1 port map( A1 => n4574, A2 => n6396, B1 => n1700, B2 => 
                           n6395, ZN => n2837);
   U1534 : OAI22_X1 port map( A1 => n4593, A2 => n6396, B1 => n1692, B2 => 
                           n6395, ZN => n2841);
   U1532 : OAI22_X1 port map( A1 => n4598, A2 => n6396, B1 => n1690, B2 => 
                           n6395, ZN => n2842);
   U1544 : OAI22_X1 port map( A1 => n4573, A2 => n6396, B1 => n1702, B2 => 
                           n6395, ZN => n2836);
   U1528 : OAI22_X1 port map( A1 => n4603, A2 => n6396, B1 => n1686, B2 => 
                           n6395, ZN => n2844);
   U1530 : OAI22_X1 port map( A1 => n4599, A2 => n6396, B1 => n1688, B2 => 
                           n6395, ZN => n2843);
   U1562 : OAI22_X1 port map( A1 => n4539, A2 => n6396, B1 => n1720, B2 => 
                           n6395, ZN => n2827);
   U1538 : OAI22_X1 port map( A1 => n4583, A2 => n6396, B1 => n1696, B2 => 
                           n6395, ZN => n2839);
   U1526 : OAI22_X1 port map( A1 => n4604, A2 => n6396, B1 => n1684, B2 => 
                           n6395, ZN => n2845);
   U1546 : OAI22_X1 port map( A1 => n4569, A2 => n6396, B1 => n1704, B2 => 
                           n6395, ZN => n2835);
   U1540 : OAI22_X1 port map( A1 => n4575, A2 => n6396, B1 => n1698, B2 => 
                           n6395, ZN => n2838);
   U1556 : OAI22_X1 port map( A1 => n4545, A2 => n6396, B1 => n1714, B2 => 
                           n6395, ZN => n2830);
   U1522 : OAI22_X1 port map( A1 => n4613, A2 => n4110, B1 => n1680, B2 => 
                           n6395, ZN => n2847);
   U1554 : OAI22_X1 port map( A1 => n4553, A2 => n6396, B1 => n1712, B2 => 
                           n6395, ZN => n2831);
   U1552 : OAI22_X1 port map( A1 => n4562, A2 => n6396, B1 => n1710, B2 => 
                           n6395, ZN => n2832);
   U1524 : OAI22_X1 port map( A1 => n4605, A2 => n6396, B1 => n1682, B2 => 
                           n6395, ZN => n2846);
   U1564 : OAI22_X1 port map( A1 => n4538, A2 => n6396, B1 => n1722, B2 => 
                           n6395, ZN => n2826);
   U1075 : OAI22_X1 port map( A1 => n4808, A2 => n6412, B1 => n1702, B2 => 
                           n6411, ZN => n3124);
   U1071 : OAI22_X1 port map( A1 => n4813, A2 => n6412, B1 => n1698, B2 => 
                           n6411, ZN => n3126);
   U1073 : OAI22_X1 port map( A1 => n4809, A2 => n6412, B1 => n1700, B2 => 
                           n6411, ZN => n3125);
   U1069 : OAI22_X1 port map( A1 => n4814, A2 => n6412, B1 => n1696, B2 => 
                           n6411, ZN => n3127);
   U1067 : OAI22_X1 port map( A1 => n4815, A2 => n6412, B1 => n1694, B2 => 
                           n6411, ZN => n3128);
   U1065 : OAI22_X1 port map( A1 => n4823, A2 => n6412, B1 => n1692, B2 => 
                           n6411, ZN => n3129);
   U1055 : OAI22_X1 port map( A1 => n4843, A2 => n6412, B1 => n1682, B2 => 
                           n6411, ZN => n3134);
   U1063 : OAI22_X1 port map( A1 => n4832, A2 => n6412, B1 => n1690, B2 => 
                           n6411, ZN => n3130);
   U1061 : OAI22_X1 port map( A1 => n4833, A2 => n6412, B1 => n1688, B2 => 
                           n6411, ZN => n3131);
   U1059 : OAI22_X1 port map( A1 => n4838, A2 => n6412, B1 => n1686, B2 => 
                           n6411, ZN => n3132);
   U1095 : OAI22_X1 port map( A1 => n4772, A2 => n6412, B1 => n1722, B2 => 
                           n6411, ZN => n3114);
   U1057 : OAI22_X1 port map( A1 => n4839, A2 => n6412, B1 => n1684, B2 => 
                           n6411, ZN => n3133);
   U1087 : OAI22_X1 port map( A1 => n4783, A2 => n6412, B1 => n1714, B2 => 
                           n6411, ZN => n3118);
   U1053 : OAI22_X1 port map( A1 => n4844, A2 => n3926, B1 => n1680, B2 => 
                           n6411, ZN => n3135);
   U1083 : OAI22_X1 port map( A1 => n4785, A2 => n6412, B1 => n1710, B2 => 
                           n6411, ZN => n3120);
   U1085 : OAI22_X1 port map( A1 => n4784, A2 => n6412, B1 => n1712, B2 => 
                           n6411, ZN => n3119);
   U1097 : OAI22_X1 port map( A1 => n4763, A2 => n6412, B1 => n1724, B2 => 
                           n6411, ZN => n3113);
   U1093 : OAI22_X1 port map( A1 => n4773, A2 => n6412, B1 => n1720, B2 => 
                           n6411, ZN => n3115);
   U667 : OAI22_X1 port map( A1 => n6290, A2 => n6425, B1 => n1694, B2 => n6424
                           , ZN => n3352);
   U653 : OAI22_X1 port map( A1 => n6297, A2 => n1956, B1 => n1680, B2 => n6424
                           , ZN => n3359);
   U657 : OAI22_X1 port map( A1 => n6295, A2 => n6425, B1 => n1684, B2 => n6424
                           , ZN => n3357);
   U655 : OAI22_X1 port map( A1 => n6296, A2 => n6425, B1 => n1682, B2 => n6424
                           , ZN => n3358);
   U659 : OAI22_X1 port map( A1 => n6294, A2 => n6425, B1 => n1686, B2 => n6424
                           , ZN => n3356);
   U753 : OAI22_X1 port map( A1 => n6093, A2 => n6423, B1 => n1714, B2 => n6422
                           , ZN => n3310);
   U661 : OAI22_X1 port map( A1 => n6293, A2 => n6425, B1 => n1688, B2 => n6424
                           , ZN => n3355);
   U669 : OAI22_X1 port map( A1 => n6289, A2 => n6425, B1 => n1696, B2 => n6424
                           , ZN => n3351);
   U671 : OAI22_X1 port map( A1 => n6288, A2 => n6425, B1 => n1698, B2 => n6424
                           , ZN => n3350);
   U739 : OAI22_X1 port map( A1 => n6100, A2 => n6423, B1 => n1700, B2 => n6422
                           , ZN => n3317);
   U663 : OAI22_X1 port map( A1 => n6292, A2 => n6425, B1 => n1690, B2 => n6424
                           , ZN => n3354);
   U763 : OAI22_X1 port map( A1 => n6088, A2 => n6423, B1 => n1724, B2 => n6422
                           , ZN => n3305);
   U761 : OAI22_X1 port map( A1 => n6089, A2 => n6423, B1 => n1722, B2 => n6422
                           , ZN => n3306);
   U759 : OAI22_X1 port map( A1 => n6090, A2 => n6423, B1 => n1720, B2 => n6422
                           , ZN => n3307);
   U721 : OAI22_X1 port map( A1 => n6109, A2 => n6423, B1 => n1682, B2 => n6422
                           , ZN => n3326);
   U719 : OAI22_X1 port map( A1 => n6110, A2 => n1990, B1 => n1680, B2 => n6422
                           , ZN => n3327);
   U675 : OAI22_X1 port map( A1 => n6286, A2 => n6425, B1 => n1702, B2 => n6424
                           , ZN => n3348);
   U697 : OAI22_X1 port map( A1 => n6275, A2 => n6425, B1 => n1724, B2 => n6424
                           , ZN => n3337);
   U665 : OAI22_X1 port map( A1 => n6291, A2 => n6425, B1 => n1692, B2 => n6424
                           , ZN => n3353);
   U693 : OAI22_X1 port map( A1 => n6277, A2 => n6425, B1 => n1720, B2 => n6424
                           , ZN => n3339);
   U687 : OAI22_X1 port map( A1 => n6280, A2 => n6425, B1 => n1714, B2 => n6424
                           , ZN => n3342);
   U685 : OAI22_X1 port map( A1 => n6281, A2 => n6425, B1 => n1712, B2 => n6424
                           , ZN => n3343);
   U683 : OAI22_X1 port map( A1 => n6282, A2 => n6425, B1 => n1710, B2 => n6424
                           , ZN => n3344);
   U737 : OAI22_X1 port map( A1 => n6101, A2 => n6423, B1 => n1698, B2 => n6422
                           , ZN => n3318);
   U735 : OAI22_X1 port map( A1 => n6102, A2 => n6423, B1 => n1696, B2 => n6422
                           , ZN => n3319);
   U733 : OAI22_X1 port map( A1 => n6103, A2 => n6423, B1 => n1694, B2 => n6422
                           , ZN => n3320);
   U731 : OAI22_X1 port map( A1 => n6104, A2 => n6423, B1 => n1692, B2 => n6422
                           , ZN => n3321);
   U727 : OAI22_X1 port map( A1 => n6106, A2 => n6423, B1 => n1688, B2 => n6422
                           , ZN => n3323);
   U729 : OAI22_X1 port map( A1 => n6105, A2 => n6423, B1 => n1690, B2 => n6422
                           , ZN => n3322);
   U673 : OAI22_X1 port map( A1 => n6287, A2 => n6425, B1 => n1700, B2 => n6424
                           , ZN => n3349);
   U725 : OAI22_X1 port map( A1 => n6107, A2 => n6423, B1 => n1686, B2 => n6422
                           , ZN => n3324);
   U749 : OAI22_X1 port map( A1 => n6095, A2 => n6423, B1 => n1710, B2 => n6422
                           , ZN => n3312);
   U723 : OAI22_X1 port map( A1 => n6108, A2 => n6423, B1 => n1684, B2 => n6422
                           , ZN => n3325);
   U695 : OAI22_X1 port map( A1 => n6276, A2 => n6425, B1 => n1722, B2 => n6424
                           , ZN => n3338);
   U751 : OAI22_X1 port map( A1 => n6094, A2 => n6423, B1 => n1712, B2 => n6422
                           , ZN => n3311);
   U741 : OAI22_X1 port map( A1 => n6099, A2 => n6423, B1 => n1702, B2 => n6422
                           , ZN => n3316);
   U617 : OAI22_X1 port map( A1 => n4904, A2 => n6427, B1 => n1710, B2 => n6426
                           , ZN => n3376);
   U605 : OAI22_X1 port map( A1 => n4929, A2 => n6427, B1 => n1698, B2 => n6426
                           , ZN => n3382);
   U603 : OAI22_X1 port map( A1 => n4933, A2 => n6427, B1 => n1696, B2 => n6426
                           , ZN => n3383);
   U627 : OAI22_X1 port map( A1 => n4892, A2 => n6427, B1 => n1720, B2 => n6426
                           , ZN => n3371);
   U607 : OAI22_X1 port map( A1 => n4928, A2 => n6427, B1 => n1700, B2 => n6426
                           , ZN => n3381);
   U609 : OAI22_X1 port map( A1 => n4923, A2 => n6427, B1 => n1702, B2 => n6426
                           , ZN => n3380);
   U591 : OAI22_X1 port map( A1 => n4958, A2 => n6427, B1 => n1684, B2 => n6426
                           , ZN => n3389);
   U619 : OAI22_X1 port map( A1 => n4903, A2 => n6427, B1 => n1712, B2 => n6426
                           , ZN => n3375);
   U621 : OAI22_X1 port map( A1 => n4899, A2 => n6427, B1 => n1714, B2 => n6426
                           , ZN => n3374);
   U587 : OAI22_X1 port map( A1 => n4963, A2 => n1921, B1 => n1680, B2 => n6426
                           , ZN => n3391);
   U629 : OAI22_X1 port map( A1 => n4883, A2 => n6427, B1 => n1722, B2 => n6426
                           , ZN => n3370);
   U631 : OAI22_X1 port map( A1 => n4875, A2 => n6427, B1 => n1724, B2 => n6426
                           , ZN => n3369);
   U597 : OAI22_X1 port map( A1 => n4943, A2 => n6427, B1 => n1690, B2 => n6426
                           , ZN => n3386);
   U589 : OAI22_X1 port map( A1 => n4959, A2 => n6427, B1 => n1682, B2 => n6426
                           , ZN => n3390);
   U593 : OAI22_X1 port map( A1 => n4953, A2 => n6427, B1 => n1686, B2 => n6426
                           , ZN => n3388);
   U595 : OAI22_X1 port map( A1 => n4952, A2 => n6427, B1 => n1688, B2 => n6426
                           , ZN => n3387);
   U601 : OAI22_X1 port map( A1 => n4934, A2 => n6427, B1 => n1694, B2 => n6426
                           , ZN => n3384);
   U599 : OAI22_X1 port map( A1 => n4935, A2 => n6427, B1 => n1692, B2 => n6426
                           , ZN => n3385);
   U1692 : OAI22_X1 port map( A1 => n4515, A2 => n6392, B1 => n1668, B2 => 
                           n6391, ZN => n2787);
   U1666 : OAI22_X1 port map( A1 => n4523, A2 => n4180, B1 => n1666, B2 => 
                           n6391, ZN => n2789);
   U1718 : OAI22_X1 port map( A1 => n4514, A2 => n6392, B1 => n1670, B2 => 
                           n6391, ZN => n2785);
   U2160 : OAI22_X1 port map( A1 => n4453, A2 => n6392, B1 => n1704, B2 => 
                           n6391, ZN => n2751);
   U1796 : OAI22_X1 port map( A1 => n4508, A2 => n6392, B1 => n1676, B2 => 
                           n6391, ZN => n2779);
   U1822 : OAI22_X1 port map( A1 => n4503, A2 => n4180, B1 => n1678, B2 => 
                           n6391, ZN => n2777);
   U1848 : OAI22_X1 port map( A1 => n4502, A2 => n4180, B1 => n1680, B2 => 
                           n6391, ZN => n2775);
   U1952 : OAI22_X1 port map( A1 => n4483, A2 => n6392, B1 => n1688, B2 => 
                           n6391, ZN => n2767);
   U1978 : OAI22_X1 port map( A1 => n4479, A2 => n6392, B1 => n1690, B2 => 
                           n6391, ZN => n2765);
   U2004 : OAI22_X1 port map( A1 => n4478, A2 => n6392, B1 => n1692, B2 => 
                           n6391, ZN => n2763);
   U2030 : OAI22_X1 port map( A1 => n4473, A2 => n6392, B1 => n1694, B2 => 
                           n6391, ZN => n2761);
   U2056 : OAI22_X1 port map( A1 => n4472, A2 => n6392, B1 => n1696, B2 => 
                           n6391, ZN => n2759);
   U2082 : OAI22_X1 port map( A1 => n4463, A2 => n6392, B1 => n1698, B2 => 
                           n6391, ZN => n2757);
   U2186 : OAI22_X1 port map( A1 => n4449, A2 => n6392, B1 => n1706, B2 => 
                           n6391, ZN => n2749);
   U2238 : OAI22_X1 port map( A1 => n4443, A2 => n6392, B1 => n1710, B2 => 
                           n6391, ZN => n2745);
   U2108 : OAI22_X1 port map( A1 => n4455, A2 => n6392, B1 => n1700, B2 => 
                           n6391, ZN => n2755);
   U2212 : OAI22_X1 port map( A1 => n4448, A2 => n6392, B1 => n1708, B2 => 
                           n6391, ZN => n2747);
   U2134 : OAI22_X1 port map( A1 => n4454, A2 => n6392, B1 => n1702, B2 => 
                           n6391, ZN => n2753);
   U1179 : OAI22_X1 port map( A1 => n525, A2 => n6408, B1 => n6407, B2 => n1684
                           , ZN => n3069);
   U1181 : OAI22_X1 port map( A1 => n527, A2 => n6408, B1 => n6407, B2 => n1688
                           , ZN => n3067);
   U1178 : OAI22_X1 port map( A1 => n524, A2 => n6408, B1 => n6407, B2 => n1682
                           , ZN => n3070);
   U1183 : OAI22_X1 port map( A1 => n529, A2 => n6408, B1 => n6407, B2 => n1692
                           , ZN => n3065);
   U1184 : OAI22_X1 port map( A1 => n530, A2 => n6408, B1 => n6407, B2 => n1694
                           , ZN => n3064);
   U1198 : OAI22_X1 port map( A1 => n544, A2 => n6408, B1 => n6407, B2 => n1722
                           , ZN => n3050);
   U1185 : OAI22_X1 port map( A1 => n531, A2 => n6408, B1 => n6407, B2 => n1696
                           , ZN => n3063);
   U1186 : OAI22_X1 port map( A1 => n532, A2 => n6408, B1 => n6407, B2 => n1698
                           , ZN => n3062);
   U1187 : OAI22_X1 port map( A1 => n533, A2 => n6408, B1 => n6407, B2 => n1700
                           , ZN => n3061);
   U1177 : OAI22_X1 port map( A1 => n523, A2 => n3994, B1 => n6407, B2 => n1680
                           , ZN => n3071);
   U1188 : OAI22_X1 port map( A1 => n534, A2 => n6408, B1 => n6407, B2 => n1702
                           , ZN => n3060);
   U1192 : OAI22_X1 port map( A1 => n538, A2 => n6408, B1 => n6407, B2 => n1710
                           , ZN => n3056);
   U1193 : OAI22_X1 port map( A1 => n539, A2 => n6408, B1 => n6407, B2 => n1712
                           , ZN => n3055);
   U1180 : OAI22_X1 port map( A1 => n526, A2 => n6408, B1 => n6407, B2 => n1686
                           , ZN => n3068);
   U1194 : OAI22_X1 port map( A1 => n540, A2 => n6408, B1 => n6407, B2 => n1714
                           , ZN => n3054);
   U1197 : OAI22_X1 port map( A1 => n543, A2 => n6408, B1 => n6407, B2 => n1720
                           , ZN => n3051);
   U1182 : OAI22_X1 port map( A1 => n528, A2 => n6408, B1 => n6407, B2 => n1690
                           , ZN => n3066);
   U1189 : OAI22_X1 port map( A1 => n535, A2 => n6408, B1 => n6407, B2 => n1704
                           , ZN => n3059);
   U783 : OAI22_X1 port map( A1 => n718, A2 => n6421, B1 => n6420, B2 => n1692,
                           ZN => n3289);
   U786 : OAI22_X1 port map( A1 => n721, A2 => n6421, B1 => n6420, B2 => n1698,
                           ZN => n3286);
   U782 : OAI22_X1 port map( A1 => n717, A2 => n6421, B1 => n6420, B2 => n1690,
                           ZN => n3290);
   U781 : OAI22_X1 port map( A1 => n716, A2 => n6421, B1 => n6420, B2 => n1688,
                           ZN => n3291);
   U780 : OAI22_X1 port map( A1 => n715, A2 => n6421, B1 => n6420, B2 => n1686,
                           ZN => n3292);
   U779 : OAI22_X1 port map( A1 => n714, A2 => n6421, B1 => n6420, B2 => n1684,
                           ZN => n3293);
   U778 : OAI22_X1 port map( A1 => n713, A2 => n6421, B1 => n6420, B2 => n1682,
                           ZN => n3294);
   U777 : OAI22_X1 port map( A1 => n712, A2 => n2023, B1 => n6420, B2 => n1680,
                           ZN => n3295);
   U788 : OAI22_X1 port map( A1 => n723, A2 => n6421, B1 => n6420, B2 => n1702,
                           ZN => n3284);
   U798 : OAI22_X1 port map( A1 => n733, A2 => n6421, B1 => n6420, B2 => n1722,
                           ZN => n3274);
   U797 : OAI22_X1 port map( A1 => n732, A2 => n6421, B1 => n6420, B2 => n1720,
                           ZN => n3275);
   U794 : OAI22_X1 port map( A1 => n729, A2 => n6421, B1 => n6420, B2 => n1714,
                           ZN => n3278);
   U793 : OAI22_X1 port map( A1 => n728, A2 => n6421, B1 => n6420, B2 => n1712,
                           ZN => n3279);
   U792 : OAI22_X1 port map( A1 => n727, A2 => n6421, B1 => n6420, B2 => n1710,
                           ZN => n3280);
   U789 : OAI22_X1 port map( A1 => n724, A2 => n6421, B1 => n6420, B2 => n1704,
                           ZN => n3283);
   U785 : OAI22_X1 port map( A1 => n720, A2 => n6421, B1 => n6420, B2 => n1696,
                           ZN => n3287);
   U787 : OAI22_X1 port map( A1 => n722, A2 => n6421, B1 => n6420, B2 => n1700,
                           ZN => n3285);
   U784 : OAI22_X1 port map( A1 => n719, A2 => n6421, B1 => n6420, B2 => n1694,
                           ZN => n3288);
   U1609 : OAI22_X1 port map( A1 => n6193, A2 => n6394, B1 => n1700, B2 => 
                           n6393, ZN => n2805);
   U1629 : OAI22_X1 port map( A1 => n6183, A2 => n6394, B1 => n1720, B2 => 
                           n6393, ZN => n2795);
   U1619 : OAI22_X1 port map( A1 => n6188, A2 => n6394, B1 => n1710, B2 => 
                           n6393, ZN => n2800);
   U1605 : OAI22_X1 port map( A1 => n6195, A2 => n6394, B1 => n1696, B2 => 
                           n6393, ZN => n2807);
   U1603 : OAI22_X1 port map( A1 => n6196, A2 => n6394, B1 => n1694, B2 => 
                           n6393, ZN => n2808);
   U1601 : OAI22_X1 port map( A1 => n6197, A2 => n6394, B1 => n1692, B2 => 
                           n6393, ZN => n2809);
   U1595 : OAI22_X1 port map( A1 => n6200, A2 => n6394, B1 => n1686, B2 => 
                           n6393, ZN => n2812);
   U1631 : OAI22_X1 port map( A1 => n6182, A2 => n6394, B1 => n1722, B2 => 
                           n6393, ZN => n2794);
   U1621 : OAI22_X1 port map( A1 => n6187, A2 => n6394, B1 => n1712, B2 => 
                           n6393, ZN => n2799);
   U1607 : OAI22_X1 port map( A1 => n6194, A2 => n6394, B1 => n1698, B2 => 
                           n6393, ZN => n2806);
   U1613 : OAI22_X1 port map( A1 => n6191, A2 => n6394, B1 => n1704, B2 => 
                           n6393, ZN => n2803);
   U1599 : OAI22_X1 port map( A1 => n6198, A2 => n6394, B1 => n1690, B2 => 
                           n6393, ZN => n2810);
   U1597 : OAI22_X1 port map( A1 => n6199, A2 => n6394, B1 => n1688, B2 => 
                           n6393, ZN => n2811);
   U1593 : OAI22_X1 port map( A1 => n6201, A2 => n6394, B1 => n1684, B2 => 
                           n6393, ZN => n2813);
   U1611 : OAI22_X1 port map( A1 => n6192, A2 => n6394, B1 => n1702, B2 => 
                           n6393, ZN => n2804);
   U1591 : OAI22_X1 port map( A1 => n6202, A2 => n6394, B1 => n1682, B2 => 
                           n6393, ZN => n2814);
   U1623 : OAI22_X1 port map( A1 => n6186, A2 => n6394, B1 => n1714, B2 => 
                           n6393, ZN => n2798);
   U1589 : OAI22_X1 port map( A1 => n6203, A2 => n4145, B1 => n1680, B2 => 
                           n6393, ZN => n2815);
   U1163 : OAI22_X1 port map( A1 => n4652, A2 => n6410, B1 => n1724, B2 => 
                           n6409, ZN => n3081);
   U1109 : OAI22_X1 port map( A1 => n4749, A2 => n6410, B1 => n1670, B2 => 
                           n6409, ZN => n3108);
   U1165 : OAI22_X1 port map( A1 => n6340, A2 => n6410, B1 => n1726, B2 => 
                           n6409, ZN => n3080);
   U1113 : OAI22_X1 port map( A1 => n4743, A2 => n6410, B1 => n1674, B2 => 
                           n6409, ZN => n3106);
   U1151 : OAI22_X1 port map( A1 => n4665, A2 => n6410, B1 => n1712, B2 => 
                           n6409, ZN => n3087);
   U1137 : OAI22_X1 port map( A1 => n4694, A2 => n6410, B1 => n1698, B2 => 
                           n6409, ZN => n3094);
   U1135 : OAI22_X1 port map( A1 => n4695, A2 => n6410, B1 => n1696, B2 => 
                           n6409, ZN => n3095);
   U1155 : OAI22_X1 port map( A1 => n4663, A2 => n6410, B1 => n1716, B2 => 
                           n6409, ZN => n3085);
   U1139 : OAI22_X1 port map( A1 => n4693, A2 => n6410, B1 => n1700, B2 => 
                           n6409, ZN => n3093);
   U1157 : OAI22_X1 port map( A1 => n4659, A2 => n6410, B1 => n1718, B2 => 
                           n6409, ZN => n3084);
   U1159 : OAI22_X1 port map( A1 => n4658, A2 => n6410, B1 => n1720, B2 => 
                           n6409, ZN => n3083);
   U1161 : OAI22_X1 port map( A1 => n4653, A2 => n6410, B1 => n1722, B2 => 
                           n6409, ZN => n3082);
   U1125 : OAI22_X1 port map( A1 => n4719, A2 => n6410, B1 => n1686, B2 => 
                           n6409, ZN => n3100);
   U1149 : OAI22_X1 port map( A1 => n4673, A2 => n6410, B1 => n1710, B2 => 
                           n6409, ZN => n3088);
   U1153 : OAI22_X1 port map( A1 => n4664, A2 => n6410, B1 => n1714, B2 => 
                           n6409, ZN => n3086);
   U1145 : OAI22_X1 port map( A1 => n4683, A2 => n6410, B1 => n1706, B2 => 
                           n6409, ZN => n3090);
   U1143 : OAI22_X1 port map( A1 => n4688, A2 => n6410, B1 => n1704, B2 => 
                           n6409, ZN => n3091);
   U1127 : OAI22_X1 port map( A1 => n4718, A2 => n6410, B1 => n1688, B2 => 
                           n6409, ZN => n3099);
   U1147 : OAI22_X1 port map( A1 => n4682, A2 => n6410, B1 => n1708, B2 => 
                           n6409, ZN => n3089);
   U1490 : OAI22_X1 port map( A1 => n564, A2 => n6398, B1 => n6397, B2 => n1700
                           , ZN => n2869);
   U1489 : OAI22_X1 port map( A1 => n563, A2 => n6398, B1 => n6397, B2 => n1698
                           , ZN => n2870);
   U1487 : OAI22_X1 port map( A1 => n561, A2 => n6398, B1 => n6397, B2 => n1694
                           , ZN => n2872);
   U1486 : OAI22_X1 port map( A1 => n560, A2 => n6398, B1 => n6397, B2 => n1692
                           , ZN => n2873);
   U1500 : OAI22_X1 port map( A1 => n574, A2 => n6398, B1 => n6397, B2 => n1720
                           , ZN => n2859);
   U1488 : OAI22_X1 port map( A1 => n562, A2 => n6398, B1 => n6397, B2 => n1696
                           , ZN => n2871);
   U1483 : OAI22_X1 port map( A1 => n557, A2 => n6398, B1 => n6397, B2 => n1686
                           , ZN => n2876);
   U1482 : OAI22_X1 port map( A1 => n556, A2 => n6398, B1 => n6397, B2 => n1684
                           , ZN => n2877);
   U1481 : OAI22_X1 port map( A1 => n555, A2 => n6398, B1 => n6397, B2 => n1682
                           , ZN => n2878);
   U1480 : OAI22_X1 port map( A1 => n554, A2 => n4106, B1 => n6397, B2 => n1680
                           , ZN => n2879);
   U1491 : OAI22_X1 port map( A1 => n565, A2 => n6398, B1 => n6397, B2 => n1702
                           , ZN => n2868);
   U1485 : OAI22_X1 port map( A1 => n559, A2 => n6398, B1 => n6397, B2 => n1690
                           , ZN => n2874);
   U1502 : OAI22_X1 port map( A1 => n576, A2 => n6398, B1 => n6397, B2 => n1724
                           , ZN => n2857);
   U1501 : OAI22_X1 port map( A1 => n575, A2 => n6398, B1 => n6397, B2 => n1722
                           , ZN => n2858);
   U1495 : OAI22_X1 port map( A1 => n569, A2 => n6398, B1 => n6397, B2 => n1710
                           , ZN => n2864);
   U1499 : OAI22_X1 port map( A1 => n573, A2 => n6398, B1 => n6397, B2 => n1718
                           , ZN => n2860);
   U1496 : OAI22_X1 port map( A1 => n570, A2 => n6398, B1 => n6397, B2 => n1712
                           , ZN => n2863);
   U1484 : OAI22_X1 port map( A1 => n558, A2 => n6398, B1 => n6397, B2 => n1688
                           , ZN => n2875);
   U1373 : OAI22_X1 port map( A1 => n2245, A2 => n6401, B1 => n3886, B2 => 
                           n1670, ZN => n2948);
   U1389 : OAI22_X1 port map( A1 => n2229, A2 => n6401, B1 => n3886, B2 => 
                           n1702, ZN => n2932);
   U1383 : OAI22_X1 port map( A1 => n2235, A2 => n6401, B1 => n3886, B2 => 
                           n1690, ZN => n2938);
   U1380 : OAI22_X1 port map( A1 => n2238, A2 => n6401, B1 => n3886, B2 => 
                           n1684, ZN => n2941);
   U1377 : OAI22_X1 port map( A1 => n2241, A2 => n4068, B1 => n3886, B2 => 
                           n1678, ZN => n2944);
   U1378 : OAI22_X1 port map( A1 => n2240, A2 => n4068, B1 => n3886, B2 => 
                           n1680, ZN => n2943);
   U1384 : OAI22_X1 port map( A1 => n2234, A2 => n6401, B1 => n3886, B2 => 
                           n1692, ZN => n2937);
   U1385 : OAI22_X1 port map( A1 => n2233, A2 => n6401, B1 => n3886, B2 => 
                           n1694, ZN => n2936);
   U1379 : OAI22_X1 port map( A1 => n2239, A2 => n6401, B1 => n3886, B2 => 
                           n1682, ZN => n2942);
   U1387 : OAI22_X1 port map( A1 => n2231, A2 => n6401, B1 => n3886, B2 => 
                           n1698, ZN => n2934);
   U1375 : OAI22_X1 port map( A1 => n2243, A2 => n4068, B1 => n3886, B2 => 
                           n1674, ZN => n2946);
   U1386 : OAI22_X1 port map( A1 => n2232, A2 => n6401, B1 => n3886, B2 => 
                           n1696, ZN => n2935);
   U1381 : OAI22_X1 port map( A1 => n2237, A2 => n6401, B1 => n3886, B2 => 
                           n1686, ZN => n2940);
   U1382 : OAI22_X1 port map( A1 => n2236, A2 => n6401, B1 => n3886, B2 => 
                           n1688, ZN => n2939);
   U1388 : OAI22_X1 port map( A1 => n2230, A2 => n6401, B1 => n3886, B2 => 
                           n1700, ZN => n2933);
   U383 : OAI22_X1 port map( A1 => n2653, A2 => n6434, B1 => n3881, B2 => n1686
                           , ZN => n3516);
   U379 : OAI22_X1 port map( A1 => n2657, A2 => n1847, B1 => n3881, B2 => n1678
                           , ZN => n3520);
   U382 : OAI22_X1 port map( A1 => n2654, A2 => n6434, B1 => n3881, B2 => n1684
                           , ZN => n3517);
   U380 : OAI22_X1 port map( A1 => n2656, A2 => n1847, B1 => n3881, B2 => n1680
                           , ZN => n3519);
   U384 : OAI22_X1 port map( A1 => n2652, A2 => n6434, B1 => n3881, B2 => n1688
                           , ZN => n3515);
   U385 : OAI22_X1 port map( A1 => n2651, A2 => n6434, B1 => n3881, B2 => n1690
                           , ZN => n3514);
   U377 : OAI22_X1 port map( A1 => n2659, A2 => n1847, B1 => n3881, B2 => n1674
                           , ZN => n3522);
   U388 : OAI22_X1 port map( A1 => n2648, A2 => n6434, B1 => n3881, B2 => n1696
                           , ZN => n3511);
   U389 : OAI22_X1 port map( A1 => n2647, A2 => n6434, B1 => n3881, B2 => n1698
                           , ZN => n3510);
   U386 : OAI22_X1 port map( A1 => n2650, A2 => n6434, B1 => n3881, B2 => n1692
                           , ZN => n3513);
   U381 : OAI22_X1 port map( A1 => n2655, A2 => n6434, B1 => n3881, B2 => n1682
                           , ZN => n3518);
   U375 : OAI22_X1 port map( A1 => n2661, A2 => n6434, B1 => n3881, B2 => n1670
                           , ZN => n3524);
   U387 : OAI22_X1 port map( A1 => n2649, A2 => n6434, B1 => n3881, B2 => n1694
                           , ZN => n3512);
   U390 : OAI22_X1 port map( A1 => n2646, A2 => n6434, B1 => n3881, B2 => n1700
                           , ZN => n3509);
   U391 : OAI22_X1 port map( A1 => n2645, A2 => n6434, B1 => n3881, B2 => n1702
                           , ZN => n3508);
   U1400 : OAI22_X1 port map( A1 => n6243, A2 => n6401, B1 => n1724, B2 => 
                           n3886, ZN => n2921);
   U1402 : OAI22_X1 port map( A1 => n4167, A2 => n6401, B1 => n1726, B2 => 
                           n3886, ZN => n2920);
   U403 : OAI22_X1 port map( A1 => n4169, A2 => n6434, B1 => n1726, B2 => n3881
                           , ZN => n3496);
   U1348 : OAI22_X1 port map( A1 => n6158, A2 => n6403, B1 => n1708, B2 => 
                           n4036, ZN => n2961);
   U1304 : OAI22_X1 port map( A1 => n6180, A2 => n4035, B1 => n1663, B2 => 
                           n4036, ZN => n2983);
   U1306 : OAI22_X1 port map( A1 => n6179, A2 => n4035, B1 => n1666, B2 => 
                           n4036, ZN => n2982);
   U1312 : OAI22_X1 port map( A1 => n6176, A2 => n6403, B1 => n1672, B2 => 
                           n4036, ZN => n2979);
   U1356 : OAI22_X1 port map( A1 => n6154, A2 => n6403, B1 => n1716, B2 => 
                           n4036, ZN => n2957);
   U1406 : OAI22_X1 port map( A1 => n6242, A2 => n4073, B1 => n1663, B2 => 
                           n4074, ZN => n2919);
   U1346 : OAI22_X1 port map( A1 => n6159, A2 => n6403, B1 => n1706, B2 => 
                           n4036, ZN => n2962);
   U1344 : OAI22_X1 port map( A1 => n6160, A2 => n6403, B1 => n1704, B2 => 
                           n4036, ZN => n2963);
   U1318 : OAI22_X1 port map( A1 => n6173, A2 => n4035, B1 => n1678, B2 => 
                           n4036, ZN => n2976);
   U1316 : OAI22_X1 port map( A1 => n6174, A2 => n4035, B1 => n1676, B2 => 
                           n4036, ZN => n2977);
   U1314 : OAI22_X1 port map( A1 => n6175, A2 => n6403, B1 => n1674, B2 => 
                           n4036, ZN => n2978);
   U1366 : OAI22_X1 port map( A1 => n6339, A2 => n6403, B1 => n1726, B2 => 
                           n4036, ZN => n2952);
   U1358 : OAI22_X1 port map( A1 => n6153, A2 => n6403, B1 => n1718, B2 => 
                           n4036, ZN => n2956);
   U1418 : OAI22_X1 port map( A1 => n6236, A2 => n4073, B1 => n1676, B2 => 
                           n4074, ZN => n2913);
   U1420 : OAI22_X1 port map( A1 => n6235, A2 => n4073, B1 => n1678, B2 => 
                           n4074, ZN => n2912);
   U1446 : OAI22_X1 port map( A1 => n6222, A2 => n6400, B1 => n1704, B2 => 
                           n4074, ZN => n2899);
   U1448 : OAI22_X1 port map( A1 => n6221, A2 => n6400, B1 => n1706, B2 => 
                           n4074, ZN => n2898);
   U1450 : OAI22_X1 port map( A1 => n6220, A2 => n6400, B1 => n1708, B2 => 
                           n4074, ZN => n2897);
   U1458 : OAI22_X1 port map( A1 => n6216, A2 => n6400, B1 => n1716, B2 => 
                           n4074, ZN => n2893);
   U1460 : OAI22_X1 port map( A1 => n6215, A2 => n6400, B1 => n1718, B2 => 
                           n4074, ZN => n2892);
   U1468 : OAI22_X1 port map( A1 => n6348, A2 => n6400, B1 => n1726, B2 => 
                           n4074, ZN => n2888);
   U1310 : OAI22_X1 port map( A1 => n6177, A2 => n6403, B1 => n1670, B2 => 
                           n4036, ZN => n2980);
   U1308 : OAI22_X1 port map( A1 => n6178, A2 => n6403, B1 => n1668, B2 => 
                           n4036, ZN => n2981);
   U1408 : OAI22_X1 port map( A1 => n6241, A2 => n4073, B1 => n1666, B2 => 
                           n4074, ZN => n2918);
   U1410 : OAI22_X1 port map( A1 => n6240, A2 => n6400, B1 => n1668, B2 => 
                           n4074, ZN => n2917);
   U1412 : OAI22_X1 port map( A1 => n6239, A2 => n6400, B1 => n1670, B2 => 
                           n4074, ZN => n2916);
   U1414 : OAI22_X1 port map( A1 => n6238, A2 => n6400, B1 => n1672, B2 => 
                           n4074, ZN => n2915);
   U1416 : OAI22_X1 port map( A1 => n6237, A2 => n6400, B1 => n1674, B2 => 
                           n4074, ZN => n2914);
   U1250 : OAI22_X1 port map( A1 => n6143, A2 => n4000, B1 => n1676, B2 => 
                           n4001, ZN => n3009);
   U1252 : OAI22_X1 port map( A1 => n6142, A2 => n4000, B1 => n1678, B2 => 
                           n4001, ZN => n3008);
   U1278 : OAI22_X1 port map( A1 => n6129, A2 => n6405, B1 => n1704, B2 => 
                           n4001, ZN => n2995);
   U1238 : OAI22_X1 port map( A1 => n6149, A2 => n4000, B1 => n1663, B2 => 
                           n4001, ZN => n3015);
   U1240 : OAI22_X1 port map( A1 => n6148, A2 => n4000, B1 => n1666, B2 => 
                           n4001, ZN => n3014);
   U1242 : OAI22_X1 port map( A1 => n6147, A2 => n6405, B1 => n1668, B2 => 
                           n4001, ZN => n3013);
   U1244 : OAI22_X1 port map( A1 => n6146, A2 => n6405, B1 => n1670, B2 => 
                           n4001, ZN => n3012);
   U1246 : OAI22_X1 port map( A1 => n6145, A2 => n6405, B1 => n1672, B2 => 
                           n4001, ZN => n3011);
   U1248 : OAI22_X1 port map( A1 => n6144, A2 => n6405, B1 => n1674, B2 => 
                           n4001, ZN => n3010);
   U1282 : OAI22_X1 port map( A1 => n6127, A2 => n6405, B1 => n1708, B2 => 
                           n4001, ZN => n2993);
   U1290 : OAI22_X1 port map( A1 => n6123, A2 => n6405, B1 => n1716, B2 => 
                           n4001, ZN => n2989);
   U1280 : OAI22_X1 port map( A1 => n6128, A2 => n6405, B1 => n1706, B2 => 
                           n4001, ZN => n2994);
   U1292 : OAI22_X1 port map( A1 => n6122, A2 => n6405, B1 => n1718, B2 => 
                           n4001, ZN => n2988);
   U1298 : OAI22_X1 port map( A1 => n6119, A2 => n6405, B1 => n1724, B2 => 
                           n4001, ZN => n2985);
   U1391 : OAI22_X1 port map( A1 => n2227, A2 => n6401, B1 => n3886, B2 => 
                           n1706, ZN => n2930);
   U1374 : OAI22_X1 port map( A1 => n2244, A2 => n6401, B1 => n3886, B2 => 
                           n1672, ZN => n2947);
   U1390 : OAI22_X1 port map( A1 => n2228, A2 => n6401, B1 => n3886, B2 => 
                           n1704, ZN => n2931);
   U1394 : OAI22_X1 port map( A1 => n2224, A2 => n6401, B1 => n3886, B2 => 
                           n1712, ZN => n2927);
   U1372 : OAI22_X1 port map( A1 => n2246, A2 => n6401, B1 => n3886, B2 => 
                           n1668, ZN => n2949);
   U1396 : OAI22_X1 port map( A1 => n2222, A2 => n6401, B1 => n3886, B2 => 
                           n1716, ZN => n2925);
   U1397 : OAI22_X1 port map( A1 => n2221, A2 => n6401, B1 => n3886, B2 => 
                           n1718, ZN => n2924);
   U1398 : OAI22_X1 port map( A1 => n2220, A2 => n6401, B1 => n3886, B2 => 
                           n1720, ZN => n2923);
   U1399 : OAI22_X1 port map( A1 => n2219, A2 => n6401, B1 => n3886, B2 => 
                           n1722, ZN => n2922);
   U1392 : OAI22_X1 port map( A1 => n2226, A2 => n6401, B1 => n3886, B2 => 
                           n1708, ZN => n2929);
   U1393 : OAI22_X1 port map( A1 => n2225, A2 => n6401, B1 => n3886, B2 => 
                           n1710, ZN => n2928);
   U1395 : OAI22_X1 port map( A1 => n2223, A2 => n6401, B1 => n3886, B2 => 
                           n1714, ZN => n2926);
   U374 : OAI22_X1 port map( A1 => n2662, A2 => n6434, B1 => n3881, B2 => n1668
                           , ZN => n3525);
   U376 : OAI22_X1 port map( A1 => n2660, A2 => n6434, B1 => n3881, B2 => n1672
                           , ZN => n3523);
   U401 : OAI22_X1 port map( A1 => n2635, A2 => n6434, B1 => n3881, B2 => n1722
                           , ZN => n3498);
   U402 : OAI22_X1 port map( A1 => n2634, A2 => n6434, B1 => n3881, B2 => n1724
                           , ZN => n3497);
   U395 : OAI22_X1 port map( A1 => n2641, A2 => n6434, B1 => n3881, B2 => n1710
                           , ZN => n3504);
   U396 : OAI22_X1 port map( A1 => n2640, A2 => n6434, B1 => n3881, B2 => n1712
                           , ZN => n3503);
   U397 : OAI22_X1 port map( A1 => n2639, A2 => n6434, B1 => n3881, B2 => n1714
                           , ZN => n3502);
   U398 : OAI22_X1 port map( A1 => n2638, A2 => n6434, B1 => n3881, B2 => n1716
                           , ZN => n3501);
   U399 : OAI22_X1 port map( A1 => n2637, A2 => n6434, B1 => n3881, B2 => n1718
                           , ZN => n3500);
   U392 : OAI22_X1 port map( A1 => n2644, A2 => n6434, B1 => n3881, B2 => n1704
                           , ZN => n3507);
   U393 : OAI22_X1 port map( A1 => n2643, A2 => n6434, B1 => n3881, B2 => n1706
                           , ZN => n3506);
   U394 : OAI22_X1 port map( A1 => n2642, A2 => n6434, B1 => n3881, B2 => n1708
                           , ZN => n3505);
   U400 : OAI22_X1 port map( A1 => n2636, A2 => n6434, B1 => n3881, B2 => n1720
                           , ZN => n3499);
   U429 : OAI22_X1 port map( A1 => n5933, A2 => n6433, B1 => n1686, B2 => n1853
                           , ZN => n3484);
   U490 : OAI22_X1 port map( A1 => n5078, A2 => n1885, B1 => n1682, B2 => n1886
                           , ZN => n3454);
   U528 : OAI22_X1 port map( A1 => n5003, A2 => n6431, B1 => n1720, B2 => n1886
                           , ZN => n3435);
   U427 : OAI22_X1 port map( A1 => n5965, A2 => n6433, B1 => n1684, B2 => n1853
                           , ZN => n3485);
   U488 : OAI22_X1 port map( A1 => n5079, A2 => n6431, B1 => n1680, B2 => n1886
                           , ZN => n3455);
   U520 : OAI22_X1 port map( A1 => n5019, A2 => n6431, B1 => n1712, B2 => n1886
                           , ZN => n3439);
   U522 : OAI22_X1 port map( A1 => n5018, A2 => n6431, B1 => n1714, B2 => n1886
                           , ZN => n3438);
   U524 : OAI22_X1 port map( A1 => n5013, A2 => n6431, B1 => n1716, B2 => n1886
                           , ZN => n3437);
   U526 : OAI22_X1 port map( A1 => n5012, A2 => n6431, B1 => n1718, B2 => n1886
                           , ZN => n3436);
   U494 : OAI22_X1 port map( A1 => n5072, A2 => n6431, B1 => n1686, B2 => n1886
                           , ZN => n3452);
   U492 : OAI22_X1 port map( A1 => n5073, A2 => n6431, B1 => n1684, B2 => n1886
                           , ZN => n3453);
   U457 : OAI22_X1 port map( A1 => n5134, A2 => n6433, B1 => n1714, B2 => n1853
                           , ZN => n3470);
   U425 : OAI22_X1 port map( A1 => n5970, A2 => n1852, B1 => n1682, B2 => n1853
                           , ZN => n3486);
   U407 : OAI22_X1 port map( A1 => n5993, A2 => n6433, B1 => n1663, B2 => n1853
                           , ZN => n3495);
   U530 : OAI22_X1 port map( A1 => n4995, A2 => n6431, B1 => n1722, B2 => n1886
                           , ZN => n3434);
   U482 : OAI22_X1 port map( A1 => n5085, A2 => n6431, B1 => n1674, B2 => n1886
                           , ZN => n3458);
   U480 : OAI22_X1 port map( A1 => n5093, A2 => n6431, B1 => n1672, B2 => n1886
                           , ZN => n3459);
   U532 : OAI22_X1 port map( A1 => n4994, A2 => n6431, B1 => n1724, B2 => n1886
                           , ZN => n3433);
   U417 : OAI22_X1 port map( A1 => n5988, A2 => n6433, B1 => n1674, B2 => n1853
                           , ZN => n3490);
   U467 : OAI22_X1 port map( A1 => n5113, A2 => n6433, B1 => n1724, B2 => n1853
                           , ZN => n3465);
   U472 : OAI22_X1 port map( A1 => n5109, A2 => n6431, B1 => n1663, B2 => n1886
                           , ZN => n3463);
   U463 : OAI22_X1 port map( A1 => n5115, A2 => n6433, B1 => n1720, B2 => n1853
                           , ZN => n3467);
   U461 : OAI22_X1 port map( A1 => n5123, A2 => n6433, B1 => n1718, B2 => n1853
                           , ZN => n3468);
   U465 : OAI22_X1 port map( A1 => n5114, A2 => n6433, B1 => n1722, B2 => n1853
                           , ZN => n3466);
   U423 : OAI22_X1 port map( A1 => n5985, A2 => n6433, B1 => n1680, B2 => n1853
                           , ZN => n3487);
   U455 : OAI22_X1 port map( A1 => n5139, A2 => n6433, B1 => n1712, B2 => n1853
                           , ZN => n3471);
   U459 : OAI22_X1 port map( A1 => n5133, A2 => n6433, B1 => n1716, B2 => n1853
                           , ZN => n3469);
   U415 : OAI22_X1 port map( A1 => n5989, A2 => n6433, B1 => n1672, B2 => n1853
                           , ZN => n3491);
   U563 : OAI22_X1 port map( A1 => n508, A2 => n6429, B1 => n1918, B2 => n1716,
                           ZN => n3405);
   U540 : OAI22_X1 port map( A1 => n485, A2 => n6429, B1 => n1918, B2 => n1670,
                           ZN => n3428);
   U539 : OAI22_X1 port map( A1 => n484, A2 => n6429, B1 => n1918, B2 => n1668,
                           ZN => n3429);
   U558 : OAI22_X1 port map( A1 => n503, A2 => n6429, B1 => n1918, B2 => n1706,
                           ZN => n3410);
   U537 : OAI22_X1 port map( A1 => n482, A2 => n1917, B1 => n1918, B2 => n1663,
                           ZN => n3431);
   U538 : OAI22_X1 port map( A1 => n483, A2 => n1917, B1 => n1918, B2 => n1666,
                           ZN => n3430);
   U544 : OAI22_X1 port map( A1 => n489, A2 => n1917, B1 => n1918, B2 => n1678,
                           ZN => n3424);
   U568 : OAI22_X1 port map( A1 => n639, A2 => n6429, B1 => n1918, B2 => n1726,
                           ZN => n3400);
   U541 : OAI22_X1 port map( A1 => n486, A2 => n6429, B1 => n1918, B2 => n1672,
                           ZN => n3427);
   U559 : OAI22_X1 port map( A1 => n504, A2 => n6429, B1 => n1918, B2 => n1708,
                           ZN => n3409);
   U564 : OAI22_X1 port map( A1 => n509, A2 => n6429, B1 => n1918, B2 => n1718,
                           ZN => n3404);
   U543 : OAI22_X1 port map( A1 => n488, A2 => n1917, B1 => n1918, B2 => n1676,
                           ZN => n3425);
   U542 : OAI22_X1 port map( A1 => n487, A2 => n6429, B1 => n1918, B2 => n1674,
                           ZN => n3426);
   U567 : OAI22_X1 port map( A1 => n512, A2 => n6429, B1 => n1918, B2 => n1724,
                           ZN => n3401);
   U345 : OAI22_X1 port map( A1 => n616, A2 => n1843, B1 => n3883, B2 => n1680,
                           ZN => n3551);
   U348 : OAI22_X1 port map( A1 => n619, A2 => n6435, B1 => n3883, B2 => n1686,
                           ZN => n3548);
   U347 : OAI22_X1 port map( A1 => n618, A2 => n6435, B1 => n3883, B2 => n1684,
                           ZN => n3549);
   U351 : OAI22_X1 port map( A1 => n622, A2 => n6435, B1 => n3883, B2 => n1692,
                           ZN => n3545);
   U353 : OAI22_X1 port map( A1 => n624, A2 => n6435, B1 => n3883, B2 => n1696,
                           ZN => n3543);
   U346 : OAI22_X1 port map( A1 => n617, A2 => n6435, B1 => n3883, B2 => n1682,
                           ZN => n3550);
   U355 : OAI22_X1 port map( A1 => n626, A2 => n6435, B1 => n3883, B2 => n1700,
                           ZN => n3541);
   U356 : OAI22_X1 port map( A1 => n627, A2 => n6435, B1 => n3883, B2 => n1702,
                           ZN => n3540);
   U349 : OAI22_X1 port map( A1 => n620, A2 => n6435, B1 => n3883, B2 => n1688,
                           ZN => n3547);
   U350 : OAI22_X1 port map( A1 => n621, A2 => n6435, B1 => n3883, B2 => n1690,
                           ZN => n3546);
   U340 : OAI22_X1 port map( A1 => n611, A2 => n6435, B1 => n3883, B2 => n1670,
                           ZN => n3556);
   U352 : OAI22_X1 port map( A1 => n623, A2 => n6435, B1 => n3883, B2 => n1694,
                           ZN => n3544);
   U342 : OAI22_X1 port map( A1 => n613, A2 => n1843, B1 => n3883, B2 => n1674,
                           ZN => n3554);
   U354 : OAI22_X1 port map( A1 => n625, A2 => n6435, B1 => n3883, B2 => n1698,
                           ZN => n3542);
   U344 : OAI22_X1 port map( A1 => n615, A2 => n1843, B1 => n3883, B2 => n1678,
                           ZN => n3552);
   U250 : OAI22_X1 port map( A1 => n3771, A2 => n6438, B1 => n3882, B2 => n1690
                           , ZN => n3610);
   U245 : OAI22_X1 port map( A1 => n3776, A2 => n1807, B1 => n3882, B2 => n1680
                           , ZN => n3615);
   U246 : OAI22_X1 port map( A1 => n3775, A2 => n6438, B1 => n3882, B2 => n1682
                           , ZN => n3614);
   U247 : OAI22_X1 port map( A1 => n3774, A2 => n6438, B1 => n3882, B2 => n1684
                           , ZN => n3613);
   U248 : OAI22_X1 port map( A1 => n3773, A2 => n6438, B1 => n3882, B2 => n1686
                           , ZN => n3612);
   U249 : OAI22_X1 port map( A1 => n3772, A2 => n6438, B1 => n3882, B2 => n1688
                           , ZN => n3611);
   U253 : OAI22_X1 port map( A1 => n3768, A2 => n6438, B1 => n3882, B2 => n1696
                           , ZN => n3607);
   U251 : OAI22_X1 port map( A1 => n3770, A2 => n6438, B1 => n3882, B2 => n1692
                           , ZN => n3609);
   U252 : OAI22_X1 port map( A1 => n3769, A2 => n6438, B1 => n3882, B2 => n1694
                           , ZN => n3608);
   U256 : OAI22_X1 port map( A1 => n3765, A2 => n6438, B1 => n3882, B2 => n1702
                           , ZN => n3604);
   U254 : OAI22_X1 port map( A1 => n3767, A2 => n6438, B1 => n3882, B2 => n1698
                           , ZN => n3606);
   U255 : OAI22_X1 port map( A1 => n3766, A2 => n6438, B1 => n3882, B2 => n1700
                           , ZN => n3605);
   U240 : OAI22_X1 port map( A1 => n3781, A2 => n6438, B1 => n3882, B2 => n1670
                           , ZN => n3620);
   U244 : OAI22_X1 port map( A1 => n3777, A2 => n1807, B1 => n3882, B2 => n1678
                           , ZN => n3616);
   U242 : OAI22_X1 port map( A1 => n3779, A2 => n1807, B1 => n3882, B2 => n1674
                           , ZN => n3618);
   U368 : OAI22_X1 port map( A1 => n6343, A2 => n6435, B1 => n1726, B2 => n3883
                           , ZN => n3528);
   U55 : OAI22_X1 port map( A1 => n6029, A2 => n6445, B1 => n1716, B2 => n1664,
                           ZN => n3725);
   U3 : OAI22_X1 port map( A1 => n6055, A2 => n1662, B1 => n1663, B2 => n1664, 
                           ZN => n3751);
   U17 : OAI22_X1 port map( A1 => n6048, A2 => n1662, B1 => n1678, B2 => n1664,
                           ZN => n3744);
   U47 : OAI22_X1 port map( A1 => n6033, A2 => n6445, B1 => n1708, B2 => n1664,
                           ZN => n3729);
   U43 : OAI22_X1 port map( A1 => n6035, A2 => n6445, B1 => n1704, B2 => n1664,
                           ZN => n3731);
   U7 : OAI22_X1 port map( A1 => n6053, A2 => n6445, B1 => n1668, B2 => n1664, 
                           ZN => n3749);
   U9 : OAI22_X1 port map( A1 => n6052, A2 => n6445, B1 => n1670, B2 => n1664, 
                           ZN => n3748);
   U45 : OAI22_X1 port map( A1 => n6034, A2 => n6445, B1 => n1706, B2 => n1664,
                           ZN => n3730);
   U65 : OAI22_X1 port map( A1 => n6346, A2 => n6445, B1 => n1726, B2 => n1664,
                           ZN => n3720);
   U5 : OAI22_X1 port map( A1 => n6054, A2 => n1662, B1 => n1666, B2 => n1664, 
                           ZN => n3750);
   U57 : OAI22_X1 port map( A1 => n6028, A2 => n6445, B1 => n1718, B2 => n1664,
                           ZN => n3724);
   U11 : OAI22_X1 port map( A1 => n6051, A2 => n6445, B1 => n1672, B2 => n1664,
                           ZN => n3747);
   U15 : OAI22_X1 port map( A1 => n6049, A2 => n1662, B1 => n1676, B2 => n1664,
                           ZN => n3745);
   U13 : OAI22_X1 port map( A1 => n6050, A2 => n6445, B1 => n1674, B2 => n1664,
                           ZN => n3746);
   U1220 : OAI22_X1 port map( A1 => n689, A2 => n6406, B1 => n3887, B2 => n1698
                           , ZN => n3030);
   U1221 : OAI22_X1 port map( A1 => n690, A2 => n6406, B1 => n3887, B2 => n1700
                           , ZN => n3029);
   U1222 : OAI22_X1 port map( A1 => n691, A2 => n6406, B1 => n3887, B2 => n1702
                           , ZN => n3028);
   U1217 : OAI22_X1 port map( A1 => n686, A2 => n6406, B1 => n3887, B2 => n1692
                           , ZN => n3033);
   U1206 : OAI22_X1 port map( A1 => n675, A2 => n6406, B1 => n3887, B2 => n1670
                           , ZN => n3044);
   U1218 : OAI22_X1 port map( A1 => n687, A2 => n6406, B1 => n3887, B2 => n1694
                           , ZN => n3032);
   U1214 : OAI22_X1 port map( A1 => n683, A2 => n6406, B1 => n3887, B2 => n1686
                           , ZN => n3036);
   U1213 : OAI22_X1 port map( A1 => n682, A2 => n6406, B1 => n3887, B2 => n1684
                           , ZN => n3037);
   U1212 : OAI22_X1 port map( A1 => n681, A2 => n6406, B1 => n3887, B2 => n1682
                           , ZN => n3038);
   U1211 : OAI22_X1 port map( A1 => n680, A2 => n3996, B1 => n3887, B2 => n1680
                           , ZN => n3039);
   U1210 : OAI22_X1 port map( A1 => n679, A2 => n3996, B1 => n3887, B2 => n1678
                           , ZN => n3040);
   U1208 : OAI22_X1 port map( A1 => n677, A2 => n3996, B1 => n3887, B2 => n1674
                           , ZN => n3042);
   U1216 : OAI22_X1 port map( A1 => n685, A2 => n6406, B1 => n3887, B2 => n1690
                           , ZN => n3034);
   U1215 : OAI22_X1 port map( A1 => n684, A2 => n6406, B1 => n3887, B2 => n1688
                           , ZN => n3035);
   U1219 : OAI22_X1 port map( A1 => n688, A2 => n6406, B1 => n3887, B2 => n1696
                           , ZN => n3031);
   U268 : OAI22_X1 port map( A1 => n6344, A2 => n6438, B1 => n1726, B2 => n3882
                           , ZN => n3592);
   U920 : OAI22_X1 port map( A1 => n4175, A2 => n6417, B1 => n1714, B2 => n6416
                           , ZN => n3214);
   U926 : OAI22_X1 port map( A1 => n4172, A2 => n6417, B1 => n1720, B2 => n6416
                           , ZN => n3211);
   U928 : OAI22_X1 port map( A1 => n4171, A2 => n6417, B1 => n1722, B2 => n6416
                           , ZN => n3210);
   U930 : OAI22_X1 port map( A1 => n4170, A2 => n6417, B1 => n1724, B2 => n6416
                           , ZN => n3209);
   U898 : OAI22_X1 port map( A1 => n4242, A2 => n6417, B1 => n1692, B2 => n6416
                           , ZN => n3225);
   U900 : OAI22_X1 port map( A1 => n4230, A2 => n6417, B1 => n1694, B2 => n6416
                           , ZN => n3224);
   U892 : OAI22_X1 port map( A1 => n4253, A2 => n6417, B1 => n1686, B2 => n6416
                           , ZN => n3228);
   U894 : OAI22_X1 port map( A1 => n4245, A2 => n6417, B1 => n1688, B2 => n6416
                           , ZN => n3227);
   U906 : OAI22_X1 port map( A1 => n4213, A2 => n6417, B1 => n1700, B2 => n6416
                           , ZN => n3221);
   U904 : OAI22_X1 port map( A1 => n4222, A2 => n2062, B1 => n1698, B2 => n6416
                           , ZN => n3222);
   U918 : OAI22_X1 port map( A1 => n4176, A2 => n6417, B1 => n1712, B2 => n6416
                           , ZN => n3215);
   U886 : OAI22_X1 port map( A1 => n4268, A2 => n2062, B1 => n1680, B2 => n6416
                           , ZN => n3231);
   U888 : OAI22_X1 port map( A1 => n4263, A2 => n6417, B1 => n1682, B2 => n6416
                           , ZN => n3230);
   U890 : OAI22_X1 port map( A1 => n4262, A2 => n6417, B1 => n1684, B2 => n6416
                           , ZN => n3229);
   U908 : OAI22_X1 port map( A1 => n4206, A2 => n6417, B1 => n1702, B2 => n6416
                           , ZN => n3220);
   U902 : OAI22_X1 port map( A1 => n4227, A2 => n6417, B1 => n1696, B2 => n6416
                           , ZN => n3223);
   U884 : OAI22_X1 port map( A1 => n4269, A2 => n2062, B1 => n1678, B2 => n6416
                           , ZN => n3232);
   U896 : OAI22_X1 port map( A1 => n4244, A2 => n2062, B1 => n1690, B2 => n6416
                           , ZN => n3226);
   U838 : OAI22_X1 port map( A1 => n6257, A2 => n6419, B1 => n1698, B2 => n6418
                           , ZN => n3254);
   U824 : OAI22_X1 port map( A1 => n6264, A2 => n6419, B1 => n1684, B2 => n6418
                           , ZN => n3261);
   U822 : OAI22_X1 port map( A1 => n6265, A2 => n6419, B1 => n1682, B2 => n6418
                           , ZN => n3262);
   U836 : OAI22_X1 port map( A1 => n6258, A2 => n6419, B1 => n1696, B2 => n6418
                           , ZN => n3255);
   U860 : OAI22_X1 port map( A1 => n6246, A2 => n6419, B1 => n1720, B2 => n6418
                           , ZN => n3243);
   U826 : OAI22_X1 port map( A1 => n6263, A2 => n6419, B1 => n1686, B2 => n6418
                           , ZN => n3260);
   U818 : OAI22_X1 port map( A1 => n6267, A2 => n2027, B1 => n1678, B2 => n6418
                           , ZN => n3264);
   U864 : OAI22_X1 port map( A1 => n6244, A2 => n6419, B1 => n1724, B2 => n6418
                           , ZN => n3241);
   U840 : OAI22_X1 port map( A1 => n6256, A2 => n2027, B1 => n1700, B2 => n6418
                           , ZN => n3253);
   U820 : OAI22_X1 port map( A1 => n6266, A2 => n6419, B1 => n1680, B2 => n6418
                           , ZN => n3263);
   U862 : OAI22_X1 port map( A1 => n6245, A2 => n6419, B1 => n1722, B2 => n6418
                           , ZN => n3242);
   U834 : OAI22_X1 port map( A1 => n6259, A2 => n6419, B1 => n1694, B2 => n6418
                           , ZN => n3256);
   U832 : OAI22_X1 port map( A1 => n6260, A2 => n6419, B1 => n1692, B2 => n6418
                           , ZN => n3257);
   U854 : OAI22_X1 port map( A1 => n6249, A2 => n6419, B1 => n1714, B2 => n6418
                           , ZN => n3246);
   U828 : OAI22_X1 port map( A1 => n6262, A2 => n6419, B1 => n1688, B2 => n6418
                           , ZN => n3259);
   U830 : OAI22_X1 port map( A1 => n6261, A2 => n2027, B1 => n1690, B2 => n6418
                           , ZN => n3258);
   U842 : OAI22_X1 port map( A1 => n6255, A2 => n2027, B1 => n1702, B2 => n6418
                           , ZN => n3252);
   U852 : OAI22_X1 port map( A1 => n6250, A2 => n6419, B1 => n1712, B2 => n6418
                           , ZN => n3247);
   U223 : OAI22_X1 port map( A1 => n4313, A2 => n6440, B1 => n1716, B2 => n1773
                           , ZN => n3629);
   U173 : OAI22_X1 port map( A1 => n4412, A2 => n1772, B1 => n1666, B2 => n1773
                           , ZN => n3654);
   U179 : OAI22_X1 port map( A1 => n4394, A2 => n6440, B1 => n1672, B2 => n1773
                           , ZN => n3651);
   U231 : OAI22_X1 port map( A1 => n4299, A2 => n6440, B1 => n1724, B2 => n1773
                           , ZN => n3625);
   U183 : OAI22_X1 port map( A1 => n4389, A2 => n6440, B1 => n1676, B2 => n1773
                           , ZN => n3649);
   U181 : OAI22_X1 port map( A1 => n4393, A2 => n1772, B1 => n1674, B2 => n1773
                           , ZN => n3650);
   U171 : OAI22_X1 port map( A1 => n4413, A2 => n1772, B1 => n1663, B2 => n1773
                           , ZN => n3655);
   U177 : OAI22_X1 port map( A1 => n4395, A2 => n6440, B1 => n1670, B2 => n1773
                           , ZN => n3652);
   U211 : OAI22_X1 port map( A1 => n4334, A2 => n6440, B1 => n1704, B2 => n1773
                           , ZN => n3635);
   U175 : OAI22_X1 port map( A1 => n4403, A2 => n6440, B1 => n1668, B2 => n1773
                           , ZN => n3653);
   U225 : OAI22_X1 port map( A1 => n4305, A2 => n6440, B1 => n1718, B2 => n1773
                           , ZN => n3628);
   U215 : OAI22_X1 port map( A1 => n4329, A2 => n6440, B1 => n1708, B2 => n1773
                           , ZN => n3633);
   U213 : OAI22_X1 port map( A1 => n4333, A2 => n6440, B1 => n1706, B2 => n1773
                           , ZN => n3634);
   U185 : OAI22_X1 port map( A1 => n4388, A2 => n1772, B1 => n1678, B2 => n1773
                           , ZN => n3648);
   U358 : OAI22_X1 port map( A1 => n629, A2 => n6435, B1 => n3883, B2 => n1706,
                           ZN => n3538);
   U362 : OAI22_X1 port map( A1 => n633, A2 => n6435, B1 => n3883, B2 => n1714,
                           ZN => n3534);
   U363 : OAI22_X1 port map( A1 => n634, A2 => n6435, B1 => n3883, B2 => n1716,
                           ZN => n3533);
   U360 : OAI22_X1 port map( A1 => n631, A2 => n6435, B1 => n3883, B2 => n1710,
                           ZN => n3536);
   U359 : OAI22_X1 port map( A1 => n630, A2 => n6435, B1 => n3883, B2 => n1708,
                           ZN => n3537);
   U357 : OAI22_X1 port map( A1 => n628, A2 => n6435, B1 => n3883, B2 => n1704,
                           ZN => n3539);
   U361 : OAI22_X1 port map( A1 => n632, A2 => n6435, B1 => n3883, B2 => n1712,
                           ZN => n3535);
   U339 : OAI22_X1 port map( A1 => n610, A2 => n6435, B1 => n3883, B2 => n1668,
                           ZN => n3557);
   U341 : OAI22_X1 port map( A1 => n612, A2 => n6435, B1 => n3883, B2 => n1672,
                           ZN => n3555);
   U366 : OAI22_X1 port map( A1 => n637, A2 => n6435, B1 => n3883, B2 => n1722,
                           ZN => n3530);
   U365 : OAI22_X1 port map( A1 => n636, A2 => n6435, B1 => n3883, B2 => n1720,
                           ZN => n3531);
   U367 : OAI22_X1 port map( A1 => n638, A2 => n6435, B1 => n3883, B2 => n1724,
                           ZN => n3529);
   U364 : OAI22_X1 port map( A1 => n635, A2 => n6435, B1 => n3883, B2 => n1718,
                           ZN => n3532);
   U257 : OAI22_X1 port map( A1 => n3764, A2 => n6438, B1 => n3882, B2 => n1704
                           , ZN => n3603);
   U259 : OAI22_X1 port map( A1 => n3762, A2 => n6438, B1 => n3882, B2 => n1708
                           , ZN => n3601);
   U258 : OAI22_X1 port map( A1 => n3763, A2 => n6438, B1 => n3882, B2 => n1706
                           , ZN => n3602);
   U267 : OAI22_X1 port map( A1 => n3754, A2 => n6438, B1 => n3882, B2 => n1724
                           , ZN => n3593);
   U263 : OAI22_X1 port map( A1 => n3758, A2 => n6438, B1 => n3882, B2 => n1716
                           , ZN => n3597);
   U265 : OAI22_X1 port map( A1 => n3756, A2 => n6438, B1 => n3882, B2 => n1720
                           , ZN => n3595);
   U264 : OAI22_X1 port map( A1 => n3757, A2 => n6438, B1 => n3882, B2 => n1718
                           , ZN => n3596);
   U260 : OAI22_X1 port map( A1 => n3761, A2 => n6438, B1 => n3882, B2 => n1710
                           , ZN => n3600);
   U239 : OAI22_X1 port map( A1 => n3782, A2 => n6438, B1 => n3882, B2 => n1668
                           , ZN => n3621);
   U262 : OAI22_X1 port map( A1 => n3759, A2 => n6438, B1 => n3882, B2 => n1714
                           , ZN => n3598);
   U261 : OAI22_X1 port map( A1 => n3760, A2 => n6438, B1 => n3882, B2 => n1712
                           , ZN => n3599);
   U241 : OAI22_X1 port map( A1 => n3780, A2 => n6438, B1 => n3882, B2 => n1672
                           , ZN => n3619);
   U266 : OAI22_X1 port map( A1 => n3755, A2 => n6438, B1 => n3882, B2 => n1722
                           , ZN => n3594);
   U1558 : OAI22_X1 port map( A1 => n4544, A2 => n6396, B1 => n1716, B2 => 
                           n4111, ZN => n2829);
   U1510 : OAI22_X1 port map( A1 => n4634, A2 => n6396, B1 => n1668, B2 => 
                           n4111, ZN => n2853);
   U1508 : OAI22_X1 port map( A1 => n4635, A2 => n4110, B1 => n1666, B2 => 
                           n4111, ZN => n2854);
   U1568 : OAI22_X1 port map( A1 => n6338, A2 => n6396, B1 => n1726, B2 => 
                           n4111, ZN => n2824);
   U1566 : OAI22_X1 port map( A1 => n4533, A2 => n6396, B1 => n1724, B2 => 
                           n4111, ZN => n2825);
   U1520 : OAI22_X1 port map( A1 => n4622, A2 => n4110, B1 => n1678, B2 => 
                           n4111, ZN => n2848);
   U1518 : OAI22_X1 port map( A1 => n4623, A2 => n4110, B1 => n1676, B2 => 
                           n4111, ZN => n2849);
   U1516 : OAI22_X1 port map( A1 => n4628, A2 => n6396, B1 => n1674, B2 => 
                           n4111, ZN => n2850);
   U1514 : OAI22_X1 port map( A1 => n4629, A2 => n6396, B1 => n1672, B2 => 
                           n4111, ZN => n2851);
   U1506 : OAI22_X1 port map( A1 => n4643, A2 => n4110, B1 => n1663, B2 => 
                           n4111, ZN => n2855);
   U1550 : OAI22_X1 port map( A1 => n4563, A2 => n6396, B1 => n1708, B2 => 
                           n4111, ZN => n2833);
   U1548 : OAI22_X1 port map( A1 => n4568, A2 => n6396, B1 => n1706, B2 => 
                           n4111, ZN => n2834);
   U1560 : OAI22_X1 port map( A1 => n4543, A2 => n6396, B1 => n1718, B2 => 
                           n4111, ZN => n2828);
   U1512 : OAI22_X1 port map( A1 => n4633, A2 => n6396, B1 => n1670, B2 => 
                           n4111, ZN => n2852);
   U1234 : OAI22_X1 port map( A1 => n6350, A2 => n6406, B1 => n1726, B2 => 
                           n3887, ZN => n3016);
   U332 : OAI22_X1 port map( A1 => n6306, A2 => n6437, B1 => n1724, B2 => n1812
                           , ZN => n3561);
   U330 : OAI22_X1 port map( A1 => n6307, A2 => n6437, B1 => n1722, B2 => n1812
                           , ZN => n3562);
   U328 : OAI22_X1 port map( A1 => n6308, A2 => n6437, B1 => n1720, B2 => n1812
                           , ZN => n3563);
   U326 : OAI22_X1 port map( A1 => n6309, A2 => n6437, B1 => n1718, B2 => n1812
                           , ZN => n3564);
   U324 : OAI22_X1 port map( A1 => n6310, A2 => n6437, B1 => n1716, B2 => n1812
                           , ZN => n3565);
   U322 : OAI22_X1 port map( A1 => n6311, A2 => n6437, B1 => n1714, B2 => n1812
                           , ZN => n3566);
   U320 : OAI22_X1 port map( A1 => n6312, A2 => n6437, B1 => n1712, B2 => n1812
                           , ZN => n3567);
   U280 : OAI22_X1 port map( A1 => n6332, A2 => n6437, B1 => n1672, B2 => n1812
                           , ZN => n3587);
   U282 : OAI22_X1 port map( A1 => n6331, A2 => n6437, B1 => n1674, B2 => n1812
                           , ZN => n3586);
   U288 : OAI22_X1 port map( A1 => n6328, A2 => n6437, B1 => n1680, B2 => n1812
                           , ZN => n3583);
   U290 : OAI22_X1 port map( A1 => n6327, A2 => n1811, B1 => n1682, B2 => n1812
                           , ZN => n3582);
   U1079 : OAI22_X1 port map( A1 => n4802, A2 => n6412, B1 => n1706, B2 => 
                           n3927, ZN => n3122);
   U1081 : OAI22_X1 port map( A1 => n4793, A2 => n6412, B1 => n1708, B2 => 
                           n3927, ZN => n3121);
   U1089 : OAI22_X1 port map( A1 => n4779, A2 => n6412, B1 => n1716, B2 => 
                           n3927, ZN => n3117);
   U1091 : OAI22_X1 port map( A1 => n4778, A2 => n6412, B1 => n1718, B2 => 
                           n3927, ZN => n3116);
   U1099 : OAI22_X1 port map( A1 => n6341, A2 => n6412, B1 => n1726, B2 => 
                           n3927, ZN => n3112);
   U1039 : OAI22_X1 port map( A1 => n4873, A2 => n3926, B1 => n1666, B2 => 
                           n3927, ZN => n3142);
   U1077 : OAI22_X1 port map( A1 => n4803, A2 => n6412, B1 => n1704, B2 => 
                           n3927, ZN => n3123);
   U1041 : OAI22_X1 port map( A1 => n4869, A2 => n6412, B1 => n1668, B2 => 
                           n3927, ZN => n3141);
   U1043 : OAI22_X1 port map( A1 => n4868, A2 => n6412, B1 => n1670, B2 => 
                           n3927, ZN => n3140);
   U1047 : OAI22_X1 port map( A1 => n4862, A2 => n6412, B1 => n1674, B2 => 
                           n3927, ZN => n3138);
   U1049 : OAI22_X1 port map( A1 => n4853, A2 => n3926, B1 => n1676, B2 => 
                           n3927, ZN => n3137);
   U294 : OAI22_X1 port map( A1 => n6325, A2 => n6437, B1 => n1686, B2 => n1812
                           , ZN => n3580);
   U272 : OAI22_X1 port map( A1 => n6336, A2 => n6437, B1 => n1663, B2 => n1812
                           , ZN => n3591);
   U1045 : OAI22_X1 port map( A1 => n4863, A2 => n6412, B1 => n1672, B2 => 
                           n3927, ZN => n3139);
   U1051 : OAI22_X1 port map( A1 => n4845, A2 => n3926, B1 => n1678, B2 => 
                           n3927, ZN => n3136);
   U292 : OAI22_X1 port map( A1 => n6326, A2 => n6437, B1 => n1684, B2 => n1812
                           , ZN => n3581);
   U1037 : OAI22_X1 port map( A1 => n4874, A2 => n3926, B1 => n1663, B2 => 
                           n3927, ZN => n3143);
   U128 : OAI22_X1 port map( A1 => n6012, A2 => n6442, B1 => n1688, B2 => n6441
                           , ZN => n3675);
   U122 : OAI22_X1 port map( A1 => n6015, A2 => n6442, B1 => n1682, B2 => n6441
                           , ZN => n3678);
   U124 : OAI22_X1 port map( A1 => n6014, A2 => n6442, B1 => n1684, B2 => n6441
                           , ZN => n3677);
   U120 : OAI22_X1 port map( A1 => n6016, A2 => n6442, B1 => n1680, B2 => n6441
                           , ZN => n3679);
   U152 : OAI22_X1 port map( A1 => n6000, A2 => n6442, B1 => n1712, B2 => n6441
                           , ZN => n3663);
   U134 : OAI22_X1 port map( A1 => n6009, A2 => n6442, B1 => n1694, B2 => n6441
                           , ZN => n3672);
   U126 : OAI22_X1 port map( A1 => n6013, A2 => n1735, B1 => n1686, B2 => n6441
                           , ZN => n3676);
   U160 : OAI22_X1 port map( A1 => n5996, A2 => n6442, B1 => n1720, B2 => n6441
                           , ZN => n3659);
   U136 : OAI22_X1 port map( A1 => n6008, A2 => n1735, B1 => n1696, B2 => n6441
                           , ZN => n3671);
   U162 : OAI22_X1 port map( A1 => n5995, A2 => n6442, B1 => n1722, B2 => n6441
                           , ZN => n3658);
   U154 : OAI22_X1 port map( A1 => n5999, A2 => n6442, B1 => n1714, B2 => n6441
                           , ZN => n3662);
   U138 : OAI22_X1 port map( A1 => n6007, A2 => n6442, B1 => n1698, B2 => n6441
                           , ZN => n3670);
   U118 : OAI22_X1 port map( A1 => n6017, A2 => n6442, B1 => n1678, B2 => n6441
                           , ZN => n3680);
   U130 : OAI22_X1 port map( A1 => n6011, A2 => n6442, B1 => n1690, B2 => n6441
                           , ZN => n3674);
   U132 : OAI22_X1 port map( A1 => n6010, A2 => n6442, B1 => n1692, B2 => n6441
                           , ZN => n3673);
   U140 : OAI22_X1 port map( A1 => n6006, A2 => n1735, B1 => n1700, B2 => n6441
                           , ZN => n3669);
   U164 : OAI22_X1 port map( A1 => n5994, A2 => n6442, B1 => n1724, B2 => n6441
                           , ZN => n3657);
   U142 : OAI22_X1 port map( A1 => n6005, A2 => n1735, B1 => n1702, B2 => n6441
                           , ZN => n3668);
   U715 : OAI22_X1 port map( A1 => n6112, A2 => n1990, B1 => n1676, B2 => n1991
                           , ZN => n3329);
   U699 : OAI22_X1 port map( A1 => n6352, A2 => n6425, B1 => n1726, B2 => n1957
                           , ZN => n3336);
   U677 : OAI22_X1 port map( A1 => n6285, A2 => n6425, B1 => n1704, B2 => n1957
                           , ZN => n3347);
   U717 : OAI22_X1 port map( A1 => n6111, A2 => n1990, B1 => n1678, B2 => n1991
                           , ZN => n3328);
   U641 : OAI22_X1 port map( A1 => n6303, A2 => n6425, B1 => n1668, B2 => n1957
                           , ZN => n3365);
   U639 : OAI22_X1 port map( A1 => n6304, A2 => n1956, B1 => n1666, B2 => n1957
                           , ZN => n3366);
   U681 : OAI22_X1 port map( A1 => n6283, A2 => n6425, B1 => n1708, B2 => n1957
                           , ZN => n3345);
   U689 : OAI22_X1 port map( A1 => n6279, A2 => n6425, B1 => n1716, B2 => n1957
                           , ZN => n3341);
   U691 : OAI22_X1 port map( A1 => n6278, A2 => n6425, B1 => n1718, B2 => n1957
                           , ZN => n3340);
   U679 : OAI22_X1 port map( A1 => n6284, A2 => n6425, B1 => n1706, B2 => n1957
                           , ZN => n3346);
   U705 : OAI22_X1 port map( A1 => n6117, A2 => n1990, B1 => n1666, B2 => n1991
                           , ZN => n3334);
   U713 : OAI22_X1 port map( A1 => n6113, A2 => n6423, B1 => n1674, B2 => n1991
                           , ZN => n3330);
   U709 : OAI22_X1 port map( A1 => n6115, A2 => n6423, B1 => n1670, B2 => n1991
                           , ZN => n3332);
   U711 : OAI22_X1 port map( A1 => n6114, A2 => n6423, B1 => n1672, B2 => n1991
                           , ZN => n3331);
   U743 : OAI22_X1 port map( A1 => n6098, A2 => n6423, B1 => n1704, B2 => n1991
                           , ZN => n3315);
   U745 : OAI22_X1 port map( A1 => n6097, A2 => n6423, B1 => n1706, B2 => n1991
                           , ZN => n3314);
   U747 : OAI22_X1 port map( A1 => n6096, A2 => n6423, B1 => n1708, B2 => n1991
                           , ZN => n3313);
   U765 : OAI22_X1 port map( A1 => n6087, A2 => n6423, B1 => n1726, B2 => n1991
                           , ZN => n3304);
   U643 : OAI22_X1 port map( A1 => n6302, A2 => n6425, B1 => n1670, B2 => n1957
                           , ZN => n3364);
   U651 : OAI22_X1 port map( A1 => n6298, A2 => n1956, B1 => n1678, B2 => n1957
                           , ZN => n3360);
   U755 : OAI22_X1 port map( A1 => n6092, A2 => n6423, B1 => n1716, B2 => n1991
                           , ZN => n3309);
   U757 : OAI22_X1 port map( A1 => n6091, A2 => n6423, B1 => n1718, B2 => n1991
                           , ZN => n3308);
   U649 : OAI22_X1 port map( A1 => n6299, A2 => n1956, B1 => n1676, B2 => n1957
                           , ZN => n3361);
   U647 : OAI22_X1 port map( A1 => n6300, A2 => n6425, B1 => n1674, B2 => n1957
                           , ZN => n3362);
   U645 : OAI22_X1 port map( A1 => n6301, A2 => n6425, B1 => n1672, B2 => n1957
                           , ZN => n3363);
   U637 : OAI22_X1 port map( A1 => n6305, A2 => n1956, B1 => n1663, B2 => n1957
                           , ZN => n3367);
   U707 : OAI22_X1 port map( A1 => n6116, A2 => n6423, B1 => n1668, B2 => n1991
                           , ZN => n3333);
   U703 : OAI22_X1 port map( A1 => n6118, A2 => n1990, B1 => n1663, B2 => n1991
                           , ZN => n3335);
   U613 : OAI22_X1 port map( A1 => n4913, A2 => n6427, B1 => n1706, B2 => n1922
                           , ZN => n3378);
   U573 : OAI22_X1 port map( A1 => n4989, A2 => n1921, B1 => n1666, B2 => n1922
                           , ZN => n3398);
   U575 : OAI22_X1 port map( A1 => n4988, A2 => n6427, B1 => n1668, B2 => n1922
                           , ZN => n3397);
   U623 : OAI22_X1 port map( A1 => n4898, A2 => n6427, B1 => n1716, B2 => n1922
                           , ZN => n3373);
   U611 : OAI22_X1 port map( A1 => n4922, A2 => n6427, B1 => n1704, B2 => n1922
                           , ZN => n3379);
   U585 : OAI22_X1 port map( A1 => n4964, A2 => n1921, B1 => n1678, B2 => n1922
                           , ZN => n3392);
   U625 : OAI22_X1 port map( A1 => n4893, A2 => n6427, B1 => n1718, B2 => n1922
                           , ZN => n3372);
   U615 : OAI22_X1 port map( A1 => n4905, A2 => n6427, B1 => n1708, B2 => n1922
                           , ZN => n3377);
   U579 : OAI22_X1 port map( A1 => n4982, A2 => n6427, B1 => n1672, B2 => n1922
                           , ZN => n3395);
   U577 : OAI22_X1 port map( A1 => n4983, A2 => n6427, B1 => n1670, B2 => n1922
                           , ZN => n3396);
   U633 : OAI22_X1 port map( A1 => n6342, A2 => n6427, B1 => n1726, B2 => n1922
                           , ZN => n3368);
   U583 : OAI22_X1 port map( A1 => n4965, A2 => n1921, B1 => n1676, B2 => n1922
                           , ZN => n3393);
   U571 : OAI22_X1 port map( A1 => n4993, A2 => n1921, B1 => n1663, B2 => n1922
                           , ZN => n3399);
   U581 : OAI22_X1 port map( A1 => n4973, A2 => n6427, B1 => n1674, B2 => n1922
                           , ZN => n3394);
   U1225 : OAI22_X1 port map( A1 => n694, A2 => n6406, B1 => n3887, B2 => n1708
                           , ZN => n3025);
   U1224 : OAI22_X1 port map( A1 => n693, A2 => n6406, B1 => n3887, B2 => n1706
                           , ZN => n3026);
   U1233 : OAI22_X1 port map( A1 => n702, A2 => n6406, B1 => n3887, B2 => n1724
                           , ZN => n3017);
   U1232 : OAI22_X1 port map( A1 => n701, A2 => n6406, B1 => n3887, B2 => n1722
                           , ZN => n3018);
   U1207 : OAI22_X1 port map( A1 => n676, A2 => n6406, B1 => n3887, B2 => n1672
                           , ZN => n3043);
   U1205 : OAI22_X1 port map( A1 => n674, A2 => n6406, B1 => n3887, B2 => n1668
                           , ZN => n3045);
   U1223 : OAI22_X1 port map( A1 => n692, A2 => n6406, B1 => n3887, B2 => n1704
                           , ZN => n3027);
   U1227 : OAI22_X1 port map( A1 => n696, A2 => n6406, B1 => n3887, B2 => n1712
                           , ZN => n3023);
   U1231 : OAI22_X1 port map( A1 => n700, A2 => n6406, B1 => n3887, B2 => n1720
                           , ZN => n3019);
   U1230 : OAI22_X1 port map( A1 => n699, A2 => n6406, B1 => n3887, B2 => n1718
                           , ZN => n3020);
   U1229 : OAI22_X1 port map( A1 => n698, A2 => n6406, B1 => n3887, B2 => n1716
                           , ZN => n3021);
   U1226 : OAI22_X1 port map( A1 => n695, A2 => n6406, B1 => n3887, B2 => n1710
                           , ZN => n3024);
   U1228 : OAI22_X1 port map( A1 => n697, A2 => n6406, B1 => n3887, B2 => n1714
                           , ZN => n3022);
   U2448 : OAI22_X1 port map( A1 => n2087, A2 => n6392, B1 => n4181, B2 => 
                           n1726, ZN => n2729);
   U1770 : OAI22_X1 port map( A1 => n4509, A2 => n4180, B1 => n1674, B2 => 
                           n4181, ZN => n2781);
   U2420 : OAI22_X1 port map( A1 => n4418, A2 => n6392, B1 => n1724, B2 => 
                           n4181, ZN => n2731);
   U1874 : OAI22_X1 port map( A1 => n4493, A2 => n6392, B1 => n1682, B2 => 
                           n4181, ZN => n2773);
   U1744 : OAI22_X1 port map( A1 => n4513, A2 => n6392, B1 => n1672, B2 => 
                           n4181, ZN => n2783);
   U1640 : OAI22_X1 port map( A1 => n4532, A2 => n4180, B1 => n1663, B2 => 
                           n4181, ZN => n2791);
   U2264 : OAI22_X1 port map( A1 => n4442, A2 => n6392, B1 => n1712, B2 => 
                           n4181, ZN => n2743);
   U1900 : OAI22_X1 port map( A1 => n4485, A2 => n6392, B1 => n1684, B2 => 
                           n4181, ZN => n2771);
   U1926 : OAI22_X1 port map( A1 => n4484, A2 => n6392, B1 => n1686, B2 => 
                           n4181, ZN => n2769);
   U2316 : OAI22_X1 port map( A1 => n4425, A2 => n6392, B1 => n1716, B2 => 
                           n4181, ZN => n2739);
   U2394 : OAI22_X1 port map( A1 => n4419, A2 => n6392, B1 => n1722, B2 => 
                           n4181, ZN => n2733);
   U2290 : OAI22_X1 port map( A1 => n4433, A2 => n6392, B1 => n1714, B2 => 
                           n4181, ZN => n2741);
   U2368 : OAI22_X1 port map( A1 => n4423, A2 => n6392, B1 => n1720, B2 => 
                           n4181, ZN => n2735);
   U2342 : OAI22_X1 port map( A1 => n4424, A2 => n6392, B1 => n1718, B2 => 
                           n4181, ZN => n2737);
   U1627 : OAI22_X1 port map( A1 => n6184, A2 => n6394, B1 => n1718, B2 => 
                           n4146, ZN => n2796);
   U1583 : OAI22_X1 port map( A1 => n6206, A2 => n4145, B1 => n1674, B2 => 
                           n4146, ZN => n2818);
   U1587 : OAI22_X1 port map( A1 => n6204, A2 => n4145, B1 => n1678, B2 => 
                           n4146, ZN => n2816);
   U1617 : OAI22_X1 port map( A1 => n6189, A2 => n6394, B1 => n1708, B2 => 
                           n4146, ZN => n2801);
   U1615 : OAI22_X1 port map( A1 => n6190, A2 => n6394, B1 => n1706, B2 => 
                           n4146, ZN => n2802);
   U1573 : OAI22_X1 port map( A1 => n6211, A2 => n4145, B1 => n1663, B2 => 
                           n4146, ZN => n2823);
   U1625 : OAI22_X1 port map( A1 => n6185, A2 => n6394, B1 => n1716, B2 => 
                           n4146, ZN => n2797);
   U1577 : OAI22_X1 port map( A1 => n6209, A2 => n6394, B1 => n1668, B2 => 
                           n4146, ZN => n2821);
   U1581 : OAI22_X1 port map( A1 => n6207, A2 => n6394, B1 => n1672, B2 => 
                           n4146, ZN => n2819);
   U1635 : OAI22_X1 port map( A1 => n6347, A2 => n6394, B1 => n1726, B2 => 
                           n4146, ZN => n2792);
   U1579 : OAI22_X1 port map( A1 => n6208, A2 => n6394, B1 => n1670, B2 => 
                           n4146, ZN => n2820);
   U1633 : OAI22_X1 port map( A1 => n6181, A2 => n6394, B1 => n1724, B2 => 
                           n4146, ZN => n2793);
   U1585 : OAI22_X1 port map( A1 => n6205, A2 => n6394, B1 => n1676, B2 => 
                           n4146, ZN => n2817);
   U1575 : OAI22_X1 port map( A1 => n6210, A2 => n4145, B1 => n1666, B2 => 
                           n4146, ZN => n2822);
   U1195 : OAI22_X1 port map( A1 => n541, A2 => n6408, B1 => n3995, B2 => n1716
                           , ZN => n3053);
   U1190 : OAI22_X1 port map( A1 => n536, A2 => n6408, B1 => n3995, B2 => n1706
                           , ZN => n3058);
   U1170 : OAI22_X1 port map( A1 => n516, A2 => n3994, B1 => n3995, B2 => n1666
                           , ZN => n3078);
   U1200 : OAI22_X1 port map( A1 => n671, A2 => n6408, B1 => n3995, B2 => n1726
                           , ZN => n3048);
   U1173 : OAI22_X1 port map( A1 => n519, A2 => n6408, B1 => n3995, B2 => n1672
                           , ZN => n3075);
   U1174 : OAI22_X1 port map( A1 => n520, A2 => n6408, B1 => n3995, B2 => n1674
                           , ZN => n3074);
   U1199 : OAI22_X1 port map( A1 => n545, A2 => n6408, B1 => n3995, B2 => n1724
                           , ZN => n3049);
   U1171 : OAI22_X1 port map( A1 => n517, A2 => n6408, B1 => n3995, B2 => n1668
                           , ZN => n3077);
   U1172 : OAI22_X1 port map( A1 => n518, A2 => n6408, B1 => n3995, B2 => n1670
                           , ZN => n3076);
   U1196 : OAI22_X1 port map( A1 => n542, A2 => n6408, B1 => n3995, B2 => n1718
                           , ZN => n3052);
   U1191 : OAI22_X1 port map( A1 => n537, A2 => n6408, B1 => n3995, B2 => n1708
                           , ZN => n3057);
   U1176 : OAI22_X1 port map( A1 => n522, A2 => n3994, B1 => n3995, B2 => n1678
                           , ZN => n3072);
   U1169 : OAI22_X1 port map( A1 => n515, A2 => n3994, B1 => n3995, B2 => n1663
                           , ZN => n3079);
   U1175 : OAI22_X1 port map( A1 => n521, A2 => n3994, B1 => n3995, B2 => n1676
                           , ZN => n3073);
   U773 : OAI22_X1 port map( A1 => n708, A2 => n6421, B1 => n2024, B2 => n1672,
                           ZN => n3299);
   U791 : OAI22_X1 port map( A1 => n726, A2 => n6421, B1 => n2024, B2 => n1708,
                           ZN => n3281);
   U790 : OAI22_X1 port map( A1 => n725, A2 => n6421, B1 => n2024, B2 => n1706,
                           ZN => n3282);
   U770 : OAI22_X1 port map( A1 => n705, A2 => n2023, B1 => n2024, B2 => n1666,
                           ZN => n3302);
   U776 : OAI22_X1 port map( A1 => n711, A2 => n2023, B1 => n2024, B2 => n1678,
                           ZN => n3296);
   U795 : OAI22_X1 port map( A1 => n730, A2 => n6421, B1 => n2024, B2 => n1716,
                           ZN => n3277);
   U774 : OAI22_X1 port map( A1 => n709, A2 => n6421, B1 => n2024, B2 => n1674,
                           ZN => n3298);
   U772 : OAI22_X1 port map( A1 => n707, A2 => n6421, B1 => n2024, B2 => n1670,
                           ZN => n3300);
   U771 : OAI22_X1 port map( A1 => n706, A2 => n6421, B1 => n2024, B2 => n1668,
                           ZN => n3301);
   U796 : OAI22_X1 port map( A1 => n731, A2 => n6421, B1 => n2024, B2 => n1718,
                           ZN => n3276);
   U769 : OAI22_X1 port map( A1 => n704, A2 => n2023, B1 => n2024, B2 => n1663,
                           ZN => n3303);
   U799 : OAI22_X1 port map( A1 => n734, A2 => n6421, B1 => n2024, B2 => n1724,
                           ZN => n3273);
   U800 : OAI22_X1 port map( A1 => n513, A2 => n6421, B1 => n2024, B2 => n1726,
                           ZN => n3272);
   U775 : OAI22_X1 port map( A1 => n710, A2 => n2023, B1 => n2024, B2 => n1676,
                           ZN => n3297);
   U1129 : OAI22_X1 port map( A1 => n4713, A2 => n6410, B1 => n1690, B2 => 
                           n3962, ZN => n3098);
   U1121 : OAI22_X1 port map( A1 => n4724, A2 => n6410, B1 => n1682, B2 => 
                           n3962, ZN => n3102);
   U1103 : OAI22_X1 port map( A1 => n4755, A2 => n3961, B1 => n1663, B2 => 
                           n3962, ZN => n3111);
   U1107 : OAI22_X1 port map( A1 => n4753, A2 => n6410, B1 => n1668, B2 => 
                           n3962, ZN => n3109);
   U1117 : OAI22_X1 port map( A1 => n4733, A2 => n3961, B1 => n1678, B2 => 
                           n3962, ZN => n3104);
   U1133 : OAI22_X1 port map( A1 => n4703, A2 => n6410, B1 => n1694, B2 => 
                           n3962, ZN => n3096);
   U1141 : OAI22_X1 port map( A1 => n4689, A2 => n6410, B1 => n1702, B2 => 
                           n3962, ZN => n3092);
   U1123 : OAI22_X1 port map( A1 => n4723, A2 => n6410, B1 => n1684, B2 => 
                           n3962, ZN => n3101);
   U1105 : OAI22_X1 port map( A1 => n4754, A2 => n3961, B1 => n1666, B2 => 
                           n3962, ZN => n3110);
   U1115 : OAI22_X1 port map( A1 => n4742, A2 => n3961, B1 => n1676, B2 => 
                           n3962, ZN => n3105);
   U1131 : OAI22_X1 port map( A1 => n4712, A2 => n6410, B1 => n1692, B2 => 
                           n3962, ZN => n3097);
   U1119 : OAI22_X1 port map( A1 => n4725, A2 => n3961, B1 => n1680, B2 => 
                           n3962, ZN => n3103);
   U1111 : OAI22_X1 port map( A1 => n4748, A2 => n6410, B1 => n1672, B2 => 
                           n3962, ZN => n3107);
   U1474 : OAI22_X1 port map( A1 => n548, A2 => n6398, B1 => n4107, B2 => n1668
                           , ZN => n2885);
   U1473 : OAI22_X1 port map( A1 => n547, A2 => n6398, B1 => n4107, B2 => n1666
                           , ZN => n2886);
   U1475 : OAI22_X1 port map( A1 => n549, A2 => n6398, B1 => n4107, B2 => n1670
                           , ZN => n2884);
   U1498 : OAI22_X1 port map( A1 => n572, A2 => n6398, B1 => n4107, B2 => n1716
                           , ZN => n2861);
   U1477 : OAI22_X1 port map( A1 => n551, A2 => n6398, B1 => n4107, B2 => n1674
                           , ZN => n2882);
   U1497 : OAI22_X1 port map( A1 => n571, A2 => n6398, B1 => n4107, B2 => n1714
                           , ZN => n2862);
   U1503 : OAI22_X1 port map( A1 => n703, A2 => n6398, B1 => n4107, B2 => n1726
                           , ZN => n2856);
   U1479 : OAI22_X1 port map( A1 => n553, A2 => n4106, B1 => n4107, B2 => n1678
                           , ZN => n2880);
   U1492 : OAI22_X1 port map( A1 => n566, A2 => n4106, B1 => n4107, B2 => n1704
                           , ZN => n2867);
   U1472 : OAI22_X1 port map( A1 => n546, A2 => n4106, B1 => n4107, B2 => n1663
                           , ZN => n2887);
   U1476 : OAI22_X1 port map( A1 => n550, A2 => n6398, B1 => n4107, B2 => n1672
                           , ZN => n2883);
   U1494 : OAI22_X1 port map( A1 => n568, A2 => n6398, B1 => n4107, B2 => n1708
                           , ZN => n2865);
   U1493 : OAI22_X1 port map( A1 => n567, A2 => n6398, B1 => n4107, B2 => n1706
                           , ZN => n2866);
   U1478 : OAI22_X1 port map( A1 => n552, A2 => n4106, B1 => n4107, B2 => n1676
                           , ZN => n2881);
   U1017 : OAI22_X1 port map( A1 => n6063, A2 => n3892, B1 => n1710, B2 => 
                           n6413, ZN => n3152);
   U1009 : OAI22_X1 port map( A1 => n6067, A2 => n6414, B1 => n1702, B2 => 
                           n6413, ZN => n3156);
   U1007 : OAI22_X1 port map( A1 => n6068, A2 => n6414, B1 => n1700, B2 => 
                           n6413, ZN => n3157);
   U973 : OAI22_X1 port map( A1 => n6085, A2 => n6414, B1 => n1666, B2 => n6413
                           , ZN => n3174);
   U1015 : OAI22_X1 port map( A1 => n6064, A2 => n3892, B1 => n1708, B2 => 
                           n6413, ZN => n3153);
   U1013 : OAI22_X1 port map( A1 => n6065, A2 => n3892, B1 => n1706, B2 => 
                           n6413, ZN => n3154);
   U1005 : OAI22_X1 port map( A1 => n6069, A2 => n6414, B1 => n1698, B2 => 
                           n6413, ZN => n3158);
   U999 : OAI22_X1 port map( A1 => n6072, A2 => n6414, B1 => n1692, B2 => n6413
                           , ZN => n3161);
   U997 : OAI22_X1 port map( A1 => n6073, A2 => n6414, B1 => n1690, B2 => n6413
                           , ZN => n3162);
   U995 : OAI22_X1 port map( A1 => n6074, A2 => n6414, B1 => n1688, B2 => n6413
                           , ZN => n3163);
   U1003 : OAI22_X1 port map( A1 => n6070, A2 => n6414, B1 => n1696, B2 => 
                           n6413, ZN => n3159);
   U1001 : OAI22_X1 port map( A1 => n6071, A2 => n6414, B1 => n1694, B2 => 
                           n6413, ZN => n3160);
   U985 : OAI22_X1 port map( A1 => n6079, A2 => n6414, B1 => n1678, B2 => n6413
                           , ZN => n3168);
   U983 : OAI22_X1 port map( A1 => n6080, A2 => n6414, B1 => n1676, B2 => n6413
                           , ZN => n3169);
   U977 : OAI22_X1 port map( A1 => n6083, A2 => n6414, B1 => n1670, B2 => n6413
                           , ZN => n3172);
   U1011 : OAI22_X1 port map( A1 => n6066, A2 => n6414, B1 => n1704, B2 => 
                           n6413, ZN => n3155);
   U975 : OAI22_X1 port map( A1 => n6084, A2 => n6414, B1 => n1668, B2 => n6413
                           , ZN => n3173);
   U1033 : OAI22_X1 port map( A1 => n514, A2 => n6414, B1 => n6413, B2 => n1726
                           , ZN => n3144);
   U943 : OAI22_X1 port map( A1 => n647, A2 => n3888, B1 => n3884, B2 => n1678,
                           ZN => n3200);
   U953 : OAI22_X1 port map( A1 => n657, A2 => n3888, B1 => n3884, B2 => n1698,
                           ZN => n3190);
   U950 : OAI22_X1 port map( A1 => n654, A2 => n3888, B1 => n3884, B2 => n1692,
                           ZN => n3193);
   U941 : OAI22_X1 port map( A1 => n645, A2 => n3888, B1 => n3884, B2 => n1674,
                           ZN => n3202);
   U954 : OAI22_X1 port map( A1 => n658, A2 => n3888, B1 => n3884, B2 => n1700,
                           ZN => n3189);
   U949 : OAI22_X1 port map( A1 => n653, A2 => n3888, B1 => n3884, B2 => n1690,
                           ZN => n3194);
   U955 : OAI22_X1 port map( A1 => n659, A2 => n3888, B1 => n3884, B2 => n1702,
                           ZN => n3188);
   U951 : OAI22_X1 port map( A1 => n655, A2 => n6415, B1 => n3884, B2 => n1694,
                           ZN => n3192);
   U946 : OAI22_X1 port map( A1 => n650, A2 => n6415, B1 => n3884, B2 => n1684,
                           ZN => n3197);
   U947 : OAI22_X1 port map( A1 => n651, A2 => n3888, B1 => n3884, B2 => n1686,
                           ZN => n3196);
   U944 : OAI22_X1 port map( A1 => n648, A2 => n3888, B1 => n3884, B2 => n1680,
                           ZN => n3199);
   U945 : OAI22_X1 port map( A1 => n649, A2 => n3888, B1 => n3884, B2 => n1682,
                           ZN => n3198);
   U948 : OAI22_X1 port map( A1 => n652, A2 => n3888, B1 => n3884, B2 => n1688,
                           ZN => n3195);
   U952 : OAI22_X1 port map( A1 => n656, A2 => n6415, B1 => n3884, B2 => n1696,
                           ZN => n3191);
   U967 : OAI22_X1 port map( A1 => n6337, A2 => n6415, B1 => n1726, B2 => n3884
                           , ZN => n3176);
   U81 : OAI22_X1 port map( A1 => n589, A2 => n1730, B1 => n3885, B2 => n1688, 
                           ZN => n3707);
   U84 : OAI22_X1 port map( A1 => n592, A2 => n1730, B1 => n3885, B2 => n1694, 
                           ZN => n3704);
   U85 : OAI22_X1 port map( A1 => n593, A2 => n1730, B1 => n3885, B2 => n1696, 
                           ZN => n3703);
   U78 : OAI22_X1 port map( A1 => n586, A2 => n1730, B1 => n3885, B2 => n1682, 
                           ZN => n3710);
   U83 : OAI22_X1 port map( A1 => n591, A2 => n1730, B1 => n3885, B2 => n1692, 
                           ZN => n3705);
   U80 : OAI22_X1 port map( A1 => n588, A2 => n1730, B1 => n3885, B2 => n1686, 
                           ZN => n3708);
   U74 : OAI22_X1 port map( A1 => n582, A2 => n1730, B1 => n3885, B2 => n1674, 
                           ZN => n3714);
   U88 : OAI22_X1 port map( A1 => n596, A2 => n6443, B1 => n3885, B2 => n1702, 
                           ZN => n3700);
   U87 : OAI22_X1 port map( A1 => n595, A2 => n6443, B1 => n3885, B2 => n1700, 
                           ZN => n3701);
   U77 : OAI22_X1 port map( A1 => n585, A2 => n1730, B1 => n3885, B2 => n1680, 
                           ZN => n3711);
   U82 : OAI22_X1 port map( A1 => n590, A2 => n1730, B1 => n3885, B2 => n1690, 
                           ZN => n3706);
   U79 : OAI22_X1 port map( A1 => n587, A2 => n1730, B1 => n3885, B2 => n1684, 
                           ZN => n3709);
   U86 : OAI22_X1 port map( A1 => n594, A2 => n1730, B1 => n3885, B2 => n1698, 
                           ZN => n3702);
   U76 : OAI22_X1 port map( A1 => n584, A2 => n6443, B1 => n3885, B2 => n1678, 
                           ZN => n3712);
   U963 : OAI22_X1 port map( A1 => n667, A2 => n6415, B1 => n3884, B2 => n1718,
                           ZN => n3180);
   U958 : OAI22_X1 port map( A1 => n662, A2 => n6415, B1 => n3884, B2 => n1708,
                           ZN => n3185);
   U961 : OAI22_X1 port map( A1 => n665, A2 => n6415, B1 => n3884, B2 => n1714,
                           ZN => n3182);
   U962 : OAI22_X1 port map( A1 => n666, A2 => n6415, B1 => n3884, B2 => n1716,
                           ZN => n3181);
   U956 : OAI22_X1 port map( A1 => n660, A2 => n6415, B1 => n3884, B2 => n1704,
                           ZN => n3187);
   U966 : OAI22_X1 port map( A1 => n670, A2 => n6415, B1 => n3884, B2 => n1724,
                           ZN => n3177);
   U957 : OAI22_X1 port map( A1 => n661, A2 => n6415, B1 => n3884, B2 => n1706,
                           ZN => n3186);
   U964 : OAI22_X1 port map( A1 => n668, A2 => n6415, B1 => n3884, B2 => n1720,
                           ZN => n3179);
   U959 : OAI22_X1 port map( A1 => n663, A2 => n6415, B1 => n3884, B2 => n1710,
                           ZN => n3184);
   U940 : OAI22_X1 port map( A1 => n644, A2 => n6415, B1 => n3884, B2 => n1672,
                           ZN => n3203);
   U960 : OAI22_X1 port map( A1 => n664, A2 => n6415, B1 => n3884, B2 => n1712,
                           ZN => n3183);
   U965 : OAI22_X1 port map( A1 => n669, A2 => n6415, B1 => n3884, B2 => n1722,
                           ZN => n3178);
   U100 : OAI22_X1 port map( A1 => n6345, A2 => n6443, B1 => n1726, B2 => n3885
                           , ZN => n3688);
   U73 : OAI22_X1 port map( A1 => n581, A2 => n6443, B1 => n3885, B2 => n1672, 
                           ZN => n3715);
   U98 : OAI22_X1 port map( A1 => n606, A2 => n6443, B1 => n3885, B2 => n1722, 
                           ZN => n3690);
   U90 : OAI22_X1 port map( A1 => n598, A2 => n6443, B1 => n3885, B2 => n1706, 
                           ZN => n3698);
   U95 : OAI22_X1 port map( A1 => n603, A2 => n6443, B1 => n3885, B2 => n1716, 
                           ZN => n3693);
   U96 : OAI22_X1 port map( A1 => n604, A2 => n6443, B1 => n3885, B2 => n1718, 
                           ZN => n3692);
   U89 : OAI22_X1 port map( A1 => n597, A2 => n6443, B1 => n3885, B2 => n1704, 
                           ZN => n3699);
   U94 : OAI22_X1 port map( A1 => n602, A2 => n6443, B1 => n3885, B2 => n1714, 
                           ZN => n3694);
   U97 : OAI22_X1 port map( A1 => n605, A2 => n6443, B1 => n3885, B2 => n1720, 
                           ZN => n3691);
   U99 : OAI22_X1 port map( A1 => n607, A2 => n6443, B1 => n3885, B2 => n1724, 
                           ZN => n3689);
   U92 : OAI22_X1 port map( A1 => n600, A2 => n6443, B1 => n3885, B2 => n1710, 
                           ZN => n3696);
   U91 : OAI22_X1 port map( A1 => n599, A2 => n6443, B1 => n3885, B2 => n1708, 
                           ZN => n3697);
   U93 : OAI22_X1 port map( A1 => n601, A2 => n6443, B1 => n3885, B2 => n1712, 
                           ZN => n3695);
   U870 : OAI22_X1 port map( A1 => n4298, A2 => n2062, B1 => n1663, B2 => n2063
                           , ZN => n3239);
   U912 : OAI22_X1 port map( A1 => n4191, A2 => n6417, B1 => n1706, B2 => n2063
                           , ZN => n3218);
   U910 : OAI22_X1 port map( A1 => n4193, A2 => n6417, B1 => n1704, B2 => n2063
                           , ZN => n3219);
   U922 : OAI22_X1 port map( A1 => n4174, A2 => n6417, B1 => n1716, B2 => n2063
                           , ZN => n3213);
   U872 : OAI22_X1 port map( A1 => n4293, A2 => n2062, B1 => n1666, B2 => n2063
                           , ZN => n3238);
   U874 : OAI22_X1 port map( A1 => n4292, A2 => n2062, B1 => n1668, B2 => n2063
                           , ZN => n3237);
   U932 : OAI22_X1 port map( A1 => n4168, A2 => n6417, B1 => n1726, B2 => n2063
                           , ZN => n3208);
   U882 : OAI22_X1 port map( A1 => n4273, A2 => n2062, B1 => n1676, B2 => n2063
                           , ZN => n3233);
   U916 : OAI22_X1 port map( A1 => n4177, A2 => n6417, B1 => n1710, B2 => n2063
                           , ZN => n3216);
   U914 : OAI22_X1 port map( A1 => n4179, A2 => n6417, B1 => n1708, B2 => n2063
                           , ZN => n3217);
   U876 : OAI22_X1 port map( A1 => n4283, A2 => n2062, B1 => n1670, B2 => n2063
                           , ZN => n3236);
   U924 : OAI22_X1 port map( A1 => n4173, A2 => n6417, B1 => n1718, B2 => n2063
                           , ZN => n3212);
   U880 : OAI22_X1 port map( A1 => n4274, A2 => n2062, B1 => n1674, B2 => n2063
                           , ZN => n3234);
   U878 : OAI22_X1 port map( A1 => n4275, A2 => n2062, B1 => n1672, B2 => n2063
                           , ZN => n3235);
   U844 : OAI22_X1 port map( A1 => n6254, A2 => n2027, B1 => n1704, B2 => n2028
                           , ZN => n3251);
   U850 : OAI22_X1 port map( A1 => n6251, A2 => n6419, B1 => n1710, B2 => n2028
                           , ZN => n3248);
   U848 : OAI22_X1 port map( A1 => n6252, A2 => n6419, B1 => n1708, B2 => n2028
                           , ZN => n3249);
   U846 : OAI22_X1 port map( A1 => n6253, A2 => n6419, B1 => n1706, B2 => n2028
                           , ZN => n3250);
   U816 : OAI22_X1 port map( A1 => n6268, A2 => n6419, B1 => n1676, B2 => n2028
                           , ZN => n3265);
   U814 : OAI22_X1 port map( A1 => n6269, A2 => n2027, B1 => n1674, B2 => n2028
                           , ZN => n3266);
   U812 : OAI22_X1 port map( A1 => n6270, A2 => n2027, B1 => n1672, B2 => n2028
                           , ZN => n3267);
   U866 : OAI22_X1 port map( A1 => n6351, A2 => n6419, B1 => n1726, B2 => n2028
                           , ZN => n3240);
   U808 : OAI22_X1 port map( A1 => n6272, A2 => n2027, B1 => n1668, B2 => n2028
                           , ZN => n3269);
   U806 : OAI22_X1 port map( A1 => n6273, A2 => n2027, B1 => n1666, B2 => n2028
                           , ZN => n3270);
   U804 : OAI22_X1 port map( A1 => n6274, A2 => n2027, B1 => n1663, B2 => n2028
                           , ZN => n3271);
   U856 : OAI22_X1 port map( A1 => n6248, A2 => n6419, B1 => n1716, B2 => n2028
                           , ZN => n3245);
   U858 : OAI22_X1 port map( A1 => n6247, A2 => n6419, B1 => n1718, B2 => n2028
                           , ZN => n3244);
   U810 : OAI22_X1 port map( A1 => n6271, A2 => n2027, B1 => n1670, B2 => n2028
                           , ZN => n3268);
   U110 : OAI22_X1 port map( A1 => n6021, A2 => n1735, B1 => n1670, B2 => n1736
                           , ZN => n3684);
   U144 : OAI22_X1 port map( A1 => n6004, A2 => n6442, B1 => n1704, B2 => n1736
                           , ZN => n3667);
   U158 : OAI22_X1 port map( A1 => n5997, A2 => n6442, B1 => n1718, B2 => n1736
                           , ZN => n3660);
   U156 : OAI22_X1 port map( A1 => n5998, A2 => n6442, B1 => n1716, B2 => n1736
                           , ZN => n3661);
   U146 : OAI22_X1 port map( A1 => n6003, A2 => n6442, B1 => n1706, B2 => n1736
                           , ZN => n3666);
   U116 : OAI22_X1 port map( A1 => n6018, A2 => n1735, B1 => n1676, B2 => n1736
                           , ZN => n3681);
   U166 : OAI22_X1 port map( A1 => n6354, A2 => n6442, B1 => n1726, B2 => n1736
                           , ZN => n3656);
   U150 : OAI22_X1 port map( A1 => n6001, A2 => n6442, B1 => n1710, B2 => n1736
                           , ZN => n3664);
   U148 : OAI22_X1 port map( A1 => n6002, A2 => n6442, B1 => n1708, B2 => n1736
                           , ZN => n3665);
   U108 : OAI22_X1 port map( A1 => n6022, A2 => n1735, B1 => n1668, B2 => n1736
                           , ZN => n3685);
   U106 : OAI22_X1 port map( A1 => n6023, A2 => n1735, B1 => n1666, B2 => n1736
                           , ZN => n3686);
   U114 : OAI22_X1 port map( A1 => n6019, A2 => n1735, B1 => n1674, B2 => n1736
                           , ZN => n3682);
   U112 : OAI22_X1 port map( A1 => n6020, A2 => n1735, B1 => n1672, B2 => n1736
                           , ZN => n3683);
   U104 : OAI22_X1 port map( A1 => n6024, A2 => n1735, B1 => n1663, B2 => n1736
                           , ZN => n3687);
   U1376 : OAI22_X1 port map( A1 => n2242, A2 => n6401, B1 => n4069, B2 => 
                           n1676, ZN => n2945);
   U1370 : OAI22_X1 port map( A1 => n2248, A2 => n4068, B1 => n4069, B2 => 
                           n1663, ZN => n2951);
   U1371 : OAI22_X1 port map( A1 => n2247, A2 => n4068, B1 => n4069, B2 => 
                           n1666, ZN => n2950);
   U372 : OAI22_X1 port map( A1 => n2664, A2 => n1847, B1 => n1848, B2 => n1663
                           , ZN => n3527);
   U373 : OAI22_X1 port map( A1 => n2663, A2 => n1847, B1 => n1848, B2 => n1666
                           , ZN => n3526);
   U378 : OAI22_X1 port map( A1 => n2658, A2 => n6434, B1 => n1848, B2 => n1676
                           , ZN => n3521);
   U338 : OAI22_X1 port map( A1 => n609, A2 => n1843, B1 => n1844, B2 => n1666,
                           ZN => n3558);
   U337 : OAI22_X1 port map( A1 => n608, A2 => n1843, B1 => n1844, B2 => n1663,
                           ZN => n3559);
   U343 : OAI22_X1 port map( A1 => n614, A2 => n6435, B1 => n1844, B2 => n1676,
                           ZN => n3553);
   U237 : OAI22_X1 port map( A1 => n3784, A2 => n1807, B1 => n1808, B2 => n1663
                           , ZN => n3623);
   U243 : OAI22_X1 port map( A1 => n3778, A2 => n6438, B1 => n1808, B2 => n1676
                           , ZN => n3617);
   U238 : OAI22_X1 port map( A1 => n3783, A2 => n1807, B1 => n1808, B2 => n1666
                           , ZN => n3622);
   U1204 : OAI22_X1 port map( A1 => n673, A2 => n3996, B1 => n3997, B2 => n1666
                           , ZN => n3046);
   U1209 : OAI22_X1 port map( A1 => n678, A2 => n6406, B1 => n3997, B2 => n1676
                           , ZN => n3041);
   U1203 : OAI22_X1 port map( A1 => n672, A2 => n3996, B1 => n3997, B2 => n1663
                           , ZN => n3047);
   U979 : OAI22_X1 port map( A1 => n6082, A2 => n6414, B1 => n1672, B2 => n3893
                           , ZN => n3171);
   U1021 : OAI22_X1 port map( A1 => n6061, A2 => n6414, B1 => n1714, B2 => 
                           n3893, ZN => n3150);
   U1031 : OAI22_X1 port map( A1 => n6056, A2 => n6414, B1 => n1724, B2 => 
                           n3893, ZN => n3145);
   U991 : OAI22_X1 port map( A1 => n6076, A2 => n6414, B1 => n1684, B2 => n3893
                           , ZN => n3165);
   U1025 : OAI22_X1 port map( A1 => n6059, A2 => n6414, B1 => n1718, B2 => 
                           n3893, ZN => n3148);
   U971 : OAI22_X1 port map( A1 => n6086, A2 => n6414, B1 => n1663, B2 => n3893
                           , ZN => n3175);
   U1019 : OAI22_X1 port map( A1 => n6062, A2 => n6414, B1 => n1712, B2 => 
                           n3893, ZN => n3151);
   U987 : OAI22_X1 port map( A1 => n6078, A2 => n6414, B1 => n1680, B2 => n3893
                           , ZN => n3167);
   U1027 : OAI22_X1 port map( A1 => n6058, A2 => n6414, B1 => n1720, B2 => 
                           n3893, ZN => n3147);
   U1029 : OAI22_X1 port map( A1 => n6057, A2 => n6414, B1 => n1722, B2 => 
                           n3893, ZN => n3146);
   U989 : OAI22_X1 port map( A1 => n6077, A2 => n6414, B1 => n1682, B2 => n3893
                           , ZN => n3166);
   U1023 : OAI22_X1 port map( A1 => n6060, A2 => n6414, B1 => n1716, B2 => 
                           n3893, ZN => n3149);
   U981 : OAI22_X1 port map( A1 => n6081, A2 => n6414, B1 => n1674, B2 => n3893
                           , ZN => n3170);
   U993 : OAI22_X1 port map( A1 => n6075, A2 => n6414, B1 => n1686, B2 => n3893
                           , ZN => n3164);
   U937 : OAI22_X1 port map( A1 => n641, A2 => n6415, B1 => n3889, B2 => n1666,
                           ZN => n3206);
   U939 : OAI22_X1 port map( A1 => n643, A2 => n6415, B1 => n3889, B2 => n1670,
                           ZN => n3204);
   U942 : OAI22_X1 port map( A1 => n646, A2 => n6415, B1 => n3889, B2 => n1676,
                           ZN => n3201);
   U936 : OAI22_X1 port map( A1 => n640, A2 => n6415, B1 => n3889, B2 => n1663,
                           ZN => n3207);
   U938 : OAI22_X1 port map( A1 => n642, A2 => n6415, B1 => n3889, B2 => n1668,
                           ZN => n3205);
   U72 : OAI22_X1 port map( A1 => n580, A2 => n6443, B1 => n1731, B2 => n1670, 
                           ZN => n3716);
   U75 : OAI22_X1 port map( A1 => n583, A2 => n6443, B1 => n1731, B2 => n1676, 
                           ZN => n3713);
   U70 : OAI22_X1 port map( A1 => n578, A2 => n6443, B1 => n1731, B2 => n1666, 
                           ZN => n3718);
   U71 : OAI22_X1 port map( A1 => n579, A2 => n6443, B1 => n1731, B2 => n1668, 
                           ZN => n3717);
   U69 : OAI22_X1 port map( A1 => n577, A2 => n6443, B1 => n1731, B2 => n1663, 
                           ZN => n3719);
   U3540 : NOR2_X2 port map( A1 => n5953, A2 => n5939, ZN => n5264);
   U3536 : NOR2_X2 port map( A1 => n5949, A2 => n5936, ZN => n5262);
   U3515 : NOR2_X2 port map( A1 => n5938, A2 => n5936, ZN => n5213);
   U3508 : NOR2_X2 port map( A1 => n5950, A2 => n5960, ZN => n5249);
   U3507 : NOR2_X2 port map( A1 => n5959, A2 => n5951, ZN => n5248);
   U3501 : NOR2_X2 port map( A1 => n5952, A2 => n5935, ZN => n5245);
   U3500 : NOR2_X2 port map( A1 => n5953, A2 => n5951, ZN => n5244);
   U3493 : NOR2_X2 port map( A1 => n5952, A2 => n5938, ZN => n5237);
   U3492 : NOR2_X2 port map( A1 => n5952, A2 => n5953, ZN => n5236);
   U2522 : NOR2_X2 port map( A1 => n5173, A2 => n5159, ZN => n4241);
   U2518 : NOR2_X2 port map( A1 => n5169, A2 => n5156, ZN => n4240);
   U2509 : NOR2_X2 port map( A1 => n5168, A2 => n5185, ZN => n4237);
   U2498 : NOR2_X2 port map( A1 => n5158, A2 => n5156, ZN => n4186);
   U2485 : NOR2_X2 port map( A1 => n5172, A2 => n5155, ZN => n4220);
   U3542 : NAND2_X1 port map( A1 => n5964, A2 => ADD_RD1(1), ZN => n5960);
   U3538 : NAND2_X1 port map( A1 => ADD_RD1(1), A2 => ADD_RD1(2), ZN => n5951);
   U3528 : NAND2_X1 port map( A1 => ADD_RD1(2), A2 => n5963, ZN => n5948);
   U2524 : NAND2_X1 port map( A1 => n5186, A2 => ADD_RD2(1), ZN => n5182);
   U2520 : NAND2_X1 port map( A1 => ADD_RD2(2), A2 => ADD_RD2(1), ZN => n5171);
   U2511 : NAND2_X1 port map( A1 => ADD_RD2(2), A2 => n5187, ZN => n5168);
   U3547 : NOR2_X1 port map( A1 => n5206, A2 => n5981, ZN => n5977);
   U3570 : NAND3_X1 port map( A1 => ADD_WR(3), A2 => ADD_WR(2), A3 => n1770, ZN
                           => n1954);
   U2454 : INV_X1 port map( A => WR, ZN => n2025);
   U3569 : NAND3_X1 port map( A1 => ADD_WR(3), A2 => n1770, A3 => n1919, ZN => 
                           n1850);
   U3568 : NAND3_X1 port map( A1 => ADD_WR(2), A2 => n1770, A3 => n1846, ZN => 
                           n1806);
   U3573 : NAND3_X1 port map( A1 => ADD_WR(3), A2 => ADD_WR(2), A3 => n3924, ZN
                           => n4108);
   U1036 : NAND2_X1 port map( A1 => n1769, A2 => n3924, ZN => n2060);
   U536 : OAI21_X1 port map( B1 => n1733, B2 => n1850, A => n6446, ZN => n1885)
                           ;
   U471 : OAI21_X1 port map( B1 => n1728, B2 => n1850, A => n6446, ZN => n1852)
                           ;
   U3572 : NAND3_X1 port map( A1 => ADD_WR(3), A2 => n3924, A3 => n1919, ZN => 
                           n4033);
   U570 : OAI21_X1 port map( B1 => n1768, B2 => n1850, A => n6446, ZN => n1917)
                           ;
   U3571 : NAND3_X1 port map( A1 => ADD_WR(2), A2 => n3924, A3 => n1846, ZN => 
                           n3959);
   U701 : OAI21_X1 port map( B1 => n1728, B2 => n1954, A => n6446, ZN => n1956)
                           ;
   U635 : OAI21_X1 port map( B1 => n1805, B2 => n1954, A => n6446, ZN => n1921)
                           ;
   U802 : OAI21_X1 port map( B1 => n1768, B2 => n1954, A => n6446, ZN => n2023)
                           ;
   U2453 : NOR2_X1 port map( A1 => n2025, A2 => n5146, ZN => n3924);
   U3560 : INV_X1 port map( A => ADD_RD1(0), ZN => n5966);
   U3563 : INV_X1 port map( A => ADD_RD1(3), ZN => n5971);
   U3566 : INV_X1 port map( A => ADD_RD1(1), ZN => n5963);
   U3567 : INV_X1 port map( A => ADD_RD1(4), ZN => n5967);
   U3543 : INV_X1 port map( A => ADD_RD1(2), ZN => n5964);
   U2535 : INV_X1 port map( A => ADD_RD2(2), ZN => n5186);
   U2521 : INV_X1 port map( A => ADD_RD2(3), ZN => n5194);
   U2533 : INV_X1 port map( A => ADD_RD2(1), ZN => n5187);
   U2538 : INV_X1 port map( A => ADD_RD2(4), ZN => n5190);
   U2537 : INV_X1 port map( A => ADD_RD2(0), ZN => n5189);
   U3551 : INV_X1 port map( A => ADD_WR(2), ZN => n1919);
   U2451 : OAI21_X1 port map( B1 => n1768, B2 => n4108, A => n6446, ZN => n4180
                           );
   U1637 : OAI21_X1 port map( B1 => n4108, B2 => n1733, A => n6446, ZN => n4145
                           );
   U336 : OAI21_X1 port map( B1 => n1733, B2 => n1806, A => n6446, ZN => n1811)
                           ;
   U1202 : OAI21_X1 port map( B1 => n1733, B2 => n3959, A => n6446, ZN => n3994
                           );
   U370 : OAI21_X1 port map( B1 => n1768, B2 => n1806, A => n6446, ZN => n1843)
                           ;
   U1236 : OAI21_X1 port map( B1 => n1768, B2 => n3959, A => n6446, ZN => n3996
                           );
   U1470 : OAI21_X1 port map( B1 => n1768, B2 => n4033, A => n6446, ZN => n4073
                           );
   U767 : OAI21_X1 port map( B1 => n1733, B2 => n1954, A => n6446, ZN => n1990)
                           ;
   U1404 : OAI21_X1 port map( B1 => n1733, B2 => n4033, A => n6446, ZN => n4068
                           );
   U1035 : OAI21_X1 port map( B1 => n1768, B2 => n2060, A => n6446, ZN => n3892
                           );
   U3556 : NAND2_X1 port map( A1 => n4143, A2 => n4178, ZN => n1805);
   U1167 : OAI21_X1 port map( B1 => n1728, B2 => n3959, A => n6446, ZN => n3961
                           );
   U235 : OAI21_X1 port map( B1 => n1805, B2 => n1806, A => n6446, ZN => n1772)
                           ;
   U1101 : OAI21_X1 port map( B1 => n1805, B2 => n3959, A => n6446, ZN => n3926
                           );
   U405 : OAI21_X1 port map( B1 => n1805, B2 => n1850, A => n6446, ZN => n1847)
                           ;
   U1505 : OAI21_X1 port map( B1 => n1805, B2 => n4108, A => n6446, ZN => n4106
                           );
   U3555 : INV_X1 port map( A => n1805, ZN => n5984);
   U1570 : OAI21_X1 port map( B1 => n4108, B2 => n1728, A => n6446, ZN => n4110
                           );
   U270 : OAI21_X1 port map( B1 => n1728, B2 => n1806, A => n6446, ZN => n1807)
                           ;
   U1368 : OAI21_X1 port map( B1 => n1728, B2 => n4033, A => n6446, ZN => n4035
                           );
   U67 : OAI21_X1 port map( B1 => n1728, B2 => n1729, A => n6446, ZN => n1662);
   U1302 : OAI21_X1 port map( B1 => n1805, B2 => n4033, A => n6446, ZN => n4000
                           );
   U2526 : AOI211_X1 port map( C1 => n5205, C2 => n5200, A => Rst, B => n5197, 
                           ZN => n4199);
   U3545 : AOI211_X1 port map( C1 => n5980, C2 => n5977, A => Rst, B => n5974, 
                           ZN => n5225);
   U2512 : INV_X2 port map( A => n5197, ZN => n4235);
   U2523 : OR2_X1 port map( A1 => n6387, A2 => n5182, ZN => n5159);
   U2497 : OR2_X1 port map( A1 => n6387, A2 => n5170, ZN => n5184);
   U2519 : OR2_X1 port map( A1 => n6387, A2 => n5171, ZN => n5156);
   U2510 : OR2_X1 port map( A1 => n6387, A2 => n5181, ZN => n5185);
   U3514 : OR2_X1 port map( A1 => n6371, A2 => n5950, ZN => n5961);
   U3541 : OR2_X1 port map( A1 => n6371, A2 => n5960, ZN => n5939);
   U3527 : OR2_X1 port map( A1 => n6371, A2 => n5959, ZN => n5962);
   U3537 : OR2_X1 port map( A1 => n6371, A2 => n5951, ZN => n5936);
   U3474 : NOR2_X1 port map( A1 => n5935, A2 => n5936, ZN => n5219);
   U2460 : NOR2_X1 port map( A1 => n5155, A2 => n5156, ZN => n4192);
   U3510 : NOR2_X1 port map( A1 => n5961, A2 => n5952, ZN => n5251);
   U3511 : NOR2_X1 port map( A1 => n5952, A2 => n5962, ZN => n5250);
   U2515 : NOR2_X1 port map( A1 => n5157, A2 => n5159, ZN => n4239);
   U3533 : NOR2_X1 port map( A1 => n5949, A2 => n5939, ZN => n5263);
   U2516 : NOR2_X1 port map( A1 => n5169, A2 => n5159, ZN => n4243);
   U3532 : NOR2_X1 port map( A1 => n5937, A2 => n5939, ZN => n5261);
   U3526 : NOR2_X1 port map( A1 => n5948, A2 => n5962, ZN => n5259);
   U2493 : NOR2_X1 port map( A1 => n5184, A2 => n5172, ZN => n4228);
   U2494 : NOR2_X1 port map( A1 => n5172, A2 => n5185, ZN => n4229);
   U4 : INV_X4 port map( A => n5142, ZN => n4233);
   U6 : INV_X4 port map( A => n5124, ZN => n4189);
   U8 : INV_X4 port map( A => n5910, ZN => n5216);
   U10 : INV_X4 port map( A => n5925, ZN => n5256);
   U12 : INV_X4 port map( A => Rst, ZN => n6446);
   U14 : BUF_X1 port map( A => n4243, Z => n6375);
   U16 : BUF_X2 port map( A => n4229, Z => n3880);
   U18 : BUF_X1 port map( A => n1664, Z => n6444);
   U20 : BUF_X1 port map( A => n1773, Z => n6439);
   U22 : BUF_X1 port map( A => n4111, Z => n6395);
   U24 : BUF_X1 port map( A => n4181, Z => n6391);
   U26 : BUF_X2 port map( A => n1848, Z => n3881);
   U28 : BUF_X1 port map( A => n1991, Z => n6422);
   U30 : BUF_X2 port map( A => n1808, Z => n3882);
   U32 : BUF_X1 port map( A => n4146, Z => n6393);
   U34 : BUF_X2 port map( A => n1844, Z => n3883);
   U36 : BUF_X2 port map( A => n3889, Z => n3884);
   U38 : BUF_X2 port map( A => n1731, Z => n3885);
   U40 : BUF_X2 port map( A => n4069, Z => n3886);
   U42 : BUF_X2 port map( A => n3997, Z => n3887);
   U44 : INV_X2 port map( A => DATAIN(6), ZN => n1714);
   U46 : INV_X2 port map( A => DATAIN(5), ZN => n1716);
   U48 : INV_X2 port map( A => DATAIN(26), ZN => n1674);
   U50 : INV_X2 port map( A => DATAIN(4), ZN => n1718);
   U52 : INV_X2 port map( A => DATAIN(3), ZN => n1720);
   U54 : INV_X2 port map( A => DATAIN(2), ZN => n1722);
   U56 : INV_X2 port map( A => DATAIN(1), ZN => n1724);
   U58 : INV_X2 port map( A => DATAIN(0), ZN => n1726);
   U60 : INV_X2 port map( A => DATAIN(27), ZN => n1672);
   U62 : INV_X2 port map( A => DATAIN(28), ZN => n1670);
   U64 : INV_X2 port map( A => DATAIN(29), ZN => n1668);
   U66 : INV_X2 port map( A => DATAIN(21), ZN => n1684);
   U68 : INV_X2 port map( A => DATAIN(20), ZN => n1686);
   U101 : INV_X2 port map( A => DATAIN(19), ZN => n1688);
   U102 : INV_X2 port map( A => DATAIN(18), ZN => n1690);
   U103 : INV_X2 port map( A => DATAIN(22), ZN => n1682);
   U105 : INV_X2 port map( A => DATAIN(17), ZN => n1692);
   U107 : INV_X2 port map( A => DATAIN(16), ZN => n1694);
   U109 : INV_X2 port map( A => DATAIN(15), ZN => n1696);
   U111 : INV_X2 port map( A => DATAIN(23), ZN => n1680);
   U113 : INV_X2 port map( A => DATAIN(14), ZN => n1698);
   U115 : INV_X2 port map( A => DATAIN(13), ZN => n1700);
   U117 : INV_X2 port map( A => DATAIN(24), ZN => n1678);
   U119 : INV_X2 port map( A => DATAIN(12), ZN => n1702);
   U121 : INV_X2 port map( A => DATAIN(11), ZN => n1704);
   U123 : INV_X2 port map( A => DATAIN(10), ZN => n1706);
   U125 : INV_X2 port map( A => DATAIN(9), ZN => n1708);
   U127 : INV_X2 port map( A => DATAIN(8), ZN => n1710);
   U129 : INV_X2 port map( A => DATAIN(7), ZN => n1712);
   U131 : INV_X2 port map( A => DATAIN(25), ZN => n1676);
   U133 : INV_X2 port map( A => DATAIN(31), ZN => n1663);
   U135 : INV_X2 port map( A => DATAIN(30), ZN => n1666);
   U137 : BUF_X1 port map( A => n4221, Z => n3891);
   U139 : BUF_X1 port map( A => n4212, Z => n3903);
   U141 : BUF_X2 port map( A => n5259, Z => n6360);
   U143 : BUF_X2 port map( A => n5250, Z => n6363);
   U145 : BUF_X2 port map( A => n5261, Z => n6358);
   U147 : BUF_X2 port map( A => n5263, Z => n6356);
   U149 : BUF_X2 port map( A => n4239, Z => n6378);
   U151 : OR2_X1 port map( A1 => n5155, A2 => n5159, ZN => n3950);
   U153 : OR2_X1 port map( A1 => n5935, A2 => n5939, ZN => n3952);
   U155 : OR2_X1 port map( A1 => n5938, A2 => n5939, ZN => n3953);
   U157 : OR2_X1 port map( A1 => n5158, A2 => n5159, ZN => n3951);
   U159 : INV_X1 port map( A => n4199, ZN => n6387);
   U161 : INV_X1 port map( A => n5225, ZN => n6371);
   U163 : NOR2_X1 port map( A1 => ENABLE, A2 => Rst, ZN => n5197);
   U165 : NOR2_X1 port map( A1 => ENABLE, A2 => Rst, ZN => n5974);
   U167 : BUF_X1 port map( A => n4036, Z => n6402);
   U168 : BUF_X1 port map( A => n4001, Z => n6404);
   U170 : BUF_X1 port map( A => n2063, Z => n6416);
   U172 : BUF_X1 port map( A => n4107, Z => n6397);
   U174 : BUF_X1 port map( A => n3962, Z => n6409);
   U176 : BUF_X1 port map( A => n3927, Z => n6411);
   U178 : BUF_X1 port map( A => n4074, Z => n6399);
   U180 : NAND2_X1 port map( A1 => n6446, A2 => n6410, ZN => n3962);
   U182 : BUF_X1 port map( A => n1736, Z => n6441);
   U184 : NAND2_X1 port map( A1 => n6446, A2 => n6438, ZN => n1808);
   U186 : NAND2_X1 port map( A1 => n6446, A2 => n6434, ZN => n1848);
   U188 : NAND2_X1 port map( A1 => n6446, A2 => n6405, ZN => n4001);
   U190 : NAND2_X1 port map( A1 => n6446, A2 => n6412, ZN => n3927);
   U192 : NAND2_X1 port map( A1 => n6446, A2 => n6396, ZN => n4111);
   U194 : BUF_X1 port map( A => n1812, Z => n6436);
   U196 : NAND2_X1 port map( A1 => n6446, A2 => n6440, ZN => n1773);
   U198 : NAND2_X1 port map( A1 => n6446, A2 => n6398, ZN => n4107);
   U200 : NAND2_X1 port map( A1 => n6446, A2 => n6417, ZN => n2063);
   U202 : NAND2_X1 port map( A1 => n6446, A2 => n6403, ZN => n4036);
   U204 : BUF_X1 port map( A => n3995, Z => n6407);
   U206 : NAND2_X1 port map( A1 => n6446, A2 => n6445, ZN => n1664);
   U208 : NAND2_X1 port map( A1 => n6446, A2 => n6419, ZN => n2028);
   U210 : BUF_X2 port map( A => n1772, Z => n6440);
   U212 : BUF_X2 port map( A => n4110, Z => n6396);
   U214 : BUF_X2 port map( A => n1662, Z => n6445);
   U216 : BUF_X2 port map( A => n1956, Z => n6425);
   U218 : NAND2_X1 port map( A1 => n6446, A2 => n6401, ZN => n4069);
   U220 : BUF_X2 port map( A => n4106, Z => n6398);
   U222 : BUF_X2 port map( A => n4035, Z => n6403);
   U224 : BUF_X2 port map( A => n3926, Z => n6412);
   U226 : NAND2_X1 port map( A1 => n6446, A2 => n6392, ZN => n4181);
   U228 : NAND2_X1 port map( A1 => n6446, A2 => n6437, ZN => n1812);
   U230 : NAND2_X1 port map( A1 => n6446, A2 => n6408, ZN => n3995);
   U232 : BUF_X2 port map( A => n1852, Z => n6433);
   U234 : BUF_X2 port map( A => n4000, Z => n6405);
   U236 : BUF_X2 port map( A => n1807, Z => n6438);
   U269 : NAND2_X1 port map( A1 => n6446, A2 => n6423, ZN => n1991);
   U271 : BUF_X1 port map( A => n2062, Z => n6417);
   U273 : BUF_X2 port map( A => n1921, Z => n6427);
   U275 : BUF_X2 port map( A => n3961, Z => n6410);
   U277 : NAND2_X1 port map( A1 => n6446, A2 => n6415, ZN => n3889);
   U279 : NAND2_X1 port map( A1 => n6446, A2 => n6400, ZN => n4074);
   U281 : NAND2_X1 port map( A1 => n6446, A2 => n6435, ZN => n1844);
   U283 : BUF_X2 port map( A => n1847, Z => n6434);
   U285 : NAND2_X1 port map( A1 => n6446, A2 => n6442, ZN => n1736);
   U287 : NAND2_X1 port map( A1 => n6446, A2 => n6443, ZN => n1731);
   U289 : NAND2_X1 port map( A1 => n6446, A2 => n6394, ZN => n4146);
   U291 : NAND2_X1 port map( A1 => n6446, A2 => n6406, ZN => n3997);
   U293 : BUF_X2 port map( A => n3892, Z => n6414);
   U295 : NAND2_X1 port map( A1 => n6446, A2 => n3892, ZN => n3893);
   U297 : BUF_X2 port map( A => n1885, Z => n6431);
   U299 : BUF_X2 port map( A => n1990, Z => n6423);
   U301 : BUF_X2 port map( A => n3994, Z => n6408);
   U303 : BUF_X2 port map( A => n1917, Z => n6429);
   U305 : BUF_X2 port map( A => n3996, Z => n6406);
   U307 : BUF_X2 port map( A => n2023, Z => n6421);
   U309 : BUF_X2 port map( A => n1843, Z => n6435);
   U311 : BUF_X1 port map( A => n1735, Z => n6442);
   U313 : BUF_X2 port map( A => n4180, Z => n6392);
   U315 : BUF_X2 port map( A => n4145, Z => n6394);
   U317 : BUF_X2 port map( A => n4073, Z => n6400);
   U319 : BUF_X2 port map( A => n4068, Z => n6401);
   U321 : BUF_X2 port map( A => n1811, Z => n6437);
   U323 : INV_X1 port map( A => ADD_WR(1), ZN => n4143);
   U325 : BUF_X2 port map( A => n4204, Z => n6385);
   U327 : INV_X1 port map( A => ADD_WR(0), ZN => n4178);
   U329 : INV_X1 port map( A => ADD_WR(3), ZN => n1846);
   U331 : BUF_X2 port map( A => n4218, Z => n3890);
   U333 : BUF_X2 port map( A => n4224, Z => n3894);
   U335 : BUF_X2 port map( A => n4223, Z => n3895);
   U369 : BUF_X2 port map( A => n4226, Z => n3896);
   U371 : BUF_X2 port map( A => n4219, Z => n3897);
   U404 : BUF_X2 port map( A => n4205, Z => n3898);
   U406 : BUF_X2 port map( A => n4208, Z => n3899);
   U408 : BUF_X2 port map( A => n4207, Z => n3900);
   U410 : BUF_X2 port map( A => n4210, Z => n3901);
   U412 : BUF_X2 port map( A => n4209, Z => n3902);
   U414 : BUF_X2 port map( A => n4211, Z => n3904);
   U416 : BUF_X2 port map( A => n5231, Z => n3905);
   U418 : BUF_X2 port map( A => n5230, Z => n3906);
   U420 : BUF_X2 port map( A => n5233, Z => n3907);
   U422 : BUF_X2 port map( A => n5232, Z => n3908);
   U424 : BUF_X2 port map( A => n5235, Z => n3909);
   U426 : BUF_X2 port map( A => n5234, Z => n3910);
   U428 : BUF_X2 port map( A => n5246, Z => n3911);
   U430 : BUF_X2 port map( A => n5247, Z => n3912);
   U432 : BUF_X2 port map( A => n5242, Z => n3913);
   U434 : BUF_X2 port map( A => n5243, Z => n3914);
   U436 : NOR2_X2 port map( A1 => n5181, A2 => n5171, ZN => n4225);
   U438 : BUF_X2 port map( A => n5260, Z => n6359);
   U440 : BUF_X2 port map( A => n4238, Z => n6379);
   U442 : NAND2_X1 port map( A1 => n6446, A2 => n6433, ZN => n1853);
   U444 : NAND2_X1 port map( A1 => n6446, A2 => n6431, ZN => n1886);
   U446 : NAND2_X1 port map( A1 => n6446, A2 => n6429, ZN => n1918);
   U448 : NAND2_X1 port map( A1 => n6446, A2 => n6427, ZN => n1922);
   U450 : NAND2_X1 port map( A1 => n6446, A2 => n6425, ZN => n1957);
   U452 : NAND2_X1 port map( A1 => n6446, A2 => n6421, ZN => n2024);
   U454 : BUF_X2 port map( A => n4228, Z => n6382);
   U456 : BUF_X1 port map( A => n1730, Z => n6443);
   U458 : BUF_X1 port map( A => n3888, Z => n6415);
   U460 : BUF_X1 port map( A => n3893, Z => n6413);
   U462 : BUF_X1 port map( A => n2028, Z => n6418);
   U464 : BUF_X1 port map( A => n2024, Z => n6420);
   U466 : BUF_X1 port map( A => n1922, Z => n6426);
   U468 : BUF_X1 port map( A => n1957, Z => n6424);
   U470 : BUF_X1 port map( A => n1918, Z => n6428);
   U473 : BUF_X1 port map( A => n1853, Z => n6432);
   U475 : BUF_X1 port map( A => n1886, Z => n6430);
   U477 : BUF_X1 port map( A => n4240, Z => n6377);
   U479 : OAI21_X1 port map( B1 => n1768, B2 => n1729, A => n6446, ZN => n1735)
                           ;
   U481 : OAI21_X1 port map( B1 => n1728, B2 => n2060, A => n6446, ZN => n2062)
                           ;
   U483 : NAND2_X1 port map( A1 => ADD_WR(0), A2 => n4143, ZN => n1728);
   U485 : BUF_X1 port map( A => n4241, Z => n6376);
   U487 : BUF_X1 port map( A => n4192, Z => n6388);
   U489 : OAI21_X1 port map( B1 => n1733, B2 => n1729, A => n6446, ZN => n1730)
                           ;
   U491 : OAI21_X1 port map( B1 => n1733, B2 => n2060, A => n6446, ZN => n3888)
                           ;
   U493 : NAND2_X1 port map( A1 => ADD_WR(1), A2 => ADD_WR(0), ZN => n1768);
   U495 : NAND2_X1 port map( A1 => ADD_WR(1), A2 => n4178, ZN => n1733);
   U497 : BUF_X1 port map( A => n5219, Z => n6372);
   U499 : BUF_X1 port map( A => n5262, Z => n6357);
   U501 : BUF_X1 port map( A => n5264, Z => n6355);
   U503 : BUF_X1 port map( A => n4186, Z => n6390);
   U505 : BUF_X1 port map( A => n2027, Z => n6419);
   U507 : NOR2_X1 port map( A1 => ADD_WR(4), A2 => n2025, ZN => n1770);
   U509 : INV_X2 port map( A => n3950, ZN => n6381);
   U511 : BUF_X1 port map( A => n5213, Z => n6374);
   U513 : INV_X1 port map( A => ADD_WR(4), ZN => n5146);
   U515 : NOR2_X1 port map( A1 => ADD_WR(3), A2 => ADD_WR(2), ZN => n1769);
   U517 : INV_X2 port map( A => n3952, ZN => n6361);
   U519 : OAI21_X1 port map( B1 => n1805, B2 => n2060, A => n6446, ZN => n2027)
                           ;
   U521 : INV_X2 port map( A => n3951, ZN => n6389);
   U523 : BUF_X1 port map( A => n4225, Z => n6383);
   U525 : BUF_X1 port map( A => n4237, Z => n6380);
   U527 : BUF_X1 port map( A => n5236, Z => n6369);
   U529 : BUF_X1 port map( A => n5244, Z => n6367);
   U531 : BUF_X1 port map( A => n5248, Z => n6365);
   U533 : INV_X2 port map( A => n3953, ZN => n6373);
   U535 : INV_X2 port map( A => n6387, ZN => n6386);
   U569 : BUF_X1 port map( A => n4220, Z => n6384);
   U572 : OR2_X2 port map( A1 => n5168, A2 => n5184, ZN => n4194);
   U574 : OR2_X2 port map( A1 => n5179, A2 => n5156, ZN => n4234);
   U576 : INV_X2 port map( A => n6371, ZN => n6370);
   U578 : BUF_X1 port map( A => n5237, Z => n6368);
   U580 : BUF_X1 port map( A => n5245, Z => n6366);
   U582 : BUF_X1 port map( A => n5249, Z => n6364);
   U584 : BUF_X1 port map( A => n5251, Z => n6362);
   U586 : OR2_X2 port map( A1 => n5948, A2 => n5961, ZN => n5220);
   U588 : OR2_X2 port map( A1 => n5958, A2 => n5936, ZN => n5255);
   U590 : INV_X2 port map( A => n5974, ZN => n5257);
   U592 : NOR2_X1 port map( A1 => n5172, A2 => n5173, ZN => n4211);
   U594 : NOR2_X1 port map( A1 => n5948, A2 => n5937, ZN => n5230);
   U596 : NOR2_X1 port map( A1 => n5172, A2 => n5157, ZN => n4207);
   U598 : NOR2_X1 port map( A1 => n5168, A2 => n5158, ZN => n4209);
   U600 : NOR2_X1 port map( A1 => n5172, A2 => n5179, ZN => n4219);
   U602 : NOR2_X1 port map( A1 => n5168, A2 => n5179, ZN => n4223);
   U604 : NOR2_X1 port map( A1 => n5173, A2 => n5171, ZN => n4221);
   U606 : NOR2_X1 port map( A1 => n5172, A2 => n5158, ZN => n4212);
   U608 : NOR2_X1 port map( A1 => n5952, A2 => n5937, ZN => n5232);
   U610 : NOR2_X1 port map( A1 => n5948, A2 => n5938, ZN => n5234);
   U612 : NOR2_X1 port map( A1 => n5948, A2 => n5958, ZN => n5246);
   U614 : NOR2_X1 port map( A1 => n5948, A2 => n5935, ZN => n5242);
   U616 : NOR2_X1 port map( A1 => n5948, A2 => n5949, ZN => n5231);
   U618 : NOR2_X1 port map( A1 => n5170, A2 => n5182, ZN => n4226);
   U620 : NOR2_X1 port map( A1 => n5168, A2 => n5157, ZN => n4205);
   U622 : NOR2_X1 port map( A1 => n5168, A2 => n5173, ZN => n4210);
   U624 : NOR2_X1 port map( A1 => n5168, A2 => n5155, ZN => n4218);
   U626 : NOR2_X1 port map( A1 => n5181, A2 => n5182, ZN => n4224);
   U628 : NOR2_X1 port map( A1 => n5170, A2 => n5171, ZN => n4208);
   U630 : NOR2_X1 port map( A1 => n5948, A2 => n5953, ZN => n5235);
   U632 : NOR2_X1 port map( A1 => n5959, A2 => n5960, ZN => n5247);
   U634 : NOR2_X1 port map( A1 => n5952, A2 => n5958, ZN => n5243);
   U636 : NOR2_X1 port map( A1 => n5950, A2 => n5951, ZN => n5233);
   U638 : OAI21_X1 port map( B1 => ADD_WR(4), B2 => n5983, A => WR, ZN => n5206
                           );
   U640 : AOI22_X1 port map( A1 => ADD_WR(1), A2 => ADD_RD1(1), B1 => n5963, B2
                           => n4143, ZN => n5979);
   U642 : AOI22_X1 port map( A1 => ADD_WR(1), A2 => ADD_RD2(1), B1 => n5187, B2
                           => n4143, ZN => n5201);
   U644 : AOI22_X1 port map( A1 => ADD_WR(0), A2 => ADD_RD1(0), B1 => n5966, B2
                           => n4178, ZN => n5978);
   U646 : AOI22_X1 port map( A1 => ADD_WR(0), A2 => ADD_RD2(0), B1 => n5189, B2
                           => n4178, ZN => n5202);
   U648 : AOI22_X1 port map( A1 => ADD_WR(3), A2 => ADD_RD1(3), B1 => n5971, B2
                           => n1846, ZN => n5973);

end SYN_A;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity 
   dlx_cu_MICROCODE_MEM_SIZE64_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE13 is

   port( Clk, Rst : in std_logic;  IR_IN : in std_logic_vector (31 downto 0);  
         stall_exe_i, mispredict_i : in std_logic;  D1_i, D2_i : in 
         std_logic_vector (4 downto 0);  S1_LATCH_EN, S2_LATCH_EN, S3_LATCH_EN 
         : out std_logic;  S_MUX_PC_BUS : out std_logic_vector (1 downto 0);  
         S_EXT, S_EXT_SIGN, S_EQ_NEQ : out std_logic;  S_MUX_DEST : out 
         std_logic_vector (1 downto 0);  S_MUX_LINK, S_MEM_W_R, S_MEM_EN, 
         S_RF_W_wb, S_RF_W_mem, S_RF_W_exe, S_MUX_ALUIN, stall_exe_o, 
         stall_dec_o, stall_fetch_o, stall_btb_o, was_branch_o, was_jmp_o : out
         std_logic;  ALU_WORD_o : out std_logic_vector (12 downto 0);  
         ALU_OPCODE : out std_logic_vector (0 to 4);  S_MUX_MEM_BAR : out 
         std_logic);

end dlx_cu_MICROCODE_MEM_SIZE64_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE13;

architecture SYN_dlx_cu_hw of 
   dlx_cu_MICROCODE_MEM_SIZE64_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE13 is

   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFS_X1
      port( D, CK, SN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFR_X2
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component alu_ctrl
      port( OP : in std_logic_vector (0 to 4);  ALU_WORD : out std_logic_vector
            (12 downto 0));
   end component;
   
   component cw_mem_MICROCODE_MEM_SIZE64_OP_CODE_SIZE6_CW_SIZE13
      port( OPCODE_IN : in std_logic_vector (5 downto 0);  CW_OUT : out 
            std_logic_vector (12 downto 0));
   end component;
   
   component stall_logic_FUNC_SIZE11_OP_CODE_SIZE6
      port( OPCODE_i : in std_logic_vector (5 downto 0);  FUNC_i : in 
            std_logic_vector (10 downto 0);  rA_i, rB_i, D1_i, D2_i : in 
            std_logic_vector (4 downto 0);  S_mem_LOAD_i, S_exe_LOAD_i : in 
            std_logic;  S_MUX_PC_BUS_i : in std_logic_vector (1 downto 0);  
            mispredict_i : in std_logic;  bubble_dec_o, bubble_exe_o, 
            stall_exe_o, stall_dec_o, stall_btb_o, stall_fetch_o : out 
            std_logic;  S_exe_WRITE_i_BAR : in std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal S_MUX_PC_BUS_1_port, S_MUX_PC_BUS_0_port, S_MEM_W_R_port, S_MEM_LOAD,
      S_EXE_LOAD, next_bubble_dec, stall_fetch_o_TEMP, cw_from_mem_12_port, 
      cw_from_mem_11_port, cw_from_mem_10_port, cw_from_mem_9_port, 
      cw_from_mem_8_port, cw_from_mem_7_port, cw_from_mem_6_port, 
      cw_from_mem_4_port, cw_from_mem_3_port, cw_from_mem_2_port, 
      cw_from_mem_1_port, cw_from_mem_0_port, aluOpcode_d_4_port, 
      aluOpcode_d_3_port, aluOpcode_d_2_port, aluOpcode_d_1_port, 
      aluOpcode_d_0_port, N29, N30, N31, N32, n138, n139, n140, n143, n150, 
      n151, n152, n153, n154, n155, n156, n157, n159, n2, n119, n123, net644354
      , net644355, net644356, n35, n36, n37, n38, n39, n40, n41, n42, n49, n50,
      n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65
      , n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, 
      n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94
      , n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107
      , n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n124,
      n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, 
      n137, n141, n149, n158, n160, n161, n162, n163, n164, n165, n166, n167, 
      n168, n169, n170, n171, n172, n142, n144, n147, stall_btb_o_port, n173, 
      n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, 
      n186, n187, n188, net684159, net684160, net684161, net684162, net684163, 
      net684164, net684165, net684166, net684167, net684168 : std_logic;

begin
   S_MUX_PC_BUS <= ( S_MUX_PC_BUS_1_port, S_MUX_PC_BUS_0_port );
   S_MEM_W_R <= S_MEM_W_R_port;
   stall_exe_o <= stall_exe_i;
   stall_dec_o <= stall_btb_o_port;
   stall_fetch_o <= stall_btb_o_port;
   stall_btb_o <= stall_btb_o_port;
   
   bubble_dec_reg : DFF_X1 port map( D => n157, CK => Clk, Q => n119, QN => 
                           n173);
   cw_e_reg_0_inst : DFFR_X1 port map( D => n156, CK => Clk, RN => n175, Q => 
                           net684168, QN => n123);
   cw_e_reg_5_inst : DFFR_X1 port map( D => n154, CK => Clk, RN => n175, Q => 
                           S_MUX_DEST(1), QN => n139);
   cw_e_reg_4_inst : DFFR_X1 port map( D => n153, CK => Clk, RN => n175, Q => 
                           S_MUX_DEST(0), QN => n138);
   cw_e_reg_3_inst : DFFR_X1 port map( D => n152, CK => Clk, RN => n175, Q => 
                           net684167, QN => n2);
   cw_e_reg_2_inst : DFFR_X1 port map( D => n151, CK => Clk, RN => n175, Q => 
                           net644356, QN => net684166);
   cw_e_reg_1_inst : DFFR_X1 port map( D => n150, CK => Clk, RN => n175, Q => 
                           net644355, QN => net684165);
   cw_m_reg_2_inst : DFFR_X1 port map( D => N31, CK => Clk, RN => n175, Q => 
                           S_MEM_W_R_port, QN => net644354);
   cw_m_reg_3_inst : DFFR_X1 port map( D => N32, CK => Clk, RN => n175, Q => 
                           S_MEM_EN, QN => n159);
   cw_m_reg_0_inst : DFFR_X1 port map( D => N29, CK => Clk, RN => n175, Q => 
                           S_RF_W_mem, QN => n143);
   U145 : XOR2_X1 port map( A => S_MUX_PC_BUS_1_port, B => S_MUX_PC_BUS_0_port,
                           Z => was_jmp_o);
   U146 : MUX2_X1 port map( A => next_bubble_dec, B => n119, S => Rst, Z => 
                           n157);
   U147 : NAND3_X1 port map( A1 => n174, A2 => n67, A3 => n68, ZN => n66);
   U148 : NAND3_X1 port map( A1 => IR_IN(5), A2 => IR_IN(0), A3 => IR_IN(4), ZN
                           => n80);
   U149 : NAND3_X1 port map( A1 => n137, A2 => n77, A3 => n100, ZN => n72);
   U150 : NAND3_X1 port map( A1 => IR_IN(30), A2 => n174, A3 => n93, ZN => n164
                           );
   U151 : NAND3_X1 port map( A1 => n116, A2 => n117, A3 => n141, ZN => n167);
   U152 : NAND3_X1 port map( A1 => IR_IN(1), A2 => IR_IN(3), A3 => n75, ZN => 
                           n62);
   U153 : NAND3_X1 port map( A1 => IR_IN(5), A2 => IR_IN(4), A3 => n100, ZN => 
                           n61);
   STALL_L : stall_logic_FUNC_SIZE11_OP_CODE_SIZE6 port map( OPCODE_i(5) => 
                           IR_IN(31), OPCODE_i(4) => IR_IN(30), OPCODE_i(3) => 
                           IR_IN(29), OPCODE_i(2) => n174, OPCODE_i(1) => n147,
                           OPCODE_i(0) => IR_IN(26), FUNC_i(10) => n176, 
                           FUNC_i(9) => n177, FUNC_i(8) => n178, FUNC_i(7) => 
                           n179, FUNC_i(6) => n180, FUNC_i(5) => n181, 
                           FUNC_i(4) => n182, FUNC_i(3) => n183, FUNC_i(2) => 
                           n184, FUNC_i(1) => n185, FUNC_i(0) => n186, rA_i(4) 
                           => IR_IN(25), rA_i(3) => IR_IN(24), rA_i(2) => 
                           IR_IN(23), rA_i(1) => IR_IN(22), rA_i(0) => 
                           IR_IN(21), rB_i(4) => IR_IN(20), rB_i(3) => 
                           IR_IN(19), rB_i(2) => IR_IN(18), rB_i(1) => 
                           IR_IN(17), rB_i(0) => IR_IN(16), D1_i(4) => D1_i(4),
                           D1_i(3) => D1_i(3), D1_i(2) => D1_i(2), D1_i(1) => 
                           D1_i(1), D1_i(0) => D1_i(0), D2_i(4) => D2_i(4), 
                           D2_i(3) => D2_i(3), D2_i(2) => D2_i(2), D2_i(1) => 
                           D2_i(1), D2_i(0) => D2_i(0), S_mem_LOAD_i => 
                           S_MEM_LOAD, S_exe_LOAD_i => S_EXE_LOAD, 
                           S_MUX_PC_BUS_i(1) => n187, S_MUX_PC_BUS_i(0) => n188
                           , mispredict_i => mispredict_i, bubble_dec_o => 
                           next_bubble_dec, bubble_exe_o => net684161, 
                           stall_exe_o => net684162, stall_dec_o => net684163, 
                           stall_btb_o => net684164, stall_fetch_o => 
                           stall_fetch_o_TEMP, S_exe_WRITE_i_BAR => n123);
   CWM : cw_mem_MICROCODE_MEM_SIZE64_OP_CODE_SIZE6_CW_SIZE13 port map( 
                           OPCODE_IN(5) => IR_IN(31), OPCODE_IN(4) => IR_IN(30)
                           , OPCODE_IN(3) => IR_IN(29), OPCODE_IN(2) => 
                           IR_IN(28), OPCODE_IN(1) => IR_IN(27), OPCODE_IN(0) 
                           => IR_IN(26), CW_OUT(12) => cw_from_mem_12_port, 
                           CW_OUT(11) => cw_from_mem_11_port, CW_OUT(10) => 
                           cw_from_mem_10_port, CW_OUT(9) => cw_from_mem_9_port
                           , CW_OUT(8) => cw_from_mem_8_port, CW_OUT(7) => 
                           cw_from_mem_7_port, CW_OUT(6) => cw_from_mem_6_port,
                           CW_OUT(5) => net684160, CW_OUT(4) => 
                           cw_from_mem_4_port, CW_OUT(3) => cw_from_mem_3_port,
                           CW_OUT(2) => cw_from_mem_2_port, CW_OUT(1) => 
                           cw_from_mem_1_port, CW_OUT(0) => cw_from_mem_0_port)
                           ;
   ALU_C : alu_ctrl port map( OP(0) => aluOpcode_d_4_port, OP(1) => 
                           aluOpcode_d_3_port, OP(2) => aluOpcode_d_2_port, 
                           OP(3) => aluOpcode_d_1_port, OP(4) => 
                           aluOpcode_d_0_port, ALU_WORD(12) => ALU_WORD_o(12), 
                           ALU_WORD(11) => ALU_WORD_o(11), ALU_WORD(10) => 
                           ALU_WORD_o(10), ALU_WORD(9) => ALU_WORD_o(9), 
                           ALU_WORD(8) => ALU_WORD_o(8), ALU_WORD(7) => 
                           ALU_WORD_o(7), ALU_WORD(6) => ALU_WORD_o(6), 
                           ALU_WORD(5) => ALU_WORD_o(5), ALU_WORD(4) => 
                           ALU_WORD_o(4), ALU_WORD(3) => ALU_WORD_o(3), 
                           ALU_WORD(2) => ALU_WORD_o(2), ALU_WORD(1) => 
                           ALU_WORD_o(1), ALU_WORD(0) => ALU_WORD_o(0));
   cw_m_reg_1_inst : DFFR_X1 port map( D => N30, CK => Clk, RN => n175, Q => 
                           net684159, QN => S_MUX_MEM_BAR);
   U137 : AND2_X1 port map( A1 => cw_from_mem_8_port, A2 => n173, ZN => 
                           S_EQ_NEQ);
   U116 : NOR4_X1 port map( A1 => IR_IN(7), A2 => IR_IN(9), A3 => IR_IN(8), A4 
                           => IR_IN(6), ZN => n169);
   U112 : NAND4_X1 port map( A1 => n169, A2 => n170, A3 => n106, A4 => n165, ZN
                           => n168);
   U37 : NAND2_X1 port map( A1 => IR_IN(5), A2 => IR_IN(4), ZN => n50);
   U70 : NAND2_X1 port map( A1 => IR_IN(5), A2 => IR_IN(0), ZN => n54);
   U77 : NAND4_X1 port map( A1 => IR_IN(2), A2 => n59, A3 => IR_IN(3), A4 => 
                           n99, ZN => n55);
   U36 : NOR2_X1 port map( A1 => n61, A2 => n62, ZN => n60);
   U52 : NAND2_X1 port map( A1 => IR_IN(26), A2 => n82, ZN => n57);
   U34 : OAI211_X1 port map( C1 => n54, C2 => n55, A => n56, B => n57, ZN => 
                           n52);
   U106 : NOR2_X1 port map( A1 => IR_IN(0), A2 => n99, ZN => n116);
   U102 : NOR3_X1 port map( A1 => n124, A2 => n168, A3 => n75, ZN => n117);
   U101 : NOR3_X1 port map( A1 => IR_IN(5), A2 => n166, A3 => n167, ZN => n83);
   U64 : NAND2_X1 port map( A1 => n59, A2 => n76, ZN => n114);
   U128 : NOR2_X1 port map( A1 => IR_IN(5), A2 => IR_IN(4), ZN => n115);
   U63 : NAND4_X1 port map( A1 => IR_IN(3), A2 => n115, A3 => n116, A4 => n117,
                           ZN => n94);
   U62 : OAI21_X1 port map( B1 => n62, B2 => n114, A => n94, ZN => n84);
   U45 : OAI221_X1 port map( B1 => n55, B2 => n61, C1 => n55, C2 => n80, A => 
                           n81, ZN => n53);
   U33 : NOR2_X1 port map( A1 => n52, A2 => n53, ZN => n51);
   U59 : NAND2_X1 port map( A1 => n106, A2 => n107, ZN => n86);
   U79 : NAND2_X1 port map( A1 => n82, A2 => n124, ZN => n64);
   U127 : NAND2_X1 port map( A1 => IR_IN(0), A2 => IR_IN(1), ZN => n78);
   U43 : AOI22_X1 port map( A1 => IR_IN(1), A2 => n76, B1 => n77, B2 => n78, ZN
                           => n74);
   U42 : NOR3_X1 port map( A1 => IR_IN(3), A2 => n74, A3 => n75, ZN => n69);
   U108 : NAND2_X1 port map( A1 => n77, A2 => n75, ZN => n96);
   U107 : NOR2_X1 port map( A1 => n141, A2 => n96, ZN => n73);
   U85 : NOR3_X1 port map( A1 => IR_IN(1), A2 => n75, A3 => n141, ZN => n137);
   U40 : OAI211_X1 port map( C1 => n61, C2 => n62, A => n71, B => n72, ZN => 
                           n70);
   U39 : OAI21_X1 port map( B1 => n69, B2 => n70, A => n59, ZN => n65);
   U38 : NAND4_X1 port map( A1 => n63, A2 => n64, A3 => n65, A4 => n66, ZN => 
                           aluOpcode_d_3_port);
   U124 : NAND2_X1 port map( A1 => n100, A2 => n99, ZN => n133);
   U84 : NAND2_X1 port map( A1 => n59, A2 => n73, ZN => n128);
   U81 : OAI21_X1 port map( B1 => n105, B2 => n87, A => n107, ZN => n134);
   U78 : OAI211_X1 port map( C1 => n133, C2 => n128, A => n134, B => n64, ZN =>
                           n131);
   U76 : AOI221_X1 port map( B1 => n99, B2 => n55, C1 => n49, C2 => n55, A => 
                           n61, ZN => n132);
   U75 : AOI211_X1 port map( C1 => n59, C2 => n104, A => n131, B => n132, ZN =>
                           n108);
   U73 : NOR2_X1 port map( A1 => n128, A2 => n78, ZN => n127);
   U69 : OAI21_X1 port map( B1 => IR_IN(5), B2 => IR_IN(2), A => n54, ZN => 
                           n118);
   U68 : NOR3_X1 port map( A1 => n118, A2 => IR_IN(4), A3 => n99, ZN => n112);
   U66 : NOR2_X1 port map( A1 => IR_IN(1), A2 => n80, ZN => n103);
   U61 : AOI221_X1 port map( B1 => n112, B2 => n113, C1 => n103, C2 => n113, A 
                           => n84, ZN => n111);
   U60 : NAND4_X1 port map( A1 => n108, A2 => n109, A3 => n110, A4 => n111, ZN 
                           => aluOpcode_d_1_port);
   U122 : AOI21_X1 port map( B1 => n78, B2 => n133, A => n75, ZN => n171);
   U121 : NOR2_X1 port map( A1 => IR_IN(1), A2 => n100, ZN => n172);
   U117 : AOI221_X1 port map( B1 => n115, B2 => n171, C1 => n172, C2 => n77, A 
                           => n97, ZN => n129);
   U105 : NAND2_X1 port map( A1 => n73, A2 => n116, ZN => n102);
   U104 : OAI21_X1 port map( B1 => n62, B2 => n61, A => n102, ZN => n149);
   U96 : NAND2_X1 port map( A1 => n67, A2 => n165, ZN => n160);
   U88 : AOI21_X1 port map( B1 => n162, B2 => n126, A => n163, ZN => n161);
   U87 : OAI221_X1 port map( B1 => n124, B2 => n160, C1 => IR_IN(26), C2 => n85
                           , A => n161, ZN => n158);
   U86 : AOI211_X1 port map( C1 => n59, C2 => n149, A => n83, B => n158, ZN => 
                           n130);
   U74 : OAI211_X1 port map( C1 => n129, C2 => n49, A => n130, B => n108, ZN =>
                           aluOpcode_d_0_port);
   U57 : AOI21_X1 port map( B1 => IR_IN(2), B2 => n103, A => n104, ZN => n101);
   U56 : OAI211_X1 port map( C1 => n96, C2 => n100, A => n101, B => n102, ZN =>
                           n90);
   U55 : NOR2_X1 port map( A1 => n99, A2 => n80, ZN => n98);
   U54 : AOI22_X1 port map( A1 => IR_IN(2), A2 => n97, B1 => n98, B2 => n75, ZN
                           => n95);
   U53 : AOI21_X1 port map( B1 => n95, B2 => n96, A => n49, ZN => n91);
   U50 : AOI211_X1 port map( C1 => n59, C2 => n90, A => n91, B => n92, ZN => 
                           n89);
   U19 : NOR2_X1 port map( A1 => n119, A2 => stall_btb_o_port, ZN => n37);
   U18 : AOI22_X1 port map( A1 => stall_exe_i, A2 => net644355, B1 => n37, B2 
                           => cw_from_mem_1_port, ZN => n42);
   U16 : AOI22_X1 port map( A1 => stall_exe_i, A2 => net644356, B1 => n37, B2 
                           => cw_from_mem_2_port, ZN => n41);
   U143 : INV_X1 port map( A => stall_exe_i, ZN => n35);
   U10 : NAND2_X1 port map( A1 => n37, A2 => cw_from_mem_6_port, ZN => n38);
   U8 : OAI21_X1 port map( B1 => n140, B2 => n35, A => n38, ZN => n155);
   U9 : OAI21_X1 port map( B1 => n139, B2 => n35, A => n38, ZN => n154);
   U14 : NAND2_X1 port map( A1 => n37, A2 => cw_from_mem_3_port, ZN => n40);
   U13 : OAI21_X1 port map( B1 => n35, B2 => n2, A => n40, ZN => n152);
   U12 : NAND2_X1 port map( A1 => n37, A2 => cw_from_mem_4_port, ZN => n39);
   U11 : OAI21_X1 port map( B1 => n35, B2 => n138, A => n39, ZN => n153);
   U7 : NAND2_X1 port map( A1 => n37, A2 => cw_from_mem_0_port, ZN => n36);
   U6 : OAI21_X1 port map( B1 => n35, B2 => n123, A => n36, ZN => n156);
   U140 : NOR2_X1 port map( A1 => stall_exe_i, A2 => n2, ZN => N32);
   U144 : NOR2_X1 port map( A1 => stall_exe_i, A2 => n123, ZN => N29);
   U131 : AND2_X2 port map( A1 => cw_from_mem_7_port, A2 => n173, ZN => 
                           S_MUX_LINK);
   U111 : NOR2_X1 port map( A1 => IR_IN(26), A2 => n168, ZN => n59);
   U109 : NAND2_X1 port map( A1 => n59, A2 => n141, ZN => n49);
   U103 : INV_X1 port map( A => IR_IN(26), ZN => n124);
   U32 : OAI21_X1 port map( B1 => n49, B2 => n50, A => n51, ZN => 
                           aluOpcode_d_4_port);
   U49 : OAI211_X1 port map( C1 => n87, C2 => n86, A => n88, B => n89, ZN => 
                           aluOpcode_d_2_port);
   U136 : NOR2_X1 port map( A1 => net644356, A2 => n2, ZN => S_EXE_LOAD);
   cw_e_reg_6_inst : DFFR_X2 port map( D => n155, CK => Clk, RN => n175, Q => 
                           S_MUX_ALUIN, QN => n140);
   U120 : INV_X1 port map( A => IR_IN(4), ZN => n166);
   U126 : INV_X1 port map( A => IR_IN(0), ZN => n100);
   U125 : INV_X1 port map( A => IR_IN(1), ZN => n99);
   U123 : INV_X1 port map( A => IR_IN(2), ZN => n75);
   U110 : INV_X1 port map( A => IR_IN(3), ZN => n141);
   U65 : INV_X1 port map( A => n80, ZN => n76);
   U119 : AND2_X1 port map( A1 => n166, A2 => IR_IN(5), ZN => n77);
   U97 : AND2_X1 port map( A1 => n135, A2 => n107, ZN => n67);
   U118 : INV_X1 port map( A => n61, ZN => n97);
   U92 : INV_X1 port map( A => n68, ZN => n162);
   U48 : INV_X1 port map( A => n86, ZN => n79);
   U47 : INV_X1 port map( A => n85, ZN => n58);
   U41 : INV_X1 port map( A => n73, ZN => n71);
   U67 : INV_X1 port map( A => n49, ZN => n113);
   U141 : AND2_X1 port map( A1 => n35, A2 => net644356, ZN => N31);
   U5 : AND2_X1 port map( A1 => S_MUX_PC_BUS_1_port, A2 => S_MUX_PC_BUS_0_port,
                           ZN => was_branch_o);
   U17 : INV_X1 port map( A => n42, ZN => n150);
   U15 : INV_X1 port map( A => n41, ZN => n151);
   cw_w_reg_0_inst : DFFS_X1 port map( D => n143, CK => Clk, SN => n175, Q => 
                           n144, QN => S_RF_W_wb);
   U3 : OAI21_X1 port map( B1 => n78, B2 => n142, A => n72, ZN => n104);
   U4 : OR2_X1 port map( A1 => n96, A2 => IR_IN(3), ZN => n142);
   U20 : AND2_X1 port map( A1 => n173, A2 => cw_from_mem_10_port, ZN => S_EXT);
   U21 : AND2_X1 port map( A1 => n173, A2 => cw_from_mem_11_port, ZN => 
                           S_MUX_PC_BUS_0_port);
   U22 : NOR2_X1 port map( A1 => n159, A2 => S_MEM_W_R_port, ZN => S_MEM_LOAD);
   U23 : OR2_X2 port map( A1 => stall_exe_i, A2 => stall_fetch_o_TEMP, ZN => 
                           stall_btb_o_port);
   U24 : INV_X1 port map( A => n165, ZN => n147);
   U25 : INV_X1 port map( A => n174, ZN => n106);
   U26 : INV_X1 port map( A => Rst, ZN => n175);
   U27 : AND2_X2 port map( A1 => cw_from_mem_9_port, A2 => n173, ZN => 
                           S_EXT_SIGN);
   U28 : AND2_X1 port map( A1 => net644355, A2 => n35, ZN => N30);
   U29 : INV_X1 port map( A => IR_IN(27), ZN => n165);
   U30 : INV_X1 port map( A => IR_IN(30), ZN => n135);
   U31 : AND2_X1 port map( A1 => cw_from_mem_12_port, A2 => n173, ZN => 
                           S_MUX_PC_BUS_1_port);
   U35 : BUF_X1 port map( A => IR_IN(28), Z => n174);
   U44 : NOR2_X1 port map( A1 => IR_IN(29), A2 => n164, ZN => n126);
   U46 : INV_X1 port map( A => IR_IN(29), ZN => n136);
   U51 : AOI21_X1 port map( B1 => n105, B2 => IR_IN(31), A => n83, ZN => n88);
   U58 : AOI22_X1 port map( A1 => IR_IN(31), A2 => n58, B1 => n59, B2 => n60, 
                           ZN => n56);
   U71 : OAI221_X1 port map( B1 => IR_IN(31), B2 => n64, C1 => n93, C2 => n57, 
                           A => n94, ZN => n92);
   U72 : NOR2_X1 port map( A1 => IR_IN(31), A2 => n136, ZN => n107);
   U80 : AOI211_X1 port map( C1 => n82, C2 => IR_IN(31), A => n83, B => n84, ZN
                           => n81);
   U82 : INV_X1 port map( A => IR_IN(31), ZN => n93);
   U83 : AOI211_X1 port map( C1 => IR_IN(30), C2 => n79, A => n58, B => n53, ZN
                           => n63);
   U89 : NOR4_X1 port map( A1 => IR_IN(10), A2 => IR_IN(31), A3 => IR_IN(29), 
                           A4 => IR_IN(30), ZN => n170);
   U90 : NOR3_X1 port map( A1 => n174, A2 => n135, A3 => n136, ZN => n125);
   U91 : NOR3_X1 port map( A1 => IR_IN(30), A2 => n174, A3 => n68, ZN => n105);
   U93 : AOI21_X1 port map( B1 => n147, B2 => n126, A => n127, ZN => n109);
   U94 : OAI221_X1 port map( B1 => n124, B2 => n125, C1 => IR_IN(26), C2 => n67
                           , A => n147, ZN => n110);
   U95 : NOR3_X1 port map( A1 => n164, A2 => IR_IN(26), A3 => n147, ZN => n163)
                           ;
   U98 : NAND2_X1 port map( A1 => n147, A2 => n125, ZN => n85);
   U99 : NOR3_X1 port map( A1 => IR_IN(26), A2 => n147, A3 => n135, ZN => n87);
   U100 : NAND2_X1 port map( A1 => IR_IN(26), A2 => n147, ZN => n68);
   U113 : NOR4_X1 port map( A1 => n147, A2 => n135, A3 => n136, A4 => n106, ZN 
                           => n82);
   n176 <= '0';
   n177 <= '0';
   n178 <= '0';
   n179 <= '0';
   n180 <= '0';
   n181 <= '0';
   n182 <= '0';
   n183 <= '0';
   n184 <= '0';
   n185 <= '0';
   n186 <= '0';
   n187 <= '0';
   n188 <= '0';

end SYN_dlx_cu_hw;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity jump_logic is

   port( NPCF_i, IR_i, A_i : in std_logic_vector (31 downto 0);  A_o : out 
         std_logic_vector (31 downto 0);  rA_o, rB_o, rC_o : out 
         std_logic_vector (4 downto 0);  branch_target_o, sum_addr_o, 
         extended_imm : out std_logic_vector (31 downto 0);  taken_o : out 
         std_logic;  FW_X_i, FW_W_i : in std_logic_vector (31 downto 0);  
         S_FW_Adec_i : in std_logic_vector (1 downto 0);  S_EXT_i, S_EXT_SIGN_i
         , S_MUX_LINK_i, S_EQ_NEQ_i : in std_logic);

end jump_logic;

architecture SYN_struct of jump_logic is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component mux41_MUX_SIZE32
      port( IN0, IN1, IN2, IN3 : in std_logic_vector (31 downto 0);  CTRL : in 
            std_logic_vector (1 downto 0);  OUT1 : out std_logic_vector (31 
            downto 0));
   end component;
   
   component mux21_4
      port( IN0, IN1 : in std_logic_vector (31 downto 0);  CTRL : in std_logic;
            OUT1 : out std_logic_vector (31 downto 0));
   end component;
   
   component zerocheck
      port( IN0 : in std_logic_vector (31 downto 0);  CTRL : in std_logic;  
            OUT1 : out std_logic);
   end component;
   
   component mux21_2
      port( IN0, IN1 : in std_logic_vector (31 downto 0);  CTRL : in std_logic;
            OUT1 : out std_logic_vector (31 downto 0));
   end component;
   
   component p4add_N32_logN5_0
      port( A, B : in std_logic_vector (31 downto 0);  Cin, sign : in std_logic
            ;  S : out std_logic_vector (31 downto 0);  Cout : out std_logic);
   end component;
   
   component extender_32
      port( IN1 : in std_logic_vector (31 downto 0);  CTRL, SIGN : in std_logic
            ;  OUT1 : out std_logic_vector (31 downto 0));
   end component;
   
   signal X_Logic0_port, A_o_31_port, A_o_30_port, A_o_29_port, A_o_28_port, 
      A_o_27_port, A_o_26_port, A_o_25_port, A_o_24_port, A_o_23_port, 
      A_o_22_port, A_o_21_port, A_o_20_port, A_o_19_port, A_o_18_port, 
      A_o_17_port, A_o_16_port, A_o_15_port, A_o_14_port, A_o_13_port, 
      A_o_12_port, A_o_11_port, A_o_10_port, A_o_9_port, A_o_8_port, A_o_7_port
      , A_o_6_port, A_o_5_port, A_o_4_port, A_o_3_port, A_o_2_port, A_o_1_port,
      A_o_0_port, sum_addr_o_31_port, sum_addr_o_30_port, sum_addr_o_29_port, 
      sum_addr_o_28_port, sum_addr_o_27_port, sum_addr_o_26_port, 
      sum_addr_o_25_port, sum_addr_o_24_port, sum_addr_o_23_port, 
      sum_addr_o_22_port, sum_addr_o_21_port, sum_addr_o_20_port, 
      sum_addr_o_19_port, sum_addr_o_18_port, sum_addr_o_17_port, 
      sum_addr_o_16_port, sum_addr_o_15_port, sum_addr_o_14_port, 
      sum_addr_o_13_port, sum_addr_o_12_port, sum_addr_o_11_port, 
      sum_addr_o_10_port, sum_addr_o_9_port, sum_addr_o_8_port, 
      sum_addr_o_7_port, sum_addr_o_6_port, sum_addr_o_5_port, 
      sum_addr_o_4_port, sum_addr_o_3_port, sum_addr_o_2_port, 
      sum_addr_o_1_port, sum_addr_o_0_port, ext_imm_31_port, ext_imm_30_port, 
      ext_imm_29_port, ext_imm_28_port, ext_imm_27_port, ext_imm_26_port, 
      ext_imm_25_port, ext_imm_24_port, ext_imm_23_port, ext_imm_22_port, 
      ext_imm_21_port, ext_imm_20_port, ext_imm_18_port, ext_imm_17_port, 
      ext_imm_16_port, ext_imm_15_port, ext_imm_14_port, ext_imm_13_port, 
      ext_imm_12_port, ext_imm_11_port, ext_imm_10_port, ext_imm_9_port, 
      ext_imm_8_port, ext_imm_7_port, ext_imm_6_port, ext_imm_5_port, 
      ext_imm_4_port, ext_imm_3_port, ext_imm_2_port, ext_imm_1_port, 
      ext_imm_0_port, branch_sel, n1, n2, n4, n5, n6, n7, n8, n9, net684158 : 
      std_logic;

begin
   A_o <= ( A_o_31_port, A_o_30_port, A_o_29_port, A_o_28_port, A_o_27_port, 
      A_o_26_port, A_o_25_port, A_o_24_port, A_o_23_port, A_o_22_port, 
      A_o_21_port, A_o_20_port, A_o_19_port, A_o_18_port, A_o_17_port, 
      A_o_16_port, A_o_15_port, A_o_14_port, A_o_13_port, A_o_12_port, 
      A_o_11_port, A_o_10_port, A_o_9_port, A_o_8_port, A_o_7_port, A_o_6_port,
      A_o_5_port, A_o_4_port, A_o_3_port, A_o_2_port, A_o_1_port, A_o_0_port );
   rA_o <= ( IR_i(25), IR_i(24), IR_i(23), IR_i(22), IR_i(21) );
   rB_o <= ( IR_i(20), IR_i(19), IR_i(18), IR_i(17), IR_i(16) );
   rC_o <= ( IR_i(15), IR_i(14), IR_i(13), IR_i(12), IR_i(11) );
   sum_addr_o <= ( sum_addr_o_31_port, sum_addr_o_30_port, sum_addr_o_29_port, 
      sum_addr_o_28_port, sum_addr_o_27_port, sum_addr_o_26_port, 
      sum_addr_o_25_port, sum_addr_o_24_port, sum_addr_o_23_port, 
      sum_addr_o_22_port, sum_addr_o_21_port, sum_addr_o_20_port, 
      sum_addr_o_19_port, sum_addr_o_18_port, sum_addr_o_17_port, 
      sum_addr_o_16_port, sum_addr_o_15_port, sum_addr_o_14_port, 
      sum_addr_o_13_port, sum_addr_o_12_port, sum_addr_o_11_port, 
      sum_addr_o_10_port, sum_addr_o_9_port, sum_addr_o_8_port, 
      sum_addr_o_7_port, sum_addr_o_6_port, sum_addr_o_5_port, 
      sum_addr_o_4_port, sum_addr_o_3_port, sum_addr_o_2_port, 
      sum_addr_o_1_port, sum_addr_o_0_port );
   
   X_Logic0_port <= '0';
   EXTENDER : extender_32 port map( IN1(31) => n4, IN1(30) => n5, IN1(29) => n6
                           , IN1(28) => n7, IN1(27) => n8, IN1(26) => n9, 
                           IN1(25) => IR_i(25), IN1(24) => IR_i(24), IN1(23) =>
                           IR_i(23), IN1(22) => IR_i(22), IN1(21) => IR_i(21), 
                           IN1(20) => IR_i(20), IN1(19) => IR_i(19), IN1(18) =>
                           IR_i(18), IN1(17) => IR_i(17), IN1(16) => IR_i(16), 
                           IN1(15) => IR_i(15), IN1(14) => IR_i(14), IN1(13) =>
                           IR_i(13), IN1(12) => IR_i(12), IN1(11) => IR_i(11), 
                           IN1(10) => IR_i(10), IN1(9) => IR_i(9), IN1(8) => 
                           IR_i(8), IN1(7) => IR_i(7), IN1(6) => IR_i(6), 
                           IN1(5) => IR_i(5), IN1(4) => IR_i(4), IN1(3) => 
                           IR_i(3), IN1(2) => IR_i(2), IN1(1) => IR_i(1), 
                           IN1(0) => IR_i(0), CTRL => S_EXT_i, SIGN => 
                           S_EXT_SIGN_i, OUT1(31) => ext_imm_31_port, OUT1(30) 
                           => ext_imm_30_port, OUT1(29) => ext_imm_29_port, 
                           OUT1(28) => ext_imm_28_port, OUT1(27) => 
                           ext_imm_27_port, OUT1(26) => ext_imm_26_port, 
                           OUT1(25) => ext_imm_25_port, OUT1(24) => 
                           ext_imm_24_port, OUT1(23) => ext_imm_23_port, 
                           OUT1(22) => ext_imm_22_port, OUT1(21) => 
                           ext_imm_21_port, OUT1(20) => ext_imm_20_port, 
                           OUT1(19) => n1, OUT1(18) => ext_imm_18_port, 
                           OUT1(17) => ext_imm_17_port, OUT1(16) => 
                           ext_imm_16_port, OUT1(15) => ext_imm_15_port, 
                           OUT1(14) => ext_imm_14_port, OUT1(13) => 
                           ext_imm_13_port, OUT1(12) => ext_imm_12_port, 
                           OUT1(11) => ext_imm_11_port, OUT1(10) => 
                           ext_imm_10_port, OUT1(9) => ext_imm_9_port, OUT1(8) 
                           => ext_imm_8_port, OUT1(7) => ext_imm_7_port, 
                           OUT1(6) => ext_imm_6_port, OUT1(5) => ext_imm_5_port
                           , OUT1(4) => ext_imm_4_port, OUT1(3) => 
                           ext_imm_3_port, OUT1(2) => ext_imm_2_port, OUT1(1) 
                           => ext_imm_1_port, OUT1(0) => ext_imm_0_port);
   JUMPADDER : p4add_N32_logN5_0 port map( A(31) => NPCF_i(31), A(30) => 
                           NPCF_i(30), A(29) => NPCF_i(29), A(28) => NPCF_i(28)
                           , A(27) => NPCF_i(27), A(26) => NPCF_i(26), A(25) =>
                           NPCF_i(25), A(24) => NPCF_i(24), A(23) => NPCF_i(23)
                           , A(22) => NPCF_i(22), A(21) => NPCF_i(21), A(20) =>
                           NPCF_i(20), A(19) => NPCF_i(19), A(18) => NPCF_i(18)
                           , A(17) => NPCF_i(17), A(16) => NPCF_i(16), A(15) =>
                           NPCF_i(15), A(14) => NPCF_i(14), A(13) => NPCF_i(13)
                           , A(12) => NPCF_i(12), A(11) => NPCF_i(11), A(10) =>
                           NPCF_i(10), A(9) => NPCF_i(9), A(8) => NPCF_i(8), 
                           A(7) => NPCF_i(7), A(6) => NPCF_i(6), A(5) => 
                           NPCF_i(5), A(4) => NPCF_i(4), A(3) => NPCF_i(3), 
                           A(2) => NPCF_i(2), A(1) => NPCF_i(1), A(0) => 
                           NPCF_i(0), B(31) => ext_imm_31_port, B(30) => 
                           ext_imm_30_port, B(29) => ext_imm_29_port, B(28) => 
                           ext_imm_28_port, B(27) => ext_imm_27_port, B(26) => 
                           ext_imm_26_port, B(25) => ext_imm_25_port, B(24) => 
                           ext_imm_24_port, B(23) => ext_imm_23_port, B(22) => 
                           ext_imm_22_port, B(21) => ext_imm_21_port, B(20) => 
                           ext_imm_20_port, B(19) => n1, B(18) => 
                           ext_imm_18_port, B(17) => ext_imm_17_port, B(16) => 
                           ext_imm_16_port, B(15) => ext_imm_15_port, B(14) => 
                           ext_imm_14_port, B(13) => ext_imm_13_port, B(12) => 
                           ext_imm_12_port, B(11) => ext_imm_11_port, B(10) => 
                           ext_imm_10_port, B(9) => ext_imm_9_port, B(8) => 
                           ext_imm_8_port, B(7) => ext_imm_7_port, B(6) => 
                           ext_imm_6_port, B(5) => ext_imm_5_port, B(4) => 
                           ext_imm_4_port, B(3) => ext_imm_3_port, B(2) => 
                           ext_imm_2_port, B(1) => ext_imm_1_port, B(0) => 
                           ext_imm_0_port, Cin => X_Logic0_port, sign => 
                           X_Logic0_port, S(31) => sum_addr_o_31_port, S(30) =>
                           sum_addr_o_30_port, S(29) => sum_addr_o_29_port, 
                           S(28) => sum_addr_o_28_port, S(27) => 
                           sum_addr_o_27_port, S(26) => sum_addr_o_26_port, 
                           S(25) => sum_addr_o_25_port, S(24) => 
                           sum_addr_o_24_port, S(23) => sum_addr_o_23_port, 
                           S(22) => sum_addr_o_22_port, S(21) => 
                           sum_addr_o_21_port, S(20) => sum_addr_o_20_port, 
                           S(19) => sum_addr_o_19_port, S(18) => 
                           sum_addr_o_18_port, S(17) => sum_addr_o_17_port, 
                           S(16) => sum_addr_o_16_port, S(15) => 
                           sum_addr_o_15_port, S(14) => sum_addr_o_14_port, 
                           S(13) => sum_addr_o_13_port, S(12) => 
                           sum_addr_o_12_port, S(11) => sum_addr_o_11_port, 
                           S(10) => sum_addr_o_10_port, S(9) => 
                           sum_addr_o_9_port, S(8) => sum_addr_o_8_port, S(7) 
                           => sum_addr_o_7_port, S(6) => sum_addr_o_6_port, 
                           S(5) => sum_addr_o_5_port, S(4) => sum_addr_o_4_port
                           , S(3) => sum_addr_o_3_port, S(2) => 
                           sum_addr_o_2_port, S(1) => sum_addr_o_1_port, S(0) 
                           => sum_addr_o_0_port, Cout => net684158);
   BRANCHMUX : mux21_2 port map( IN0(31) => sum_addr_o_31_port, IN0(30) => 
                           sum_addr_o_30_port, IN0(29) => sum_addr_o_29_port, 
                           IN0(28) => sum_addr_o_28_port, IN0(27) => 
                           sum_addr_o_27_port, IN0(26) => sum_addr_o_26_port, 
                           IN0(25) => sum_addr_o_25_port, IN0(24) => 
                           sum_addr_o_24_port, IN0(23) => sum_addr_o_23_port, 
                           IN0(22) => sum_addr_o_22_port, IN0(21) => 
                           sum_addr_o_21_port, IN0(20) => sum_addr_o_20_port, 
                           IN0(19) => sum_addr_o_19_port, IN0(18) => 
                           sum_addr_o_18_port, IN0(17) => sum_addr_o_17_port, 
                           IN0(16) => sum_addr_o_16_port, IN0(15) => 
                           sum_addr_o_15_port, IN0(14) => sum_addr_o_14_port, 
                           IN0(13) => sum_addr_o_13_port, IN0(12) => 
                           sum_addr_o_12_port, IN0(11) => sum_addr_o_11_port, 
                           IN0(10) => sum_addr_o_10_port, IN0(9) => 
                           sum_addr_o_9_port, IN0(8) => sum_addr_o_8_port, 
                           IN0(7) => sum_addr_o_7_port, IN0(6) => 
                           sum_addr_o_6_port, IN0(5) => sum_addr_o_5_port, 
                           IN0(4) => sum_addr_o_4_port, IN0(3) => 
                           sum_addr_o_3_port, IN0(2) => sum_addr_o_2_port, 
                           IN0(1) => sum_addr_o_1_port, IN0(0) => 
                           sum_addr_o_0_port, IN1(31) => NPCF_i(31), IN1(30) =>
                           NPCF_i(30), IN1(29) => NPCF_i(29), IN1(28) => 
                           NPCF_i(28), IN1(27) => NPCF_i(27), IN1(26) => 
                           NPCF_i(26), IN1(25) => NPCF_i(25), IN1(24) => 
                           NPCF_i(24), IN1(23) => NPCF_i(23), IN1(22) => 
                           NPCF_i(22), IN1(21) => NPCF_i(21), IN1(20) => 
                           NPCF_i(20), IN1(19) => NPCF_i(19), IN1(18) => 
                           NPCF_i(18), IN1(17) => NPCF_i(17), IN1(16) => 
                           NPCF_i(16), IN1(15) => NPCF_i(15), IN1(14) => 
                           NPCF_i(14), IN1(13) => NPCF_i(13), IN1(12) => 
                           NPCF_i(12), IN1(11) => NPCF_i(11), IN1(10) => 
                           NPCF_i(10), IN1(9) => NPCF_i(9), IN1(8) => NPCF_i(8)
                           , IN1(7) => NPCF_i(7), IN1(6) => NPCF_i(6), IN1(5) 
                           => NPCF_i(5), IN1(4) => NPCF_i(4), IN1(3) => 
                           NPCF_i(3), IN1(2) => NPCF_i(2), IN1(1) => NPCF_i(1),
                           IN1(0) => NPCF_i(0), CTRL => branch_sel, OUT1(31) =>
                           branch_target_o(31), OUT1(30) => branch_target_o(30)
                           , OUT1(29) => branch_target_o(29), OUT1(28) => 
                           branch_target_o(28), OUT1(27) => branch_target_o(27)
                           , OUT1(26) => branch_target_o(26), OUT1(25) => 
                           branch_target_o(25), OUT1(24) => branch_target_o(24)
                           , OUT1(23) => branch_target_o(23), OUT1(22) => 
                           branch_target_o(22), OUT1(21) => branch_target_o(21)
                           , OUT1(20) => branch_target_o(20), OUT1(19) => 
                           branch_target_o(19), OUT1(18) => branch_target_o(18)
                           , OUT1(17) => branch_target_o(17), OUT1(16) => 
                           branch_target_o(16), OUT1(15) => branch_target_o(15)
                           , OUT1(14) => branch_target_o(14), OUT1(13) => 
                           branch_target_o(13), OUT1(12) => branch_target_o(12)
                           , OUT1(11) => branch_target_o(11), OUT1(10) => 
                           branch_target_o(10), OUT1(9) => branch_target_o(9), 
                           OUT1(8) => branch_target_o(8), OUT1(7) => 
                           branch_target_o(7), OUT1(6) => branch_target_o(6), 
                           OUT1(5) => branch_target_o(5), OUT1(4) => 
                           branch_target_o(4), OUT1(3) => branch_target_o(3), 
                           OUT1(2) => branch_target_o(2), OUT1(1) => 
                           branch_target_o(1), OUT1(0) => branch_target_o(0));
   ZC : zerocheck port map( IN0(31) => A_o_31_port, IN0(30) => A_o_30_port, 
                           IN0(29) => A_o_29_port, IN0(28) => A_o_28_port, 
                           IN0(27) => A_o_27_port, IN0(26) => A_o_26_port, 
                           IN0(25) => A_o_25_port, IN0(24) => A_o_24_port, 
                           IN0(23) => A_o_23_port, IN0(22) => A_o_22_port, 
                           IN0(21) => A_o_21_port, IN0(20) => A_o_20_port, 
                           IN0(19) => A_o_19_port, IN0(18) => A_o_18_port, 
                           IN0(17) => A_o_17_port, IN0(16) => A_o_16_port, 
                           IN0(15) => A_o_15_port, IN0(14) => A_o_14_port, 
                           IN0(13) => A_o_13_port, IN0(12) => A_o_12_port, 
                           IN0(11) => A_o_11_port, IN0(10) => A_o_10_port, 
                           IN0(9) => A_o_9_port, IN0(8) => A_o_8_port, IN0(7) 
                           => A_o_7_port, IN0(6) => A_o_6_port, IN0(5) => 
                           A_o_5_port, IN0(4) => A_o_4_port, IN0(3) => 
                           A_o_3_port, IN0(2) => A_o_2_port, IN0(1) => 
                           A_o_1_port, IN0(0) => A_o_0_port, CTRL => S_EQ_NEQ_i
                           , OUT1 => branch_sel);
   MUXLINK : mux21_4 port map( IN0(31) => ext_imm_31_port, IN0(30) => 
                           ext_imm_30_port, IN0(29) => ext_imm_29_port, IN0(28)
                           => ext_imm_28_port, IN0(27) => ext_imm_31_port, 
                           IN0(26) => ext_imm_26_port, IN0(25) => 
                           ext_imm_25_port, IN0(24) => ext_imm_24_port, IN0(23)
                           => ext_imm_23_port, IN0(22) => ext_imm_22_port, 
                           IN0(21) => ext_imm_21_port, IN0(20) => 
                           ext_imm_20_port, IN0(19) => n1, IN0(18) => 
                           ext_imm_18_port, IN0(17) => ext_imm_17_port, IN0(16)
                           => ext_imm_16_port, IN0(15) => ext_imm_15_port, 
                           IN0(14) => ext_imm_14_port, IN0(13) => 
                           ext_imm_13_port, IN0(12) => ext_imm_12_port, IN0(11)
                           => ext_imm_11_port, IN0(10) => ext_imm_10_port, 
                           IN0(9) => ext_imm_9_port, IN0(8) => ext_imm_8_port, 
                           IN0(7) => ext_imm_7_port, IN0(6) => ext_imm_6_port, 
                           IN0(5) => ext_imm_5_port, IN0(4) => ext_imm_4_port, 
                           IN0(3) => ext_imm_3_port, IN0(2) => ext_imm_2_port, 
                           IN0(1) => ext_imm_1_port, IN0(0) => ext_imm_0_port, 
                           IN1(31) => NPCF_i(31), IN1(30) => NPCF_i(30), 
                           IN1(29) => NPCF_i(29), IN1(28) => NPCF_i(28), 
                           IN1(27) => NPCF_i(27), IN1(26) => NPCF_i(26), 
                           IN1(25) => NPCF_i(25), IN1(24) => NPCF_i(24), 
                           IN1(23) => NPCF_i(23), IN1(22) => NPCF_i(22), 
                           IN1(21) => NPCF_i(21), IN1(20) => NPCF_i(20), 
                           IN1(19) => NPCF_i(19), IN1(18) => NPCF_i(18), 
                           IN1(17) => NPCF_i(17), IN1(16) => NPCF_i(16), 
                           IN1(15) => NPCF_i(15), IN1(14) => NPCF_i(14), 
                           IN1(13) => NPCF_i(13), IN1(12) => NPCF_i(12), 
                           IN1(11) => NPCF_i(11), IN1(10) => NPCF_i(10), IN1(9)
                           => NPCF_i(9), IN1(8) => NPCF_i(8), IN1(7) => 
                           NPCF_i(7), IN1(6) => NPCF_i(6), IN1(5) => NPCF_i(5),
                           IN1(4) => NPCF_i(4), IN1(3) => NPCF_i(3), IN1(2) => 
                           NPCF_i(2), IN1(1) => NPCF_i(1), IN1(0) => NPCF_i(0),
                           CTRL => S_MUX_LINK_i, OUT1(31) => extended_imm(31), 
                           OUT1(30) => extended_imm(30), OUT1(29) => 
                           extended_imm(29), OUT1(28) => extended_imm(28), 
                           OUT1(27) => extended_imm(27), OUT1(26) => 
                           extended_imm(26), OUT1(25) => extended_imm(25), 
                           OUT1(24) => extended_imm(24), OUT1(23) => 
                           extended_imm(23), OUT1(22) => extended_imm(22), 
                           OUT1(21) => extended_imm(21), OUT1(20) => 
                           extended_imm(20), OUT1(19) => extended_imm(19), 
                           OUT1(18) => extended_imm(18), OUT1(17) => 
                           extended_imm(17), OUT1(16) => extended_imm(16), 
                           OUT1(15) => extended_imm(15), OUT1(14) => 
                           extended_imm(14), OUT1(13) => extended_imm(13), 
                           OUT1(12) => extended_imm(12), OUT1(11) => 
                           extended_imm(11), OUT1(10) => extended_imm(10), 
                           OUT1(9) => extended_imm(9), OUT1(8) => 
                           extended_imm(8), OUT1(7) => extended_imm(7), OUT1(6)
                           => extended_imm(6), OUT1(5) => extended_imm(5), 
                           OUT1(4) => extended_imm(4), OUT1(3) => 
                           extended_imm(3), OUT1(2) => extended_imm(2), OUT1(1)
                           => extended_imm(1), OUT1(0) => extended_imm(0));
   MUX_FWA : mux41_MUX_SIZE32 port map( IN0(31) => A_i(31), IN0(30) => A_i(30),
                           IN0(29) => A_i(29), IN0(28) => A_i(28), IN0(27) => 
                           A_i(27), IN0(26) => A_i(26), IN0(25) => A_i(25), 
                           IN0(24) => A_i(24), IN0(23) => A_i(23), IN0(22) => 
                           A_i(22), IN0(21) => A_i(21), IN0(20) => A_i(20), 
                           IN0(19) => A_i(19), IN0(18) => A_i(18), IN0(17) => 
                           A_i(17), IN0(16) => A_i(16), IN0(15) => A_i(15), 
                           IN0(14) => A_i(14), IN0(13) => A_i(13), IN0(12) => 
                           A_i(12), IN0(11) => A_i(11), IN0(10) => A_i(10), 
                           IN0(9) => A_i(9), IN0(8) => A_i(8), IN0(7) => A_i(7)
                           , IN0(6) => A_i(6), IN0(5) => A_i(5), IN0(4) => 
                           A_i(4), IN0(3) => A_i(3), IN0(2) => A_i(2), IN0(1) 
                           => A_i(1), IN0(0) => A_i(0), IN1(31) => FW_X_i(31), 
                           IN1(30) => FW_X_i(30), IN1(29) => FW_X_i(29), 
                           IN1(28) => FW_X_i(28), IN1(27) => FW_X_i(27), 
                           IN1(26) => FW_X_i(26), IN1(25) => FW_X_i(25), 
                           IN1(24) => FW_X_i(24), IN1(23) => FW_X_i(23), 
                           IN1(22) => FW_X_i(22), IN1(21) => FW_X_i(21), 
                           IN1(20) => FW_X_i(20), IN1(19) => FW_X_i(19), 
                           IN1(18) => FW_X_i(18), IN1(17) => FW_X_i(17), 
                           IN1(16) => FW_X_i(16), IN1(15) => FW_X_i(15), 
                           IN1(14) => FW_X_i(14), IN1(13) => FW_X_i(13), 
                           IN1(12) => FW_X_i(12), IN1(11) => FW_X_i(11), 
                           IN1(10) => FW_X_i(10), IN1(9) => FW_X_i(9), IN1(8) 
                           => FW_X_i(8), IN1(7) => FW_X_i(7), IN1(6) => 
                           FW_X_i(6), IN1(5) => FW_X_i(5), IN1(4) => FW_X_i(4),
                           IN1(3) => FW_X_i(3), IN1(2) => FW_X_i(2), IN1(1) => 
                           FW_X_i(1), IN1(0) => FW_X_i(0), IN2(31) => 
                           FW_W_i(31), IN2(30) => FW_W_i(30), IN2(29) => 
                           FW_W_i(29), IN2(28) => FW_W_i(28), IN2(27) => 
                           FW_W_i(27), IN2(26) => FW_W_i(26), IN2(25) => 
                           FW_W_i(25), IN2(24) => FW_W_i(24), IN2(23) => 
                           FW_W_i(23), IN2(22) => FW_W_i(22), IN2(21) => 
                           FW_W_i(21), IN2(20) => FW_W_i(20), IN2(19) => 
                           FW_W_i(19), IN2(18) => FW_W_i(18), IN2(17) => 
                           FW_W_i(17), IN2(16) => FW_W_i(16), IN2(15) => 
                           FW_W_i(15), IN2(14) => FW_W_i(14), IN2(13) => 
                           FW_W_i(13), IN2(12) => FW_W_i(12), IN2(11) => 
                           FW_W_i(11), IN2(10) => FW_W_i(10), IN2(9) => 
                           FW_W_i(9), IN2(8) => FW_W_i(8), IN2(7) => FW_W_i(7),
                           IN2(6) => FW_W_i(6), IN2(5) => FW_W_i(5), IN2(4) => 
                           FW_W_i(4), IN2(3) => FW_W_i(3), IN2(2) => FW_W_i(2),
                           IN2(1) => FW_W_i(1), IN2(0) => FW_W_i(0), IN3(31) =>
                           X_Logic0_port, IN3(30) => X_Logic0_port, IN3(29) => 
                           X_Logic0_port, IN3(28) => X_Logic0_port, IN3(27) => 
                           X_Logic0_port, IN3(26) => X_Logic0_port, IN3(25) => 
                           X_Logic0_port, IN3(24) => X_Logic0_port, IN3(23) => 
                           X_Logic0_port, IN3(22) => X_Logic0_port, IN3(21) => 
                           X_Logic0_port, IN3(20) => X_Logic0_port, IN3(19) => 
                           X_Logic0_port, IN3(18) => X_Logic0_port, IN3(17) => 
                           X_Logic0_port, IN3(16) => X_Logic0_port, IN3(15) => 
                           X_Logic0_port, IN3(14) => X_Logic0_port, IN3(13) => 
                           X_Logic0_port, IN3(12) => X_Logic0_port, IN3(11) => 
                           X_Logic0_port, IN3(10) => X_Logic0_port, IN3(9) => 
                           X_Logic0_port, IN3(8) => X_Logic0_port, IN3(7) => 
                           X_Logic0_port, IN3(6) => X_Logic0_port, IN3(5) => 
                           X_Logic0_port, IN3(4) => X_Logic0_port, IN3(3) => 
                           X_Logic0_port, IN3(2) => X_Logic0_port, IN3(1) => 
                           X_Logic0_port, IN3(0) => X_Logic0_port, CTRL(1) => 
                           S_FW_Adec_i(1), CTRL(0) => S_FW_Adec_i(0), OUT1(31) 
                           => A_o_31_port, OUT1(30) => A_o_30_port, OUT1(29) =>
                           A_o_29_port, OUT1(28) => A_o_28_port, OUT1(27) => 
                           A_o_27_port, OUT1(26) => A_o_26_port, OUT1(25) => 
                           A_o_25_port, OUT1(24) => A_o_24_port, OUT1(23) => 
                           A_o_23_port, OUT1(22) => A_o_22_port, OUT1(21) => 
                           A_o_21_port, OUT1(20) => A_o_20_port, OUT1(19) => 
                           A_o_19_port, OUT1(18) => A_o_18_port, OUT1(17) => 
                           A_o_17_port, OUT1(16) => A_o_16_port, OUT1(15) => 
                           A_o_15_port, OUT1(14) => A_o_14_port, OUT1(13) => 
                           A_o_13_port, OUT1(12) => A_o_12_port, OUT1(11) => 
                           A_o_11_port, OUT1(10) => A_o_10_port, OUT1(9) => 
                           A_o_9_port, OUT1(8) => A_o_8_port, OUT1(7) => 
                           A_o_7_port, OUT1(6) => A_o_6_port, OUT1(5) => 
                           A_o_5_port, OUT1(4) => A_o_4_port, OUT1(3) => 
                           A_o_3_port, OUT1(2) => A_o_2_port, OUT1(1) => 
                           A_o_1_port, OUT1(0) => A_o_0_port);
   U2 : CLKBUF_X1 port map( A => branch_sel, Z => n2);
   U3 : INV_X1 port map( A => n2, ZN => taken_o);
   n4 <= '0';
   n5 <= '0';
   n6 <= '0';
   n7 <= '0';
   n8 <= '0';
   n9 <= '0';

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity fetch_regs is

   port( NPCF_i, IR_i : in std_logic_vector (31 downto 0);  NPCF_o, IR_o : out 
         std_logic_vector (31 downto 0);  stall_i, clk, rst : in std_logic);

end fetch_regs;

architecture SYN_struct of fetch_regs is

   component INV_X4
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component ff32_en_IR
      port( D : in std_logic_vector (31 downto 0);  en, clk, rst : in std_logic
            ;  Q : out std_logic_vector (31 downto 0));
   end component;
   
   component ff32_en_1
      port( D : in std_logic_vector (31 downto 0);  en, clk, rst : in std_logic
            ;  Q : out std_logic_vector (31 downto 0));
   end component;
   
   signal n2 : std_logic;

begin
   
   NPCF : ff32_en_1 port map( D(31) => NPCF_i(31), D(30) => NPCF_i(30), D(29) 
                           => NPCF_i(29), D(28) => NPCF_i(28), D(27) => 
                           NPCF_i(27), D(26) => NPCF_i(26), D(25) => NPCF_i(25)
                           , D(24) => NPCF_i(24), D(23) => NPCF_i(23), D(22) =>
                           NPCF_i(22), D(21) => NPCF_i(21), D(20) => NPCF_i(20)
                           , D(19) => NPCF_i(19), D(18) => NPCF_i(18), D(17) =>
                           NPCF_i(17), D(16) => NPCF_i(16), D(15) => NPCF_i(15)
                           , D(14) => NPCF_i(14), D(13) => NPCF_i(13), D(12) =>
                           NPCF_i(12), D(11) => NPCF_i(11), D(10) => NPCF_i(10)
                           , D(9) => NPCF_i(9), D(8) => NPCF_i(8), D(7) => 
                           NPCF_i(7), D(6) => NPCF_i(6), D(5) => NPCF_i(5), 
                           D(4) => NPCF_i(4), D(3) => NPCF_i(3), D(2) => 
                           NPCF_i(2), D(1) => NPCF_i(1), D(0) => NPCF_i(0), en 
                           => n2, clk => clk, rst => rst, Q(31) => NPCF_o(31), 
                           Q(30) => NPCF_o(30), Q(29) => NPCF_o(29), Q(28) => 
                           NPCF_o(28), Q(27) => NPCF_o(27), Q(26) => NPCF_o(26)
                           , Q(25) => NPCF_o(25), Q(24) => NPCF_o(24), Q(23) =>
                           NPCF_o(23), Q(22) => NPCF_o(22), Q(21) => NPCF_o(21)
                           , Q(20) => NPCF_o(20), Q(19) => NPCF_o(19), Q(18) =>
                           NPCF_o(18), Q(17) => NPCF_o(17), Q(16) => NPCF_o(16)
                           , Q(15) => NPCF_o(15), Q(14) => NPCF_o(14), Q(13) =>
                           NPCF_o(13), Q(12) => NPCF_o(12), Q(11) => NPCF_o(11)
                           , Q(10) => NPCF_o(10), Q(9) => NPCF_o(9), Q(8) => 
                           NPCF_o(8), Q(7) => NPCF_o(7), Q(6) => NPCF_o(6), 
                           Q(5) => NPCF_o(5), Q(4) => NPCF_o(4), Q(3) => 
                           NPCF_o(3), Q(2) => NPCF_o(2), Q(1) => NPCF_o(1), 
                           Q(0) => NPCF_o(0));
   IR : ff32_en_IR port map( D(31) => IR_i(31), D(30) => IR_i(30), D(29) => 
                           IR_i(29), D(28) => IR_i(28), D(27) => IR_i(27), 
                           D(26) => IR_i(26), D(25) => IR_i(25), D(24) => 
                           IR_i(24), D(23) => IR_i(23), D(22) => IR_i(22), 
                           D(21) => IR_i(21), D(20) => IR_i(20), D(19) => 
                           IR_i(19), D(18) => IR_i(18), D(17) => IR_i(17), 
                           D(16) => IR_i(16), D(15) => IR_i(15), D(14) => 
                           IR_i(14), D(13) => IR_i(13), D(12) => IR_i(12), 
                           D(11) => IR_i(11), D(10) => IR_i(10), D(9) => 
                           IR_i(9), D(8) => IR_i(8), D(7) => IR_i(7), D(6) => 
                           IR_i(6), D(5) => IR_i(5), D(4) => IR_i(4), D(3) => 
                           IR_i(3), D(2) => IR_i(2), D(1) => IR_i(1), D(0) => 
                           IR_i(0), en => n2, clk => clk, rst => rst, Q(31) => 
                           IR_o(31), Q(30) => IR_o(30), Q(29) => IR_o(29), 
                           Q(28) => IR_o(28), Q(27) => IR_o(27), Q(26) => 
                           IR_o(26), Q(25) => IR_o(25), Q(24) => IR_o(24), 
                           Q(23) => IR_o(23), Q(22) => IR_o(22), Q(21) => 
                           IR_o(21), Q(20) => IR_o(20), Q(19) => IR_o(19), 
                           Q(18) => IR_o(18), Q(17) => IR_o(17), Q(16) => 
                           IR_o(16), Q(15) => IR_o(15), Q(14) => IR_o(14), 
                           Q(13) => IR_o(13), Q(12) => IR_o(12), Q(11) => 
                           IR_o(11), Q(10) => IR_o(10), Q(9) => IR_o(9), Q(8) 
                           => IR_o(8), Q(7) => IR_o(7), Q(6) => IR_o(6), Q(5) 
                           => IR_o(5), Q(4) => IR_o(4), Q(3) => IR_o(3), Q(2) 
                           => IR_o(2), Q(1) => IR_o(1), Q(0) => IR_o(0));
   U1 : INV_X4 port map( A => stall_i, ZN => n2);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity btb_N_LINES4_SIZE32 is

   port( clock, reset, stall_i : in std_logic;  TAG_i : in std_logic_vector (3 
         downto 0);  target_PC_i : in std_logic_vector (31 downto 0);  
         was_taken_i : in std_logic;  predicted_next_PC_o : out 
         std_logic_vector (31 downto 0);  taken_o, mispredict_o : out std_logic
         );

end btb_N_LINES4_SIZE32;

architecture SYN_bhe of btb_N_LINES4_SIZE32 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component predictor_2_1
      port( clock, reset, enable, taken_i : in std_logic;  prediction_o : out 
            std_logic);
   end component;
   
   component predictor_2_2
      port( clock, reset, enable, taken_i : in std_logic;  prediction_o : out 
            std_logic);
   end component;
   
   component predictor_2_3
      port( clock, reset, enable, taken_i : in std_logic;  prediction_o : out 
            std_logic);
   end component;
   
   component predictor_2_4
      port( clock, reset, enable, taken_i : in std_logic;  prediction_o : out 
            std_logic);
   end component;
   
   component predictor_2_5
      port( clock, reset, enable, taken_i : in std_logic;  prediction_o : out 
            std_logic);
   end component;
   
   component predictor_2_6
      port( clock, reset, enable, taken_i : in std_logic;  prediction_o : out 
            std_logic);
   end component;
   
   component predictor_2_7
      port( clock, reset, enable, taken_i : in std_logic;  prediction_o : out 
            std_logic);
   end component;
   
   component predictor_2_8
      port( clock, reset, enable, taken_i : in std_logic;  prediction_o : out 
            std_logic);
   end component;
   
   component predictor_2_9
      port( clock, reset, enable, taken_i : in std_logic;  prediction_o : out 
            std_logic);
   end component;
   
   component predictor_2_10
      port( clock, reset, enable, taken_i : in std_logic;  prediction_o : out 
            std_logic);
   end component;
   
   component predictor_2_11
      port( clock, reset, enable, taken_i : in std_logic;  prediction_o : out 
            std_logic);
   end component;
   
   component predictor_2_12
      port( clock, reset, enable, taken_i : in std_logic;  prediction_o : out 
            std_logic);
   end component;
   
   component predictor_2_13
      port( clock, reset, enable, taken_i : in std_logic;  prediction_o : out 
            std_logic);
   end component;
   
   component predictor_2_14
      port( clock, reset, enable, taken_i : in std_logic;  prediction_o : out 
            std_logic);
   end component;
   
   component predictor_2_15
      port( clock, reset, enable, taken_i : in std_logic;  prediction_o : out 
            std_logic);
   end component;
   
   component predictor_2_0
      port( clock, reset, enable, taken_i : in std_logic;  prediction_o : out 
            std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal predicted_next_PC_o_31_port, predicted_next_PC_o_30_port, 
      predicted_next_PC_o_29_port, predicted_next_PC_o_28_port, 
      predicted_next_PC_o_27_port, predicted_next_PC_o_26_port, 
      predicted_next_PC_o_25_port, predicted_next_PC_o_24_port, 
      predicted_next_PC_o_23_port, predicted_next_PC_o_22_port, 
      predicted_next_PC_o_21_port, predicted_next_PC_o_20_port, 
      predicted_next_PC_o_19_port, predicted_next_PC_o_18_port, 
      predicted_next_PC_o_17_port, predicted_next_PC_o_16_port, 
      predicted_next_PC_o_15_port, predicted_next_PC_o_14_port, 
      predicted_next_PC_o_13_port, predicted_next_PC_o_12_port, 
      predicted_next_PC_o_11_port, predicted_next_PC_o_10_port, 
      predicted_next_PC_o_9_port, predicted_next_PC_o_8_port, 
      predicted_next_PC_o_7_port, predicted_next_PC_o_6_port, 
      predicted_next_PC_o_5_port, predicted_next_PC_o_4_port, 
      predicted_next_PC_o_3_port, predicted_next_PC_o_2_port, 
      predicted_next_PC_o_1_port, predicted_next_PC_o_0_port, taken_o_port, 
      mispredict_o_port, taken_15_port, taken_14_port, taken_13_port, 
      taken_12_port, taken_11_port, taken_10_port, taken_9_port, taken_8_port, 
      taken_7_port, taken_6_port, taken_5_port, taken_4_port, taken_3_port, 
      taken_2_port, taken_1_port, taken_0_port, write_enable_15_port, 
      write_enable_14_port, write_enable_13_port, write_enable_12_port, 
      write_enable_11_port, write_enable_10_port, write_enable_9_port, 
      write_enable_8_port, write_enable_7_port, write_enable_6_port, 
      write_enable_5_port, write_enable_4_port, write_enable_3_port, 
      write_enable_2_port, write_enable_1_port, write_enable_0_port, 
      predict_PC_0_31_port, predict_PC_0_30_port, predict_PC_0_29_port, 
      predict_PC_0_28_port, predict_PC_0_27_port, predict_PC_0_26_port, 
      predict_PC_0_25_port, predict_PC_0_24_port, predict_PC_0_23_port, 
      predict_PC_0_22_port, predict_PC_0_21_port, predict_PC_0_20_port, 
      predict_PC_0_19_port, predict_PC_0_18_port, predict_PC_0_17_port, 
      predict_PC_0_16_port, predict_PC_0_15_port, predict_PC_0_14_port, 
      predict_PC_0_13_port, predict_PC_0_12_port, predict_PC_0_11_port, 
      predict_PC_0_10_port, predict_PC_0_9_port, predict_PC_0_8_port, 
      predict_PC_0_7_port, predict_PC_0_6_port, predict_PC_0_5_port, 
      predict_PC_0_4_port, predict_PC_0_3_port, predict_PC_0_2_port, 
      predict_PC_0_1_port, predict_PC_0_0_port, predict_PC_1_31_port, 
      predict_PC_1_30_port, predict_PC_1_29_port, predict_PC_1_28_port, 
      predict_PC_1_27_port, predict_PC_1_26_port, predict_PC_1_25_port, 
      predict_PC_1_24_port, predict_PC_1_23_port, predict_PC_1_22_port, 
      predict_PC_1_21_port, predict_PC_1_20_port, predict_PC_1_19_port, 
      predict_PC_1_18_port, predict_PC_1_17_port, predict_PC_1_16_port, 
      predict_PC_1_15_port, predict_PC_1_14_port, predict_PC_1_13_port, 
      predict_PC_1_12_port, predict_PC_1_11_port, predict_PC_1_10_port, 
      predict_PC_1_9_port, predict_PC_1_8_port, predict_PC_1_7_port, 
      predict_PC_1_6_port, predict_PC_1_5_port, predict_PC_1_4_port, 
      predict_PC_1_3_port, predict_PC_1_2_port, predict_PC_1_1_port, 
      predict_PC_1_0_port, predict_PC_2_31_port, predict_PC_2_30_port, 
      predict_PC_2_29_port, predict_PC_2_28_port, predict_PC_2_27_port, 
      predict_PC_2_26_port, predict_PC_2_25_port, predict_PC_2_24_port, 
      predict_PC_2_23_port, predict_PC_2_22_port, predict_PC_2_21_port, 
      predict_PC_2_20_port, predict_PC_2_19_port, predict_PC_2_18_port, 
      predict_PC_2_17_port, predict_PC_2_16_port, predict_PC_2_15_port, 
      predict_PC_2_14_port, predict_PC_2_13_port, predict_PC_2_12_port, 
      predict_PC_2_11_port, predict_PC_2_10_port, predict_PC_2_9_port, 
      predict_PC_2_8_port, predict_PC_2_7_port, predict_PC_2_6_port, 
      predict_PC_2_5_port, predict_PC_2_4_port, predict_PC_2_3_port, 
      predict_PC_2_2_port, predict_PC_2_1_port, predict_PC_2_0_port, 
      predict_PC_3_31_port, predict_PC_3_30_port, predict_PC_3_29_port, 
      predict_PC_3_28_port, predict_PC_3_27_port, predict_PC_3_26_port, 
      predict_PC_3_25_port, predict_PC_3_24_port, predict_PC_3_23_port, 
      predict_PC_3_22_port, predict_PC_3_21_port, predict_PC_3_20_port, 
      predict_PC_3_19_port, predict_PC_3_18_port, predict_PC_3_17_port, 
      predict_PC_3_16_port, predict_PC_3_15_port, predict_PC_3_14_port, 
      predict_PC_3_13_port, predict_PC_3_12_port, predict_PC_3_11_port, 
      predict_PC_3_10_port, predict_PC_3_9_port, predict_PC_3_8_port, 
      predict_PC_3_7_port, predict_PC_3_6_port, predict_PC_3_5_port, 
      predict_PC_3_4_port, predict_PC_3_3_port, predict_PC_3_2_port, 
      predict_PC_3_1_port, predict_PC_3_0_port, predict_PC_4_31_port, 
      predict_PC_4_30_port, predict_PC_4_29_port, predict_PC_4_28_port, 
      predict_PC_4_27_port, predict_PC_4_26_port, predict_PC_4_25_port, 
      predict_PC_4_24_port, predict_PC_4_23_port, predict_PC_4_22_port, 
      predict_PC_4_21_port, predict_PC_4_20_port, predict_PC_4_19_port, 
      predict_PC_4_18_port, predict_PC_4_17_port, predict_PC_4_16_port, 
      predict_PC_4_15_port, predict_PC_4_14_port, predict_PC_4_13_port, 
      predict_PC_4_12_port, predict_PC_4_11_port, predict_PC_4_10_port, 
      predict_PC_4_9_port, predict_PC_4_8_port, predict_PC_4_7_port, 
      predict_PC_4_6_port, predict_PC_4_5_port, predict_PC_4_4_port, 
      predict_PC_4_3_port, predict_PC_4_2_port, predict_PC_4_1_port, 
      predict_PC_4_0_port, predict_PC_5_31_port, predict_PC_5_30_port, 
      predict_PC_5_29_port, predict_PC_5_28_port, predict_PC_5_27_port, 
      predict_PC_5_26_port, predict_PC_5_25_port, predict_PC_5_24_port, 
      predict_PC_5_23_port, predict_PC_5_22_port, predict_PC_5_21_port, 
      predict_PC_5_20_port, predict_PC_5_19_port, predict_PC_5_18_port, 
      predict_PC_5_17_port, predict_PC_5_16_port, predict_PC_5_15_port, 
      predict_PC_5_14_port, predict_PC_5_13_port, predict_PC_5_12_port, 
      predict_PC_5_11_port, predict_PC_5_10_port, predict_PC_5_9_port, 
      predict_PC_5_8_port, predict_PC_5_7_port, predict_PC_5_6_port, 
      predict_PC_5_5_port, predict_PC_5_4_port, predict_PC_5_3_port, 
      predict_PC_5_2_port, predict_PC_5_1_port, predict_PC_5_0_port, 
      predict_PC_6_31_port, predict_PC_6_30_port, predict_PC_6_29_port, 
      predict_PC_6_28_port, predict_PC_6_27_port, predict_PC_6_26_port, 
      predict_PC_6_25_port, predict_PC_6_24_port, predict_PC_6_23_port, 
      predict_PC_6_22_port, predict_PC_6_21_port, predict_PC_6_20_port, 
      predict_PC_6_19_port, predict_PC_6_18_port, predict_PC_6_17_port, 
      predict_PC_6_16_port, predict_PC_6_15_port, predict_PC_6_14_port, 
      predict_PC_6_13_port, predict_PC_6_12_port, predict_PC_6_11_port, 
      predict_PC_6_10_port, predict_PC_6_9_port, predict_PC_6_8_port, 
      predict_PC_6_7_port, predict_PC_6_6_port, predict_PC_6_5_port, 
      predict_PC_6_4_port, predict_PC_6_3_port, predict_PC_6_2_port, 
      predict_PC_6_1_port, predict_PC_6_0_port, predict_PC_7_31_port, 
      predict_PC_7_30_port, predict_PC_7_29_port, predict_PC_7_28_port, 
      predict_PC_7_27_port, predict_PC_7_26_port, predict_PC_7_25_port, 
      predict_PC_7_24_port, predict_PC_7_23_port, predict_PC_7_22_port, 
      predict_PC_7_21_port, predict_PC_7_20_port, predict_PC_7_19_port, 
      predict_PC_7_18_port, predict_PC_7_17_port, predict_PC_7_16_port, 
      predict_PC_7_15_port, predict_PC_7_14_port, predict_PC_7_13_port, 
      predict_PC_7_12_port, predict_PC_7_11_port, predict_PC_7_10_port, 
      predict_PC_7_9_port, predict_PC_7_8_port, predict_PC_7_7_port, 
      predict_PC_7_6_port, predict_PC_7_5_port, predict_PC_7_4_port, 
      predict_PC_7_3_port, predict_PC_7_2_port, predict_PC_7_1_port, 
      predict_PC_7_0_port, predict_PC_8_31_port, predict_PC_8_30_port, 
      predict_PC_8_29_port, predict_PC_8_28_port, predict_PC_8_27_port, 
      predict_PC_8_26_port, predict_PC_8_25_port, predict_PC_8_24_port, 
      predict_PC_8_23_port, predict_PC_8_22_port, predict_PC_8_21_port, 
      predict_PC_8_20_port, predict_PC_8_19_port, predict_PC_8_18_port, 
      predict_PC_8_17_port, predict_PC_8_16_port, predict_PC_8_15_port, 
      predict_PC_8_14_port, predict_PC_8_13_port, predict_PC_8_12_port, 
      predict_PC_8_11_port, predict_PC_8_10_port, predict_PC_8_9_port, 
      predict_PC_8_8_port, predict_PC_8_7_port, predict_PC_8_6_port, 
      predict_PC_8_5_port, predict_PC_8_4_port, predict_PC_8_3_port, 
      predict_PC_8_2_port, predict_PC_8_1_port, predict_PC_8_0_port, 
      predict_PC_9_31_port, predict_PC_9_30_port, predict_PC_9_29_port, 
      predict_PC_9_28_port, predict_PC_9_27_port, predict_PC_9_26_port, 
      predict_PC_9_25_port, predict_PC_9_24_port, predict_PC_9_23_port, 
      predict_PC_9_22_port, predict_PC_9_21_port, predict_PC_9_20_port, 
      predict_PC_9_19_port, predict_PC_9_18_port, predict_PC_9_17_port, 
      predict_PC_9_16_port, predict_PC_9_15_port, predict_PC_9_14_port, 
      predict_PC_9_13_port, predict_PC_9_12_port, predict_PC_9_11_port, 
      predict_PC_9_10_port, predict_PC_9_9_port, predict_PC_9_8_port, 
      predict_PC_9_7_port, predict_PC_9_6_port, predict_PC_9_5_port, 
      predict_PC_9_4_port, predict_PC_9_3_port, predict_PC_9_2_port, 
      predict_PC_9_1_port, predict_PC_9_0_port, predict_PC_10_31_port, 
      predict_PC_10_30_port, predict_PC_10_29_port, predict_PC_10_28_port, 
      predict_PC_10_27_port, predict_PC_10_26_port, predict_PC_10_25_port, 
      predict_PC_10_24_port, predict_PC_10_23_port, predict_PC_10_22_port, 
      predict_PC_10_21_port, predict_PC_10_20_port, predict_PC_10_19_port, 
      predict_PC_10_18_port, predict_PC_10_17_port, predict_PC_10_16_port, 
      predict_PC_10_15_port, predict_PC_10_14_port, predict_PC_10_13_port, 
      predict_PC_10_12_port, predict_PC_10_11_port, predict_PC_10_10_port, 
      predict_PC_10_9_port, predict_PC_10_8_port, predict_PC_10_7_port, 
      predict_PC_10_6_port, predict_PC_10_5_port, predict_PC_10_4_port, 
      predict_PC_10_3_port, predict_PC_10_2_port, predict_PC_10_1_port, 
      predict_PC_10_0_port, predict_PC_11_31_port, predict_PC_11_30_port, 
      predict_PC_11_29_port, predict_PC_11_28_port, predict_PC_11_27_port, 
      predict_PC_11_26_port, predict_PC_11_25_port, predict_PC_11_24_port, 
      predict_PC_11_23_port, predict_PC_11_22_port, predict_PC_11_21_port, 
      predict_PC_11_20_port, predict_PC_11_19_port, predict_PC_11_18_port, 
      predict_PC_11_17_port, predict_PC_11_16_port, predict_PC_11_15_port, 
      predict_PC_11_14_port, predict_PC_11_13_port, predict_PC_11_12_port, 
      predict_PC_11_11_port, predict_PC_11_10_port, predict_PC_11_9_port, 
      predict_PC_11_8_port, predict_PC_11_7_port, predict_PC_11_6_port, 
      predict_PC_11_5_port, predict_PC_11_4_port, predict_PC_11_3_port, 
      predict_PC_11_2_port, predict_PC_11_1_port, predict_PC_11_0_port, 
      predict_PC_12_31_port, predict_PC_12_30_port, predict_PC_12_29_port, 
      predict_PC_12_28_port, predict_PC_12_27_port, predict_PC_12_26_port, 
      predict_PC_12_25_port, predict_PC_12_24_port, predict_PC_12_23_port, 
      predict_PC_12_22_port, predict_PC_12_21_port, predict_PC_12_20_port, 
      predict_PC_12_19_port, predict_PC_12_18_port, predict_PC_12_17_port, 
      predict_PC_12_16_port, predict_PC_12_15_port, predict_PC_12_14_port, 
      predict_PC_12_13_port, predict_PC_12_12_port, predict_PC_12_11_port, 
      predict_PC_12_10_port, predict_PC_12_9_port, predict_PC_12_8_port, 
      predict_PC_12_7_port, predict_PC_12_6_port, predict_PC_12_5_port, 
      predict_PC_12_4_port, predict_PC_12_3_port, predict_PC_12_2_port, 
      predict_PC_12_1_port, predict_PC_12_0_port, predict_PC_13_31_port, 
      predict_PC_13_30_port, predict_PC_13_29_port, predict_PC_13_28_port, 
      predict_PC_13_27_port, predict_PC_13_26_port, predict_PC_13_25_port, 
      predict_PC_13_24_port, predict_PC_13_23_port, predict_PC_13_22_port, 
      predict_PC_13_21_port, predict_PC_13_20_port, predict_PC_13_19_port, 
      predict_PC_13_18_port, predict_PC_13_17_port, predict_PC_13_16_port, 
      predict_PC_13_15_port, predict_PC_13_14_port, predict_PC_13_13_port, 
      predict_PC_13_12_port, predict_PC_13_11_port, predict_PC_13_10_port, 
      predict_PC_13_9_port, predict_PC_13_8_port, predict_PC_13_7_port, 
      predict_PC_13_6_port, predict_PC_13_5_port, predict_PC_13_4_port, 
      predict_PC_13_3_port, predict_PC_13_2_port, predict_PC_13_1_port, 
      predict_PC_13_0_port, predict_PC_14_31_port, predict_PC_14_30_port, 
      predict_PC_14_29_port, predict_PC_14_28_port, predict_PC_14_27_port, 
      predict_PC_14_26_port, predict_PC_14_25_port, predict_PC_14_24_port, 
      predict_PC_14_23_port, predict_PC_14_22_port, predict_PC_14_21_port, 
      predict_PC_14_20_port, predict_PC_14_19_port, predict_PC_14_18_port, 
      predict_PC_14_17_port, predict_PC_14_16_port, predict_PC_14_15_port, 
      predict_PC_14_14_port, predict_PC_14_13_port, predict_PC_14_12_port, 
      predict_PC_14_11_port, predict_PC_14_10_port, predict_PC_14_9_port, 
      predict_PC_14_8_port, predict_PC_14_7_port, predict_PC_14_6_port, 
      predict_PC_14_5_port, predict_PC_14_4_port, predict_PC_14_3_port, 
      predict_PC_14_2_port, predict_PC_14_1_port, predict_PC_14_0_port, 
      predict_PC_15_31_port, predict_PC_15_30_port, predict_PC_15_29_port, 
      predict_PC_15_28_port, predict_PC_15_27_port, predict_PC_15_26_port, 
      predict_PC_15_25_port, predict_PC_15_24_port, predict_PC_15_23_port, 
      predict_PC_15_22_port, predict_PC_15_21_port, predict_PC_15_20_port, 
      predict_PC_15_19_port, predict_PC_15_18_port, predict_PC_15_17_port, 
      predict_PC_15_16_port, predict_PC_15_15_port, predict_PC_15_14_port, 
      predict_PC_15_13_port, predict_PC_15_12_port, predict_PC_15_11_port, 
      predict_PC_15_10_port, predict_PC_15_9_port, predict_PC_15_8_port, 
      predict_PC_15_7_port, predict_PC_15_6_port, predict_PC_15_5_port, 
      predict_PC_15_4_port, predict_PC_15_3_port, predict_PC_15_2_port, 
      predict_PC_15_1_port, predict_PC_15_0_port, n1535, n1536, n1537, n1538, 
      n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, 
      n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, 
      n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, 
      n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, 
      n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, 
      n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, 
      n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, 
      n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, 
      n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, 
      n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, 
      n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, 
      n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, 
      n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, 
      n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, 
      n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, 
      n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, 
      n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, 
      n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, 
      n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, 
      n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, 
      n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, 
      n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, 
      n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, 
      n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, 
      n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, 
      n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, 
      n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, 
      n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, 
      n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, 
      n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, 
      n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, 
      n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, 
      n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, 
      n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, 
      n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, 
      n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, 
      n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, 
      n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, 
      n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, 
      n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, 
      n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, 
      n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, 
      n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, 
      n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, 
      n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, 
      n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, 
      n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, 
      n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, 
      n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, 
      n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, 
      n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, 
      n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, 
      n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, 
      n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, 
      n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, 
      n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, 
      n2099, n2100, n6, n7, n8, n9, n588, n589, n590, n591, n592, n593, n598, 
      n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, 
      n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, 
      n623, n624, net643832, net643833, net643834, net643835, net643836, 
      net643837, net643838, net643839, net643840, net643841, net643842, 
      net643843, net643844, net643845, net643846, net643847, net643848, 
      net643849, net643850, net643851, net643852, net643853, net643854, 
      net643855, net643856, net643857, net643858, net643859, net643860, 
      net643861, net643862, net643863, net643864, net643865, net643866, 
      net643867, net643868, net643869, net643870, net643871, net643872, 
      net643873, net643874, net643875, net643876, net643877, net643878, 
      net643879, net643880, net643881, net643882, net643883, net643884, 
      net643885, net643886, net643887, net643888, net643889, net643890, 
      net643891, net643892, net643893, net643894, net643895, net643896, 
      net643897, net643898, net643899, net643900, net643901, net643902, 
      net643903, net643904, net643905, net643906, net643907, net643908, 
      net643909, net643910, net643911, net643912, net643913, net643914, 
      net643915, net643916, net643917, net643918, net643919, net643920, 
      net643921, net643922, net643923, net643924, net643925, net643926, 
      net643927, net643928, net643929, net643930, net643931, net643932, 
      net643933, net643934, net643935, net643936, net643937, net643938, 
      net643939, net643940, net643941, net643942, net643943, net643944, 
      net643945, net643946, net643947, net643948, net643949, net643950, 
      net643951, net643952, net643953, net643954, net643955, net643956, 
      net643957, net643958, net643959, net643960, net643961, net643962, 
      net643963, net643964, net643965, net643966, net643967, net643968, 
      net643969, net643970, net643971, net643972, net643973, net643974, 
      net643975, net643976, net643977, net643978, net643979, net643980, 
      net643981, net643982, net643983, net643984, net643985, net643986, 
      net643987, net643988, net643989, net643990, net643991, net643992, 
      net643993, net643994, net643995, net643996, net643997, net643998, 
      net643999, net644000, net644001, net644002, net644003, net644004, 
      net644005, net644006, net644007, net644008, net644009, net644010, 
      net644011, net644012, net644013, net644014, net644015, net644016, 
      net644017, net644018, net644019, net644020, net644021, net644022, 
      net644023, net644024, net644025, net644026, net644027, net644028, 
      net644029, net644030, net644031, net644032, net644033, net644034, 
      net644035, net644036, net644037, net644038, net644039, net644040, 
      net644041, net644042, net644043, net644044, net644045, net644046, 
      net644047, net644048, net644049, net644050, net644051, net644052, 
      net644053, net644054, net644055, net644056, net644057, net644058, 
      net644059, net644060, net644061, net644062, net644063, net644064, 
      net644065, net644066, net644067, net644068, net644069, net644070, 
      net644071, net644072, net644073, net644074, net644075, net644076, 
      net644077, net644078, net644079, net644080, net644081, net644082, 
      net644083, net644084, net644085, net644086, net644087, net644088, 
      net644089, net644090, net644091, net644092, net644093, net644094, 
      net644095, net644096, net644097, net644098, net644099, net644100, 
      net644101, net644102, net644103, net644104, net644105, net644106, 
      net644107, net644108, net644109, net644110, net644111, net644112, 
      net644113, net644114, net644115, net644116, net644117, net644118, 
      net644119, net644120, net644121, net644122, net644123, net644124, 
      net644125, net644126, net644127, net644128, net644129, net644130, 
      net644131, net644132, net644133, net644134, net644135, net644136, 
      net644137, net644138, net644139, net644140, net644141, net644142, 
      net644143, net644144, net644145, net644146, net644147, net644148, 
      net644149, net644150, net644151, net644152, net644153, net644154, 
      net644155, net644156, net644157, net644158, net644159, net644160, 
      net644161, net644162, net644163, net644164, net644165, net644166, 
      net644167, net644168, net644169, net644170, net644171, net644172, 
      net644173, net644174, net644175, net644176, net644177, net644178, 
      net644179, net644180, net644181, net644182, net644183, net644184, 
      net644185, net644186, net644187, net644188, net644189, net644190, 
      net644191, net644192, net644193, net644194, net644195, net644196, 
      net644197, net644198, net644199, net644200, net644201, net644202, 
      net644203, net644204, net644205, net644206, net644207, net644208, 
      net644209, net644210, net644211, net644212, net644213, net644214, 
      net644215, net644216, net644217, net644218, net644219, net644220, 
      net644221, net644222, net644223, net644224, net644225, net644226, 
      net644227, net644228, net644229, net644230, net644231, net644232, 
      net644233, net644234, net644235, net644236, net644237, net644238, 
      net644239, net644240, net644241, net644242, net644243, net644244, 
      net644245, net644246, net644247, net644248, net644249, net644250, 
      net644251, net644252, net644253, net644254, net644255, net644256, 
      net644257, net644258, net644259, net644260, net644261, net644262, 
      net644263, net644264, net644265, net644266, net644267, net644268, 
      net644269, net644270, net644271, net644272, net644273, net644274, 
      net644275, net644276, net644277, net644278, net644279, net644280, 
      net644281, net644282, net644283, net644284, net644285, net644286, 
      net644287, net644288, net644289, net644290, net644291, net644292, 
      net644293, net644294, net644295, net644296, net644297, net644298, 
      net644299, net644300, net644301, net644302, net644303, net644304, 
      net644305, net644306, net644307, net644308, net644309, net644310, 
      net644311, net644312, net644313, net644314, net644315, net644316, 
      net644317, net644318, net644319, net644320, net644321, net644322, 
      net644323, net644324, net644325, net644326, net644327, net644328, 
      net644329, net644330, net644331, net644332, net644333, net644334, 
      net644335, net644336, net644337, net644338, net644339, net644340, 
      net644341, net644342, net644343, net644344, n666, n667, n668, n669, n670,
      n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, 
      n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n696, 
      n697, n699, n701, n703, n736, n738, n739, n740, n741, n742, n743, n744, 
      n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, 
      n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, 
      n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, 
      n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, 
      n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, 
      n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, 
      n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, 
      n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, 
      n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, 
      n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, 
      n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, 
      n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, 
      n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, 
      n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, 
      n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, 
      n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, 
      n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, 
      n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, 
      n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, 
      n973, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, 
      n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, 
      n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, 
      n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, 
      n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, 
      n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, 
      n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, 
      n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, 
      n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, 
      n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, 
      n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, 
      n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, 
      n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, 
      n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, 
      n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, 
      n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, 
      n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, 
      n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, 
      n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, 
      n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, 
      n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, 
      n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, 
      n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, 
      n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, 
      n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, 
      n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, 
      n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, 
      n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, 
      n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, 
      n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, 
      n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, 
      n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, 
      n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, 
      n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, 
      n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, 
      n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, 
      n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, 
      n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, 
      n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, 
      n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, 
      n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, 
      n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, 
      n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, 
      n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, 
      n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, 
      n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, 
      n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, 
      n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, 
      n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, 
      n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, 
      n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, 
      n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, 
      n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, 
      n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, 
      n1531, n1532, n1533, n1534, n2101, n2102, n2103, n2104, n2105, n2106, 
      n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, 
      n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, 
      n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, 
      n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, 
      n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, 
      n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, 
      n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, 
      n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, 
      n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, 
      n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, 
      n2207, n2208, n2209, n2210, n2221, n2222, n2224, n2225, n2252, n2251, 
      n2250, n2249, n2248, n2247, n2246, n2245, n2244, n2243, n2242, n2241, 
      n2240, n2239, n2238, n2237, n2236, n2235, n2234, n2233, n2232, n2231, 
      n2230, n2229, n2228, n2227, n2226, n2223, n2220, n2219, n2218, n2217, 
      n2212, n2211, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
      n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, 
      n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, 
      n664, n665, n694, n695, n698, n700, n702, n704, n705, n706, n707, n708, 
      n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, 
      n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, 
      n733, n734, n735, n737, n974, n975, n976, n977, n978, n979, n980, n981, 
      n982, n983, n984, n985, n986, n987, n988, n989, n2213, n2214, n2215, 
      n2216, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, 
      n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, 
      n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, 
      n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, 
      n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, 
      n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, 
      net684125, net684126, net684127, net684128, net684129, net684130, 
      net684131, net684132, net684133, net684134, net684135, net684136, 
      net684137, net684138, net684139, net684140, net684141, net684142, 
      net684143, net684144, net684145, net684146, net684147, net684148, 
      net684149, net684150, net684151, net684152, net684153, net684154, 
      net684155, net684156, net684157 : std_logic;

begin
   predicted_next_PC_o <= ( predicted_next_PC_o_31_port, 
      predicted_next_PC_o_30_port, predicted_next_PC_o_29_port, 
      predicted_next_PC_o_28_port, predicted_next_PC_o_27_port, 
      predicted_next_PC_o_26_port, predicted_next_PC_o_25_port, 
      predicted_next_PC_o_24_port, predicted_next_PC_o_23_port, 
      predicted_next_PC_o_22_port, predicted_next_PC_o_21_port, 
      predicted_next_PC_o_20_port, predicted_next_PC_o_19_port, 
      predicted_next_PC_o_18_port, predicted_next_PC_o_17_port, 
      predicted_next_PC_o_16_port, predicted_next_PC_o_15_port, 
      predicted_next_PC_o_14_port, predicted_next_PC_o_13_port, 
      predicted_next_PC_o_12_port, predicted_next_PC_o_11_port, 
      predicted_next_PC_o_10_port, predicted_next_PC_o_9_port, 
      predicted_next_PC_o_8_port, predicted_next_PC_o_7_port, 
      predicted_next_PC_o_6_port, predicted_next_PC_o_5_port, 
      predicted_next_PC_o_4_port, predicted_next_PC_o_3_port, 
      predicted_next_PC_o_2_port, predicted_next_PC_o_1_port, 
      predicted_next_PC_o_0_port );
   taken_o <= taken_o_port;
   mispredict_o <= mispredict_o_port;
   
   last_TAG_reg_3_inst : DFFR_X1 port map( D => n2100, CK => clock, RN => n2288
                           , Q => n591, QN => n664);
   last_TAG_reg_2_inst : DFFR_X1 port map( D => n2099, CK => clock, RN => n2303
                           , Q => n590, QN => n661);
   last_TAG_reg_1_inst : DFFR_X1 port map( D => n2098, CK => clock, RN => n2291
                           , Q => n589, QN => n662);
   last_TAG_reg_0_inst : DFFR_X1 port map( D => n2097, CK => clock, RN => n2299
                           , Q => n588, QN => n660);
   write_enable_reg_15_inst : DFFR_X1 port map( D => n2096, CK => clock, RN => 
                           n2305, Q => write_enable_15_port, QN => n713);
   write_enable_reg_14_inst : DFFR_X1 port map( D => n2095, CK => clock, RN => 
                           n2310, Q => write_enable_14_port, QN => n712);
   write_enable_reg_13_inst : DFFR_X1 port map( D => n2094, CK => clock, RN => 
                           n2300, Q => write_enable_13_port, QN => n711);
   write_enable_reg_12_inst : DFFR_X1 port map( D => n2093, CK => clock, RN => 
                           n2307, Q => write_enable_12_port, QN => n710);
   write_enable_reg_11_inst : DFFR_X1 port map( D => n2092, CK => clock, RN => 
                           n2309, Q => write_enable_11_port, QN => n709);
   write_enable_reg_10_inst : DFFR_X1 port map( D => n2091, CK => clock, RN => 
                           n2310, Q => write_enable_10_port, QN => n708);
   write_enable_reg_9_inst : DFFR_X1 port map( D => n2090, CK => clock, RN => 
                           n2296, Q => write_enable_9_port, QN => n707);
   write_enable_reg_8_inst : DFFR_X1 port map( D => n2089, CK => clock, RN => 
                           n2290, Q => write_enable_8_port, QN => n706);
   write_enable_reg_7_inst : DFFR_X1 port map( D => n2088, CK => clock, RN => 
                           n2309, Q => write_enable_7_port, QN => n705);
   write_enable_reg_6_inst : DFFR_X1 port map( D => n2087, CK => clock, RN => 
                           n2310, Q => write_enable_6_port, QN => n704);
   write_enable_reg_5_inst : DFFR_X1 port map( D => n2086, CK => clock, RN => 
                           n2296, Q => write_enable_5_port, QN => n702);
   write_enable_reg_4_inst : DFFR_X1 port map( D => n2085, CK => clock, RN => 
                           n2299, Q => write_enable_4_port, QN => n700);
   write_enable_reg_3_inst : DFFR_X1 port map( D => n2084, CK => clock, RN => 
                           n2305, Q => write_enable_3_port, QN => n698);
   write_enable_reg_2_inst : DFFR_X1 port map( D => n2083, CK => clock, RN => 
                           n2302, Q => write_enable_2_port, QN => n695);
   write_enable_reg_1_inst : DFFR_X1 port map( D => n2082, CK => clock, RN => 
                           n2307, Q => write_enable_1_port, QN => n694);
   write_enable_reg_0_inst : DFFR_X1 port map( D => n2081, CK => clock, RN => 
                           n2289, Q => write_enable_0_port, QN => n665);
   last_taken_reg : DFF_X1 port map( D => n2080, CK => clock, Q => n663, QN => 
                           net644344);
   predict_PC_reg_0_31_inst : DFFR_X1 port map( D => n2079, CK => clock, RN => 
                           n2308, Q => predict_PC_0_31_port, QN => net644343);
   predict_PC_reg_0_30_inst : DFFR_X1 port map( D => n2078, CK => clock, RN => 
                           n2298, Q => predict_PC_0_30_port, QN => net644342);
   predict_PC_reg_0_29_inst : DFFR_X1 port map( D => n2077, CK => clock, RN => 
                           n2303, Q => predict_PC_0_29_port, QN => net644341);
   predict_PC_reg_0_28_inst : DFFR_X1 port map( D => n2076, CK => clock, RN => 
                           n2308, Q => predict_PC_0_28_port, QN => net644340);
   predict_PC_reg_0_27_inst : DFFR_X1 port map( D => n2075, CK => clock, RN => 
                           n2302, Q => predict_PC_0_27_port, QN => net644339);
   predict_PC_reg_0_26_inst : DFFR_X1 port map( D => n2074, CK => clock, RN => 
                           n2301, Q => predict_PC_0_26_port, QN => net644338);
   predict_PC_reg_0_25_inst : DFFR_X1 port map( D => n2073, CK => clock, RN => 
                           n2309, Q => predict_PC_0_25_port, QN => net644337);
   predict_PC_reg_0_24_inst : DFFR_X1 port map( D => n2072, CK => clock, RN => 
                           n2308, Q => predict_PC_0_24_port, QN => net644336);
   predict_PC_reg_0_23_inst : DFFR_X1 port map( D => n2071, CK => clock, RN => 
                           n2308, Q => predict_PC_0_23_port, QN => net644335);
   predict_PC_reg_0_22_inst : DFFR_X1 port map( D => n2070, CK => clock, RN => 
                           n2292, Q => predict_PC_0_22_port, QN => net644334);
   predict_PC_reg_0_21_inst : DFFR_X1 port map( D => n2069, CK => clock, RN => 
                           n2292, Q => predict_PC_0_21_port, QN => net644333);
   predict_PC_reg_0_20_inst : DFFR_X1 port map( D => n2068, CK => clock, RN => 
                           n2292, Q => predict_PC_0_20_port, QN => net644332);
   predict_PC_reg_0_19_inst : DFFR_X1 port map( D => n2067, CK => clock, RN => 
                           n2292, Q => predict_PC_0_19_port, QN => net644331);
   predict_PC_reg_0_18_inst : DFFR_X1 port map( D => n2066, CK => clock, RN => 
                           n2307, Q => predict_PC_0_18_port, QN => net644330);
   predict_PC_reg_0_17_inst : DFFR_X1 port map( D => n2065, CK => clock, RN => 
                           n2292, Q => predict_PC_0_17_port, QN => net644329);
   predict_PC_reg_0_16_inst : DFFR_X1 port map( D => n2064, CK => clock, RN => 
                           n2292, Q => predict_PC_0_16_port, QN => net644328);
   predict_PC_reg_0_15_inst : DFFR_X1 port map( D => n2063, CK => clock, RN => 
                           n2292, Q => predict_PC_0_15_port, QN => net644327);
   predict_PC_reg_0_14_inst : DFFR_X1 port map( D => n2062, CK => clock, RN => 
                           n2292, Q => predict_PC_0_14_port, QN => net644326);
   predict_PC_reg_0_13_inst : DFFR_X1 port map( D => n2061, CK => clock, RN => 
                           n2292, Q => predict_PC_0_13_port, QN => net644325);
   predict_PC_reg_0_12_inst : DFFR_X1 port map( D => n2060, CK => clock, RN => 
                           n2292, Q => predict_PC_0_12_port, QN => net644324);
   predict_PC_reg_0_11_inst : DFFR_X1 port map( D => n2059, CK => clock, RN => 
                           n2292, Q => predict_PC_0_11_port, QN => net644323);
   predict_PC_reg_0_10_inst : DFFR_X1 port map( D => n2058, CK => clock, RN => 
                           n2298, Q => predict_PC_0_10_port, QN => net644322);
   predict_PC_reg_0_9_inst : DFFR_X1 port map( D => n2057, CK => clock, RN => 
                           n2297, Q => predict_PC_0_9_port, QN => net644321);
   predict_PC_reg_0_8_inst : DFFR_X1 port map( D => n2056, CK => clock, RN => 
                           n2301, Q => predict_PC_0_8_port, QN => net644320);
   predict_PC_reg_0_7_inst : DFFR_X1 port map( D => n2055, CK => clock, RN => 
                           n2303, Q => predict_PC_0_7_port, QN => net644319);
   predict_PC_reg_0_6_inst : DFFR_X1 port map( D => n2054, CK => clock, RN => 
                           n2294, Q => predict_PC_0_6_port, QN => net644318);
   predict_PC_reg_0_5_inst : DFFR_X1 port map( D => n2053, CK => clock, RN => 
                           n2306, Q => predict_PC_0_5_port, QN => net644317);
   predict_PC_reg_0_4_inst : DFFR_X1 port map( D => n2052, CK => clock, RN => 
                           n2300, Q => predict_PC_0_4_port, QN => net644316);
   predict_PC_reg_0_3_inst : DFFR_X1 port map( D => n2051, CK => clock, RN => 
                           n2308, Q => predict_PC_0_3_port, QN => net644315);
   predict_PC_reg_0_2_inst : DFFR_X1 port map( D => n2050, CK => clock, RN => 
                           n2295, Q => predict_PC_0_2_port, QN => net644314);
   predict_PC_reg_0_1_inst : DFFR_X1 port map( D => n2049, CK => clock, RN => 
                           n2295, Q => predict_PC_0_1_port, QN => net644313);
   predict_PC_reg_0_0_inst : DFFR_X1 port map( D => n2048, CK => clock, RN => 
                           n2306, Q => predict_PC_0_0_port, QN => net644312);
   predict_PC_reg_1_31_inst : DFFR_X1 port map( D => n2047, CK => clock, RN => 
                           n2307, Q => predict_PC_1_31_port, QN => net644311);
   predict_PC_reg_1_30_inst : DFFR_X1 port map( D => n2046, CK => clock, RN => 
                           n2298, Q => predict_PC_1_30_port, QN => net644310);
   predict_PC_reg_1_29_inst : DFFR_X1 port map( D => n2045, CK => clock, RN => 
                           n2303, Q => predict_PC_1_29_port, QN => net644309);
   predict_PC_reg_1_28_inst : DFFR_X1 port map( D => n2044, CK => clock, RN => 
                           n2307, Q => predict_PC_1_28_port, QN => net644308);
   predict_PC_reg_1_27_inst : DFFR_X1 port map( D => n2043, CK => clock, RN => 
                           n2302, Q => predict_PC_1_27_port, QN => net644307);
   predict_PC_reg_1_26_inst : DFFR_X1 port map( D => n2042, CK => clock, RN => 
                           n2301, Q => predict_PC_1_26_port, QN => net644306);
   predict_PC_reg_1_25_inst : DFFR_X1 port map( D => n2041, CK => clock, RN => 
                           n2299, Q => predict_PC_1_25_port, QN => net644305);
   predict_PC_reg_1_24_inst : DFFR_X1 port map( D => n2040, CK => clock, RN => 
                           n2310, Q => predict_PC_1_24_port, QN => net644304);
   predict_PC_reg_1_23_inst : DFFR_X1 port map( D => n2039, CK => clock, RN => 
                           n2302, Q => predict_PC_1_23_port, QN => net644303);
   predict_PC_reg_1_22_inst : DFFR_X1 port map( D => n2038, CK => clock, RN => 
                           n2301, Q => predict_PC_1_22_port, QN => net644302);
   predict_PC_reg_1_21_inst : DFFR_X1 port map( D => n2037, CK => clock, RN => 
                           n2303, Q => predict_PC_1_21_port, QN => net644301);
   predict_PC_reg_1_20_inst : DFFR_X1 port map( D => n2036, CK => clock, RN => 
                           n2294, Q => predict_PC_1_20_port, QN => net644300);
   predict_PC_reg_1_19_inst : DFFR_X1 port map( D => n2035, CK => clock, RN => 
                           n2298, Q => predict_PC_1_19_port, QN => net644299);
   predict_PC_reg_1_18_inst : DFFR_X1 port map( D => n2034, CK => clock, RN => 
                           n2300, Q => predict_PC_1_18_port, QN => net644298);
   predict_PC_reg_1_17_inst : DFFR_X1 port map( D => n2033, CK => clock, RN => 
                           n2308, Q => predict_PC_1_17_port, QN => net644297);
   predict_PC_reg_1_16_inst : DFFR_X1 port map( D => n2032, CK => clock, RN => 
                           n2294, Q => predict_PC_1_16_port, QN => net644296);
   predict_PC_reg_1_15_inst : DFFR_X1 port map( D => n2031, CK => clock, RN => 
                           n2294, Q => predict_PC_1_15_port, QN => net644295);
   predict_PC_reg_1_14_inst : DFFR_X1 port map( D => n2030, CK => clock, RN => 
                           n2294, Q => predict_PC_1_14_port, QN => net644294);
   predict_PC_reg_1_13_inst : DFFR_X1 port map( D => n2029, CK => clock, RN => 
                           n2294, Q => predict_PC_1_13_port, QN => net644293);
   predict_PC_reg_1_12_inst : DFFR_X1 port map( D => n2028, CK => clock, RN => 
                           n2294, Q => predict_PC_1_12_port, QN => net644292);
   predict_PC_reg_1_11_inst : DFFR_X1 port map( D => n2027, CK => clock, RN => 
                           n2294, Q => predict_PC_1_11_port, QN => net644291);
   predict_PC_reg_1_10_inst : DFFR_X1 port map( D => n2026, CK => clock, RN => 
                           n2294, Q => predict_PC_1_10_port, QN => net644290);
   predict_PC_reg_1_9_inst : DFFR_X1 port map( D => n2025, CK => clock, RN => 
                           n2304, Q => predict_PC_1_9_port, QN => net644289);
   predict_PC_reg_1_8_inst : DFFR_X1 port map( D => n2024, CK => clock, RN => 
                           n2294, Q => predict_PC_1_8_port, QN => net644288);
   predict_PC_reg_1_7_inst : DFFR_X1 port map( D => n2023, CK => clock, RN => 
                           n2294, Q => predict_PC_1_7_port, QN => net644287);
   predict_PC_reg_1_6_inst : DFFR_X1 port map( D => n2022, CK => clock, RN => 
                           n2297, Q => predict_PC_1_6_port, QN => net644286);
   predict_PC_reg_1_5_inst : DFFR_X1 port map( D => n2021, CK => clock, RN => 
                           n2306, Q => predict_PC_1_5_port, QN => net644285);
   predict_PC_reg_1_4_inst : DFFR_X1 port map( D => n2020, CK => clock, RN => 
                           n2306, Q => predict_PC_1_4_port, QN => net644284);
   predict_PC_reg_1_3_inst : DFFR_X1 port map( D => n2019, CK => clock, RN => 
                           n2306, Q => predict_PC_1_3_port, QN => net644283);
   predict_PC_reg_1_2_inst : DFFR_X1 port map( D => n2018, CK => clock, RN => 
                           n2307, Q => predict_PC_1_2_port, QN => net644282);
   predict_PC_reg_1_1_inst : DFFR_X1 port map( D => n2017, CK => clock, RN => 
                           n2295, Q => predict_PC_1_1_port, QN => net644281);
   predict_PC_reg_1_0_inst : DFFR_X1 port map( D => n2016, CK => clock, RN => 
                           n2307, Q => predict_PC_1_0_port, QN => net644280);
   predict_PC_reg_2_31_inst : DFFR_X1 port map( D => n2015, CK => clock, RN => 
                           n2302, Q => predict_PC_2_31_port, QN => net644279);
   predict_PC_reg_2_30_inst : DFFR_X1 port map( D => n2014, CK => clock, RN => 
                           n2303, Q => predict_PC_2_30_port, QN => net644278);
   predict_PC_reg_2_29_inst : DFFR_X1 port map( D => n2013, CK => clock, RN => 
                           n2302, Q => predict_PC_2_29_port, QN => net644277);
   predict_PC_reg_2_28_inst : DFFR_X1 port map( D => n2012, CK => clock, RN => 
                           n2302, Q => predict_PC_2_28_port, QN => net644276);
   predict_PC_reg_2_27_inst : DFFR_X1 port map( D => n2011, CK => clock, RN => 
                           n2302, Q => predict_PC_2_27_port, QN => net644275);
   predict_PC_reg_2_26_inst : DFFR_X1 port map( D => n2010, CK => clock, RN => 
                           n2289, Q => predict_PC_2_26_port, QN => net644274);
   predict_PC_reg_2_25_inst : DFFR_X1 port map( D => n2009, CK => clock, RN => 
                           n2299, Q => predict_PC_2_25_port, QN => net644273);
   predict_PC_reg_2_24_inst : DFFR_X1 port map( D => n2008, CK => clock, RN => 
                           n2289, Q => predict_PC_2_24_port, QN => net644272);
   predict_PC_reg_2_23_inst : DFFR_X1 port map( D => n2007, CK => clock, RN => 
                           n2288, Q => predict_PC_2_23_port, QN => net644271);
   predict_PC_reg_2_22_inst : DFFR_X1 port map( D => n2006, CK => clock, RN => 
                           n2288, Q => predict_PC_2_22_port, QN => net644270);
   predict_PC_reg_2_21_inst : DFFR_X1 port map( D => n2005, CK => clock, RN => 
                           n2311, Q => predict_PC_2_21_port, QN => net644269);
   predict_PC_reg_2_20_inst : DFFR_X1 port map( D => n2004, CK => clock, RN => 
                           n2288, Q => predict_PC_2_20_port, QN => net644268);
   predict_PC_reg_2_19_inst : DFFR_X1 port map( D => n2003, CK => clock, RN => 
                           n2311, Q => predict_PC_2_19_port, QN => net644267);
   predict_PC_reg_2_18_inst : DFFR_X1 port map( D => n2002, CK => clock, RN => 
                           n2298, Q => predict_PC_2_18_port, QN => net644266);
   predict_PC_reg_2_17_inst : DFFR_X1 port map( D => n2001, CK => clock, RN => 
                           n2301, Q => predict_PC_2_17_port, QN => net644265);
   predict_PC_reg_2_16_inst : DFFR_X1 port map( D => n2000, CK => clock, RN => 
                           n2288, Q => predict_PC_2_16_port, QN => net644264);
   predict_PC_reg_2_15_inst : DFFR_X1 port map( D => n1999, CK => clock, RN => 
                           n2310, Q => predict_PC_2_15_port, QN => net644263);
   predict_PC_reg_2_14_inst : DFFR_X1 port map( D => n1998, CK => clock, RN => 
                           n2289, Q => predict_PC_2_14_port, QN => net644262);
   predict_PC_reg_2_13_inst : DFFR_X1 port map( D => n1997, CK => clock, RN => 
                           n2310, Q => predict_PC_2_13_port, QN => net644261);
   predict_PC_reg_2_12_inst : DFFR_X1 port map( D => n1996, CK => clock, RN => 
                           n2311, Q => predict_PC_2_12_port, QN => net644260);
   predict_PC_reg_2_11_inst : DFFR_X1 port map( D => n1995, CK => clock, RN => 
                           n2311, Q => predict_PC_2_11_port, QN => net644259);
   predict_PC_reg_2_10_inst : DFFR_X1 port map( D => n1994, CK => clock, RN => 
                           n2311, Q => predict_PC_2_10_port, QN => net644258);
   predict_PC_reg_2_9_inst : DFFR_X1 port map( D => n1993, CK => clock, RN => 
                           n2304, Q => predict_PC_2_9_port, QN => net644257);
   predict_PC_reg_2_8_inst : DFFR_X1 port map( D => n1992, CK => clock, RN => 
                           n2311, Q => predict_PC_2_8_port, QN => net644256);
   predict_PC_reg_2_7_inst : DFFR_X1 port map( D => n1991, CK => clock, RN => 
                           n2289, Q => predict_PC_2_7_port, QN => net644255);
   predict_PC_reg_2_6_inst : DFFR_X1 port map( D => n1990, CK => clock, RN => 
                           n2295, Q => predict_PC_2_6_port, QN => net644254);
   predict_PC_reg_2_5_inst : DFFR_X1 port map( D => n1989, CK => clock, RN => 
                           n2306, Q => predict_PC_2_5_port, QN => net644253);
   predict_PC_reg_2_4_inst : DFFR_X1 port map( D => n1988, CK => clock, RN => 
                           n2311, Q => predict_PC_2_4_port, QN => net644252);
   predict_PC_reg_2_3_inst : DFFR_X1 port map( D => n1987, CK => clock, RN => 
                           n2311, Q => predict_PC_2_3_port, QN => net644251);
   predict_PC_reg_2_2_inst : DFFR_X1 port map( D => n1986, CK => clock, RN => 
                           n2300, Q => predict_PC_2_2_port, QN => net644250);
   predict_PC_reg_2_1_inst : DFFR_X1 port map( D => n1985, CK => clock, RN => 
                           n2295, Q => predict_PC_2_1_port, QN => net644249);
   predict_PC_reg_2_0_inst : DFFR_X1 port map( D => n1984, CK => clock, RN => 
                           n2311, Q => predict_PC_2_0_port, QN => net644248);
   predict_PC_reg_3_31_inst : DFFR_X1 port map( D => n1983, CK => clock, RN => 
                           n2309, Q => predict_PC_3_31_port, QN => net644247);
   predict_PC_reg_3_30_inst : DFFR_X1 port map( D => n1982, CK => clock, RN => 
                           n2303, Q => predict_PC_3_30_port, QN => net644246);
   predict_PC_reg_3_29_inst : DFFR_X1 port map( D => n1981, CK => clock, RN => 
                           n2302, Q => predict_PC_3_29_port, QN => net644245);
   predict_PC_reg_3_28_inst : DFFR_X1 port map( D => n1980, CK => clock, RN => 
                           n2297, Q => predict_PC_3_28_port, QN => net644244);
   predict_PC_reg_3_27_inst : DFFR_X1 port map( D => n1979, CK => clock, RN => 
                           n2302, Q => predict_PC_3_27_port, QN => net644243);
   predict_PC_reg_3_26_inst : DFFR_X1 port map( D => n1978, CK => clock, RN => 
                           n2299, Q => predict_PC_3_26_port, QN => net644242);
   predict_PC_reg_3_25_inst : DFFR_X1 port map( D => n1977, CK => clock, RN => 
                           n2299, Q => predict_PC_3_25_port, QN => net644241);
   predict_PC_reg_3_24_inst : DFFR_X1 port map( D => n1976, CK => clock, RN => 
                           n2299, Q => predict_PC_3_24_port, QN => net644240);
   predict_PC_reg_3_23_inst : DFFR_X1 port map( D => n1975, CK => clock, RN => 
                           n2306, Q => predict_PC_3_23_port, QN => net644239);
   predict_PC_reg_3_22_inst : DFFR_X1 port map( D => n1974, CK => clock, RN => 
                           n2295, Q => predict_PC_3_22_port, QN => net644238);
   predict_PC_reg_3_21_inst : DFFR_X1 port map( D => n1973, CK => clock, RN => 
                           n2308, Q => predict_PC_3_21_port, QN => net644237);
   predict_PC_reg_3_20_inst : DFFR_X1 port map( D => n1972, CK => clock, RN => 
                           n2295, Q => predict_PC_3_20_port, QN => net644236);
   predict_PC_reg_3_19_inst : DFFR_X1 port map( D => n1971, CK => clock, RN => 
                           n2291, Q => predict_PC_3_19_port, QN => net644235);
   predict_PC_reg_3_18_inst : DFFR_X1 port map( D => n1970, CK => clock, RN => 
                           n2300, Q => predict_PC_3_18_port, QN => net644234);
   predict_PC_reg_3_17_inst : DFFR_X1 port map( D => n1969, CK => clock, RN => 
                           n2290, Q => predict_PC_3_17_port, QN => net644233);
   predict_PC_reg_3_16_inst : DFFR_X1 port map( D => n1968, CK => clock, RN => 
                           n2290, Q => predict_PC_3_16_port, QN => net644232);
   predict_PC_reg_3_15_inst : DFFR_X1 port map( D => n1967, CK => clock, RN => 
                           n2290, Q => predict_PC_3_15_port, QN => net644231);
   predict_PC_reg_3_14_inst : DFFR_X1 port map( D => n1966, CK => clock, RN => 
                           n2290, Q => predict_PC_3_14_port, QN => net644230);
   predict_PC_reg_3_13_inst : DFFR_X1 port map( D => n1965, CK => clock, RN => 
                           n2290, Q => predict_PC_3_13_port, QN => net644229);
   predict_PC_reg_3_12_inst : DFFR_X1 port map( D => n1964, CK => clock, RN => 
                           n2290, Q => predict_PC_3_12_port, QN => net644228);
   predict_PC_reg_3_11_inst : DFFR_X1 port map( D => n1963, CK => clock, RN => 
                           n2290, Q => predict_PC_3_11_port, QN => net644227);
   predict_PC_reg_3_10_inst : DFFR_X1 port map( D => n1962, CK => clock, RN => 
                           n2290, Q => predict_PC_3_10_port, QN => net644226);
   predict_PC_reg_3_9_inst : DFFR_X1 port map( D => n1961, CK => clock, RN => 
                           n2304, Q => predict_PC_3_9_port, QN => net644225);
   predict_PC_reg_3_8_inst : DFFR_X1 port map( D => n1960, CK => clock, RN => 
                           n2290, Q => predict_PC_3_8_port, QN => net644224);
   predict_PC_reg_3_7_inst : DFFR_X1 port map( D => n1959, CK => clock, RN => 
                           n2309, Q => predict_PC_3_7_port, QN => net644223);
   predict_PC_reg_3_6_inst : DFFR_X1 port map( D => n1958, CK => clock, RN => 
                           n2309, Q => predict_PC_3_6_port, QN => net644222);
   predict_PC_reg_3_5_inst : DFFR_X1 port map( D => n1957, CK => clock, RN => 
                           n2306, Q => predict_PC_3_5_port, QN => net644221);
   predict_PC_reg_3_4_inst : DFFR_X1 port map( D => n1956, CK => clock, RN => 
                           n2309, Q => predict_PC_3_4_port, QN => net644220);
   predict_PC_reg_3_3_inst : DFFR_X1 port map( D => n1955, CK => clock, RN => 
                           n2309, Q => predict_PC_3_3_port, QN => net644219);
   predict_PC_reg_3_2_inst : DFFR_X1 port map( D => n1954, CK => clock, RN => 
                           n2309, Q => predict_PC_3_2_port, QN => net644218);
   predict_PC_reg_3_1_inst : DFFR_X1 port map( D => n1953, CK => clock, RN => 
                           n2295, Q => predict_PC_3_1_port, QN => net644217);
   predict_PC_reg_3_0_inst : DFFR_X1 port map( D => n1952, CK => clock, RN => 
                           n2309, Q => predict_PC_3_0_port, QN => net644216);
   predict_PC_reg_4_31_inst : DFFR_X1 port map( D => n1951, CK => clock, RN => 
                           n2297, Q => predict_PC_4_31_port, QN => net644215);
   predict_PC_reg_4_30_inst : DFFR_X1 port map( D => n1950, CK => clock, RN => 
                           n2303, Q => predict_PC_4_30_port, QN => net644214);
   predict_PC_reg_4_29_inst : DFFR_X1 port map( D => n1949, CK => clock, RN => 
                           n2302, Q => predict_PC_4_29_port, QN => net644213);
   predict_PC_reg_4_28_inst : DFFR_X1 port map( D => n1948, CK => clock, RN => 
                           n2309, Q => predict_PC_4_28_port, QN => net644212);
   predict_PC_reg_4_27_inst : DFFR_X1 port map( D => n1947, CK => clock, RN => 
                           n2302, Q => predict_PC_4_27_port, QN => net644211);
   predict_PC_reg_4_26_inst : DFFR_X1 port map( D => n1946, CK => clock, RN => 
                           n2299, Q => predict_PC_4_26_port, QN => net644210);
   predict_PC_reg_4_25_inst : DFFR_X1 port map( D => n1945, CK => clock, RN => 
                           n2300, Q => predict_PC_4_25_port, QN => net644209);
   predict_PC_reg_4_24_inst : DFFR_X1 port map( D => n1944, CK => clock, RN => 
                           n2302, Q => predict_PC_4_24_port, QN => net644208);
   predict_PC_reg_4_23_inst : DFFR_X1 port map( D => n1943, CK => clock, RN => 
                           n2293, Q => predict_PC_4_23_port, QN => net644207);
   predict_PC_reg_4_22_inst : DFFR_X1 port map( D => n1942, CK => clock, RN => 
                           n2293, Q => predict_PC_4_22_port, QN => net644206);
   predict_PC_reg_4_21_inst : DFFR_X1 port map( D => n1941, CK => clock, RN => 
                           n2293, Q => predict_PC_4_21_port, QN => net644205);
   predict_PC_reg_4_20_inst : DFFR_X1 port map( D => n1940, CK => clock, RN => 
                           n2293, Q => predict_PC_4_20_port, QN => net644204);
   predict_PC_reg_4_19_inst : DFFR_X1 port map( D => n1939, CK => clock, RN => 
                           n2293, Q => predict_PC_4_19_port, QN => net644203);
   predict_PC_reg_4_18_inst : DFFR_X1 port map( D => n1938, CK => clock, RN => 
                           n2290, Q => predict_PC_4_18_port, QN => net644202);
   predict_PC_reg_4_17_inst : DFFR_X1 port map( D => n1937, CK => clock, RN => 
                           n2293, Q => predict_PC_4_17_port, QN => net644201);
   predict_PC_reg_4_16_inst : DFFR_X1 port map( D => n1936, CK => clock, RN => 
                           n2293, Q => predict_PC_4_16_port, QN => net644200);
   predict_PC_reg_4_15_inst : DFFR_X1 port map( D => n1935, CK => clock, RN => 
                           n2293, Q => predict_PC_4_15_port, QN => net644199);
   predict_PC_reg_4_14_inst : DFFR_X1 port map( D => n1934, CK => clock, RN => 
                           n2293, Q => predict_PC_4_14_port, QN => net644198);
   predict_PC_reg_4_13_inst : DFFR_X1 port map( D => n1933, CK => clock, RN => 
                           n2293, Q => predict_PC_4_13_port, QN => net644197);
   predict_PC_reg_4_12_inst : DFFR_X1 port map( D => n1932, CK => clock, RN => 
                           n2293, Q => predict_PC_4_12_port, QN => net644196);
   predict_PC_reg_4_11_inst : DFFR_X1 port map( D => n1931, CK => clock, RN => 
                           n2292, Q => predict_PC_4_11_port, QN => net644195);
   predict_PC_reg_4_10_inst : DFFR_X1 port map( D => n1930, CK => clock, RN => 
                           n2304, Q => predict_PC_4_10_port, QN => net644194);
   predict_PC_reg_4_9_inst : DFFR_X1 port map( D => n1929, CK => clock, RN => 
                           n2304, Q => predict_PC_4_9_port, QN => net644193);
   predict_PC_reg_4_8_inst : DFFR_X1 port map( D => n1928, CK => clock, RN => 
                           n2307, Q => predict_PC_4_8_port, QN => net644192);
   predict_PC_reg_4_7_inst : DFFR_X1 port map( D => n1927, CK => clock, RN => 
                           n2302, Q => predict_PC_4_7_port, QN => net644191);
   predict_PC_reg_4_6_inst : DFFR_X1 port map( D => n1926, CK => clock, RN => 
                           n2290, Q => predict_PC_4_6_port, QN => net644190);
   predict_PC_reg_4_5_inst : DFFR_X1 port map( D => n1925, CK => clock, RN => 
                           n2306, Q => predict_PC_4_5_port, QN => net644189);
   predict_PC_reg_4_4_inst : DFFR_X1 port map( D => n1924, CK => clock, RN => 
                           n2293, Q => predict_PC_4_4_port, QN => net644188);
   predict_PC_reg_4_3_inst : DFFR_X1 port map( D => n1923, CK => clock, RN => 
                           n2291, Q => predict_PC_4_3_port, QN => net644187);
   predict_PC_reg_4_2_inst : DFFR_X1 port map( D => n1922, CK => clock, RN => 
                           n2311, Q => predict_PC_4_2_port, QN => net644186);
   predict_PC_reg_4_1_inst : DFFR_X1 port map( D => n1921, CK => clock, RN => 
                           n2307, Q => predict_PC_4_1_port, QN => net644185);
   predict_PC_reg_4_0_inst : DFFR_X1 port map( D => n1920, CK => clock, RN => 
                           n2292, Q => predict_PC_4_0_port, QN => net644184);
   predict_PC_reg_5_31_inst : DFFR_X1 port map( D => n1919, CK => clock, RN => 
                           n2296, Q => predict_PC_5_31_port, QN => net644183);
   predict_PC_reg_5_30_inst : DFFR_X1 port map( D => n1918, CK => clock, RN => 
                           n2303, Q => predict_PC_5_30_port, QN => net644182);
   predict_PC_reg_5_29_inst : DFFR_X1 port map( D => n1917, CK => clock, RN => 
                           n2302, Q => predict_PC_5_29_port, QN => net644181);
   predict_PC_reg_5_28_inst : DFFR_X1 port map( D => n1916, CK => clock, RN => 
                           n2296, Q => predict_PC_5_28_port, QN => net644180);
   predict_PC_reg_5_27_inst : DFFR_X1 port map( D => n1915, CK => clock, RN => 
                           n2298, Q => predict_PC_5_27_port, QN => net644179);
   predict_PC_reg_5_26_inst : DFFR_X1 port map( D => n1914, CK => clock, RN => 
                           n2299, Q => predict_PC_5_26_port, QN => net644178);
   predict_PC_reg_5_25_inst : DFFR_X1 port map( D => n1913, CK => clock, RN => 
                           n2300, Q => predict_PC_5_25_port, QN => net644177);
   predict_PC_reg_5_24_inst : DFFR_X1 port map( D => n1912, CK => clock, RN => 
                           n2296, Q => predict_PC_5_24_port, QN => net644176);
   predict_PC_reg_5_23_inst : DFFR_X1 port map( D => n1911, CK => clock, RN => 
                           n2296, Q => predict_PC_5_23_port, QN => net644175);
   predict_PC_reg_5_22_inst : DFFR_X1 port map( D => n1910, CK => clock, RN => 
                           n2296, Q => predict_PC_5_22_port, QN => net644174);
   predict_PC_reg_5_21_inst : DFFR_X1 port map( D => n1909, CK => clock, RN => 
                           n2296, Q => predict_PC_5_21_port, QN => net644173);
   predict_PC_reg_5_20_inst : DFFR_X1 port map( D => n1908, CK => clock, RN => 
                           n2295, Q => predict_PC_5_20_port, QN => net644172);
   predict_PC_reg_5_19_inst : DFFR_X1 port map( D => n1907, CK => clock, RN => 
                           n2295, Q => predict_PC_5_19_port, QN => net644171);
   predict_PC_reg_5_18_inst : DFFR_X1 port map( D => n1906, CK => clock, RN => 
                           n2288, Q => predict_PC_5_18_port, QN => net644170);
   predict_PC_reg_5_17_inst : DFFR_X1 port map( D => n1905, CK => clock, RN => 
                           n2295, Q => predict_PC_5_17_port, QN => net644169);
   predict_PC_reg_5_16_inst : DFFR_X1 port map( D => n1904, CK => clock, RN => 
                           n2295, Q => predict_PC_5_16_port, QN => net644168);
   predict_PC_reg_5_15_inst : DFFR_X1 port map( D => n1903, CK => clock, RN => 
                           n2305, Q => predict_PC_5_15_port, QN => net644167);
   predict_PC_reg_5_14_inst : DFFR_X1 port map( D => n1902, CK => clock, RN => 
                           n2305, Q => predict_PC_5_14_port, QN => net644166);
   predict_PC_reg_5_13_inst : DFFR_X1 port map( D => n1901, CK => clock, RN => 
                           n2305, Q => predict_PC_5_13_port, QN => net644165);
   predict_PC_reg_5_12_inst : DFFR_X1 port map( D => n1900, CK => clock, RN => 
                           n2306, Q => predict_PC_5_12_port, QN => net644164);
   predict_PC_reg_5_11_inst : DFFR_X1 port map( D => n1899, CK => clock, RN => 
                           n2306, Q => predict_PC_5_11_port, QN => net644163);
   predict_PC_reg_5_10_inst : DFFR_X1 port map( D => n1898, CK => clock, RN => 
                           n2306, Q => predict_PC_5_10_port, QN => net644162);
   predict_PC_reg_5_9_inst : DFFR_X1 port map( D => n1897, CK => clock, RN => 
                           n2304, Q => predict_PC_5_9_port, QN => net644161);
   predict_PC_reg_5_8_inst : DFFR_X1 port map( D => n1896, CK => clock, RN => 
                           n2306, Q => predict_PC_5_8_port, QN => net644160);
   predict_PC_reg_5_7_inst : DFFR_X1 port map( D => n1895, CK => clock, RN => 
                           n2306, Q => predict_PC_5_7_port, QN => net644159);
   predict_PC_reg_5_6_inst : DFFR_X1 port map( D => n1894, CK => clock, RN => 
                           n2306, Q => predict_PC_5_6_port, QN => net644158);
   predict_PC_reg_5_5_inst : DFFR_X1 port map( D => n1893, CK => clock, RN => 
                           n2306, Q => predict_PC_5_5_port, QN => net644157);
   predict_PC_reg_5_4_inst : DFFR_X1 port map( D => n1892, CK => clock, RN => 
                           n2306, Q => predict_PC_5_4_port, QN => net644156);
   predict_PC_reg_5_3_inst : DFFR_X1 port map( D => n1891, CK => clock, RN => 
                           n2306, Q => predict_PC_5_3_port, QN => net644155);
   predict_PC_reg_5_2_inst : DFFR_X1 port map( D => n1890, CK => clock, RN => 
                           n2306, Q => predict_PC_5_2_port, QN => net644154);
   predict_PC_reg_5_1_inst : DFFR_X1 port map( D => n1889, CK => clock, RN => 
                           n2307, Q => predict_PC_5_1_port, QN => net644153);
   predict_PC_reg_5_0_inst : DFFR_X1 port map( D => n1888, CK => clock, RN => 
                           n2296, Q => predict_PC_5_0_port, QN => net644152);
   predict_PC_reg_6_31_inst : DFFR_X1 port map( D => n1887, CK => clock, RN => 
                           n2310, Q => predict_PC_6_31_port, QN => net644151);
   predict_PC_reg_6_30_inst : DFFR_X1 port map( D => n1886, CK => clock, RN => 
                           n2303, Q => predict_PC_6_30_port, QN => net644150);
   predict_PC_reg_6_29_inst : DFFR_X1 port map( D => n1885, CK => clock, RN => 
                           n2302, Q => predict_PC_6_29_port, QN => net644149);
   predict_PC_reg_6_28_inst : DFFR_X1 port map( D => n1884, CK => clock, RN => 
                           n2310, Q => predict_PC_6_28_port, QN => net644148);
   predict_PC_reg_6_27_inst : DFFR_X1 port map( D => n1883, CK => clock, RN => 
                           n2298, Q => predict_PC_6_27_port, QN => net644147);
   predict_PC_reg_6_26_inst : DFFR_X1 port map( D => n1882, CK => clock, RN => 
                           n2299, Q => predict_PC_6_26_port, QN => net644146);
   predict_PC_reg_6_25_inst : DFFR_X1 port map( D => n1881, CK => clock, RN => 
                           n2300, Q => predict_PC_6_25_port, QN => net644145);
   predict_PC_reg_6_24_inst : DFFR_X1 port map( D => n1880, CK => clock, RN => 
                           n2311, Q => predict_PC_6_24_port, QN => net644144);
   predict_PC_reg_6_23_inst : DFFR_X1 port map( D => n1879, CK => clock, RN => 
                           n2288, Q => predict_PC_6_23_port, QN => net644143);
   predict_PC_reg_6_22_inst : DFFR_X1 port map( D => n1878, CK => clock, RN => 
                           n2288, Q => predict_PC_6_22_port, QN => net644142);
   predict_PC_reg_6_21_inst : DFFR_X1 port map( D => n1877, CK => clock, RN => 
                           n2311, Q => predict_PC_6_21_port, QN => net644141);
   predict_PC_reg_6_20_inst : DFFR_X1 port map( D => n1876, CK => clock, RN => 
                           n2308, Q => predict_PC_6_20_port, QN => net644140);
   predict_PC_reg_6_19_inst : DFFR_X1 port map( D => n1875, CK => clock, RN => 
                           n2311, Q => predict_PC_6_19_port, QN => net644139);
   predict_PC_reg_6_18_inst : DFFR_X1 port map( D => n1874, CK => clock, RN => 
                           n2288, Q => predict_PC_6_18_port, QN => net644138);
   predict_PC_reg_6_17_inst : DFFR_X1 port map( D => n1873, CK => clock, RN => 
                           n2304, Q => predict_PC_6_17_port, QN => net644137);
   predict_PC_reg_6_16_inst : DFFR_X1 port map( D => n1872, CK => clock, RN => 
                           n2289, Q => predict_PC_6_16_port, QN => net644136);
   predict_PC_reg_6_15_inst : DFFR_X1 port map( D => n1871, CK => clock, RN => 
                           n2289, Q => predict_PC_6_15_port, QN => net644135);
   predict_PC_reg_6_14_inst : DFFR_X1 port map( D => n1870, CK => clock, RN => 
                           n2289, Q => predict_PC_6_14_port, QN => net644134);
   predict_PC_reg_6_13_inst : DFFR_X1 port map( D => n1869, CK => clock, RN => 
                           n2289, Q => predict_PC_6_13_port, QN => net644133);
   predict_PC_reg_6_12_inst : DFFR_X1 port map( D => n1868, CK => clock, RN => 
                           n2289, Q => predict_PC_6_12_port, QN => net644132);
   predict_PC_reg_6_11_inst : DFFR_X1 port map( D => n1867, CK => clock, RN => 
                           n2289, Q => predict_PC_6_11_port, QN => net644131);
   predict_PC_reg_6_10_inst : DFFR_X1 port map( D => n1866, CK => clock, RN => 
                           n2289, Q => predict_PC_6_10_port, QN => net644130);
   predict_PC_reg_6_9_inst : DFFR_X1 port map( D => n1865, CK => clock, RN => 
                           n2304, Q => predict_PC_6_9_port, QN => net644129);
   predict_PC_reg_6_8_inst : DFFR_X1 port map( D => n1864, CK => clock, RN => 
                           n2289, Q => predict_PC_6_8_port, QN => net644128);
   predict_PC_reg_6_7_inst : DFFR_X1 port map( D => n1863, CK => clock, RN => 
                           n2289, Q => predict_PC_6_7_port, QN => net644127);
   predict_PC_reg_6_6_inst : DFFR_X1 port map( D => n1862, CK => clock, RN => 
                           n2308, Q => predict_PC_6_6_port, QN => net644126);
   predict_PC_reg_6_5_inst : DFFR_X1 port map( D => n1861, CK => clock, RN => 
                           n2306, Q => predict_PC_6_5_port, QN => net644125);
   predict_PC_reg_6_4_inst : DFFR_X1 port map( D => n1860, CK => clock, RN => 
                           n2289, Q => predict_PC_6_4_port, QN => net644124);
   predict_PC_reg_6_3_inst : DFFR_X1 port map( D => n1859, CK => clock, RN => 
                           n2289, Q => predict_PC_6_3_port, QN => net644123);
   predict_PC_reg_6_2_inst : DFFR_X1 port map( D => n1858, CK => clock, RN => 
                           n2300, Q => predict_PC_6_2_port, QN => net644122);
   predict_PC_reg_6_1_inst : DFFR_X1 port map( D => n1857, CK => clock, RN => 
                           n2307, Q => predict_PC_6_1_port, QN => net644121);
   predict_PC_reg_6_0_inst : DFFR_X1 port map( D => n1856, CK => clock, RN => 
                           n2310, Q => predict_PC_6_0_port, QN => net644120);
   predict_PC_reg_7_31_inst : DFFR_X1 port map( D => n1855, CK => clock, RN => 
                           n2309, Q => predict_PC_7_31_port, QN => net644119);
   predict_PC_reg_7_30_inst : DFFR_X1 port map( D => n1854, CK => clock, RN => 
                           n2303, Q => predict_PC_7_30_port, QN => net644118);
   predict_PC_reg_7_29_inst : DFFR_X1 port map( D => n1853, CK => clock, RN => 
                           n2302, Q => predict_PC_7_29_port, QN => net644117);
   predict_PC_reg_7_28_inst : DFFR_X1 port map( D => n1852, CK => clock, RN => 
                           n2309, Q => predict_PC_7_28_port, QN => net644116);
   predict_PC_reg_7_27_inst : DFFR_X1 port map( D => n1851, CK => clock, RN => 
                           n2298, Q => predict_PC_7_27_port, QN => net644115);
   predict_PC_reg_7_26_inst : DFFR_X1 port map( D => n1850, CK => clock, RN => 
                           n2299, Q => predict_PC_7_26_port, QN => net644114);
   predict_PC_reg_7_25_inst : DFFR_X1 port map( D => n1849, CK => clock, RN => 
                           n2300, Q => predict_PC_7_25_port, QN => net644113);
   predict_PC_reg_7_24_inst : DFFR_X1 port map( D => n1848, CK => clock, RN => 
                           n2309, Q => predict_PC_7_24_port, QN => net644112);
   predict_PC_reg_7_23_inst : DFFR_X1 port map( D => n1847, CK => clock, RN => 
                           n2309, Q => predict_PC_7_23_port, QN => net644111);
   predict_PC_reg_7_22_inst : DFFR_X1 port map( D => n1846, CK => clock, RN => 
                           n2309, Q => predict_PC_7_22_port, QN => net644110);
   predict_PC_reg_7_21_inst : DFFR_X1 port map( D => n1845, CK => clock, RN => 
                           n2291, Q => predict_PC_7_21_port, QN => net644109);
   predict_PC_reg_7_20_inst : DFFR_X1 port map( D => n1844, CK => clock, RN => 
                           n2291, Q => predict_PC_7_20_port, QN => net644108);
   predict_PC_reg_7_19_inst : DFFR_X1 port map( D => n1843, CK => clock, RN => 
                           n2291, Q => predict_PC_7_19_port, QN => net644107);
   predict_PC_reg_7_18_inst : DFFR_X1 port map( D => n1842, CK => clock, RN => 
                           n2288, Q => predict_PC_7_18_port, QN => net644106);
   predict_PC_reg_7_17_inst : DFFR_X1 port map( D => n1841, CK => clock, RN => 
                           n2291, Q => predict_PC_7_17_port, QN => net644105);
   predict_PC_reg_7_16_inst : DFFR_X1 port map( D => n1840, CK => clock, RN => 
                           n2291, Q => predict_PC_7_16_port, QN => net644104);
   predict_PC_reg_7_15_inst : DFFR_X1 port map( D => n1839, CK => clock, RN => 
                           n2291, Q => predict_PC_7_15_port, QN => net644103);
   predict_PC_reg_7_14_inst : DFFR_X1 port map( D => n1838, CK => clock, RN => 
                           n2291, Q => predict_PC_7_14_port, QN => net644102);
   predict_PC_reg_7_13_inst : DFFR_X1 port map( D => n1837, CK => clock, RN => 
                           n2291, Q => predict_PC_7_13_port, QN => net644101);
   predict_PC_reg_7_12_inst : DFFR_X1 port map( D => n1836, CK => clock, RN => 
                           n2291, Q => predict_PC_7_12_port, QN => net644100);
   predict_PC_reg_7_11_inst : DFFR_X1 port map( D => n1835, CK => clock, RN => 
                           n2291, Q => predict_PC_7_11_port, QN => net644099);
   predict_PC_reg_7_10_inst : DFFR_X1 port map( D => n1834, CK => clock, RN => 
                           n2291, Q => predict_PC_7_10_port, QN => net644098);
   predict_PC_reg_7_9_inst : DFFR_X1 port map( D => n1833, CK => clock, RN => 
                           n2304, Q => predict_PC_7_9_port, QN => net644097);
   predict_PC_reg_7_8_inst : DFFR_X1 port map( D => n1832, CK => clock, RN => 
                           n2291, Q => predict_PC_7_8_port, QN => net644096);
   predict_PC_reg_7_7_inst : DFFR_X1 port map( D => n1831, CK => clock, RN => 
                           n2308, Q => predict_PC_7_7_port, QN => net644095);
   predict_PC_reg_7_6_inst : DFFR_X1 port map( D => n1830, CK => clock, RN => 
                           n2308, Q => predict_PC_7_6_port, QN => net644094);
   predict_PC_reg_7_5_inst : DFFR_X1 port map( D => n1829, CK => clock, RN => 
                           n2306, Q => predict_PC_7_5_port, QN => net644093);
   predict_PC_reg_7_4_inst : DFFR_X1 port map( D => n1828, CK => clock, RN => 
                           n2308, Q => predict_PC_7_4_port, QN => net644092);
   predict_PC_reg_7_3_inst : DFFR_X1 port map( D => n1827, CK => clock, RN => 
                           n2308, Q => predict_PC_7_3_port, QN => net644091);
   predict_PC_reg_7_2_inst : DFFR_X1 port map( D => n1826, CK => clock, RN => 
                           n2308, Q => predict_PC_7_2_port, QN => net644090);
   predict_PC_reg_7_1_inst : DFFR_X1 port map( D => n1825, CK => clock, RN => 
                           n2307, Q => predict_PC_7_1_port, QN => net644089);
   predict_PC_reg_7_0_inst : DFFR_X1 port map( D => n1824, CK => clock, RN => 
                           n2308, Q => predict_PC_7_0_port, QN => net644088);
   predict_PC_reg_8_31_inst : DFFR_X1 port map( D => n1823, CK => clock, RN => 
                           n2309, Q => predict_PC_8_31_port, QN => net644087);
   predict_PC_reg_8_30_inst : DFFR_X1 port map( D => n1822, CK => clock, RN => 
                           n2303, Q => predict_PC_8_30_port, QN => net644086);
   predict_PC_reg_8_29_inst : DFFR_X1 port map( D => n1821, CK => clock, RN => 
                           n2302, Q => predict_PC_8_29_port, QN => net644085);
   predict_PC_reg_8_28_inst : DFFR_X1 port map( D => n1820, CK => clock, RN => 
                           n2309, Q => predict_PC_8_28_port, QN => net644084);
   predict_PC_reg_8_27_inst : DFFR_X1 port map( D => n1819, CK => clock, RN => 
                           n2298, Q => predict_PC_8_27_port, QN => net644083);
   predict_PC_reg_8_26_inst : DFFR_X1 port map( D => n1818, CK => clock, RN => 
                           n2299, Q => predict_PC_8_26_port, QN => net644082);
   predict_PC_reg_8_25_inst : DFFR_X1 port map( D => n1817, CK => clock, RN => 
                           n2300, Q => predict_PC_8_25_port, QN => net644081);
   predict_PC_reg_8_24_inst : DFFR_X1 port map( D => n1816, CK => clock, RN => 
                           n2309, Q => predict_PC_8_24_port, QN => net644080);
   predict_PC_reg_8_23_inst : DFFR_X1 port map( D => n1815, CK => clock, RN => 
                           n2290, Q => predict_PC_8_23_port, QN => net644079);
   predict_PC_reg_8_22_inst : DFFR_X1 port map( D => n1814, CK => clock, RN => 
                           n2288, Q => predict_PC_8_22_port, QN => net644078);
   predict_PC_reg_8_21_inst : DFFR_X1 port map( D => n1813, CK => clock, RN => 
                           n2288, Q => predict_PC_8_21_port, QN => net644077);
   predict_PC_reg_8_20_inst : DFFR_X1 port map( D => n1812, CK => clock, RN => 
                           n2309, Q => predict_PC_8_20_port, QN => net644076);
   predict_PC_reg_8_19_inst : DFFR_X1 port map( D => n1811, CK => clock, RN => 
                           n2311, Q => predict_PC_8_19_port, QN => net644075);
   predict_PC_reg_8_18_inst : DFFR_X1 port map( D => n1810, CK => clock, RN => 
                           n2301, Q => predict_PC_8_18_port, QN => net644074);
   predict_PC_reg_8_17_inst : DFFR_X1 port map( D => n1809, CK => clock, RN => 
                           n2300, Q => predict_PC_8_17_port, QN => net644073);
   predict_PC_reg_8_16_inst : DFFR_X1 port map( D => n1808, CK => clock, RN => 
                           n2292, Q => predict_PC_8_16_port, QN => net644072);
   predict_PC_reg_8_15_inst : DFFR_X1 port map( D => n1807, CK => clock, RN => 
                           n2290, Q => predict_PC_8_15_port, QN => net644071);
   predict_PC_reg_8_14_inst : DFFR_X1 port map( D => n1806, CK => clock, RN => 
                           n2311, Q => predict_PC_8_14_port, QN => net644070);
   predict_PC_reg_8_13_inst : DFFR_X1 port map( D => n1805, CK => clock, RN => 
                           n2290, Q => predict_PC_8_13_port, QN => net644069);
   predict_PC_reg_8_12_inst : DFFR_X1 port map( D => n1804, CK => clock, RN => 
                           n2290, Q => predict_PC_8_12_port, QN => net644068);
   predict_PC_reg_8_11_inst : DFFR_X1 port map( D => n1803, CK => clock, RN => 
                           n2290, Q => predict_PC_8_11_port, QN => net644067);
   predict_PC_reg_8_10_inst : DFFR_X1 port map( D => n1802, CK => clock, RN => 
                           n2305, Q => predict_PC_8_10_port, QN => net644066);
   predict_PC_reg_8_9_inst : DFFR_X1 port map( D => n1801, CK => clock, RN => 
                           n2304, Q => predict_PC_8_9_port, QN => net644065);
   predict_PC_reg_8_8_inst : DFFR_X1 port map( D => n1800, CK => clock, RN => 
                           n2290, Q => predict_PC_8_8_port, QN => net644064);
   predict_PC_reg_8_7_inst : DFFR_X1 port map( D => n1799, CK => clock, RN => 
                           n2289, Q => predict_PC_8_7_port, QN => net644063);
   predict_PC_reg_8_6_inst : DFFR_X1 port map( D => n1798, CK => clock, RN => 
                           n2292, Q => predict_PC_8_6_port, QN => net644062);
   predict_PC_reg_8_5_inst : DFFR_X1 port map( D => n1797, CK => clock, RN => 
                           n2295, Q => predict_PC_8_5_port, QN => net644061);
   predict_PC_reg_8_4_inst : DFFR_X1 port map( D => n1796, CK => clock, RN => 
                           n2290, Q => predict_PC_8_4_port, QN => net644060);
   predict_PC_reg_8_3_inst : DFFR_X1 port map( D => n1795, CK => clock, RN => 
                           n2289, Q => predict_PC_8_3_port, QN => net644059);
   predict_PC_reg_8_2_inst : DFFR_X1 port map( D => n1794, CK => clock, RN => 
                           n2300, Q => predict_PC_8_2_port, QN => net644058);
   predict_PC_reg_8_1_inst : DFFR_X1 port map( D => n1793, CK => clock, RN => 
                           n2307, Q => predict_PC_8_1_port, QN => net644057);
   predict_PC_reg_8_0_inst : DFFR_X1 port map( D => n1792, CK => clock, RN => 
                           n2306, Q => predict_PC_8_0_port, QN => net644056);
   predict_PC_reg_9_31_inst : DFFR_X1 port map( D => n1791, CK => clock, RN => 
                           n2296, Q => predict_PC_9_31_port, QN => net644055);
   predict_PC_reg_9_30_inst : DFFR_X1 port map( D => n1790, CK => clock, RN => 
                           n2303, Q => predict_PC_9_30_port, QN => net644054);
   predict_PC_reg_9_29_inst : DFFR_X1 port map( D => n1789, CK => clock, RN => 
                           n2297, Q => predict_PC_9_29_port, QN => net644053);
   predict_PC_reg_9_28_inst : DFFR_X1 port map( D => n1788, CK => clock, RN => 
                           n2296, Q => predict_PC_9_28_port, QN => net644052);
   predict_PC_reg_9_27_inst : DFFR_X1 port map( D => n1787, CK => clock, RN => 
                           n2298, Q => predict_PC_9_27_port, QN => net644051);
   predict_PC_reg_9_26_inst : DFFR_X1 port map( D => n1786, CK => clock, RN => 
                           n2299, Q => predict_PC_9_26_port, QN => net644050);
   predict_PC_reg_9_25_inst : DFFR_X1 port map( D => n1785, CK => clock, RN => 
                           n2300, Q => predict_PC_9_25_port, QN => net644049);
   predict_PC_reg_9_24_inst : DFFR_X1 port map( D => n1784, CK => clock, RN => 
                           n2296, Q => predict_PC_9_24_port, QN => net644048);
   predict_PC_reg_9_23_inst : DFFR_X1 port map( D => n1783, CK => clock, RN => 
                           n2296, Q => predict_PC_9_23_port, QN => net644047);
   predict_PC_reg_9_22_inst : DFFR_X1 port map( D => n1782, CK => clock, RN => 
                           n2296, Q => predict_PC_9_22_port, QN => net644046);
   predict_PC_reg_9_21_inst : DFFR_X1 port map( D => n1781, CK => clock, RN => 
                           n2296, Q => predict_PC_9_21_port, QN => net644045);
   predict_PC_reg_9_20_inst : DFFR_X1 port map( D => n1780, CK => clock, RN => 
                           n2296, Q => predict_PC_9_20_port, QN => net644044);
   predict_PC_reg_9_19_inst : DFFR_X1 port map( D => n1779, CK => clock, RN => 
                           n2296, Q => predict_PC_9_19_port, QN => net644043);
   predict_PC_reg_9_18_inst : DFFR_X1 port map( D => n1778, CK => clock, RN => 
                           n2301, Q => predict_PC_9_18_port, QN => net644042);
   predict_PC_reg_9_17_inst : DFFR_X1 port map( D => n1777, CK => clock, RN => 
                           n2296, Q => predict_PC_9_17_port, QN => net644041);
   predict_PC_reg_9_16_inst : DFFR_X1 port map( D => n1776, CK => clock, RN => 
                           n2296, Q => predict_PC_9_16_port, QN => net644040);
   predict_PC_reg_9_15_inst : DFFR_X1 port map( D => n1775, CK => clock, RN => 
                           n2305, Q => predict_PC_9_15_port, QN => net644039);
   predict_PC_reg_9_14_inst : DFFR_X1 port map( D => n1774, CK => clock, RN => 
                           n2305, Q => predict_PC_9_14_port, QN => net644038);
   predict_PC_reg_9_13_inst : DFFR_X1 port map( D => n1773, CK => clock, RN => 
                           n2305, Q => predict_PC_9_13_port, QN => net644037);
   predict_PC_reg_9_12_inst : DFFR_X1 port map( D => n1772, CK => clock, RN => 
                           n2305, Q => predict_PC_9_12_port, QN => net644036);
   predict_PC_reg_9_11_inst : DFFR_X1 port map( D => n1771, CK => clock, RN => 
                           n2305, Q => predict_PC_9_11_port, QN => net644035);
   predict_PC_reg_9_10_inst : DFFR_X1 port map( D => n1770, CK => clock, RN => 
                           n2305, Q => predict_PC_9_10_port, QN => net644034);
   predict_PC_reg_9_9_inst : DFFR_X1 port map( D => n1769, CK => clock, RN => 
                           n2304, Q => predict_PC_9_9_port, QN => net644033);
   predict_PC_reg_9_8_inst : DFFR_X1 port map( D => n1768, CK => clock, RN => 
                           n2305, Q => predict_PC_9_8_port, QN => net644032);
   predict_PC_reg_9_7_inst : DFFR_X1 port map( D => n1767, CK => clock, RN => 
                           n2305, Q => predict_PC_9_7_port, QN => net644031);
   predict_PC_reg_9_6_inst : DFFR_X1 port map( D => n1766, CK => clock, RN => 
                           n2305, Q => predict_PC_9_6_port, QN => net644030);
   predict_PC_reg_9_5_inst : DFFR_X1 port map( D => n1765, CK => clock, RN => 
                           n2295, Q => predict_PC_9_5_port, QN => net644029);
   predict_PC_reg_9_4_inst : DFFR_X1 port map( D => n1764, CK => clock, RN => 
                           n2305, Q => predict_PC_9_4_port, QN => net644028);
   predict_PC_reg_9_3_inst : DFFR_X1 port map( D => n1763, CK => clock, RN => 
                           n2305, Q => predict_PC_9_3_port, QN => net644027);
   predict_PC_reg_9_2_inst : DFFR_X1 port map( D => n1762, CK => clock, RN => 
                           n2305, Q => predict_PC_9_2_port, QN => net644026);
   predict_PC_reg_9_1_inst : DFFR_X1 port map( D => n1761, CK => clock, RN => 
                           n2307, Q => predict_PC_9_1_port, QN => net644025);
   predict_PC_reg_9_0_inst : DFFR_X1 port map( D => n1760, CK => clock, RN => 
                           n2290, Q => predict_PC_9_0_port, QN => net644024);
   predict_PC_reg_10_31_inst : DFFR_X1 port map( D => n1759, CK => clock, RN =>
                           n2310, Q => predict_PC_10_31_port, QN => net644023);
   predict_PC_reg_10_30_inst : DFFR_X1 port map( D => n1758, CK => clock, RN =>
                           n2303, Q => predict_PC_10_30_port, QN => net644022);
   predict_PC_reg_10_29_inst : DFFR_X1 port map( D => n1757, CK => clock, RN =>
                           n2298, Q => predict_PC_10_29_port, QN => net644021);
   predict_PC_reg_10_28_inst : DFFR_X1 port map( D => n1756, CK => clock, RN =>
                           n2310, Q => predict_PC_10_28_port, QN => net644020);
   predict_PC_reg_10_27_inst : DFFR_X1 port map( D => n1755, CK => clock, RN =>
                           n2298, Q => predict_PC_10_27_port, QN => net644019);
   predict_PC_reg_10_26_inst : DFFR_X1 port map( D => n1754, CK => clock, RN =>
                           n2299, Q => predict_PC_10_26_port, QN => net644018);
   predict_PC_reg_10_25_inst : DFFR_X1 port map( D => n1753, CK => clock, RN =>
                           n2300, Q => predict_PC_10_25_port, QN => net644017);
   predict_PC_reg_10_24_inst : DFFR_X1 port map( D => n1752, CK => clock, RN =>
                           n2310, Q => predict_PC_10_24_port, QN => net644016);
   predict_PC_reg_10_23_inst : DFFR_X1 port map( D => n1751, CK => clock, RN =>
                           n2297, Q => predict_PC_10_23_port, QN => net644015);
   predict_PC_reg_10_22_inst : DFFR_X1 port map( D => n1750, CK => clock, RN =>
                           n2288, Q => predict_PC_10_22_port, QN => net644014);
   predict_PC_reg_10_21_inst : DFFR_X1 port map( D => n1749, CK => clock, RN =>
                           n2288, Q => predict_PC_10_21_port, QN => net644013);
   predict_PC_reg_10_20_inst : DFFR_X1 port map( D => n1748, CK => clock, RN =>
                           n2310, Q => predict_PC_10_20_port, QN => net644012);
   predict_PC_reg_10_19_inst : DFFR_X1 port map( D => n1747, CK => clock, RN =>
                           n2311, Q => predict_PC_10_19_port, QN => net644011);
   predict_PC_reg_10_18_inst : DFFR_X1 port map( D => n1746, CK => clock, RN =>
                           n2301, Q => predict_PC_10_18_port, QN => net644010);
   predict_PC_reg_10_17_inst : DFFR_X1 port map( D => n1745, CK => clock, RN =>
                           n2300, Q => predict_PC_10_17_port, QN => net644009);
   predict_PC_reg_10_16_inst : DFFR_X1 port map( D => n1744, CK => clock, RN =>
                           n2310, Q => predict_PC_10_16_port, QN => net644008);
   predict_PC_reg_10_15_inst : DFFR_X1 port map( D => n1743, CK => clock, RN =>
                           n2310, Q => predict_PC_10_15_port, QN => net644007);
   predict_PC_reg_10_14_inst : DFFR_X1 port map( D => n1742, CK => clock, RN =>
                           n2311, Q => predict_PC_10_14_port, QN => net644006);
   predict_PC_reg_10_13_inst : DFFR_X1 port map( D => n1741, CK => clock, RN =>
                           n2310, Q => predict_PC_10_13_port, QN => net644005);
   predict_PC_reg_10_12_inst : DFFR_X1 port map( D => n1740, CK => clock, RN =>
                           n2310, Q => predict_PC_10_12_port, QN => net644004);
   predict_PC_reg_10_11_inst : DFFR_X1 port map( D => n1739, CK => clock, RN =>
                           n2310, Q => predict_PC_10_11_port, QN => net644003);
   predict_PC_reg_10_10_inst : DFFR_X1 port map( D => n1738, CK => clock, RN =>
                           n2310, Q => predict_PC_10_10_port, QN => net644002);
   predict_PC_reg_10_9_inst : DFFR_X1 port map( D => n1737, CK => clock, RN => 
                           n2304, Q => predict_PC_10_9_port, QN => net644001);
   predict_PC_reg_10_8_inst : DFFR_X1 port map( D => n1736, CK => clock, RN => 
                           n2292, Q => predict_PC_10_8_port, QN => net644000);
   predict_PC_reg_10_7_inst : DFFR_X1 port map( D => n1735, CK => clock, RN => 
                           n2289, Q => predict_PC_10_7_port, QN => net643999);
   predict_PC_reg_10_6_inst : DFFR_X1 port map( D => n1734, CK => clock, RN => 
                           n2298, Q => predict_PC_10_6_port, QN => net643998);
   predict_PC_reg_10_5_inst : DFFR_X1 port map( D => n1733, CK => clock, RN => 
                           n2295, Q => predict_PC_10_5_port, QN => net643997);
   predict_PC_reg_10_4_inst : DFFR_X1 port map( D => n1732, CK => clock, RN => 
                           n2311, Q => predict_PC_10_4_port, QN => net643996);
   predict_PC_reg_10_3_inst : DFFR_X1 port map( D => n1731, CK => clock, RN => 
                           n2291, Q => predict_PC_10_3_port, QN => net643995);
   predict_PC_reg_10_2_inst : DFFR_X1 port map( D => n1730, CK => clock, RN => 
                           n2292, Q => predict_PC_10_2_port, QN => net643994);
   predict_PC_reg_10_1_inst : DFFR_X1 port map( D => n1729, CK => clock, RN => 
                           n2307, Q => predict_PC_10_1_port, QN => net643993);
   predict_PC_reg_10_0_inst : DFFR_X1 port map( D => n1728, CK => clock, RN => 
                           n2293, Q => predict_PC_10_0_port, QN => net643992);
   predict_PC_reg_11_31_inst : DFFR_X1 port map( D => n1727, CK => clock, RN =>
                           n2308, Q => predict_PC_11_31_port, QN => net643991);
   predict_PC_reg_11_30_inst : DFFR_X1 port map( D => n1726, CK => clock, RN =>
                           n2303, Q => predict_PC_11_30_port, QN => net643990);
   predict_PC_reg_11_29_inst : DFFR_X1 port map( D => n1725, CK => clock, RN =>
                           n2298, Q => predict_PC_11_29_port, QN => net643989);
   predict_PC_reg_11_28_inst : DFFR_X1 port map( D => n1724, CK => clock, RN =>
                           n2309, Q => predict_PC_11_28_port, QN => net643988);
   predict_PC_reg_11_27_inst : DFFR_X1 port map( D => n1723, CK => clock, RN =>
                           n2298, Q => predict_PC_11_27_port, QN => net643987);
   predict_PC_reg_11_26_inst : DFFR_X1 port map( D => n1722, CK => clock, RN =>
                           n2299, Q => predict_PC_11_26_port, QN => net643986);
   predict_PC_reg_11_25_inst : DFFR_X1 port map( D => n1721, CK => clock, RN =>
                           n2300, Q => predict_PC_11_25_port, QN => net643985);
   predict_PC_reg_11_24_inst : DFFR_X1 port map( D => n1720, CK => clock, RN =>
                           n2309, Q => predict_PC_11_24_port, QN => net643984);
   predict_PC_reg_11_23_inst : DFFR_X1 port map( D => n1719, CK => clock, RN =>
                           n2308, Q => predict_PC_11_23_port, QN => net643983);
   predict_PC_reg_11_22_inst : DFFR_X1 port map( D => n1718, CK => clock, RN =>
                           n2308, Q => predict_PC_11_22_port, QN => net643982);
   predict_PC_reg_11_21_inst : DFFR_X1 port map( D => n1717, CK => clock, RN =>
                           n2292, Q => predict_PC_11_21_port, QN => net643981);
   predict_PC_reg_11_20_inst : DFFR_X1 port map( D => n1716, CK => clock, RN =>
                           n2291, Q => predict_PC_11_20_port, QN => net643980);
   predict_PC_reg_11_19_inst : DFFR_X1 port map( D => n1715, CK => clock, RN =>
                           n2292, Q => predict_PC_11_19_port, QN => net643979);
   predict_PC_reg_11_18_inst : DFFR_X1 port map( D => n1714, CK => clock, RN =>
                           n2301, Q => predict_PC_11_18_port, QN => net643978);
   predict_PC_reg_11_17_inst : DFFR_X1 port map( D => n1713, CK => clock, RN =>
                           n2292, Q => predict_PC_11_17_port, QN => net643977);
   predict_PC_reg_11_16_inst : DFFR_X1 port map( D => n1712, CK => clock, RN =>
                           n2291, Q => predict_PC_11_16_port, QN => net643976);
   predict_PC_reg_11_15_inst : DFFR_X1 port map( D => n1711, CK => clock, RN =>
                           n2292, Q => predict_PC_11_15_port, QN => net643975);
   predict_PC_reg_11_14_inst : DFFR_X1 port map( D => n1710, CK => clock, RN =>
                           n2292, Q => predict_PC_11_14_port, QN => net643974);
   predict_PC_reg_11_13_inst : DFFR_X1 port map( D => n1709, CK => clock, RN =>
                           n2291, Q => predict_PC_11_13_port, QN => net643973);
   predict_PC_reg_11_12_inst : DFFR_X1 port map( D => n1708, CK => clock, RN =>
                           n2291, Q => predict_PC_11_12_port, QN => net643972);
   predict_PC_reg_11_11_inst : DFFR_X1 port map( D => n1707, CK => clock, RN =>
                           n2291, Q => predict_PC_11_11_port, QN => net643971);
   predict_PC_reg_11_10_inst : DFFR_X1 port map( D => n1706, CK => clock, RN =>
                           n2292, Q => predict_PC_11_10_port, QN => net643970);
   predict_PC_reg_11_9_inst : DFFR_X1 port map( D => n1705, CK => clock, RN => 
                           n2303, Q => predict_PC_11_9_port, QN => net643969);
   predict_PC_reg_11_8_inst : DFFR_X1 port map( D => n1704, CK => clock, RN => 
                           n2291, Q => predict_PC_11_8_port, QN => net643968);
   predict_PC_reg_11_7_inst : DFFR_X1 port map( D => n1703, CK => clock, RN => 
                           n2308, Q => predict_PC_11_7_port, QN => net643967);
   predict_PC_reg_11_6_inst : DFFR_X1 port map( D => n1702, CK => clock, RN => 
                           n2308, Q => predict_PC_11_6_port, QN => net643966);
   predict_PC_reg_11_5_inst : DFFR_X1 port map( D => n1701, CK => clock, RN => 
                           n2295, Q => predict_PC_11_5_port, QN => net643965);
   predict_PC_reg_11_4_inst : DFFR_X1 port map( D => n1700, CK => clock, RN => 
                           n2308, Q => predict_PC_11_4_port, QN => net643964);
   predict_PC_reg_11_3_inst : DFFR_X1 port map( D => n1699, CK => clock, RN => 
                           n2308, Q => predict_PC_11_3_port, QN => net643963);
   predict_PC_reg_11_2_inst : DFFR_X1 port map( D => n1698, CK => clock, RN => 
                           n2308, Q => predict_PC_11_2_port, QN => net643962);
   predict_PC_reg_11_1_inst : DFFR_X1 port map( D => n1697, CK => clock, RN => 
                           n2307, Q => predict_PC_11_1_port, QN => net643961);
   predict_PC_reg_11_0_inst : DFFR_X1 port map( D => n1696, CK => clock, RN => 
                           n2308, Q => predict_PC_11_0_port, QN => net643960);
   predict_PC_reg_12_31_inst : DFFR_X1 port map( D => n1695, CK => clock, RN =>
                           n2300, Q => predict_PC_12_31_port, QN => net643959);
   predict_PC_reg_12_30_inst : DFFR_X1 port map( D => n1694, CK => clock, RN =>
                           n2303, Q => predict_PC_12_30_port, QN => net643958);
   predict_PC_reg_12_29_inst : DFFR_X1 port map( D => n1693, CK => clock, RN =>
                           n2298, Q => predict_PC_12_29_port, QN => net643957);
   predict_PC_reg_12_28_inst : DFFR_X1 port map( D => n1692, CK => clock, RN =>
                           n2305, Q => predict_PC_12_28_port, QN => net643956);
   predict_PC_reg_12_27_inst : DFFR_X1 port map( D => n1691, CK => clock, RN =>
                           n2299, Q => predict_PC_12_27_port, QN => net643955);
   predict_PC_reg_12_26_inst : DFFR_X1 port map( D => n1690, CK => clock, RN =>
                           n2299, Q => predict_PC_12_26_port, QN => net643954);
   predict_PC_reg_12_25_inst : DFFR_X1 port map( D => n1689, CK => clock, RN =>
                           n2300, Q => predict_PC_12_25_port, QN => net643953);
   predict_PC_reg_12_24_inst : DFFR_X1 port map( D => n1688, CK => clock, RN =>
                           n2289, Q => predict_PC_12_24_port, QN => net643952);
   predict_PC_reg_12_23_inst : DFFR_X1 port map( D => n1687, CK => clock, RN =>
                           n2294, Q => predict_PC_12_23_port, QN => net643951);
   predict_PC_reg_12_22_inst : DFFR_X1 port map( D => n1686, CK => clock, RN =>
                           n2294, Q => predict_PC_12_22_port, QN => net643950);
   predict_PC_reg_12_21_inst : DFFR_X1 port map( D => n1685, CK => clock, RN =>
                           n2294, Q => predict_PC_12_21_port, QN => net643949);
   predict_PC_reg_12_20_inst : DFFR_X1 port map( D => n1684, CK => clock, RN =>
                           n2294, Q => predict_PC_12_20_port, QN => net643948);
   predict_PC_reg_12_19_inst : DFFR_X1 port map( D => n1683, CK => clock, RN =>
                           n2293, Q => predict_PC_12_19_port, QN => net643947);
   predict_PC_reg_12_18_inst : DFFR_X1 port map( D => n1682, CK => clock, RN =>
                           n2301, Q => predict_PC_12_18_port, QN => net643946);
   predict_PC_reg_12_17_inst : DFFR_X1 port map( D => n1681, CK => clock, RN =>
                           n2293, Q => predict_PC_12_17_port, QN => net643945);
   predict_PC_reg_12_16_inst : DFFR_X1 port map( D => n1680, CK => clock, RN =>
                           n2293, Q => predict_PC_12_16_port, QN => net643944);
   predict_PC_reg_12_15_inst : DFFR_X1 port map( D => n1679, CK => clock, RN =>
                           n2293, Q => predict_PC_12_15_port, QN => net643943);
   predict_PC_reg_12_14_inst : DFFR_X1 port map( D => n1678, CK => clock, RN =>
                           n2293, Q => predict_PC_12_14_port, QN => net643942);
   predict_PC_reg_12_13_inst : DFFR_X1 port map( D => n1677, CK => clock, RN =>
                           n2293, Q => predict_PC_12_13_port, QN => net643941);
   predict_PC_reg_12_12_inst : DFFR_X1 port map( D => n1676, CK => clock, RN =>
                           n2293, Q => predict_PC_12_12_port, QN => net643940);
   predict_PC_reg_12_11_inst : DFFR_X1 port map( D => n1675, CK => clock, RN =>
                           n2293, Q => predict_PC_12_11_port, QN => net643939);
   predict_PC_reg_12_10_inst : DFFR_X1 port map( D => n1674, CK => clock, RN =>
                           n2294, Q => predict_PC_12_10_port, QN => net643938);
   predict_PC_reg_12_9_inst : DFFR_X1 port map( D => n1673, CK => clock, RN => 
                           n2303, Q => predict_PC_12_9_port, QN => net643937);
   predict_PC_reg_12_8_inst : DFFR_X1 port map( D => n1672, CK => clock, RN => 
                           n2294, Q => predict_PC_12_8_port, QN => net643936);
   predict_PC_reg_12_7_inst : DFFR_X1 port map( D => n1671, CK => clock, RN => 
                           n2294, Q => predict_PC_12_7_port, QN => net643935);
   predict_PC_reg_12_6_inst : DFFR_X1 port map( D => n1670, CK => clock, RN => 
                           n2294, Q => predict_PC_12_6_port, QN => net643934);
   predict_PC_reg_12_5_inst : DFFR_X1 port map( D => n1669, CK => clock, RN => 
                           n2295, Q => predict_PC_12_5_port, QN => net643933);
   predict_PC_reg_12_4_inst : DFFR_X1 port map( D => n1668, CK => clock, RN => 
                           n2294, Q => predict_PC_12_4_port, QN => net643932);
   predict_PC_reg_12_3_inst : DFFR_X1 port map( D => n1667, CK => clock, RN => 
                           n2295, Q => predict_PC_12_3_port, QN => net643931);
   predict_PC_reg_12_2_inst : DFFR_X1 port map( D => n1666, CK => clock, RN => 
                           n2295, Q => predict_PC_12_2_port, QN => net643930);
   predict_PC_reg_12_1_inst : DFFR_X1 port map( D => n1665, CK => clock, RN => 
                           n2307, Q => predict_PC_12_1_port, QN => net643929);
   predict_PC_reg_12_0_inst : DFFR_X1 port map( D => n1664, CK => clock, RN => 
                           n2306, Q => predict_PC_12_0_port, QN => net643928);
   predict_PC_reg_13_31_inst : DFFR_X1 port map( D => n1663, CK => clock, RN =>
                           n2294, Q => predict_PC_13_31_port, QN => net643927);
   predict_PC_reg_13_30_inst : DFFR_X1 port map( D => n1662, CK => clock, RN =>
                           n2303, Q => predict_PC_13_30_port, QN => net643926);
   predict_PC_reg_13_29_inst : DFFR_X1 port map( D => n1661, CK => clock, RN =>
                           n2298, Q => predict_PC_13_29_port, QN => net643925);
   predict_PC_reg_13_28_inst : DFFR_X1 port map( D => n1660, CK => clock, RN =>
                           n2303, Q => predict_PC_13_28_port, QN => net643924);
   predict_PC_reg_13_27_inst : DFFR_X1 port map( D => n1659, CK => clock, RN =>
                           n2299, Q => predict_PC_13_27_port, QN => net643923);
   predict_PC_reg_13_26_inst : DFFR_X1 port map( D => n1658, CK => clock, RN =>
                           n2299, Q => predict_PC_13_26_port, QN => net643922);
   predict_PC_reg_13_25_inst : DFFR_X1 port map( D => n1657, CK => clock, RN =>
                           n2301, Q => predict_PC_13_25_port, QN => net643921);
   predict_PC_reg_13_24_inst : DFFR_X1 port map( D => n1656, CK => clock, RN =>
                           n2301, Q => predict_PC_13_24_port, QN => net643920);
   predict_PC_reg_13_23_inst : DFFR_X1 port map( D => n1655, CK => clock, RN =>
                           n2298, Q => predict_PC_13_23_port, QN => net643919);
   predict_PC_reg_13_22_inst : DFFR_X1 port map( D => n1654, CK => clock, RN =>
                           n2292, Q => predict_PC_13_22_port, QN => net643918);
   predict_PC_reg_13_21_inst : DFFR_X1 port map( D => n1653, CK => clock, RN =>
                           n2311, Q => predict_PC_13_21_port, QN => net643917);
   predict_PC_reg_13_20_inst : DFFR_X1 port map( D => n1652, CK => clock, RN =>
                           n2291, Q => predict_PC_13_20_port, QN => net643916);
   predict_PC_reg_13_19_inst : DFFR_X1 port map( D => n1651, CK => clock, RN =>
                           n2293, Q => predict_PC_13_19_port, QN => net643915);
   predict_PC_reg_13_18_inst : DFFR_X1 port map( D => n1650, CK => clock, RN =>
                           n2301, Q => predict_PC_13_18_port, QN => net643914);
   predict_PC_reg_13_17_inst : DFFR_X1 port map( D => n1649, CK => clock, RN =>
                           n2310, Q => predict_PC_13_17_port, QN => net643913);
   predict_PC_reg_13_16_inst : DFFR_X1 port map( D => n1648, CK => clock, RN =>
                           n2296, Q => predict_PC_13_16_port, QN => net643912);
   predict_PC_reg_13_15_inst : DFFR_X1 port map( D => n1647, CK => clock, RN =>
                           n2304, Q => predict_PC_13_15_port, QN => net643911);
   predict_PC_reg_13_14_inst : DFFR_X1 port map( D => n1646, CK => clock, RN =>
                           n2304, Q => predict_PC_13_14_port, QN => net643910);
   predict_PC_reg_13_13_inst : DFFR_X1 port map( D => n1645, CK => clock, RN =>
                           n2304, Q => predict_PC_13_13_port, QN => net643909);
   predict_PC_reg_13_12_inst : DFFR_X1 port map( D => n1644, CK => clock, RN =>
                           n2304, Q => predict_PC_13_12_port, QN => net643908);
   predict_PC_reg_13_11_inst : DFFR_X1 port map( D => n1643, CK => clock, RN =>
                           n2304, Q => predict_PC_13_11_port, QN => net643907);
   predict_PC_reg_13_10_inst : DFFR_X1 port map( D => n1642, CK => clock, RN =>
                           n2304, Q => predict_PC_13_10_port, QN => net643906);
   predict_PC_reg_13_9_inst : DFFR_X1 port map( D => n1641, CK => clock, RN => 
                           n2297, Q => predict_PC_13_9_port, QN => net643905);
   predict_PC_reg_13_8_inst : DFFR_X1 port map( D => n1640, CK => clock, RN => 
                           n2304, Q => predict_PC_13_8_port, QN => net643904);
   predict_PC_reg_13_7_inst : DFFR_X1 port map( D => n1639, CK => clock, RN => 
                           n2304, Q => predict_PC_13_7_port, QN => net643903);
   predict_PC_reg_13_6_inst : DFFR_X1 port map( D => n1638, CK => clock, RN => 
                           n2305, Q => predict_PC_13_6_port, QN => net643902);
   predict_PC_reg_13_5_inst : DFFR_X1 port map( D => n1637, CK => clock, RN => 
                           n2295, Q => predict_PC_13_5_port, QN => net643901);
   predict_PC_reg_13_4_inst : DFFR_X1 port map( D => n1636, CK => clock, RN => 
                           n2305, Q => predict_PC_13_4_port, QN => net643900);
   predict_PC_reg_13_3_inst : DFFR_X1 port map( D => n1635, CK => clock, RN => 
                           n2305, Q => predict_PC_13_3_port, QN => net643899);
   predict_PC_reg_13_2_inst : DFFR_X1 port map( D => n1634, CK => clock, RN => 
                           n2305, Q => predict_PC_13_2_port, QN => net643898);
   predict_PC_reg_13_1_inst : DFFR_X1 port map( D => n1633, CK => clock, RN => 
                           n2307, Q => predict_PC_13_1_port, QN => net643897);
   predict_PC_reg_13_0_inst : DFFR_X1 port map( D => n1632, CK => clock, RN => 
                           n2297, Q => predict_PC_13_0_port, QN => net643896);
   predict_PC_reg_14_31_inst : DFFR_X1 port map( D => n1631, CK => clock, RN =>
                           n2296, Q => predict_PC_14_31_port, QN => net643895);
   predict_PC_reg_14_30_inst : DFFR_X1 port map( D => n1630, CK => clock, RN =>
                           n2297, Q => predict_PC_14_30_port, QN => net643894);
   predict_PC_reg_14_29_inst : DFFR_X1 port map( D => n1629, CK => clock, RN =>
                           n2298, Q => predict_PC_14_29_port, QN => net643893);
   predict_PC_reg_14_28_inst : DFFR_X1 port map( D => n1628, CK => clock, RN =>
                           n2290, Q => predict_PC_14_28_port, QN => net643892);
   predict_PC_reg_14_27_inst : DFFR_X1 port map( D => n1627, CK => clock, RN =>
                           n2299, Q => predict_PC_14_27_port, QN => net643891);
   predict_PC_reg_14_26_inst : DFFR_X1 port map( D => n1626, CK => clock, RN =>
                           n2299, Q => predict_PC_14_26_port, QN => net643890);
   predict_PC_reg_14_25_inst : DFFR_X1 port map( D => n1625, CK => clock, RN =>
                           n2301, Q => predict_PC_14_25_port, QN => net643889);
   predict_PC_reg_14_24_inst : DFFR_X1 port map( D => n1624, CK => clock, RN =>
                           n2302, Q => predict_PC_14_24_port, QN => net643888);
   predict_PC_reg_14_23_inst : DFFR_X1 port map( D => n1623, CK => clock, RN =>
                           n2299, Q => predict_PC_14_23_port, QN => net643887);
   predict_PC_reg_14_22_inst : DFFR_X1 port map( D => n1622, CK => clock, RN =>
                           n2288, Q => predict_PC_14_22_port, QN => net643886);
   predict_PC_reg_14_21_inst : DFFR_X1 port map( D => n1621, CK => clock, RN =>
                           n2288, Q => predict_PC_14_21_port, QN => net643885);
   predict_PC_reg_14_20_inst : DFFR_X1 port map( D => n1620, CK => clock, RN =>
                           n2307, Q => predict_PC_14_20_port, QN => net643884);
   predict_PC_reg_14_19_inst : DFFR_X1 port map( D => n1619, CK => clock, RN =>
                           n2311, Q => predict_PC_14_19_port, QN => net643883);
   predict_PC_reg_14_18_inst : DFFR_X1 port map( D => n1618, CK => clock, RN =>
                           n2301, Q => predict_PC_14_18_port, QN => net643882);
   predict_PC_reg_14_17_inst : DFFR_X1 port map( D => n1617, CK => clock, RN =>
                           n2300, Q => predict_PC_14_17_port, QN => net643881);
   predict_PC_reg_14_16_inst : DFFR_X1 port map( D => n1616, CK => clock, RN =>
                           n2304, Q => predict_PC_14_16_port, QN => net643880);
   predict_PC_reg_14_15_inst : DFFR_X1 port map( D => n1615, CK => clock, RN =>
                           n2289, Q => predict_PC_14_15_port, QN => net643879);
   predict_PC_reg_14_14_inst : DFFR_X1 port map( D => n1614, CK => clock, RN =>
                           n2311, Q => predict_PC_14_14_port, QN => net643878);
   predict_PC_reg_14_13_inst : DFFR_X1 port map( D => n1613, CK => clock, RN =>
                           n2305, Q => predict_PC_14_13_port, QN => net643877);
   predict_PC_reg_14_12_inst : DFFR_X1 port map( D => n1612, CK => clock, RN =>
                           n2304, Q => predict_PC_14_12_port, QN => net643876);
   predict_PC_reg_14_11_inst : DFFR_X1 port map( D => n1611, CK => clock, RN =>
                           n2307, Q => predict_PC_14_11_port, QN => net643875);
   predict_PC_reg_14_10_inst : DFFR_X1 port map( D => n1610, CK => clock, RN =>
                           n2302, Q => predict_PC_14_10_port, QN => net643874);
   predict_PC_reg_14_9_inst : DFFR_X1 port map( D => n1609, CK => clock, RN => 
                           n2297, Q => predict_PC_14_9_port, QN => net643873);
   predict_PC_reg_14_8_inst : DFFR_X1 port map( D => n1608, CK => clock, RN => 
                           n2290, Q => predict_PC_14_8_port, QN => net643872);
   predict_PC_reg_14_7_inst : DFFR_X1 port map( D => n1607, CK => clock, RN => 
                           n2289, Q => predict_PC_14_7_port, QN => net643871);
   predict_PC_reg_14_6_inst : DFFR_X1 port map( D => n1606, CK => clock, RN => 
                           n2294, Q => predict_PC_14_6_port, QN => net643870);
   predict_PC_reg_14_5_inst : DFFR_X1 port map( D => n1605, CK => clock, RN => 
                           n2295, Q => predict_PC_14_5_port, QN => net643869);
   predict_PC_reg_14_4_inst : DFFR_X1 port map( D => n1604, CK => clock, RN => 
                           n2296, Q => predict_PC_14_4_port, QN => net643868);
   predict_PC_reg_14_3_inst : DFFR_X1 port map( D => n1603, CK => clock, RN => 
                           n2310, Q => predict_PC_14_3_port, QN => net643867);
   predict_PC_reg_14_2_inst : DFFR_X1 port map( D => n1602, CK => clock, RN => 
                           n2309, Q => predict_PC_14_2_port, QN => net643866);
   predict_PC_reg_14_1_inst : DFFR_X1 port map( D => n1601, CK => clock, RN => 
                           n2307, Q => predict_PC_14_1_port, QN => net643865);
   predict_PC_reg_14_0_inst : DFFR_X1 port map( D => n1600, CK => clock, RN => 
                           n2293, Q => predict_PC_14_0_port, QN => net643864);
   predict_PC_reg_15_31_inst : DFFR_X1 port map( D => n1599, CK => clock, RN =>
                           n2299, Q => predict_PC_15_31_port, QN => net643863);
   last_PC_reg_31_inst : DFFR_X1 port map( D => n1598, CK => clock, RN => n2297
                           , Q => net684157, QN => n593);
   predict_PC_reg_15_30_inst : DFFR_X1 port map( D => n1597, CK => clock, RN =>
                           n2297, Q => predict_PC_15_30_port, QN => net643862);
   last_PC_reg_30_inst : DFFR_X1 port map( D => n1596, CK => clock, RN => n2297
                           , Q => n6, QN => net684156);
   predict_PC_reg_15_29_inst : DFFR_X1 port map( D => n1595, CK => clock, RN =>
                           n2298, Q => predict_PC_15_29_port, QN => net643861);
   last_PC_reg_29_inst : DFFR_X1 port map( D => n1594, CK => clock, RN => n2298
                           , Q => n7, QN => net684155);
   predict_PC_reg_15_28_inst : DFFR_X1 port map( D => n1593, CK => clock, RN =>
                           n2297, Q => predict_PC_15_28_port, QN => net643860);
   last_PC_reg_28_inst : DFFR_X1 port map( D => n1592, CK => clock, RN => n2297
                           , Q => n8, QN => net684154);
   predict_PC_reg_15_27_inst : DFFR_X1 port map( D => n1591, CK => clock, RN =>
                           n2299, Q => predict_PC_15_27_port, QN => net643859);
   last_PC_reg_27_inst : DFFR_X1 port map( D => n1590, CK => clock, RN => n2303
                           , Q => n9, QN => net684153);
   predict_PC_reg_15_26_inst : DFFR_X1 port map( D => n1589, CK => clock, RN =>
                           n2302, Q => predict_PC_15_26_port, QN => net643858);
   last_PC_reg_26_inst : DFFR_X1 port map( D => n1588, CK => clock, RN => n2302
                           , Q => net684152, QN => n598);
   predict_PC_reg_15_25_inst : DFFR_X1 port map( D => n1587, CK => clock, RN =>
                           n2301, Q => predict_PC_15_25_port, QN => net643857);
   last_PC_reg_25_inst : DFFR_X1 port map( D => n1586, CK => clock, RN => n2301
                           , Q => net684151, QN => n599);
   predict_PC_reg_15_24_inst : DFFR_X1 port map( D => n1585, CK => clock, RN =>
                           n2309, Q => predict_PC_15_24_port, QN => net643856);
   last_PC_reg_24_inst : DFFR_X1 port map( D => n1584, CK => clock, RN => n2297
                           , Q => net684150, QN => n600);
   predict_PC_reg_15_23_inst : DFFR_X1 port map( D => n1583, CK => clock, RN =>
                           n2306, Q => predict_PC_15_23_port, QN => net643855);
   last_PC_reg_23_inst : DFFR_X1 port map( D => n1582, CK => clock, RN => n2301
                           , Q => net684149, QN => n601);
   predict_PC_reg_15_22_inst : DFFR_X1 port map( D => n1581, CK => clock, RN =>
                           n2288, Q => predict_PC_15_22_port, QN => net643854);
   last_PC_reg_22_inst : DFFR_X1 port map( D => n1580, CK => clock, RN => n2301
                           , Q => net684148, QN => n602);
   predict_PC_reg_15_21_inst : DFFR_X1 port map( D => n1579, CK => clock, RN =>
                           n2288, Q => predict_PC_15_21_port, QN => net643853);
   last_PC_reg_21_inst : DFFR_X1 port map( D => n1578, CK => clock, RN => n2301
                           , Q => net684147, QN => n603);
   predict_PC_reg_15_20_inst : DFFR_X1 port map( D => n1577, CK => clock, RN =>
                           n2304, Q => predict_PC_15_20_port, QN => net643852);
   last_PC_reg_20_inst : DFFR_X1 port map( D => n1576, CK => clock, RN => n2297
                           , Q => net684146, QN => n604);
   predict_PC_reg_15_19_inst : DFFR_X1 port map( D => n1575, CK => clock, RN =>
                           n2311, Q => predict_PC_15_19_port, QN => net643851);
   last_PC_reg_19_inst : DFFR_X1 port map( D => n1574, CK => clock, RN => n2301
                           , Q => net684145, QN => n605);
   predict_PC_reg_15_18_inst : DFFR_X1 port map( D => n1573, CK => clock, RN =>
                           n2300, Q => predict_PC_15_18_port, QN => net643850);
   last_PC_reg_18_inst : DFFR_X1 port map( D => n1572, CK => clock, RN => n2304
                           , Q => net684144, QN => n606);
   predict_PC_reg_15_17_inst : DFFR_X1 port map( D => n1571, CK => clock, RN =>
                           n2300, Q => predict_PC_15_17_port, QN => net643849);
   last_PC_reg_17_inst : DFFR_X1 port map( D => n1570, CK => clock, RN => n2300
                           , Q => net684143, QN => n607);
   predict_PC_reg_15_16_inst : DFFR_X1 port map( D => n1569, CK => clock, RN =>
                           n2300, Q => predict_PC_15_16_port, QN => net643848);
   last_PC_reg_16_inst : DFFR_X1 port map( D => n1568, CK => clock, RN => n2297
                           , Q => net684142, QN => n608);
   predict_PC_reg_15_15_inst : DFFR_X1 port map( D => n1567, CK => clock, RN =>
                           n2290, Q => predict_PC_15_15_port, QN => net643847);
   last_PC_reg_15_inst : DFFR_X1 port map( D => n1566, CK => clock, RN => n2303
                           , Q => net684141, QN => n609);
   predict_PC_reg_15_14_inst : DFFR_X1 port map( D => n1565, CK => clock, RN =>
                           n2311, Q => predict_PC_15_14_port, QN => net643846);
   last_PC_reg_14_inst : DFFR_X1 port map( D => n1564, CK => clock, RN => n2301
                           , Q => net684140, QN => n610);
   predict_PC_reg_15_13_inst : DFFR_X1 port map( D => n1563, CK => clock, RN =>
                           n2290, Q => predict_PC_15_13_port, QN => net643845);
   last_PC_reg_13_inst : DFFR_X1 port map( D => n1562, CK => clock, RN => n2303
                           , Q => net684139, QN => n611);
   predict_PC_reg_15_12_inst : DFFR_X1 port map( D => n1561, CK => clock, RN =>
                           n2296, Q => predict_PC_15_12_port, QN => net643844);
   last_PC_reg_12_inst : DFFR_X1 port map( D => n1560, CK => clock, RN => n2297
                           , Q => net684138, QN => n612);
   predict_PC_reg_15_11_inst : DFFR_X1 port map( D => n1559, CK => clock, RN =>
                           n2298, Q => predict_PC_15_11_port, QN => net643843);
   last_PC_reg_11_inst : DFFR_X1 port map( D => n1558, CK => clock, RN => n2298
                           , Q => net684137, QN => n613);
   predict_PC_reg_15_10_inst : DFFR_X1 port map( D => n1557, CK => clock, RN =>
                           n2310, Q => predict_PC_15_10_port, QN => net643842);
   last_PC_reg_10_inst : DFFR_X1 port map( D => n1556, CK => clock, RN => n2302
                           , Q => net684136, QN => n614);
   predict_PC_reg_15_9_inst : DFFR_X1 port map( D => n1555, CK => clock, RN => 
                           n2297, Q => predict_PC_15_9_port, QN => net643841);
   last_PC_reg_9_inst : DFFR_X1 port map( D => n1554, CK => clock, RN => n2297,
                           Q => net684135, QN => n615);
   predict_PC_reg_15_8_inst : DFFR_X1 port map( D => n1553, CK => clock, RN => 
                           n2294, Q => predict_PC_15_8_port, QN => net643840);
   last_PC_reg_8_inst : DFFR_X1 port map( D => n1552, CK => clock, RN => n2298,
                           Q => net684134, QN => n616);
   predict_PC_reg_15_7_inst : DFFR_X1 port map( D => n1551, CK => clock, RN => 
                           n2289, Q => predict_PC_15_7_port, QN => net643839);
   last_PC_reg_7_inst : DFFR_X1 port map( D => n1550, CK => clock, RN => n2301,
                           Q => net684133, QN => n617);
   predict_PC_reg_15_6_inst : DFFR_X1 port map( D => n1549, CK => clock, RN => 
                           n2303, Q => predict_PC_15_6_port, QN => net643838);
   last_PC_reg_6_inst : DFFR_X1 port map( D => n1548, CK => clock, RN => n2289,
                           Q => net684132, QN => n618);
   predict_PC_reg_15_5_inst : DFFR_X1 port map( D => n1547, CK => clock, RN => 
                           n2295, Q => predict_PC_15_5_port, QN => net643837);
   last_PC_reg_5_inst : DFFR_X1 port map( D => n1546, CK => clock, RN => n2295,
                           Q => net684131, QN => n619);
   predict_PC_reg_15_4_inst : DFFR_X1 port map( D => n1545, CK => clock, RN => 
                           n2301, Q => predict_PC_15_4_port, QN => net643836);
   last_PC_reg_4_inst : DFFR_X1 port map( D => n1544, CK => clock, RN => n2297,
                           Q => net684130, QN => n620);
   predict_PC_reg_15_3_inst : DFFR_X1 port map( D => n1543, CK => clock, RN => 
                           n2310, Q => predict_PC_15_3_port, QN => net643835);
   last_PC_reg_3_inst : DFFR_X1 port map( D => n1542, CK => clock, RN => n2302,
                           Q => net684129, QN => n621);
   predict_PC_reg_15_2_inst : DFFR_X1 port map( D => n1541, CK => clock, RN => 
                           n2297, Q => predict_PC_15_2_port, QN => net643834);
   last_PC_reg_2_inst : DFFR_X1 port map( D => n1540, CK => clock, RN => n2307,
                           Q => net684128, QN => n622);
   predict_PC_reg_15_1_inst : DFFR_X1 port map( D => n1539, CK => clock, RN => 
                           n2307, Q => predict_PC_15_1_port, QN => net643833);
   last_PC_reg_1_inst : DFFR_X1 port map( D => n1538, CK => clock, RN => n2295,
                           Q => net684127, QN => n623);
   predict_PC_reg_15_0_inst : DFFR_X1 port map( D => n1537, CK => clock, RN => 
                           n2307, Q => predict_PC_15_0_port, QN => net643832);
   last_PC_reg_0_inst : DFFR_X1 port map( D => n1536, CK => clock, RN => n2297,
                           Q => net684126, QN => n624);
   last_mispredict_reg : DFFR_X1 port map( D => n1535, CK => clock, RN => n2294
                           , Q => net684125, QN => n592);
   U1603 : MUX2_X1 port map( A => n6, B => predicted_next_PC_o_30_port, S => 
                           n2286, Z => n1596);
   U1604 : MUX2_X1 port map( A => n7, B => predicted_next_PC_o_29_port, S => 
                           n2286, Z => n1594);
   U1605 : MUX2_X1 port map( A => n8, B => predicted_next_PC_o_28_port, S => 
                           n2286, Z => n1592);
   U1606 : MUX2_X1 port map( A => n9, B => predicted_next_PC_o_27_port, S => 
                           n2286, Z => n1590);
   pred_x_0 : predictor_2_0 port map( clock => clock, reset => reset, enable =>
                           write_enable_0_port, taken_i => was_taken_i, 
                           prediction_o => taken_0_port);
   pred_x_1 : predictor_2_15 port map( clock => clock, reset => reset, enable 
                           => write_enable_1_port, taken_i => was_taken_i, 
                           prediction_o => taken_1_port);
   pred_x_2 : predictor_2_14 port map( clock => clock, reset => reset, enable 
                           => write_enable_2_port, taken_i => was_taken_i, 
                           prediction_o => taken_2_port);
   pred_x_3 : predictor_2_13 port map( clock => clock, reset => reset, enable 
                           => write_enable_3_port, taken_i => was_taken_i, 
                           prediction_o => taken_3_port);
   pred_x_4 : predictor_2_12 port map( clock => clock, reset => reset, enable 
                           => write_enable_4_port, taken_i => was_taken_i, 
                           prediction_o => taken_4_port);
   pred_x_5 : predictor_2_11 port map( clock => clock, reset => reset, enable 
                           => write_enable_5_port, taken_i => was_taken_i, 
                           prediction_o => taken_5_port);
   pred_x_6 : predictor_2_10 port map( clock => clock, reset => reset, enable 
                           => write_enable_6_port, taken_i => was_taken_i, 
                           prediction_o => taken_6_port);
   pred_x_7 : predictor_2_9 port map( clock => clock, reset => reset, enable =>
                           write_enable_7_port, taken_i => was_taken_i, 
                           prediction_o => taken_7_port);
   pred_x_8 : predictor_2_8 port map( clock => clock, reset => reset, enable =>
                           write_enable_8_port, taken_i => was_taken_i, 
                           prediction_o => taken_8_port);
   pred_x_9 : predictor_2_7 port map( clock => clock, reset => reset, enable =>
                           write_enable_9_port, taken_i => was_taken_i, 
                           prediction_o => taken_9_port);
   pred_x_10 : predictor_2_6 port map( clock => clock, reset => reset, enable 
                           => write_enable_10_port, taken_i => was_taken_i, 
                           prediction_o => taken_10_port);
   pred_x_11 : predictor_2_5 port map( clock => clock, reset => reset, enable 
                           => write_enable_11_port, taken_i => was_taken_i, 
                           prediction_o => taken_11_port);
   pred_x_12 : predictor_2_4 port map( clock => clock, reset => reset, enable 
                           => write_enable_12_port, taken_i => was_taken_i, 
                           prediction_o => taken_12_port);
   pred_x_13 : predictor_2_3 port map( clock => clock, reset => reset, enable 
                           => write_enable_13_port, taken_i => was_taken_i, 
                           prediction_o => taken_13_port);
   pred_x_14 : predictor_2_2 port map( clock => clock, reset => reset, enable 
                           => write_enable_14_port, taken_i => was_taken_i, 
                           prediction_o => taken_14_port);
   pred_x_15 : predictor_2_1 port map( clock => clock, reset => reset, enable 
                           => write_enable_15_port, taken_i => was_taken_i, 
                           prediction_o => taken_15_port);
   U1552 : NAND2_X1 port map( A1 => TAG_i(2), A2 => TAG_i(3), ZN => n2209);
   U1542 : NAND2_X1 port map( A1 => TAG_i(0), A2 => n701, ZN => n2200);
   U80 : AOI22_X1 port map( A1 => n2270, A2 => taken_12_port, B1 => n763, B2 =>
                           taken_13_port, ZN => n752);
   U1548 : NAND2_X1 port map( A1 => TAG_i(1), A2 => TAG_i(0), ZN => n2202);
   U79 : AOI22_X1 port map( A1 => n2272, A2 => taken_14_port, B1 => n761, B2 =>
                           taken_15_port, ZN => n753);
   U78 : AOI22_X1 port map( A1 => n2274, A2 => taken_10_port, B1 => n759, B2 =>
                           taken_11_port, ZN => n754);
   U77 : AOI22_X1 port map( A1 => n2276, A2 => taken_8_port, B1 => n757, B2 => 
                           taken_9_port, ZN => n755);
   U75 : AOI22_X1 port map( A1 => n2278, A2 => taken_4_port, B1 => n751, B2 => 
                           taken_5_port, ZN => n740);
   U74 : AOI22_X1 port map( A1 => n2280, A2 => taken_6_port, B1 => n749, B2 => 
                           taken_7_port, ZN => n741);
   U73 : AOI22_X1 port map( A1 => n746, A2 => taken_1_port, B1 => n2281, B2 => 
                           taken_0_port, ZN => n742);
   U72 : AOI22_X1 port map( A1 => n744, A2 => taken_3_port, B1 => n745, B2 => 
                           taken_2_port, ZN => n743);
   U1367 : AOI22_X1 port map( A1 => n2272, A2 => predict_PC_14_11_port, B1 => 
                           n2271, B2 => predict_PC_15_11_port, ZN => n1511);
   U1366 : AOI22_X1 port map( A1 => n2270, A2 => predict_PC_12_11_port, B1 => 
                           n2269, B2 => predict_PC_13_11_port, ZN => n1512);
   U1365 : AOI22_X1 port map( A1 => n2276, A2 => predict_PC_8_11_port, B1 => 
                           n2275, B2 => predict_PC_9_11_port, ZN => n1513);
   U1364 : AOI22_X1 port map( A1 => n2274, A2 => predict_PC_10_11_port, B1 => 
                           n2273, B2 => predict_PC_11_11_port, ZN => n1514);
   U1363 : NAND4_X1 port map( A1 => n1511, A2 => n1512, A3 => n1513, A4 => 
                           n1514, ZN => n1505);
   U1362 : AOI22_X1 port map( A1 => n2280, A2 => predict_PC_6_11_port, B1 => 
                           n2279, B2 => predict_PC_7_11_port, ZN => n1507);
   U1361 : AOI22_X1 port map( A1 => n2278, A2 => predict_PC_4_11_port, B1 => 
                           n2277, B2 => predict_PC_5_11_port, ZN => n1508);
   U1360 : AOI22_X1 port map( A1 => n2284, A2 => predict_PC_3_11_port, B1 => 
                           n2283, B2 => predict_PC_2_11_port, ZN => n1509);
   U1359 : AOI22_X1 port map( A1 => n2282, A2 => predict_PC_1_11_port, B1 => 
                           n2281, B2 => predict_PC_0_11_port, ZN => n1510);
   U1358 : NAND4_X1 port map( A1 => n1507, A2 => n1508, A3 => n1509, A4 => 
                           n1510, ZN => n1506);
   U1357 : NOR2_X1 port map( A1 => n1505, A2 => n1506, ZN => n691);
   U1325 : AOI22_X1 port map( A1 => n2272, A2 => predict_PC_14_14_port, B1 => 
                           n2271, B2 => predict_PC_15_14_port, ZN => n1478);
   U1324 : AOI22_X1 port map( A1 => n2270, A2 => predict_PC_12_14_port, B1 => 
                           n2269, B2 => predict_PC_13_14_port, ZN => n1479);
   U1323 : AOI22_X1 port map( A1 => n2276, A2 => predict_PC_8_14_port, B1 => 
                           n2275, B2 => predict_PC_9_14_port, ZN => n1480);
   U1322 : AOI22_X1 port map( A1 => n2274, A2 => predict_PC_10_14_port, B1 => 
                           n2273, B2 => predict_PC_11_14_port, ZN => n1481);
   U1321 : NAND4_X1 port map( A1 => n1478, A2 => n1479, A3 => n1480, A4 => 
                           n1481, ZN => n1472);
   U1320 : AOI22_X1 port map( A1 => n2280, A2 => predict_PC_6_14_port, B1 => 
                           n2279, B2 => predict_PC_7_14_port, ZN => n1474);
   U1319 : AOI22_X1 port map( A1 => n2278, A2 => predict_PC_4_14_port, B1 => 
                           n2277, B2 => predict_PC_5_14_port, ZN => n1475);
   U1318 : AOI22_X1 port map( A1 => n2284, A2 => predict_PC_3_14_port, B1 => 
                           n2283, B2 => predict_PC_2_14_port, ZN => n1476);
   U1317 : AOI22_X1 port map( A1 => n2282, A2 => predict_PC_1_14_port, B1 => 
                           n2281, B2 => predict_PC_0_14_port, ZN => n1477);
   U1316 : NAND4_X1 port map( A1 => n1474, A2 => n1475, A3 => n1476, A4 => 
                           n1477, ZN => n1473);
   U1315 : NOR2_X1 port map( A1 => n1472, A2 => n1473, ZN => n688);
   U1381 : AOI22_X1 port map( A1 => n2272, A2 => predict_PC_14_10_port, B1 => 
                           n2271, B2 => predict_PC_15_10_port, ZN => n1522);
   U1380 : AOI22_X1 port map( A1 => n2270, A2 => predict_PC_12_10_port, B1 => 
                           n2269, B2 => predict_PC_13_10_port, ZN => n1523);
   U1379 : AOI22_X1 port map( A1 => n2276, A2 => predict_PC_8_10_port, B1 => 
                           n2275, B2 => predict_PC_9_10_port, ZN => n1524);
   U1378 : AOI22_X1 port map( A1 => n2274, A2 => predict_PC_10_10_port, B1 => 
                           n2273, B2 => predict_PC_11_10_port, ZN => n1525);
   U1377 : NAND4_X1 port map( A1 => n1522, A2 => n1523, A3 => n1524, A4 => 
                           n1525, ZN => n1516);
   U1376 : AOI22_X1 port map( A1 => n2280, A2 => predict_PC_6_10_port, B1 => 
                           n2279, B2 => predict_PC_7_10_port, ZN => n1518);
   U1375 : AOI22_X1 port map( A1 => n2278, A2 => predict_PC_4_10_port, B1 => 
                           n2277, B2 => predict_PC_5_10_port, ZN => n1519);
   U1374 : AOI22_X1 port map( A1 => n2284, A2 => predict_PC_3_10_port, B1 => 
                           n2283, B2 => predict_PC_2_10_port, ZN => n1520);
   U1373 : AOI22_X1 port map( A1 => n2282, A2 => predict_PC_1_10_port, B1 => 
                           n2281, B2 => predict_PC_0_10_port, ZN => n1521);
   U1372 : NAND4_X1 port map( A1 => n1518, A2 => n1519, A3 => n1520, A4 => 
                           n1521, ZN => n1517);
   U1371 : NOR2_X1 port map( A1 => n1516, A2 => n1517, ZN => n692);
   U1091 : AOI22_X1 port map( A1 => n2272, A2 => predict_PC_14_31_port, B1 => 
                           n2271, B2 => predict_PC_15_31_port, ZN => n1291);
   U1090 : AOI22_X1 port map( A1 => n2270, A2 => predict_PC_12_31_port, B1 => 
                           n2269, B2 => predict_PC_13_31_port, ZN => n1292);
   U1089 : AOI22_X1 port map( A1 => n2276, A2 => predict_PC_8_31_port, B1 => 
                           n2275, B2 => predict_PC_9_31_port, ZN => n1293);
   U1088 : AOI22_X1 port map( A1 => n2274, A2 => predict_PC_10_31_port, B1 => 
                           n2273, B2 => predict_PC_11_31_port, ZN => n1294);
   U1087 : NAND4_X1 port map( A1 => n1291, A2 => n1292, A3 => n1293, A4 => 
                           n1294, ZN => n1285);
   U1086 : AOI22_X1 port map( A1 => n2280, A2 => predict_PC_6_31_port, B1 => 
                           n2279, B2 => predict_PC_7_31_port, ZN => n1287);
   U1085 : AOI22_X1 port map( A1 => n2278, A2 => predict_PC_4_31_port, B1 => 
                           n2277, B2 => predict_PC_5_31_port, ZN => n1288);
   U1084 : AOI22_X1 port map( A1 => n2284, A2 => predict_PC_3_31_port, B1 => 
                           n2283, B2 => predict_PC_2_31_port, ZN => n1289);
   U1083 : AOI22_X1 port map( A1 => n2282, A2 => predict_PC_1_31_port, B1 => 
                           n2281, B2 => predict_PC_0_31_port, ZN => n1290);
   U1082 : NAND4_X1 port map( A1 => n1287, A2 => n1288, A3 => n1289, A4 => 
                           n1290, ZN => n1286);
   U1081 : NOR2_X1 port map( A1 => n1285, A2 => n1286, ZN => n673);
   U1297 : AOI22_X1 port map( A1 => n760, A2 => predict_PC_14_16_port, B1 => 
                           n2271, B2 => predict_PC_15_16_port, ZN => n1456);
   U1296 : AOI22_X1 port map( A1 => n762, A2 => predict_PC_12_16_port, B1 => 
                           n2269, B2 => predict_PC_13_16_port, ZN => n1457);
   U1295 : AOI22_X1 port map( A1 => n756, A2 => predict_PC_8_16_port, B1 => 
                           n2275, B2 => predict_PC_9_16_port, ZN => n1458);
   U1294 : AOI22_X1 port map( A1 => n758, A2 => predict_PC_10_16_port, B1 => 
                           n2273, B2 => predict_PC_11_16_port, ZN => n1459);
   U1293 : NAND4_X1 port map( A1 => n1456, A2 => n1457, A3 => n1458, A4 => 
                           n1459, ZN => n1450);
   U1292 : AOI22_X1 port map( A1 => n748, A2 => predict_PC_6_16_port, B1 => 
                           n2279, B2 => predict_PC_7_16_port, ZN => n1452);
   U1291 : AOI22_X1 port map( A1 => n750, A2 => predict_PC_4_16_port, B1 => 
                           n2277, B2 => predict_PC_5_16_port, ZN => n1453);
   U1290 : AOI22_X1 port map( A1 => n2284, A2 => predict_PC_3_16_port, B1 => 
                           n2283, B2 => predict_PC_2_16_port, ZN => n1454);
   U1289 : AOI22_X1 port map( A1 => n2282, A2 => predict_PC_1_16_port, B1 => 
                           n747, B2 => predict_PC_0_16_port, ZN => n1455);
   U1288 : NAND4_X1 port map( A1 => n1452, A2 => n1453, A3 => n1454, A4 => 
                           n1455, ZN => n1451);
   U1287 : NOR2_X1 port map( A1 => n1450, A2 => n1451, ZN => n686);
   U1311 : AOI22_X1 port map( A1 => n760, A2 => predict_PC_14_15_port, B1 => 
                           n2271, B2 => predict_PC_15_15_port, ZN => n1467);
   U1310 : AOI22_X1 port map( A1 => n2270, A2 => predict_PC_12_15_port, B1 => 
                           n2269, B2 => predict_PC_13_15_port, ZN => n1468);
   U1309 : AOI22_X1 port map( A1 => n2276, A2 => predict_PC_8_15_port, B1 => 
                           n2275, B2 => predict_PC_9_15_port, ZN => n1469);
   U1308 : AOI22_X1 port map( A1 => n2274, A2 => predict_PC_10_15_port, B1 => 
                           n2273, B2 => predict_PC_11_15_port, ZN => n1470);
   U1307 : NAND4_X1 port map( A1 => n1467, A2 => n1468, A3 => n1469, A4 => 
                           n1470, ZN => n1461);
   U1306 : AOI22_X1 port map( A1 => n748, A2 => predict_PC_6_15_port, B1 => 
                           n2279, B2 => predict_PC_7_15_port, ZN => n1463);
   U1305 : AOI22_X1 port map( A1 => n750, A2 => predict_PC_4_15_port, B1 => 
                           n2277, B2 => predict_PC_5_15_port, ZN => n1464);
   U1304 : AOI22_X1 port map( A1 => n2284, A2 => predict_PC_3_15_port, B1 => 
                           n2283, B2 => predict_PC_2_15_port, ZN => n1465);
   U1303 : AOI22_X1 port map( A1 => n2282, A2 => predict_PC_1_15_port, B1 => 
                           n747, B2 => predict_PC_0_15_port, ZN => n1466);
   U1302 : NAND4_X1 port map( A1 => n1463, A2 => n1464, A3 => n1465, A4 => 
                           n1466, ZN => n1462);
   U1301 : NOR2_X1 port map( A1 => n1461, A2 => n1462, ZN => n687);
   U1269 : AOI22_X1 port map( A1 => n2272, A2 => predict_PC_14_18_port, B1 => 
                           n2271, B2 => predict_PC_15_18_port, ZN => n1434);
   U1268 : AOI22_X1 port map( A1 => n762, A2 => predict_PC_12_18_port, B1 => 
                           n2269, B2 => predict_PC_13_18_port, ZN => n1435);
   U1267 : AOI22_X1 port map( A1 => n756, A2 => predict_PC_8_18_port, B1 => 
                           n2275, B2 => predict_PC_9_18_port, ZN => n1436);
   U1266 : AOI22_X1 port map( A1 => n758, A2 => predict_PC_10_18_port, B1 => 
                           n2273, B2 => predict_PC_11_18_port, ZN => n1437);
   U1265 : NAND4_X1 port map( A1 => n1434, A2 => n1435, A3 => n1436, A4 => 
                           n1437, ZN => n1428);
   U1264 : AOI22_X1 port map( A1 => n748, A2 => predict_PC_6_18_port, B1 => 
                           n2279, B2 => predict_PC_7_18_port, ZN => n1430);
   U1263 : AOI22_X1 port map( A1 => n2278, A2 => predict_PC_4_18_port, B1 => 
                           n2277, B2 => predict_PC_5_18_port, ZN => n1431);
   U1262 : AOI22_X1 port map( A1 => n2284, A2 => predict_PC_3_18_port, B1 => 
                           n2283, B2 => predict_PC_2_18_port, ZN => n1432);
   U1261 : AOI22_X1 port map( A1 => n2282, A2 => predict_PC_1_18_port, B1 => 
                           n747, B2 => predict_PC_0_18_port, ZN => n1433);
   U1260 : NAND4_X1 port map( A1 => n1430, A2 => n1431, A3 => n1432, A4 => 
                           n1433, ZN => n1429);
   U1259 : NOR2_X1 port map( A1 => n1428, A2 => n1429, ZN => n684);
   U1283 : AOI22_X1 port map( A1 => n760, A2 => predict_PC_14_17_port, B1 => 
                           n2271, B2 => predict_PC_15_17_port, ZN => n1445);
   U1282 : AOI22_X1 port map( A1 => n762, A2 => predict_PC_12_17_port, B1 => 
                           n2269, B2 => predict_PC_13_17_port, ZN => n1446);
   U1281 : AOI22_X1 port map( A1 => n756, A2 => predict_PC_8_17_port, B1 => 
                           n2275, B2 => predict_PC_9_17_port, ZN => n1447);
   U1280 : AOI22_X1 port map( A1 => n758, A2 => predict_PC_10_17_port, B1 => 
                           n2273, B2 => predict_PC_11_17_port, ZN => n1448);
   U1279 : NAND4_X1 port map( A1 => n1445, A2 => n1446, A3 => n1447, A4 => 
                           n1448, ZN => n1439);
   U1278 : AOI22_X1 port map( A1 => n2280, A2 => predict_PC_6_17_port, B1 => 
                           n2279, B2 => predict_PC_7_17_port, ZN => n1441);
   U1277 : AOI22_X1 port map( A1 => n750, A2 => predict_PC_4_17_port, B1 => 
                           n2277, B2 => predict_PC_5_17_port, ZN => n1442);
   U1276 : AOI22_X1 port map( A1 => n2284, A2 => predict_PC_3_17_port, B1 => 
                           n2283, B2 => predict_PC_2_17_port, ZN => n1443);
   U1275 : AOI22_X1 port map( A1 => n2282, A2 => predict_PC_1_17_port, B1 => 
                           n747, B2 => predict_PC_0_17_port, ZN => n1444);
   U1274 : NAND4_X1 port map( A1 => n1441, A2 => n1442, A3 => n1443, A4 => 
                           n1444, ZN => n1440);
   U1273 : NOR2_X1 port map( A1 => n1439, A2 => n1440, ZN => n685);
   U1185 : AOI22_X1 port map( A1 => n2272, A2 => predict_PC_14_24_port, B1 => 
                           n2271, B2 => predict_PC_15_24_port, ZN => n1368);
   U1184 : AOI22_X1 port map( A1 => n2270, A2 => predict_PC_12_24_port, B1 => 
                           n2269, B2 => predict_PC_13_24_port, ZN => n1369);
   U1183 : AOI22_X1 port map( A1 => n2276, A2 => predict_PC_8_24_port, B1 => 
                           n2275, B2 => predict_PC_9_24_port, ZN => n1370);
   U1182 : AOI22_X1 port map( A1 => n2274, A2 => predict_PC_10_24_port, B1 => 
                           n2273, B2 => predict_PC_11_24_port, ZN => n1371);
   U1181 : NAND4_X1 port map( A1 => n1368, A2 => n1369, A3 => n1370, A4 => 
                           n1371, ZN => n1362);
   U1180 : AOI22_X1 port map( A1 => n2280, A2 => predict_PC_6_24_port, B1 => 
                           n2279, B2 => predict_PC_7_24_port, ZN => n1364);
   U1179 : AOI22_X1 port map( A1 => n2278, A2 => predict_PC_4_24_port, B1 => 
                           n2277, B2 => predict_PC_5_24_port, ZN => n1365);
   U1178 : AOI22_X1 port map( A1 => n2284, A2 => predict_PC_3_24_port, B1 => 
                           n2283, B2 => predict_PC_2_24_port, ZN => n1366);
   U1177 : AOI22_X1 port map( A1 => n2282, A2 => predict_PC_1_24_port, B1 => 
                           n2281, B2 => predict_PC_0_24_port, ZN => n1367);
   U1176 : NAND4_X1 port map( A1 => n1364, A2 => n1365, A3 => n1366, A4 => 
                           n1367, ZN => n1363);
   U1175 : NOR2_X1 port map( A1 => n1362, A2 => n1363, ZN => n677);
   U1143 : AOI22_X1 port map( A1 => n2272, A2 => predict_PC_14_27_port, B1 => 
                           n2271, B2 => predict_PC_15_27_port, ZN => n1335);
   U1142 : AOI22_X1 port map( A1 => n2270, A2 => predict_PC_12_27_port, B1 => 
                           n2269, B2 => predict_PC_13_27_port, ZN => n1336);
   U1141 : AOI22_X1 port map( A1 => n2276, A2 => predict_PC_8_27_port, B1 => 
                           n2275, B2 => predict_PC_9_27_port, ZN => n1337);
   U1140 : AOI22_X1 port map( A1 => n2274, A2 => predict_PC_10_27_port, B1 => 
                           n2273, B2 => predict_PC_11_27_port, ZN => n1338);
   U1139 : NAND4_X1 port map( A1 => n1335, A2 => n1336, A3 => n1337, A4 => 
                           n1338, ZN => n1329);
   U1138 : AOI22_X1 port map( A1 => n2280, A2 => predict_PC_6_27_port, B1 => 
                           n2279, B2 => predict_PC_7_27_port, ZN => n1331);
   U1137 : AOI22_X1 port map( A1 => n2278, A2 => predict_PC_4_27_port, B1 => 
                           n2277, B2 => predict_PC_5_27_port, ZN => n1332);
   U1136 : AOI22_X1 port map( A1 => n2284, A2 => predict_PC_3_27_port, B1 => 
                           n2283, B2 => predict_PC_2_27_port, ZN => n1333);
   U1135 : AOI22_X1 port map( A1 => n2282, A2 => predict_PC_1_27_port, B1 => 
                           n2281, B2 => predict_PC_0_27_port, ZN => n1334);
   U1134 : NAND4_X1 port map( A1 => n1331, A2 => n1332, A3 => n1333, A4 => 
                           n1334, ZN => n1330);
   U1213 : AOI22_X1 port map( A1 => n2272, A2 => predict_PC_14_22_port, B1 => 
                           n2271, B2 => predict_PC_15_22_port, ZN => n1390);
   U1212 : AOI22_X1 port map( A1 => n2270, A2 => predict_PC_12_22_port, B1 => 
                           n2269, B2 => predict_PC_13_22_port, ZN => n1391);
   U1211 : AOI22_X1 port map( A1 => n2276, A2 => predict_PC_8_22_port, B1 => 
                           n2275, B2 => predict_PC_9_22_port, ZN => n1392);
   U1210 : AOI22_X1 port map( A1 => n2274, A2 => predict_PC_10_22_port, B1 => 
                           n2273, B2 => predict_PC_11_22_port, ZN => n1393);
   U1209 : NAND4_X1 port map( A1 => n1390, A2 => n1391, A3 => n1392, A4 => 
                           n1393, ZN => n1384);
   U1208 : AOI22_X1 port map( A1 => n2280, A2 => predict_PC_6_22_port, B1 => 
                           n2279, B2 => predict_PC_7_22_port, ZN => n1386);
   U1207 : AOI22_X1 port map( A1 => n2278, A2 => predict_PC_4_22_port, B1 => 
                           n2277, B2 => predict_PC_5_22_port, ZN => n1387);
   U1206 : AOI22_X1 port map( A1 => n2284, A2 => predict_PC_3_22_port, B1 => 
                           n2283, B2 => predict_PC_2_22_port, ZN => n1388);
   U1205 : AOI22_X1 port map( A1 => n2282, A2 => predict_PC_1_22_port, B1 => 
                           n2281, B2 => predict_PC_0_22_port, ZN => n1389);
   U1204 : NAND4_X1 port map( A1 => n1386, A2 => n1387, A3 => n1388, A4 => 
                           n1389, ZN => n1385);
   U1203 : NOR2_X1 port map( A1 => n1384, A2 => n1385, ZN => n679);
   U1255 : AOI22_X1 port map( A1 => n2272, A2 => predict_PC_14_19_port, B1 => 
                           n2271, B2 => predict_PC_15_19_port, ZN => n1423);
   U1254 : AOI22_X1 port map( A1 => n2270, A2 => predict_PC_12_19_port, B1 => 
                           n2269, B2 => predict_PC_13_19_port, ZN => n1424);
   U1253 : AOI22_X1 port map( A1 => n2276, A2 => predict_PC_8_19_port, B1 => 
                           n2275, B2 => predict_PC_9_19_port, ZN => n1425);
   U1252 : AOI22_X1 port map( A1 => n2274, A2 => predict_PC_10_19_port, B1 => 
                           n2273, B2 => predict_PC_11_19_port, ZN => n1426);
   U1251 : NAND4_X1 port map( A1 => n1423, A2 => n1424, A3 => n1425, A4 => 
                           n1426, ZN => n1417);
   U1250 : AOI22_X1 port map( A1 => n2280, A2 => predict_PC_6_19_port, B1 => 
                           n2279, B2 => predict_PC_7_19_port, ZN => n1419);
   U1249 : AOI22_X1 port map( A1 => n2278, A2 => predict_PC_4_19_port, B1 => 
                           n2277, B2 => predict_PC_5_19_port, ZN => n1420);
   U1248 : AOI22_X1 port map( A1 => n2284, A2 => predict_PC_3_19_port, B1 => 
                           n2283, B2 => predict_PC_2_19_port, ZN => n1421);
   U1247 : AOI22_X1 port map( A1 => n2282, A2 => predict_PC_1_19_port, B1 => 
                           n2281, B2 => predict_PC_0_19_port, ZN => n1422);
   U1246 : NAND4_X1 port map( A1 => n1419, A2 => n1420, A3 => n1421, A4 => 
                           n1422, ZN => n1418);
   U1245 : NOR2_X1 port map( A1 => n1417, A2 => n1418, ZN => n683);
   U1199 : AOI22_X1 port map( A1 => n2272, A2 => predict_PC_14_23_port, B1 => 
                           n2271, B2 => predict_PC_15_23_port, ZN => n1379);
   U1198 : AOI22_X1 port map( A1 => n2270, A2 => predict_PC_12_23_port, B1 => 
                           n2269, B2 => predict_PC_13_23_port, ZN => n1380);
   U1197 : AOI22_X1 port map( A1 => n2276, A2 => predict_PC_8_23_port, B1 => 
                           n2275, B2 => predict_PC_9_23_port, ZN => n1381);
   U1196 : AOI22_X1 port map( A1 => n2274, A2 => predict_PC_10_23_port, B1 => 
                           n2273, B2 => predict_PC_11_23_port, ZN => n1382);
   U1195 : NAND4_X1 port map( A1 => n1379, A2 => n1380, A3 => n1381, A4 => 
                           n1382, ZN => n1373);
   U1194 : AOI22_X1 port map( A1 => n2280, A2 => predict_PC_6_23_port, B1 => 
                           n2279, B2 => predict_PC_7_23_port, ZN => n1375);
   U1193 : AOI22_X1 port map( A1 => n2278, A2 => predict_PC_4_23_port, B1 => 
                           n2277, B2 => predict_PC_5_23_port, ZN => n1376);
   U1192 : AOI22_X1 port map( A1 => n2284, A2 => predict_PC_3_23_port, B1 => 
                           n2283, B2 => predict_PC_2_23_port, ZN => n1377);
   U1191 : AOI22_X1 port map( A1 => n2282, A2 => predict_PC_1_23_port, B1 => 
                           n2281, B2 => predict_PC_0_23_port, ZN => n1378);
   U1190 : NAND4_X1 port map( A1 => n1375, A2 => n1376, A3 => n1377, A4 => 
                           n1378, ZN => n1374);
   U1189 : NOR2_X1 port map( A1 => n1373, A2 => n1374, ZN => n678);
   U1171 : AOI22_X1 port map( A1 => n2272, A2 => predict_PC_14_25_port, B1 => 
                           n2271, B2 => predict_PC_15_25_port, ZN => n1357);
   U1170 : AOI22_X1 port map( A1 => n2270, A2 => predict_PC_12_25_port, B1 => 
                           n2269, B2 => predict_PC_13_25_port, ZN => n1358);
   U1169 : AOI22_X1 port map( A1 => n2276, A2 => predict_PC_8_25_port, B1 => 
                           n2275, B2 => predict_PC_9_25_port, ZN => n1359);
   U1168 : AOI22_X1 port map( A1 => n2274, A2 => predict_PC_10_25_port, B1 => 
                           n2273, B2 => predict_PC_11_25_port, ZN => n1360);
   U1167 : NAND4_X1 port map( A1 => n1357, A2 => n1358, A3 => n1359, A4 => 
                           n1360, ZN => n1351);
   U1166 : AOI22_X1 port map( A1 => n2280, A2 => predict_PC_6_25_port, B1 => 
                           n2279, B2 => predict_PC_7_25_port, ZN => n1353);
   U1165 : AOI22_X1 port map( A1 => n2278, A2 => predict_PC_4_25_port, B1 => 
                           n2277, B2 => predict_PC_5_25_port, ZN => n1354);
   U1164 : AOI22_X1 port map( A1 => n2284, A2 => predict_PC_3_25_port, B1 => 
                           n2283, B2 => predict_PC_2_25_port, ZN => n1355);
   U1163 : AOI22_X1 port map( A1 => n2282, A2 => predict_PC_1_25_port, B1 => 
                           n2281, B2 => predict_PC_0_25_port, ZN => n1356);
   U1162 : NAND4_X1 port map( A1 => n1353, A2 => n1354, A3 => n1355, A4 => 
                           n1356, ZN => n1352);
   U1161 : NOR2_X1 port map( A1 => n1351, A2 => n1352, ZN => n676);
   U1157 : AOI22_X1 port map( A1 => n2272, A2 => predict_PC_14_26_port, B1 => 
                           n2271, B2 => predict_PC_15_26_port, ZN => n1346);
   U1156 : AOI22_X1 port map( A1 => n2270, A2 => predict_PC_12_26_port, B1 => 
                           n2269, B2 => predict_PC_13_26_port, ZN => n1347);
   U1155 : AOI22_X1 port map( A1 => n2276, A2 => predict_PC_8_26_port, B1 => 
                           n2275, B2 => predict_PC_9_26_port, ZN => n1348);
   U1154 : AOI22_X1 port map( A1 => n2274, A2 => predict_PC_10_26_port, B1 => 
                           n2273, B2 => predict_PC_11_26_port, ZN => n1349);
   U1153 : NAND4_X1 port map( A1 => n1346, A2 => n1347, A3 => n1348, A4 => 
                           n1349, ZN => n1340);
   U1152 : AOI22_X1 port map( A1 => n2280, A2 => predict_PC_6_26_port, B1 => 
                           n2279, B2 => predict_PC_7_26_port, ZN => n1342);
   U1151 : AOI22_X1 port map( A1 => n2278, A2 => predict_PC_4_26_port, B1 => 
                           n2277, B2 => predict_PC_5_26_port, ZN => n1343);
   U1150 : AOI22_X1 port map( A1 => n2284, A2 => predict_PC_3_26_port, B1 => 
                           n2283, B2 => predict_PC_2_26_port, ZN => n1344);
   U1149 : AOI22_X1 port map( A1 => n2282, A2 => predict_PC_1_26_port, B1 => 
                           n2281, B2 => predict_PC_0_26_port, ZN => n1345);
   U1148 : NAND4_X1 port map( A1 => n1342, A2 => n1343, A3 => n1344, A4 => 
                           n1345, ZN => n1341);
   U1147 : NOR2_X1 port map( A1 => n1340, A2 => n1341, ZN => n675);
   U1423 : AOI22_X1 port map( A1 => n760, A2 => predict_PC_14_7_port, B1 => 
                           n2271, B2 => predict_PC_15_7_port, ZN => n2121);
   U1422 : AOI22_X1 port map( A1 => n762, A2 => predict_PC_12_7_port, B1 => 
                           n2269, B2 => predict_PC_13_7_port, ZN => n2122);
   U1421 : AOI22_X1 port map( A1 => n756, A2 => predict_PC_8_7_port, B1 => 
                           n2275, B2 => predict_PC_9_7_port, ZN => n2123);
   U1420 : AOI22_X1 port map( A1 => n758, A2 => predict_PC_10_7_port, B1 => 
                           n2273, B2 => predict_PC_11_7_port, ZN => n2124);
   U1419 : NAND4_X1 port map( A1 => n2121, A2 => n2122, A3 => n2123, A4 => 
                           n2124, ZN => n2115);
   U1418 : AOI22_X1 port map( A1 => n748, A2 => predict_PC_6_7_port, B1 => 
                           n2279, B2 => predict_PC_7_7_port, ZN => n2117);
   U1417 : AOI22_X1 port map( A1 => n750, A2 => predict_PC_4_7_port, B1 => 
                           n2277, B2 => predict_PC_5_7_port, ZN => n2118);
   U1416 : AOI22_X1 port map( A1 => n2284, A2 => predict_PC_3_7_port, B1 => 
                           n2283, B2 => predict_PC_2_7_port, ZN => n2119);
   U1415 : AOI22_X1 port map( A1 => n2282, A2 => predict_PC_1_7_port, B1 => 
                           n747, B2 => predict_PC_0_7_port, ZN => n2120);
   U1414 : NAND4_X1 port map( A1 => n2117, A2 => n2118, A3 => n2119, A4 => 
                           n2120, ZN => n2116);
   U1413 : NOR2_X1 port map( A1 => n2115, A2 => n2116, ZN => n668);
   U1479 : AOI22_X1 port map( A1 => n2272, A2 => predict_PC_14_3_port, B1 => 
                           n2271, B2 => predict_PC_15_3_port, ZN => n2165);
   U1478 : AOI22_X1 port map( A1 => n2270, A2 => predict_PC_12_3_port, B1 => 
                           n2269, B2 => predict_PC_13_3_port, ZN => n2166);
   U1477 : AOI22_X1 port map( A1 => n2276, A2 => predict_PC_8_3_port, B1 => 
                           n2275, B2 => predict_PC_9_3_port, ZN => n2167);
   U1476 : AOI22_X1 port map( A1 => n2274, A2 => predict_PC_10_3_port, B1 => 
                           n2273, B2 => predict_PC_11_3_port, ZN => n2168);
   U1475 : NAND4_X1 port map( A1 => n2165, A2 => n2166, A3 => n2167, A4 => 
                           n2168, ZN => n2159);
   U1474 : AOI22_X1 port map( A1 => n2280, A2 => predict_PC_6_3_port, B1 => 
                           n2279, B2 => predict_PC_7_3_port, ZN => n2161);
   U1473 : AOI22_X1 port map( A1 => n2278, A2 => predict_PC_4_3_port, B1 => 
                           n2277, B2 => predict_PC_5_3_port, ZN => n2162);
   U1472 : AOI22_X1 port map( A1 => n2284, A2 => predict_PC_3_3_port, B1 => 
                           n2283, B2 => predict_PC_2_3_port, ZN => n2163);
   U1471 : AOI22_X1 port map( A1 => n2282, A2 => predict_PC_1_3_port, B1 => 
                           n2281, B2 => predict_PC_0_3_port, ZN => n2164);
   U1470 : NAND4_X1 port map( A1 => n2161, A2 => n2162, A3 => n2163, A4 => 
                           n2164, ZN => n2160);
   U1469 : NOR2_X1 port map( A1 => n2159, A2 => n2160, ZN => n672);
   U1227 : AOI22_X1 port map( A1 => n2272, A2 => predict_PC_14_21_port, B1 => 
                           n2271, B2 => predict_PC_15_21_port, ZN => n1401);
   U1226 : AOI22_X1 port map( A1 => n2270, A2 => predict_PC_12_21_port, B1 => 
                           n2269, B2 => predict_PC_13_21_port, ZN => n1402);
   U1225 : AOI22_X1 port map( A1 => n2276, A2 => predict_PC_8_21_port, B1 => 
                           n2275, B2 => predict_PC_9_21_port, ZN => n1403);
   U1224 : AOI22_X1 port map( A1 => n2274, A2 => predict_PC_10_21_port, B1 => 
                           n2273, B2 => predict_PC_11_21_port, ZN => n1404);
   U1223 : NAND4_X1 port map( A1 => n1401, A2 => n1402, A3 => n1403, A4 => 
                           n1404, ZN => n1395);
   U1222 : AOI22_X1 port map( A1 => n2280, A2 => predict_PC_6_21_port, B1 => 
                           n2279, B2 => predict_PC_7_21_port, ZN => n1397);
   U1221 : AOI22_X1 port map( A1 => n2278, A2 => predict_PC_4_21_port, B1 => 
                           n2277, B2 => predict_PC_5_21_port, ZN => n1398);
   U1220 : AOI22_X1 port map( A1 => n2284, A2 => predict_PC_3_21_port, B1 => 
                           n2283, B2 => predict_PC_2_21_port, ZN => n1399);
   U1219 : AOI22_X1 port map( A1 => n2282, A2 => predict_PC_1_21_port, B1 => 
                           n2281, B2 => predict_PC_0_21_port, ZN => n1400);
   U1218 : NAND4_X1 port map( A1 => n1397, A2 => n1398, A3 => n1399, A4 => 
                           n1400, ZN => n1396);
   U1217 : NOR2_X1 port map( A1 => n1395, A2 => n1396, ZN => n680);
   U1241 : AOI22_X1 port map( A1 => n2272, A2 => predict_PC_14_20_port, B1 => 
                           n2271, B2 => predict_PC_15_20_port, ZN => n1412);
   U1240 : AOI22_X1 port map( A1 => n2270, A2 => predict_PC_12_20_port, B1 => 
                           n2269, B2 => predict_PC_13_20_port, ZN => n1413);
   U1239 : AOI22_X1 port map( A1 => n2276, A2 => predict_PC_8_20_port, B1 => 
                           n2275, B2 => predict_PC_9_20_port, ZN => n1414);
   U1238 : AOI22_X1 port map( A1 => n2274, A2 => predict_PC_10_20_port, B1 => 
                           n2273, B2 => predict_PC_11_20_port, ZN => n1415);
   U1237 : NAND4_X1 port map( A1 => n1412, A2 => n1413, A3 => n1414, A4 => 
                           n1415, ZN => n1406);
   U1236 : AOI22_X1 port map( A1 => n2280, A2 => predict_PC_6_20_port, B1 => 
                           n2279, B2 => predict_PC_7_20_port, ZN => n1408);
   U1235 : AOI22_X1 port map( A1 => n2278, A2 => predict_PC_4_20_port, B1 => 
                           n2277, B2 => predict_PC_5_20_port, ZN => n1409);
   U1234 : AOI22_X1 port map( A1 => n2284, A2 => predict_PC_3_20_port, B1 => 
                           n2283, B2 => predict_PC_2_20_port, ZN => n1410);
   U1233 : AOI22_X1 port map( A1 => n2282, A2 => predict_PC_1_20_port, B1 => 
                           n2281, B2 => predict_PC_0_20_port, ZN => n1411);
   U1232 : NAND4_X1 port map( A1 => n1408, A2 => n1409, A3 => n1410, A4 => 
                           n1411, ZN => n1407);
   U1231 : NOR2_X1 port map( A1 => n1406, A2 => n1407, ZN => n681);
   U1437 : AOI22_X1 port map( A1 => n2272, A2 => predict_PC_14_6_port, B1 => 
                           n2271, B2 => predict_PC_15_6_port, ZN => n2132);
   U1436 : AOI22_X1 port map( A1 => n2270, A2 => predict_PC_12_6_port, B1 => 
                           n2269, B2 => predict_PC_13_6_port, ZN => n2133);
   U1435 : AOI22_X1 port map( A1 => n2276, A2 => predict_PC_8_6_port, B1 => 
                           n2275, B2 => predict_PC_9_6_port, ZN => n2134);
   U1434 : AOI22_X1 port map( A1 => n2274, A2 => predict_PC_10_6_port, B1 => 
                           n2273, B2 => predict_PC_11_6_port, ZN => n2135);
   U1433 : NAND4_X1 port map( A1 => n2132, A2 => n2133, A3 => n2134, A4 => 
                           n2135, ZN => n2126);
   U1432 : AOI22_X1 port map( A1 => n2280, A2 => predict_PC_6_6_port, B1 => 
                           n2279, B2 => predict_PC_7_6_port, ZN => n2128);
   U1431 : AOI22_X1 port map( A1 => n2278, A2 => predict_PC_4_6_port, B1 => 
                           n2277, B2 => predict_PC_5_6_port, ZN => n2129);
   U1430 : AOI22_X1 port map( A1 => n2284, A2 => predict_PC_3_6_port, B1 => 
                           n2283, B2 => predict_PC_2_6_port, ZN => n2130);
   U1429 : AOI22_X1 port map( A1 => n2282, A2 => predict_PC_1_6_port, B1 => 
                           n2281, B2 => predict_PC_0_6_port, ZN => n2131);
   U1428 : NAND4_X1 port map( A1 => n2128, A2 => n2129, A3 => n2130, A4 => 
                           n2131, ZN => n2127);
   U1427 : NOR2_X1 port map( A1 => n2126, A2 => n2127, ZN => n669);
   U1409 : AOI22_X1 port map( A1 => n2272, A2 => predict_PC_14_8_port, B1 => 
                           n2271, B2 => predict_PC_15_8_port, ZN => n2110);
   U1408 : AOI22_X1 port map( A1 => n2270, A2 => predict_PC_12_8_port, B1 => 
                           n2269, B2 => predict_PC_13_8_port, ZN => n2111);
   U1407 : AOI22_X1 port map( A1 => n2276, A2 => predict_PC_8_8_port, B1 => 
                           n2275, B2 => predict_PC_9_8_port, ZN => n2112);
   U1406 : AOI22_X1 port map( A1 => n2274, A2 => predict_PC_10_8_port, B1 => 
                           n2273, B2 => predict_PC_11_8_port, ZN => n2113);
   U1405 : NAND4_X1 port map( A1 => n2110, A2 => n2111, A3 => n2112, A4 => 
                           n2113, ZN => n2104);
   U1404 : AOI22_X1 port map( A1 => n2280, A2 => predict_PC_6_8_port, B1 => 
                           n2279, B2 => predict_PC_7_8_port, ZN => n2106);
   U1403 : AOI22_X1 port map( A1 => n2278, A2 => predict_PC_4_8_port, B1 => 
                           n2277, B2 => predict_PC_5_8_port, ZN => n2107);
   U1402 : AOI22_X1 port map( A1 => n2284, A2 => predict_PC_3_8_port, B1 => 
                           n2283, B2 => predict_PC_2_8_port, ZN => n2108);
   U1401 : AOI22_X1 port map( A1 => n2282, A2 => predict_PC_1_8_port, B1 => 
                           n2281, B2 => predict_PC_0_8_port, ZN => n2109);
   U1400 : NAND4_X1 port map( A1 => n2106, A2 => n2107, A3 => n2108, A4 => 
                           n2109, ZN => n2105);
   U1399 : NOR2_X1 port map( A1 => n2104, A2 => n2105, ZN => n667);
   U1395 : AOI22_X1 port map( A1 => n760, A2 => predict_PC_14_9_port, B1 => 
                           n2271, B2 => predict_PC_15_9_port, ZN => n1533);
   U1394 : AOI22_X1 port map( A1 => n762, A2 => predict_PC_12_9_port, B1 => 
                           n2269, B2 => predict_PC_13_9_port, ZN => n1534);
   U1393 : AOI22_X1 port map( A1 => n756, A2 => predict_PC_8_9_port, B1 => 
                           n2275, B2 => predict_PC_9_9_port, ZN => n2101);
   U1392 : AOI22_X1 port map( A1 => n758, A2 => predict_PC_10_9_port, B1 => 
                           n2273, B2 => predict_PC_11_9_port, ZN => n2102);
   U1391 : NAND4_X1 port map( A1 => n1533, A2 => n1534, A3 => n2101, A4 => 
                           n2102, ZN => n1527);
   U1390 : AOI22_X1 port map( A1 => n748, A2 => predict_PC_6_9_port, B1 => 
                           n2279, B2 => predict_PC_7_9_port, ZN => n1529);
   U1389 : AOI22_X1 port map( A1 => n750, A2 => predict_PC_4_9_port, B1 => 
                           n2277, B2 => predict_PC_5_9_port, ZN => n1530);
   U1388 : AOI22_X1 port map( A1 => n2284, A2 => predict_PC_3_9_port, B1 => 
                           n2283, B2 => predict_PC_2_9_port, ZN => n1531);
   U1387 : AOI22_X1 port map( A1 => n2282, A2 => predict_PC_1_9_port, B1 => 
                           n747, B2 => predict_PC_0_9_port, ZN => n1532);
   U1386 : NAND4_X1 port map( A1 => n1529, A2 => n1530, A3 => n1531, A4 => 
                           n1532, ZN => n1528);
   U1385 : NOR2_X1 port map( A1 => n1527, A2 => n1528, ZN => n666);
   U1493 : AOI22_X1 port map( A1 => n2272, A2 => predict_PC_14_2_port, B1 => 
                           n2271, B2 => predict_PC_15_2_port, ZN => n2176);
   U1492 : AOI22_X1 port map( A1 => n2270, A2 => predict_PC_12_2_port, B1 => 
                           n2269, B2 => predict_PC_13_2_port, ZN => n2177);
   U1491 : AOI22_X1 port map( A1 => n2276, A2 => predict_PC_8_2_port, B1 => 
                           n2275, B2 => predict_PC_9_2_port, ZN => n2178);
   U1490 : AOI22_X1 port map( A1 => n2274, A2 => predict_PC_10_2_port, B1 => 
                           n2273, B2 => predict_PC_11_2_port, ZN => n2179);
   U1489 : NAND4_X1 port map( A1 => n2176, A2 => n2177, A3 => n2178, A4 => 
                           n2179, ZN => n2170);
   U1488 : AOI22_X1 port map( A1 => n2280, A2 => predict_PC_6_2_port, B1 => 
                           n2279, B2 => predict_PC_7_2_port, ZN => n2172);
   U1487 : AOI22_X1 port map( A1 => n2278, A2 => predict_PC_4_2_port, B1 => 
                           n2277, B2 => predict_PC_5_2_port, ZN => n2173);
   U1486 : AOI22_X1 port map( A1 => n2284, A2 => predict_PC_3_2_port, B1 => 
                           n2283, B2 => predict_PC_2_2_port, ZN => n2174);
   U1485 : AOI22_X1 port map( A1 => n2282, A2 => predict_PC_1_2_port, B1 => 
                           n2281, B2 => predict_PC_0_2_port, ZN => n2175);
   U1484 : NAND4_X1 port map( A1 => n2172, A2 => n2173, A3 => n2174, A4 => 
                           n2175, ZN => n2171);
   U1483 : NOR2_X1 port map( A1 => n2170, A2 => n2171, ZN => n674);
   U1465 : AOI22_X1 port map( A1 => n2272, A2 => predict_PC_14_4_port, B1 => 
                           n2271, B2 => predict_PC_15_4_port, ZN => n2154);
   U1464 : AOI22_X1 port map( A1 => n2270, A2 => predict_PC_12_4_port, B1 => 
                           n2269, B2 => predict_PC_13_4_port, ZN => n2155);
   U1463 : AOI22_X1 port map( A1 => n2276, A2 => predict_PC_8_4_port, B1 => 
                           n2275, B2 => predict_PC_9_4_port, ZN => n2156);
   U1462 : AOI22_X1 port map( A1 => n2274, A2 => predict_PC_10_4_port, B1 => 
                           n2273, B2 => predict_PC_11_4_port, ZN => n2157);
   U1461 : NAND4_X1 port map( A1 => n2154, A2 => n2155, A3 => n2156, A4 => 
                           n2157, ZN => n2148);
   U1460 : AOI22_X1 port map( A1 => n2280, A2 => predict_PC_6_4_port, B1 => 
                           n2279, B2 => predict_PC_7_4_port, ZN => n2150);
   U1459 : AOI22_X1 port map( A1 => n2278, A2 => predict_PC_4_4_port, B1 => 
                           n2277, B2 => predict_PC_5_4_port, ZN => n2151);
   U1458 : AOI22_X1 port map( A1 => n2284, A2 => predict_PC_3_4_port, B1 => 
                           n2283, B2 => predict_PC_2_4_port, ZN => n2152);
   U1457 : AOI22_X1 port map( A1 => n2282, A2 => predict_PC_1_4_port, B1 => 
                           n2281, B2 => predict_PC_0_4_port, ZN => n2153);
   U1456 : NAND4_X1 port map( A1 => n2150, A2 => n2151, A3 => n2152, A4 => 
                           n2153, ZN => n2149);
   U1455 : NOR2_X1 port map( A1 => n2148, A2 => n2149, ZN => n671);
   U1117 : AOI22_X1 port map( A1 => n2272, A2 => predict_PC_14_29_port, B1 => 
                           n761, B2 => predict_PC_15_29_port, ZN => n1313);
   U1116 : AOI22_X1 port map( A1 => n2270, A2 => predict_PC_12_29_port, B1 => 
                           n2269, B2 => predict_PC_13_29_port, ZN => n1314);
   U1115 : AOI22_X1 port map( A1 => n2276, A2 => predict_PC_8_29_port, B1 => 
                           n2275, B2 => predict_PC_9_29_port, ZN => n1315);
   U1114 : AOI22_X1 port map( A1 => n2274, A2 => predict_PC_10_29_port, B1 => 
                           n2273, B2 => predict_PC_11_29_port, ZN => n1316);
   U1113 : NAND4_X1 port map( A1 => n1313, A2 => n1314, A3 => n1315, A4 => 
                           n1316, ZN => n1307);
   U1112 : AOI22_X1 port map( A1 => n2280, A2 => predict_PC_6_29_port, B1 => 
                           n2279, B2 => predict_PC_7_29_port, ZN => n1309);
   U1111 : AOI22_X1 port map( A1 => n2278, A2 => predict_PC_4_29_port, B1 => 
                           n2277, B2 => predict_PC_5_29_port, ZN => n1310);
   U1110 : AOI22_X1 port map( A1 => n2284, A2 => predict_PC_3_29_port, B1 => 
                           n2283, B2 => predict_PC_2_29_port, ZN => n1311);
   U1109 : AOI22_X1 port map( A1 => n2282, A2 => predict_PC_1_29_port, B1 => 
                           n2281, B2 => predict_PC_0_29_port, ZN => n1312);
   U1108 : NAND4_X1 port map( A1 => n1309, A2 => n1310, A3 => n1311, A4 => 
                           n1312, ZN => n1308);
   U1451 : AOI22_X1 port map( A1 => n760, A2 => predict_PC_14_5_port, B1 => 
                           n2271, B2 => predict_PC_15_5_port, ZN => n2143);
   U1450 : AOI22_X1 port map( A1 => n762, A2 => predict_PC_12_5_port, B1 => 
                           n2269, B2 => predict_PC_13_5_port, ZN => n2144);
   U1449 : AOI22_X1 port map( A1 => n756, A2 => predict_PC_8_5_port, B1 => 
                           n2275, B2 => predict_PC_9_5_port, ZN => n2145);
   U1448 : AOI22_X1 port map( A1 => n758, A2 => predict_PC_10_5_port, B1 => 
                           n2273, B2 => predict_PC_11_5_port, ZN => n2146);
   U1447 : NAND4_X1 port map( A1 => n2143, A2 => n2144, A3 => n2145, A4 => 
                           n2146, ZN => n2137);
   U1446 : AOI22_X1 port map( A1 => n748, A2 => predict_PC_6_5_port, B1 => 
                           n2279, B2 => predict_PC_7_5_port, ZN => n2139);
   U1445 : AOI22_X1 port map( A1 => n750, A2 => predict_PC_4_5_port, B1 => 
                           n2277, B2 => predict_PC_5_5_port, ZN => n2140);
   U1444 : AOI22_X1 port map( A1 => n2284, A2 => predict_PC_3_5_port, B1 => 
                           n2283, B2 => predict_PC_2_5_port, ZN => n2141);
   U1443 : AOI22_X1 port map( A1 => n2282, A2 => predict_PC_1_5_port, B1 => 
                           n747, B2 => predict_PC_0_5_port, ZN => n2142);
   U1442 : NAND4_X1 port map( A1 => n2139, A2 => n2140, A3 => n2141, A4 => 
                           n2142, ZN => n2138);
   U1441 : NOR2_X1 port map( A1 => n2137, A2 => n2138, ZN => n670);
   U1130 : AOI22_X1 port map( A1 => n2272, A2 => predict_PC_14_28_port, B1 => 
                           n761, B2 => predict_PC_15_28_port, ZN => n1324);
   U1129 : AOI22_X1 port map( A1 => n2270, A2 => predict_PC_12_28_port, B1 => 
                           n2269, B2 => predict_PC_13_28_port, ZN => n1325);
   U1128 : AOI22_X1 port map( A1 => n2276, A2 => predict_PC_8_28_port, B1 => 
                           n2275, B2 => predict_PC_9_28_port, ZN => n1326);
   U1127 : AOI22_X1 port map( A1 => n2274, A2 => predict_PC_10_28_port, B1 => 
                           n2273, B2 => predict_PC_11_28_port, ZN => n1327);
   U1126 : NAND4_X1 port map( A1 => n1324, A2 => n1325, A3 => n1326, A4 => 
                           n1327, ZN => n1318);
   U1125 : AOI22_X1 port map( A1 => n2280, A2 => predict_PC_6_28_port, B1 => 
                           n2279, B2 => predict_PC_7_28_port, ZN => n1320);
   U1124 : AOI22_X1 port map( A1 => n2278, A2 => predict_PC_4_28_port, B1 => 
                           n2277, B2 => predict_PC_5_28_port, ZN => n1321);
   U1123 : AOI22_X1 port map( A1 => n2284, A2 => predict_PC_3_28_port, B1 => 
                           n2283, B2 => predict_PC_2_28_port, ZN => n1322);
   U1122 : AOI22_X1 port map( A1 => n2282, A2 => predict_PC_1_28_port, B1 => 
                           n2281, B2 => predict_PC_0_28_port, ZN => n1323);
   U1121 : NAND4_X1 port map( A1 => n1320, A2 => n1321, A3 => n1322, A4 => 
                           n1323, ZN => n1319);
   U1546 : AOI22_X1 port map( A1 => n2272, A2 => predict_PC_14_0_port, B1 => 
                           n2271, B2 => predict_PC_15_0_port, ZN => n2204);
   U1540 : AOI22_X1 port map( A1 => n2270, A2 => predict_PC_12_0_port, B1 => 
                           n2269, B2 => predict_PC_13_0_port, ZN => n2205);
   U1535 : AOI22_X1 port map( A1 => n2276, A2 => predict_PC_8_0_port, B1 => 
                           n2275, B2 => predict_PC_9_0_port, ZN => n2206);
   U1532 : AOI22_X1 port map( A1 => n2274, A2 => predict_PC_10_0_port, B1 => 
                           n2273, B2 => predict_PC_11_0_port, ZN => n2207);
   U1531 : NAND4_X1 port map( A1 => n2204, A2 => n2205, A3 => n2206, A4 => 
                           n2207, ZN => n2192);
   U1526 : AOI22_X1 port map( A1 => n2280, A2 => predict_PC_6_0_port, B1 => 
                           n2279, B2 => predict_PC_7_0_port, ZN => n2194);
   U1523 : AOI22_X1 port map( A1 => n2278, A2 => predict_PC_4_0_port, B1 => 
                           n2277, B2 => predict_PC_5_0_port, ZN => n2195);
   U1519 : AOI22_X1 port map( A1 => n2284, A2 => predict_PC_3_0_port, B1 => 
                           n2283, B2 => predict_PC_2_0_port, ZN => n2196);
   U1516 : AOI22_X1 port map( A1 => n2282, A2 => predict_PC_1_0_port, B1 => 
                           n2281, B2 => predict_PC_0_0_port, ZN => n2197);
   U1515 : NAND4_X1 port map( A1 => n2194, A2 => n2195, A3 => n2196, A4 => 
                           n2197, ZN => n2193);
   U1514 : NOR2_X1 port map( A1 => n2192, A2 => n2193, ZN => n693);
   U1507 : AOI22_X1 port map( A1 => n2272, A2 => predict_PC_14_1_port, B1 => 
                           n2271, B2 => predict_PC_15_1_port, ZN => n2187);
   U1506 : AOI22_X1 port map( A1 => n2270, A2 => predict_PC_12_1_port, B1 => 
                           n2269, B2 => predict_PC_13_1_port, ZN => n2188);
   U1505 : AOI22_X1 port map( A1 => n2276, A2 => predict_PC_8_1_port, B1 => 
                           n2275, B2 => predict_PC_9_1_port, ZN => n2189);
   U1504 : AOI22_X1 port map( A1 => n2274, A2 => predict_PC_10_1_port, B1 => 
                           n2273, B2 => predict_PC_11_1_port, ZN => n2190);
   U1503 : NAND4_X1 port map( A1 => n2187, A2 => n2188, A3 => n2189, A4 => 
                           n2190, ZN => n2181);
   U1502 : AOI22_X1 port map( A1 => n2280, A2 => predict_PC_6_1_port, B1 => 
                           n2279, B2 => predict_PC_7_1_port, ZN => n2183);
   U1501 : AOI22_X1 port map( A1 => n2278, A2 => predict_PC_4_1_port, B1 => 
                           n2277, B2 => predict_PC_5_1_port, ZN => n2184);
   U1500 : AOI22_X1 port map( A1 => n2284, A2 => predict_PC_3_1_port, B1 => 
                           n2283, B2 => predict_PC_2_1_port, ZN => n2185);
   U1499 : AOI22_X1 port map( A1 => n2282, A2 => predict_PC_1_1_port, B1 => 
                           n2281, B2 => predict_PC_0_1_port, ZN => n2186);
   U1498 : NAND4_X1 port map( A1 => n2183, A2 => n2184, A3 => n2185, A4 => 
                           n2186, ZN => n2182);
   U1497 : NOR2_X1 port map( A1 => n2181, A2 => n2182, ZN => n682);
   U1104 : AOI22_X1 port map( A1 => n2272, A2 => predict_PC_14_30_port, B1 => 
                           n761, B2 => predict_PC_15_30_port, ZN => n1302);
   U1103 : AOI22_X1 port map( A1 => n2270, A2 => predict_PC_12_30_port, B1 => 
                           n2269, B2 => predict_PC_13_30_port, ZN => n1303);
   U1102 : AOI22_X1 port map( A1 => n2276, A2 => predict_PC_8_30_port, B1 => 
                           n2275, B2 => predict_PC_9_30_port, ZN => n1304);
   U1101 : AOI22_X1 port map( A1 => n2274, A2 => predict_PC_10_30_port, B1 => 
                           n2273, B2 => predict_PC_11_30_port, ZN => n1305);
   U1100 : NAND4_X1 port map( A1 => n1302, A2 => n1303, A3 => n1304, A4 => 
                           n1305, ZN => n1296);
   U1099 : AOI22_X1 port map( A1 => n2280, A2 => predict_PC_6_30_port, B1 => 
                           n2279, B2 => predict_PC_7_30_port, ZN => n1298);
   U1098 : AOI22_X1 port map( A1 => n2278, A2 => predict_PC_4_30_port, B1 => 
                           n2277, B2 => predict_PC_5_30_port, ZN => n1299);
   U1097 : AOI22_X1 port map( A1 => n2284, A2 => predict_PC_3_30_port, B1 => 
                           n2283, B2 => predict_PC_2_30_port, ZN => n1300);
   U1096 : AOI22_X1 port map( A1 => n2282, A2 => predict_PC_1_30_port, B1 => 
                           n2281, B2 => predict_PC_0_30_port, ZN => n1301);
   U1095 : NAND4_X1 port map( A1 => n1298, A2 => n1299, A3 => n1300, A4 => 
                           n1301, ZN => n1297);
   U1339 : AOI22_X1 port map( A1 => n2272, A2 => predict_PC_14_13_port, B1 => 
                           n2271, B2 => predict_PC_15_13_port, ZN => n1489);
   U1338 : AOI22_X1 port map( A1 => n2270, A2 => predict_PC_12_13_port, B1 => 
                           n2269, B2 => predict_PC_13_13_port, ZN => n1490);
   U1337 : AOI22_X1 port map( A1 => n2276, A2 => predict_PC_8_13_port, B1 => 
                           n2275, B2 => predict_PC_9_13_port, ZN => n1491);
   U1336 : AOI22_X1 port map( A1 => n2274, A2 => predict_PC_10_13_port, B1 => 
                           n2273, B2 => predict_PC_11_13_port, ZN => n1492);
   U1335 : NAND4_X1 port map( A1 => n1489, A2 => n1490, A3 => n1491, A4 => 
                           n1492, ZN => n1483);
   U1334 : AOI22_X1 port map( A1 => n2280, A2 => predict_PC_6_13_port, B1 => 
                           n2279, B2 => predict_PC_7_13_port, ZN => n1485);
   U1333 : AOI22_X1 port map( A1 => n2278, A2 => predict_PC_4_13_port, B1 => 
                           n2277, B2 => predict_PC_5_13_port, ZN => n1486);
   U1332 : AOI22_X1 port map( A1 => n2284, A2 => predict_PC_3_13_port, B1 => 
                           n2283, B2 => predict_PC_2_13_port, ZN => n1487);
   U1331 : AOI22_X1 port map( A1 => n2282, A2 => predict_PC_1_13_port, B1 => 
                           n2281, B2 => predict_PC_0_13_port, ZN => n1488);
   U1330 : NAND4_X1 port map( A1 => n1485, A2 => n1486, A3 => n1487, A4 => 
                           n1488, ZN => n1484);
   U1329 : NOR2_X1 port map( A1 => n1483, A2 => n1484, ZN => n689);
   U1353 : AOI22_X1 port map( A1 => n2272, A2 => predict_PC_14_12_port, B1 => 
                           n2271, B2 => predict_PC_15_12_port, ZN => n1500);
   U1352 : AOI22_X1 port map( A1 => n2270, A2 => predict_PC_12_12_port, B1 => 
                           n2269, B2 => predict_PC_13_12_port, ZN => n1501);
   U1351 : AOI22_X1 port map( A1 => n2276, A2 => predict_PC_8_12_port, B1 => 
                           n2275, B2 => predict_PC_9_12_port, ZN => n1502);
   U1350 : AOI22_X1 port map( A1 => n2274, A2 => predict_PC_10_12_port, B1 => 
                           n2273, B2 => predict_PC_11_12_port, ZN => n1503);
   U1349 : NAND4_X1 port map( A1 => n1500, A2 => n1501, A3 => n1502, A4 => 
                           n1503, ZN => n1494);
   U1348 : AOI22_X1 port map( A1 => n2280, A2 => predict_PC_6_12_port, B1 => 
                           n2279, B2 => predict_PC_7_12_port, ZN => n1496);
   U1347 : AOI22_X1 port map( A1 => n2278, A2 => predict_PC_4_12_port, B1 => 
                           n2277, B2 => predict_PC_5_12_port, ZN => n1497);
   U1346 : AOI22_X1 port map( A1 => n2284, A2 => predict_PC_3_12_port, B1 => 
                           n2283, B2 => predict_PC_2_12_port, ZN => n1498);
   U1345 : AOI22_X1 port map( A1 => n2282, A2 => predict_PC_1_12_port, B1 => 
                           n2281, B2 => predict_PC_0_12_port, ZN => n1499);
   U1344 : NAND4_X1 port map( A1 => n1496, A2 => n1497, A3 => n1498, A4 => 
                           n1499, ZN => n1495);
   U1343 : NOR2_X1 port map( A1 => n1494, A2 => n1495, ZN => n690);
   U1553 : AOI22_X1 port map( A1 => stall_i, A2 => n592, B1 => n2210, B2 => 
                           n2285, ZN => n1535);
   U1341 : OAI22_X1 port map( A1 => n1284, A2 => target_PC_i(12), B1 => 
                           predict_PC_15_12_port, B2 => n726, ZN => n1493);
   U1327 : OAI22_X1 port map( A1 => n1284, A2 => n651, B1 => 
                           predict_PC_15_13_port, B2 => n726, ZN => n1482);
   U1243 : OAI22_X1 port map( A1 => n1284, A2 => n645, B1 => 
                           predict_PC_15_19_port, B2 => n726, ZN => n1416);
   U1313 : OAI22_X1 port map( A1 => n1284, A2 => n630, B1 => 
                           predict_PC_15_14_port, B2 => n726, ZN => n1471);
   U1271 : OAI22_X1 port map( A1 => n1284, A2 => n631, B1 => 
                           predict_PC_15_17_port, B2 => n726, ZN => n1438);
   U1215 : OAI22_X1 port map( A1 => n1284, A2 => n642, B1 => 
                           predict_PC_15_21_port, B2 => n726, ZN => n1394);
   U1187 : OAI22_X1 port map( A1 => n1284, A2 => n643, B1 => 
                           predict_PC_15_23_port, B2 => n726, ZN => n1372);
   U1229 : OAI22_X1 port map( A1 => n1284, A2 => target_PC_i(20), B1 => 
                           predict_PC_15_20_port, B2 => n726, ZN => n1405);
   U1285 : OAI22_X1 port map( A1 => n1284, A2 => target_PC_i(16), B1 => 
                           predict_PC_15_16_port, B2 => n726, ZN => n1449);
   U1257 : OAI22_X1 port map( A1 => n1284, A2 => target_PC_i(18), B1 => 
                           predict_PC_15_18_port, B2 => n726, ZN => n1427);
   U1201 : OAI22_X1 port map( A1 => n1284, A2 => n632, B1 => 
                           predict_PC_15_22_port, B2 => n726, ZN => n1383);
   U1299 : OAI22_X1 port map( A1 => n1284, A2 => target_PC_i(15), B1 => 
                           predict_PC_15_15_port, B2 => n726, ZN => n1460);
   U914 : OAI22_X1 port map( A1 => n1184, A2 => n646, B1 => 
                           predict_PC_12_12_port, B2 => n735, ZN => n1203);
   U979 : OAI22_X1 port map( A1 => n1218, A2 => n651, B1 => 
                           predict_PC_13_13_port, B2 => n732, ZN => n1236);
   U1049 : OAI22_X1 port map( A1 => n1251, A2 => n646, B1 => 
                           predict_PC_14_12_port, B2 => n729, ZN => n1270);
   U1047 : OAI22_X1 port map( A1 => n1251, A2 => n651, B1 => 
                           predict_PC_14_13_port, B2 => n729, ZN => n1269);
   U912 : OAI22_X1 port map( A1 => n1184, A2 => n651, B1 => 
                           predict_PC_12_13_port, B2 => n735, ZN => n1202);
   U981 : OAI22_X1 port map( A1 => n1218, A2 => target_PC_i(12), B1 => 
                           predict_PC_13_12_port, B2 => n732, ZN => n1237);
   U973 : OAI22_X1 port map( A1 => n1218, A2 => n637, B1 => 
                           predict_PC_13_16_port, B2 => n732, ZN => n1233);
   U1033 : OAI22_X1 port map( A1 => n1251, A2 => n638, B1 => 
                           predict_PC_14_20_port, B2 => n729, ZN => n1262);
   U961 : OAI22_X1 port map( A1 => n1218, A2 => n632, B1 => 
                           predict_PC_13_22_port, B2 => n732, ZN => n1227);
   U1027 : OAI22_X1 port map( A1 => n1251, A2 => n643, B1 => 
                           predict_PC_14_23_port, B2 => n729, ZN => n1259);
   U1031 : OAI22_X1 port map( A1 => n1251, A2 => n642, B1 => 
                           predict_PC_14_21_port, B2 => n729, ZN => n1261);
   U959 : OAI22_X1 port map( A1 => n1218, A2 => n643, B1 => 
                           predict_PC_13_23_port, B2 => n732, ZN => n1226);
   U1039 : OAI22_X1 port map( A1 => n1251, A2 => n631, B1 => 
                           predict_PC_14_17_port, B2 => n729, ZN => n1265);
   U908 : OAI22_X1 port map( A1 => n1184, A2 => target_PC_i(15), B1 => 
                           predict_PC_12_15_port, B2 => n735, ZN => n1200);
   U906 : OAI22_X1 port map( A1 => n1184, A2 => n637, B1 => 
                           predict_PC_12_16_port, B2 => n735, ZN => n1199);
   U963 : OAI22_X1 port map( A1 => n1218, A2 => n642, B1 => 
                           predict_PC_13_21_port, B2 => n732, ZN => n1228);
   U965 : OAI22_X1 port map( A1 => n1218, A2 => n638, B1 => 
                           predict_PC_13_20_port, B2 => n732, ZN => n1229);
   U898 : OAI22_X1 port map( A1 => n1184, A2 => n638, B1 => 
                           predict_PC_12_20_port, B2 => n735, ZN => n1195);
   U1041 : OAI22_X1 port map( A1 => n1251, A2 => n637, B1 => 
                           predict_PC_14_16_port, B2 => n729, ZN => n1266);
   U975 : OAI22_X1 port map( A1 => n1218, A2 => target_PC_i(15), B1 => 
                           predict_PC_13_15_port, B2 => n732, ZN => n1234);
   U910 : OAI22_X1 port map( A1 => n1184, A2 => n630, B1 => 
                           predict_PC_12_14_port, B2 => n735, ZN => n1201);
   U904 : OAI22_X1 port map( A1 => n1184, A2 => n631, B1 => 
                           predict_PC_12_17_port, B2 => n735, ZN => n1198);
   U1037 : OAI22_X1 port map( A1 => n1251, A2 => target_PC_i(18), B1 => 
                           predict_PC_14_18_port, B2 => n729, ZN => n1264);
   U967 : OAI22_X1 port map( A1 => n1218, A2 => n645, B1 => 
                           predict_PC_13_19_port, B2 => n732, ZN => n1230);
   U892 : OAI22_X1 port map( A1 => n1184, A2 => n643, B1 => 
                           predict_PC_12_23_port, B2 => n735, ZN => n1192);
   U902 : OAI22_X1 port map( A1 => n1184, A2 => target_PC_i(18), B1 => 
                           predict_PC_12_18_port, B2 => n735, ZN => n1197);
   U1045 : OAI22_X1 port map( A1 => n1251, A2 => n630, B1 => 
                           predict_PC_14_14_port, B2 => n729, ZN => n1268);
   U900 : OAI22_X1 port map( A1 => n1184, A2 => n645, B1 => 
                           predict_PC_12_19_port, B2 => n735, ZN => n1196);
   U1035 : OAI22_X1 port map( A1 => n1251, A2 => n645, B1 => 
                           predict_PC_14_19_port, B2 => n729, ZN => n1263);
   U969 : OAI22_X1 port map( A1 => n1218, A2 => target_PC_i(18), B1 => 
                           predict_PC_13_18_port, B2 => n732, ZN => n1231);
   U1043 : OAI22_X1 port map( A1 => n1251, A2 => target_PC_i(15), B1 => 
                           predict_PC_14_15_port, B2 => n729, ZN => n1267);
   U971 : OAI22_X1 port map( A1 => n1218, A2 => n631, B1 => 
                           predict_PC_13_17_port, B2 => n732, ZN => n1232);
   U977 : OAI22_X1 port map( A1 => n1218, A2 => n630, B1 => 
                           predict_PC_13_14_port, B2 => n732, ZN => n1235);
   U1029 : OAI22_X1 port map( A1 => n1251, A2 => n632, B1 => 
                           predict_PC_14_22_port, B2 => n729, ZN => n1260);
   U896 : OAI22_X1 port map( A1 => n1184, A2 => n642, B1 => 
                           predict_PC_12_21_port, B2 => n735, ZN => n1194);
   U894 : OAI22_X1 port map( A1 => n1184, A2 => n632, B1 => 
                           predict_PC_12_22_port, B2 => n735, ZN => n1193);
   U384 : OAI22_X1 port map( A1 => n902, A2 => n646, B1 => predict_PC_4_12_port
                           , B2 => n2255, ZN => n921);
   U382 : OAI22_X1 port map( A1 => n902, A2 => n651, B1 => predict_PC_4_13_port
                           , B2 => n2255, ZN => n920);
   U845 : OAI22_X1 port map( A1 => n1151, A2 => n651, B1 => 
                           predict_PC_11_13_port, B2 => n975, ZN => n1169);
   U847 : OAI22_X1 port map( A1 => n1151, A2 => n646, B1 => 
                           predict_PC_11_12_port, B2 => n975, ZN => n1170);
   U713 : OAI22_X1 port map( A1 => n1085, A2 => target_PC_i(13), B1 => 
                           predict_PC_9_13_port, B2 => n981, ZN => n1103);
   U781 : OAI22_X1 port map( A1 => n1118, A2 => n646, B1 => 
                           predict_PC_10_12_port, B2 => n978, ZN => n1137);
   U649 : OAI22_X1 port map( A1 => n1051, A2 => n646, B1 => 
                           predict_PC_8_12_port, B2 => n984, ZN => n1070);
   U448 : OAI22_X1 port map( A1 => n936, A2 => n651, B1 => predict_PC_5_13_port
                           , B2 => n2216, ZN => n954);
   U514 : OAI22_X1 port map( A1 => n969, A2 => n651, B1 => predict_PC_6_13_port
                           , B2 => n2213, ZN => n1003);
   U779 : OAI22_X1 port map( A1 => n1118, A2 => n651, B1 => 
                           predict_PC_10_13_port, B2 => n978, ZN => n1136);
   U715 : OAI22_X1 port map( A1 => n1085, A2 => n646, B1 => 
                           predict_PC_9_12_port, B2 => n981, ZN => n1104);
   U450 : OAI22_X1 port map( A1 => n936, A2 => target_PC_i(12), B1 => 
                           predict_PC_5_12_port, B2 => n2216, ZN => n955);
   U582 : OAI22_X1 port map( A1 => n1018, A2 => n646, B1 => 
                           predict_PC_7_12_port, B2 => n987, ZN => n1037);
   U516 : OAI22_X1 port map( A1 => n969, A2 => n646, B1 => predict_PC_6_12_port
                           , B2 => n2213, ZN => n1004);
   U580 : OAI22_X1 port map( A1 => n1018, A2 => n651, B1 => 
                           predict_PC_7_13_port, B2 => n987, ZN => n1036);
   U647 : OAI22_X1 port map( A1 => n1051, A2 => n651, B1 => 
                           predict_PC_8_13_port, B2 => n984, ZN => n1069);
   U562 : OAI22_X1 port map( A1 => n1018, A2 => n632, B1 => 
                           predict_PC_7_22_port, B2 => n987, ZN => n1027);
   U366 : OAI22_X1 port map( A1 => n902, A2 => n642, B1 => predict_PC_4_21_port
                           , B2 => n2255, ZN => n912);
   U370 : OAI22_X1 port map( A1 => n902, A2 => n645, B1 => predict_PC_4_19_port
                           , B2 => n2255, ZN => n914);
   U372 : OAI22_X1 port map( A1 => n902, A2 => target_PC_i(18), B1 => 
                           predict_PC_4_18_port, B2 => n2255, ZN => n915);
   U368 : OAI22_X1 port map( A1 => n902, A2 => n638, B1 => predict_PC_4_20_port
                           , B2 => n2255, ZN => n913);
   U374 : OAI22_X1 port map( A1 => n902, A2 => n631, B1 => predict_PC_4_17_port
                           , B2 => n2255, ZN => n916);
   U576 : OAI22_X1 port map( A1 => n1018, A2 => target_PC_i(15), B1 => 
                           predict_PC_7_15_port, B2 => n987, ZN => n1034);
   U578 : OAI22_X1 port map( A1 => n1018, A2 => n630, B1 => 
                           predict_PC_7_14_port, B2 => n987, ZN => n1035);
   U572 : OAI22_X1 port map( A1 => n1018, A2 => n631, B1 => 
                           predict_PC_7_17_port, B2 => n987, ZN => n1032);
   U376 : OAI22_X1 port map( A1 => n902, A2 => n637, B1 => predict_PC_4_16_port
                           , B2 => n2255, ZN => n917);
   U564 : OAI22_X1 port map( A1 => n1018, A2 => n642, B1 => 
                           predict_PC_7_21_port, B2 => n987, ZN => n1028);
   U627 : OAI22_X1 port map( A1 => n1051, A2 => n643, B1 => 
                           predict_PC_8_23_port, B2 => n984, ZN => n1059);
   U629 : OAI22_X1 port map( A1 => n1051, A2 => n632, B1 => 
                           predict_PC_8_22_port, B2 => n984, ZN => n1060);
   U570 : OAI22_X1 port map( A1 => n1018, A2 => target_PC_i(18), B1 => 
                           predict_PC_7_18_port, B2 => n987, ZN => n1031);
   U631 : OAI22_X1 port map( A1 => n1051, A2 => n642, B1 => 
                           predict_PC_8_21_port, B2 => n984, ZN => n1061);
   U633 : OAI22_X1 port map( A1 => n1051, A2 => n638, B1 => 
                           predict_PC_8_20_port, B2 => n984, ZN => n1062);
   U635 : OAI22_X1 port map( A1 => n1051, A2 => n645, B1 => 
                           predict_PC_8_19_port, B2 => n984, ZN => n1063);
   U380 : OAI22_X1 port map( A1 => n902, A2 => n630, B1 => predict_PC_4_14_port
                           , B2 => n2255, ZN => n919);
   U637 : OAI22_X1 port map( A1 => n1051, A2 => target_PC_i(18), B1 => 
                           predict_PC_8_18_port, B2 => n984, ZN => n1064);
   U639 : OAI22_X1 port map( A1 => n1051, A2 => n631, B1 => 
                           predict_PC_8_17_port, B2 => n984, ZN => n1065);
   U641 : OAI22_X1 port map( A1 => n1051, A2 => n637, B1 => 
                           predict_PC_8_16_port, B2 => n984, ZN => n1066);
   U643 : OAI22_X1 port map( A1 => n1051, A2 => target_PC_i(15), B1 => 
                           predict_PC_8_15_port, B2 => n984, ZN => n1067);
   U645 : OAI22_X1 port map( A1 => n1051, A2 => n630, B1 => 
                           predict_PC_8_14_port, B2 => n984, ZN => n1068);
   U378 : OAI22_X1 port map( A1 => n902, A2 => target_PC_i(15), B1 => 
                           predict_PC_4_15_port, B2 => n2255, ZN => n918);
   U364 : OAI22_X1 port map( A1 => n902, A2 => n632, B1 => predict_PC_4_22_port
                           , B2 => n2255, ZN => n911);
   U560 : OAI22_X1 port map( A1 => n1018, A2 => n643, B1 => 
                           predict_PC_7_23_port, B2 => n987, ZN => n1026);
   U362 : OAI22_X1 port map( A1 => n902, A2 => n643, B1 => predict_PC_4_23_port
                           , B2 => n2255, ZN => n910);
   U512 : OAI22_X1 port map( A1 => n969, A2 => n630, B1 => predict_PC_6_14_port
                           , B2 => n2213, ZN => n1002);
   U574 : OAI22_X1 port map( A1 => n1018, A2 => n637, B1 => 
                           predict_PC_7_16_port, B2 => n987, ZN => n1033);
   U510 : OAI22_X1 port map( A1 => n969, A2 => target_PC_i(15), B1 => 
                           predict_PC_6_15_port, B2 => n2213, ZN => n1001);
   U693 : OAI22_X1 port map( A1 => n1085, A2 => n643, B1 => 
                           predict_PC_9_23_port, B2 => n981, ZN => n1093);
   U508 : OAI22_X1 port map( A1 => n969, A2 => n637, B1 => predict_PC_6_16_port
                           , B2 => n2213, ZN => n1000);
   U695 : OAI22_X1 port map( A1 => n1085, A2 => n632, B1 => 
                           predict_PC_9_22_port, B2 => n981, ZN => n1094);
   U506 : OAI22_X1 port map( A1 => n969, A2 => n631, B1 => predict_PC_6_17_port
                           , B2 => n2213, ZN => n999);
   U697 : OAI22_X1 port map( A1 => n1085, A2 => n642, B1 => 
                           predict_PC_9_21_port, B2 => n981, ZN => n1095);
   U504 : OAI22_X1 port map( A1 => n969, A2 => target_PC_i(18), B1 => 
                           predict_PC_6_18_port, B2 => n2213, ZN => n998);
   U699 : OAI22_X1 port map( A1 => n1085, A2 => n638, B1 => 
                           predict_PC_9_20_port, B2 => n981, ZN => n1096);
   U502 : OAI22_X1 port map( A1 => n969, A2 => n645, B1 => predict_PC_6_19_port
                           , B2 => n2213, ZN => n997);
   U701 : OAI22_X1 port map( A1 => n1085, A2 => n645, B1 => 
                           predict_PC_9_19_port, B2 => n981, ZN => n1097);
   U500 : OAI22_X1 port map( A1 => n969, A2 => n638, B1 => predict_PC_6_20_port
                           , B2 => n2213, ZN => n996);
   U703 : OAI22_X1 port map( A1 => n1085, A2 => target_PC_i(18), B1 => 
                           predict_PC_9_18_port, B2 => n981, ZN => n1098);
   U498 : OAI22_X1 port map( A1 => n969, A2 => n642, B1 => predict_PC_6_21_port
                           , B2 => n2213, ZN => n995);
   U446 : OAI22_X1 port map( A1 => n936, A2 => n630, B1 => predict_PC_5_14_port
                           , B2 => n2216, ZN => n953);
   U440 : OAI22_X1 port map( A1 => n936, A2 => n631, B1 => predict_PC_5_17_port
                           , B2 => n2216, ZN => n950);
   U767 : OAI22_X1 port map( A1 => n1118, A2 => n645, B1 => 
                           predict_PC_10_19_port, B2 => n978, ZN => n1130);
   U442 : OAI22_X1 port map( A1 => n936, A2 => n637, B1 => predict_PC_5_16_port
                           , B2 => n2216, ZN => n951);
   U839 : OAI22_X1 port map( A1 => n1151, A2 => n637, B1 => 
                           predict_PC_11_16_port, B2 => n975, ZN => n1166);
   U769 : OAI22_X1 port map( A1 => n1118, A2 => target_PC_i(18), B1 => 
                           predict_PC_10_18_port, B2 => n978, ZN => n1131);
   U432 : OAI22_X1 port map( A1 => n936, A2 => n642, B1 => predict_PC_5_21_port
                           , B2 => n2216, ZN => n946);
   U705 : OAI22_X1 port map( A1 => n1085, A2 => n631, B1 => 
                           predict_PC_9_17_port, B2 => n981, ZN => n1099);
   U833 : OAI22_X1 port map( A1 => n1151, A2 => n645, B1 => 
                           predict_PC_11_19_port, B2 => n975, ZN => n1163);
   U428 : OAI22_X1 port map( A1 => n936, A2 => n643, B1 => predict_PC_5_23_port
                           , B2 => n2216, ZN => n944);
   U496 : OAI22_X1 port map( A1 => n969, A2 => n632, B1 => predict_PC_6_22_port
                           , B2 => n2213, ZN => n994);
   U707 : OAI22_X1 port map( A1 => n1085, A2 => n637, B1 => 
                           predict_PC_9_16_port, B2 => n981, ZN => n1100);
   U494 : OAI22_X1 port map( A1 => n969, A2 => n643, B1 => predict_PC_6_23_port
                           , B2 => n2213, ZN => n993);
   U430 : OAI22_X1 port map( A1 => n936, A2 => target_PC_i(22), B1 => 
                           predict_PC_5_22_port, B2 => n2216, ZN => n945);
   U709 : OAI22_X1 port map( A1 => n1085, A2 => target_PC_i(15), B1 => 
                           predict_PC_9_15_port, B2 => n981, ZN => n1101);
   U711 : OAI22_X1 port map( A1 => n1085, A2 => n630, B1 => 
                           predict_PC_9_14_port, B2 => n981, ZN => n1102);
   U825 : OAI22_X1 port map( A1 => n1151, A2 => n643, B1 => 
                           predict_PC_11_23_port, B2 => n975, ZN => n1159);
   U777 : OAI22_X1 port map( A1 => n1118, A2 => target_PC_i(14), B1 => 
                           predict_PC_10_14_port, B2 => n978, ZN => n1135);
   U566 : OAI22_X1 port map( A1 => n1018, A2 => n638, B1 => 
                           predict_PC_7_20_port, B2 => n987, ZN => n1029);
   U568 : OAI22_X1 port map( A1 => n1018, A2 => n645, B1 => 
                           predict_PC_7_19_port, B2 => n987, ZN => n1030);
   U759 : OAI22_X1 port map( A1 => n1118, A2 => n643, B1 => 
                           predict_PC_10_23_port, B2 => n978, ZN => n1126);
   U761 : OAI22_X1 port map( A1 => n1118, A2 => n632, B1 => 
                           predict_PC_10_22_port, B2 => n978, ZN => n1127);
   U763 : OAI22_X1 port map( A1 => n1118, A2 => n642, B1 => 
                           predict_PC_10_21_port, B2 => n978, ZN => n1128);
   U843 : OAI22_X1 port map( A1 => n1151, A2 => n630, B1 => 
                           predict_PC_11_14_port, B2 => n975, ZN => n1168);
   U765 : OAI22_X1 port map( A1 => n1118, A2 => n638, B1 => 
                           predict_PC_10_20_port, B2 => n978, ZN => n1129);
   U841 : OAI22_X1 port map( A1 => n1151, A2 => target_PC_i(15), B1 => 
                           predict_PC_11_15_port, B2 => n975, ZN => n1167);
   U775 : OAI22_X1 port map( A1 => n1118, A2 => target_PC_i(15), B1 => 
                           predict_PC_10_15_port, B2 => n978, ZN => n1134);
   U438 : OAI22_X1 port map( A1 => n936, A2 => target_PC_i(18), B1 => 
                           predict_PC_5_18_port, B2 => n2216, ZN => n949);
   U827 : OAI22_X1 port map( A1 => n1151, A2 => n632, B1 => 
                           predict_PC_11_22_port, B2 => n975, ZN => n1160);
   U444 : OAI22_X1 port map( A1 => n936, A2 => target_PC_i(15), B1 => 
                           predict_PC_5_15_port, B2 => n2216, ZN => n952);
   U773 : OAI22_X1 port map( A1 => n1118, A2 => target_PC_i(16), B1 => 
                           predict_PC_10_16_port, B2 => n978, ZN => n1133);
   U837 : OAI22_X1 port map( A1 => n1151, A2 => target_PC_i(17), B1 => 
                           predict_PC_11_17_port, B2 => n975, ZN => n1165);
   U771 : OAI22_X1 port map( A1 => n1118, A2 => n631, B1 => 
                           predict_PC_10_17_port, B2 => n978, ZN => n1132);
   U835 : OAI22_X1 port map( A1 => n1151, A2 => target_PC_i(18), B1 => 
                           predict_PC_11_18_port, B2 => n975, ZN => n1164);
   U434 : OAI22_X1 port map( A1 => n936, A2 => n638, B1 => predict_PC_5_20_port
                           , B2 => n2216, ZN => n947);
   U829 : OAI22_X1 port map( A1 => n1151, A2 => n642, B1 => 
                           predict_PC_11_21_port, B2 => n975, ZN => n1161);
   U831 : OAI22_X1 port map( A1 => n1151, A2 => target_PC_i(20), B1 => 
                           predict_PC_11_20_port, B2 => n975, ZN => n1162);
   U436 : OAI22_X1 port map( A1 => n936, A2 => n645, B1 => predict_PC_5_19_port
                           , B2 => n2216, ZN => n948);
   U1355 : OAI22_X1 port map( A1 => n1284, A2 => n644, B1 => 
                           predict_PC_15_11_port, B2 => n725, ZN => n1504);
   U1439 : OAI22_X1 port map( A1 => n1284, A2 => target_PC_i(5), B1 => 
                           predict_PC_15_5_port, B2 => n725, ZN => n2136);
   U1481 : OAI22_X1 port map( A1 => n1284, A2 => target_PC_i(2), B1 => 
                           predict_PC_15_2_port, B2 => n725, ZN => n2169);
   U1495 : OAI22_X1 port map( A1 => n1284, A2 => n633, B1 => 
                           predict_PC_15_1_port, B2 => n725, ZN => n2180);
   U1467 : OAI22_X1 port map( A1 => n1284, A2 => n652, B1 => 
                           predict_PC_15_3_port, B2 => n725, ZN => n2158);
   U1425 : OAI22_X1 port map( A1 => n1284, A2 => target_PC_i(6), B1 => 
                           predict_PC_15_6_port, B2 => n725, ZN => n2125);
   U1453 : OAI22_X1 port map( A1 => n1284, A2 => n641, B1 => 
                           predict_PC_15_4_port, B2 => n725, ZN => n2147);
   U1397 : OAI22_X1 port map( A1 => n1284, A2 => n639, B1 => 
                           predict_PC_15_8_port, B2 => n725, ZN => n2103);
   U1369 : OAI22_X1 port map( A1 => n1284, A2 => n640, B1 => 
                           predict_PC_15_10_port, B2 => n725, ZN => n1515);
   U118 : OAI22_X1 port map( A1 => n765, A2 => target_PC_i(13), B1 => 
                           predict_PC_0_13_port, B2 => n2267, ZN => n783);
   U186 : OAI22_X1 port map( A1 => n800, A2 => n646, B1 => predict_PC_1_12_port
                           , B2 => n2264, ZN => n819);
   U250 : OAI22_X1 port map( A1 => n834, A2 => n651, B1 => predict_PC_2_13_port
                           , B2 => n2261, ZN => n852);
   U316 : OAI22_X1 port map( A1 => n868, A2 => n651, B1 => predict_PC_3_13_port
                           , B2 => n2258, ZN => n886);
   U318 : OAI22_X1 port map( A1 => n868, A2 => n646, B1 => predict_PC_3_12_port
                           , B2 => n2258, ZN => n887);
   U184 : OAI22_X1 port map( A1 => n800, A2 => target_PC_i(13), B1 => 
                           predict_PC_1_13_port, B2 => n2264, ZN => n818);
   U252 : OAI22_X1 port map( A1 => n834, A2 => n646, B1 => predict_PC_2_12_port
                           , B2 => n2261, ZN => n853);
   U120 : OAI22_X1 port map( A1 => n765, A2 => n646, B1 => predict_PC_0_12_port
                           , B2 => n2267, ZN => n784);
   U302 : OAI22_X1 port map( A1 => n868, A2 => n638, B1 => predict_PC_3_20_port
                           , B2 => n2258, ZN => n879);
   U238 : OAI22_X1 port map( A1 => n834, A2 => n645, B1 => predict_PC_2_19_port
                           , B2 => n2261, ZN => n846);
   U102 : OAI22_X1 port map( A1 => n765, A2 => n642, B1 => predict_PC_0_21_port
                           , B2 => n2267, ZN => n775);
   U240 : OAI22_X1 port map( A1 => n834, A2 => target_PC_i(18), B1 => 
                           predict_PC_2_18_port, B2 => n2261, ZN => n847);
   U242 : OAI22_X1 port map( A1 => n834, A2 => n631, B1 => predict_PC_2_17_port
                           , B2 => n2261, ZN => n848);
   U244 : OAI22_X1 port map( A1 => n834, A2 => n637, B1 => predict_PC_2_16_port
                           , B2 => n2261, ZN => n849);
   U100 : OAI22_X1 port map( A1 => n765, A2 => n632, B1 => predict_PC_0_22_port
                           , B2 => n2267, ZN => n774);
   U246 : OAI22_X1 port map( A1 => n834, A2 => target_PC_i(15), B1 => 
                           predict_PC_2_15_port, B2 => n2261, ZN => n850);
   U104 : OAI22_X1 port map( A1 => n765, A2 => target_PC_i(20), B1 => 
                           predict_PC_0_20_port, B2 => n2267, ZN => n776);
   U98 : OAI22_X1 port map( A1 => n765, A2 => n643, B1 => predict_PC_0_23_port,
                           B2 => n2267, ZN => n773);
   U248 : OAI22_X1 port map( A1 => n834, A2 => n630, B1 => predict_PC_2_14_port
                           , B2 => n2261, ZN => n851);
   U236 : OAI22_X1 port map( A1 => n834, A2 => n638, B1 => predict_PC_2_20_port
                           , B2 => n2261, ZN => n845);
   U234 : OAI22_X1 port map( A1 => n834, A2 => n642, B1 => predict_PC_2_21_port
                           , B2 => n2261, ZN => n844);
   U232 : OAI22_X1 port map( A1 => n834, A2 => n632, B1 => predict_PC_2_22_port
                           , B2 => n2261, ZN => n843);
   U230 : OAI22_X1 port map( A1 => n834, A2 => n643, B1 => predict_PC_2_23_port
                           , B2 => n2261, ZN => n842);
   U106 : OAI22_X1 port map( A1 => n765, A2 => n645, B1 => predict_PC_0_19_port
                           , B2 => n2267, ZN => n777);
   U108 : OAI22_X1 port map( A1 => n765, A2 => target_PC_i(18), B1 => 
                           predict_PC_0_18_port, B2 => n2267, ZN => n778);
   U110 : OAI22_X1 port map( A1 => n765, A2 => n631, B1 => predict_PC_0_17_port
                           , B2 => n2267, ZN => n779);
   U112 : OAI22_X1 port map( A1 => n765, A2 => target_PC_i(16), B1 => 
                           predict_PC_0_16_port, B2 => n2267, ZN => n780);
   U114 : OAI22_X1 port map( A1 => n765, A2 => target_PC_i(15), B1 => 
                           predict_PC_0_15_port, B2 => n2267, ZN => n781);
   U170 : OAI22_X1 port map( A1 => n800, A2 => n638, B1 => predict_PC_1_20_port
                           , B2 => n2264, ZN => n811);
   U116 : OAI22_X1 port map( A1 => n765, A2 => n630, B1 => predict_PC_0_14_port
                           , B2 => n2267, ZN => n782);
   U182 : OAI22_X1 port map( A1 => n800, A2 => n630, B1 => predict_PC_1_14_port
                           , B2 => n2264, ZN => n817);
   U178 : OAI22_X1 port map( A1 => n800, A2 => n637, B1 => predict_PC_1_16_port
                           , B2 => n2264, ZN => n815);
   U180 : OAI22_X1 port map( A1 => n800, A2 => target_PC_i(15), B1 => 
                           predict_PC_1_15_port, B2 => n2264, ZN => n816);
   U164 : OAI22_X1 port map( A1 => n800, A2 => n643, B1 => predict_PC_1_23_port
                           , B2 => n2264, ZN => n808);
   U166 : OAI22_X1 port map( A1 => n800, A2 => n632, B1 => predict_PC_1_22_port
                           , B2 => n2264, ZN => n809);
   U304 : OAI22_X1 port map( A1 => n868, A2 => n645, B1 => predict_PC_3_19_port
                           , B2 => n2258, ZN => n880);
   U168 : OAI22_X1 port map( A1 => n800, A2 => n642, B1 => predict_PC_1_21_port
                           , B2 => n2264, ZN => n810);
   U312 : OAI22_X1 port map( A1 => n868, A2 => target_PC_i(15), B1 => 
                           predict_PC_3_15_port, B2 => n2258, ZN => n884);
   U174 : OAI22_X1 port map( A1 => n800, A2 => target_PC_i(18), B1 => 
                           predict_PC_1_18_port, B2 => n2264, ZN => n813);
   U314 : OAI22_X1 port map( A1 => n868, A2 => n630, B1 => predict_PC_3_14_port
                           , B2 => n2258, ZN => n885);
   U306 : OAI22_X1 port map( A1 => n868, A2 => target_PC_i(18), B1 => 
                           predict_PC_3_18_port, B2 => n2258, ZN => n881);
   U296 : OAI22_X1 port map( A1 => n868, A2 => n643, B1 => predict_PC_3_23_port
                           , B2 => n2258, ZN => n876);
   U310 : OAI22_X1 port map( A1 => n868, A2 => n637, B1 => predict_PC_3_16_port
                           , B2 => n2258, ZN => n883);
   U308 : OAI22_X1 port map( A1 => n868, A2 => n631, B1 => predict_PC_3_17_port
                           , B2 => n2258, ZN => n882);
   U298 : OAI22_X1 port map( A1 => n868, A2 => n632, B1 => predict_PC_3_22_port
                           , B2 => n2258, ZN => n877);
   U172 : OAI22_X1 port map( A1 => n800, A2 => n645, B1 => predict_PC_1_19_port
                           , B2 => n2264, ZN => n812);
   U176 : OAI22_X1 port map( A1 => n800, A2 => n631, B1 => predict_PC_1_17_port
                           , B2 => n2264, ZN => n814);
   U300 : OAI22_X1 port map( A1 => n868, A2 => n642, B1 => predict_PC_3_21_port
                           , B2 => n2258, ZN => n878);
   U1071 : OAI22_X1 port map( A1 => n1251, A2 => n633, B1 => 
                           predict_PC_14_1_port, B2 => n728, ZN => n1281);
   U995 : OAI22_X1 port map( A1 => n1218, A2 => target_PC_i(5), B1 => 
                           predict_PC_13_5_port, B2 => n731, ZN => n1244);
   U993 : OAI22_X1 port map( A1 => n1218, A2 => target_PC_i(6), B1 => 
                           predict_PC_13_6_port, B2 => n731, ZN => n1243);
   U989 : OAI22_X1 port map( A1 => n1218, A2 => n639, B1 => 
                           predict_PC_13_8_port, B2 => n731, ZN => n1241);
   U985 : OAI22_X1 port map( A1 => n1218, A2 => n640, B1 => 
                           predict_PC_13_10_port, B2 => n731, ZN => n1239);
   U1001 : OAI22_X1 port map( A1 => n1218, A2 => target_PC_i(2), B1 => 
                           predict_PC_13_2_port, B2 => n731, ZN => n1247);
   U983 : OAI22_X1 port map( A1 => n1218, A2 => n644, B1 => 
                           predict_PC_13_11_port, B2 => n731, ZN => n1238);
   U999 : OAI22_X1 port map( A1 => n1218, A2 => n652, B1 => 
                           predict_PC_13_3_port, B2 => n731, ZN => n1246);
   U997 : OAI22_X1 port map( A1 => n1218, A2 => n641, B1 => 
                           predict_PC_13_4_port, B2 => n731, ZN => n1245);
   U1057 : OAI22_X1 port map( A1 => n1251, A2 => n639, B1 => 
                           predict_PC_14_8_port, B2 => n728, ZN => n1274);
   U1003 : OAI22_X1 port map( A1 => n1218, A2 => n633, B1 => 
                           predict_PC_13_1_port, B2 => n731, ZN => n1248);
   U932 : OAI22_X1 port map( A1 => n1184, A2 => n652, B1 => 
                           predict_PC_12_3_port, B2 => n734, ZN => n1212);
   U930 : OAI22_X1 port map( A1 => n1184, A2 => n641, B1 => 
                           predict_PC_12_4_port, B2 => n734, ZN => n1211);
   U1061 : OAI22_X1 port map( A1 => n1251, A2 => target_PC_i(6), B1 => 
                           predict_PC_14_6_port, B2 => n728, ZN => n1276);
   U926 : OAI22_X1 port map( A1 => n1184, A2 => target_PC_i(6), B1 => 
                           predict_PC_12_6_port, B2 => n734, ZN => n1209);
   U918 : OAI22_X1 port map( A1 => n1184, A2 => n640, B1 => 
                           predict_PC_12_10_port, B2 => n734, ZN => n1205);
   U1051 : OAI22_X1 port map( A1 => n1251, A2 => n644, B1 => 
                           predict_PC_14_11_port, B2 => n728, ZN => n1271);
   U922 : OAI22_X1 port map( A1 => n1184, A2 => n639, B1 => 
                           predict_PC_12_8_port, B2 => n734, ZN => n1207);
   U1069 : OAI22_X1 port map( A1 => n1251, A2 => n650, B1 => 
                           predict_PC_14_2_port, B2 => n728, ZN => n1280);
   U928 : OAI22_X1 port map( A1 => n1184, A2 => target_PC_i(5), B1 => 
                           predict_PC_12_5_port, B2 => n734, ZN => n1210);
   U1067 : OAI22_X1 port map( A1 => n1251, A2 => n652, B1 => 
                           predict_PC_14_3_port, B2 => n728, ZN => n1279);
   U934 : OAI22_X1 port map( A1 => n1184, A2 => target_PC_i(2), B1 => 
                           predict_PC_12_2_port, B2 => n734, ZN => n1213);
   U936 : OAI22_X1 port map( A1 => n1184, A2 => n633, B1 => 
                           predict_PC_12_1_port, B2 => n734, ZN => n1214);
   U1065 : OAI22_X1 port map( A1 => n1251, A2 => n641, B1 => 
                           predict_PC_14_4_port, B2 => n728, ZN => n1278);
   U916 : OAI22_X1 port map( A1 => n1184, A2 => n644, B1 => 
                           predict_PC_12_11_port, B2 => n734, ZN => n1204);
   U1053 : OAI22_X1 port map( A1 => n1251, A2 => n640, B1 => 
                           predict_PC_14_10_port, B2 => n728, ZN => n1272);
   U1063 : OAI22_X1 port map( A1 => n1251, A2 => target_PC_i(5), B1 => 
                           predict_PC_14_5_port, B2 => n728, ZN => n1277);
   U663 : OAI22_X1 port map( A1 => n1051, A2 => target_PC_i(5), B1 => 
                           predict_PC_8_5_port, B2 => n983, ZN => n1077);
   U534 : OAI22_X1 port map( A1 => n969, A2 => n652, B1 => predict_PC_6_3_port,
                           B2 => n989, ZN => n1013);
   U520 : OAI22_X1 port map( A1 => n969, A2 => n640, B1 => predict_PC_6_10_port
                           , B2 => n989, ZN => n1006);
   U530 : OAI22_X1 port map( A1 => n969, A2 => target_PC_i(5), B1 => 
                           predict_PC_6_5_port, B2 => n989, ZN => n1011);
   U604 : OAI22_X1 port map( A1 => n1018, A2 => n633, B1 => predict_PC_7_1_port
                           , B2 => n986, ZN => n1048);
   U518 : OAI22_X1 port map( A1 => n969, A2 => n644, B1 => predict_PC_6_11_port
                           , B2 => n989, ZN => n1005);
   U532 : OAI22_X1 port map( A1 => n969, A2 => n641, B1 => predict_PC_6_4_port,
                           B2 => n989, ZN => n1012);
   U524 : OAI22_X1 port map( A1 => n969, A2 => n639, B1 => predict_PC_6_8_port,
                           B2 => n989, ZN => n1008);
   U653 : OAI22_X1 port map( A1 => n1051, A2 => n640, B1 => 
                           predict_PC_8_10_port, B2 => n983, ZN => n1072);
   U528 : OAI22_X1 port map( A1 => n969, A2 => target_PC_i(6), B1 => 
                           predict_PC_6_6_port, B2 => n989, ZN => n1010);
   U651 : OAI22_X1 port map( A1 => n1051, A2 => n644, B1 => 
                           predict_PC_8_11_port, B2 => n983, ZN => n1071);
   U657 : OAI22_X1 port map( A1 => n1051, A2 => n639, B1 => predict_PC_8_8_port
                           , B2 => n983, ZN => n1074);
   U669 : OAI22_X1 port map( A1 => n1051, A2 => n650, B1 => predict_PC_8_2_port
                           , B2 => n983, ZN => n1080);
   U661 : OAI22_X1 port map( A1 => n1051, A2 => target_PC_i(6), B1 => 
                           predict_PC_8_6_port, B2 => n983, ZN => n1076);
   U590 : OAI22_X1 port map( A1 => n1018, A2 => n639, B1 => predict_PC_7_8_port
                           , B2 => n986, ZN => n1041);
   U586 : OAI22_X1 port map( A1 => n1018, A2 => target_PC_i(10), B1 => 
                           predict_PC_7_10_port, B2 => n986, ZN => n1039);
   U602 : OAI22_X1 port map( A1 => n1018, A2 => target_PC_i(2), B1 => 
                           predict_PC_7_2_port, B2 => n986, ZN => n1047);
   U719 : OAI22_X1 port map( A1 => n1085, A2 => n640, B1 => 
                           predict_PC_9_10_port, B2 => n980, ZN => n1106);
   U723 : OAI22_X1 port map( A1 => n1085, A2 => n639, B1 => predict_PC_9_8_port
                           , B2 => n980, ZN => n1108);
   U584 : OAI22_X1 port map( A1 => n1018, A2 => n644, B1 => 
                           predict_PC_7_11_port, B2 => n986, ZN => n1038);
   U665 : OAI22_X1 port map( A1 => n1051, A2 => n641, B1 => predict_PC_8_4_port
                           , B2 => n983, ZN => n1078);
   U727 : OAI22_X1 port map( A1 => n1085, A2 => target_PC_i(6), B1 => 
                           predict_PC_9_6_port, B2 => n980, ZN => n1110);
   U594 : OAI22_X1 port map( A1 => n1018, A2 => target_PC_i(6), B1 => 
                           predict_PC_7_6_port, B2 => n986, ZN => n1043);
   U667 : OAI22_X1 port map( A1 => n1051, A2 => n652, B1 => predict_PC_8_3_port
                           , B2 => n983, ZN => n1079);
   U538 : OAI22_X1 port map( A1 => n969, A2 => n633, B1 => predict_PC_6_1_port,
                           B2 => n989, ZN => n1015);
   U729 : OAI22_X1 port map( A1 => n1085, A2 => target_PC_i(5), B1 => 
                           predict_PC_9_5_port, B2 => n980, ZN => n1111);
   U717 : OAI22_X1 port map( A1 => n1085, A2 => n644, B1 => 
                           predict_PC_9_11_port, B2 => n980, ZN => n1105);
   U731 : OAI22_X1 port map( A1 => n1085, A2 => target_PC_i(4), B1 => 
                           predict_PC_9_4_port, B2 => n980, ZN => n1112);
   U671 : OAI22_X1 port map( A1 => n1051, A2 => n633, B1 => predict_PC_8_1_port
                           , B2 => n983, ZN => n1081);
   U733 : OAI22_X1 port map( A1 => n1085, A2 => target_PC_i(3), B1 => 
                           predict_PC_9_3_port, B2 => n980, ZN => n1113);
   U600 : OAI22_X1 port map( A1 => n1018, A2 => n652, B1 => predict_PC_7_3_port
                           , B2 => n986, ZN => n1046);
   U598 : OAI22_X1 port map( A1 => n1018, A2 => n641, B1 => predict_PC_7_4_port
                           , B2 => n986, ZN => n1045);
   U536 : OAI22_X1 port map( A1 => n969, A2 => n650, B1 => predict_PC_6_2_port,
                           B2 => n989, ZN => n1014);
   U596 : OAI22_X1 port map( A1 => n1018, A2 => target_PC_i(5), B1 => 
                           predict_PC_7_5_port, B2 => n986, ZN => n1044);
   U398 : OAI22_X1 port map( A1 => n902, A2 => target_PC_i(5), B1 => 
                           predict_PC_4_5_port, B2 => n2254, ZN => n928);
   U735 : OAI22_X1 port map( A1 => n1085, A2 => n650, B1 => predict_PC_9_2_port
                           , B2 => n980, ZN => n1114);
   U737 : OAI22_X1 port map( A1 => n1085, A2 => n633, B1 => predict_PC_9_1_port
                           , B2 => n980, ZN => n1115);
   U472 : OAI22_X1 port map( A1 => n936, A2 => n633, B1 => predict_PC_5_1_port,
                           B2 => n2215, ZN => n966);
   U470 : OAI22_X1 port map( A1 => n936, A2 => n650, B1 => predict_PC_5_2_port,
                           B2 => n2215, ZN => n965);
   U468 : OAI22_X1 port map( A1 => n936, A2 => n652, B1 => predict_PC_5_3_port,
                           B2 => n2215, ZN => n964);
   U466 : OAI22_X1 port map( A1 => n936, A2 => n641, B1 => predict_PC_5_4_port,
                           B2 => n2215, ZN => n963);
   U464 : OAI22_X1 port map( A1 => n936, A2 => target_PC_i(5), B1 => 
                           predict_PC_5_5_port, B2 => n2215, ZN => n962);
   U462 : OAI22_X1 port map( A1 => n936, A2 => target_PC_i(6), B1 => 
                           predict_PC_5_6_port, B2 => n2215, ZN => n961);
   U849 : OAI22_X1 port map( A1 => n1151, A2 => n644, B1 => 
                           predict_PC_11_11_port, B2 => n974, ZN => n1171);
   U851 : OAI22_X1 port map( A1 => n1151, A2 => n640, B1 => 
                           predict_PC_11_10_port, B2 => n974, ZN => n1172);
   U855 : OAI22_X1 port map( A1 => n1151, A2 => n639, B1 => 
                           predict_PC_11_8_port, B2 => n974, ZN => n1174);
   U458 : OAI22_X1 port map( A1 => n936, A2 => n639, B1 => predict_PC_5_8_port,
                           B2 => n2215, ZN => n959);
   U783 : OAI22_X1 port map( A1 => n1118, A2 => n644, B1 => 
                           predict_PC_10_11_port, B2 => n977, ZN => n1138);
   U785 : OAI22_X1 port map( A1 => n1118, A2 => n640, B1 => 
                           predict_PC_10_10_port, B2 => n977, ZN => n1139);
   U789 : OAI22_X1 port map( A1 => n1118, A2 => n639, B1 => 
                           predict_PC_10_8_port, B2 => n977, ZN => n1141);
   U454 : OAI22_X1 port map( A1 => n936, A2 => n640, B1 => predict_PC_5_10_port
                           , B2 => n2215, ZN => n957);
   U793 : OAI22_X1 port map( A1 => n1118, A2 => target_PC_i(6), B1 => 
                           predict_PC_10_6_port, B2 => n977, ZN => n1143);
   U452 : OAI22_X1 port map( A1 => n936, A2 => n644, B1 => predict_PC_5_11_port
                           , B2 => n2215, ZN => n956);
   U795 : OAI22_X1 port map( A1 => n1118, A2 => target_PC_i(5), B1 => 
                           predict_PC_10_5_port, B2 => n977, ZN => n1144);
   U803 : OAI22_X1 port map( A1 => n1118, A2 => n633, B1 => 
                           predict_PC_10_1_port, B2 => n977, ZN => n1148);
   U402 : OAI22_X1 port map( A1 => n902, A2 => n652, B1 => predict_PC_4_3_port,
                           B2 => n2254, ZN => n930);
   U406 : OAI22_X1 port map( A1 => n902, A2 => target_PC_i(1), B1 => 
                           predict_PC_4_1_port, B2 => n2254, ZN => n932);
   U400 : OAI22_X1 port map( A1 => n902, A2 => n641, B1 => predict_PC_4_4_port,
                           B2 => n2254, ZN => n929);
   U869 : OAI22_X1 port map( A1 => n1151, A2 => n633, B1 => 
                           predict_PC_11_1_port, B2 => n974, ZN => n1181);
   U797 : OAI22_X1 port map( A1 => n1118, A2 => target_PC_i(4), B1 => 
                           predict_PC_10_4_port, B2 => n977, ZN => n1145);
   U859 : OAI22_X1 port map( A1 => n1151, A2 => target_PC_i(6), B1 => 
                           predict_PC_11_6_port, B2 => n974, ZN => n1176);
   U799 : OAI22_X1 port map( A1 => n1118, A2 => n652, B1 => 
                           predict_PC_10_3_port, B2 => n977, ZN => n1146);
   U801 : OAI22_X1 port map( A1 => n1118, A2 => target_PC_i(2), B1 => 
                           predict_PC_10_2_port, B2 => n977, ZN => n1147);
   U396 : OAI22_X1 port map( A1 => n902, A2 => target_PC_i(6), B1 => 
                           predict_PC_4_6_port, B2 => n2254, ZN => n927);
   U867 : OAI22_X1 port map( A1 => n1151, A2 => n650, B1 => 
                           predict_PC_11_2_port, B2 => n974, ZN => n1180);
   U863 : OAI22_X1 port map( A1 => n1151, A2 => n641, B1 => 
                           predict_PC_11_4_port, B2 => n974, ZN => n1178);
   U865 : OAI22_X1 port map( A1 => n1151, A2 => n652, B1 => 
                           predict_PC_11_3_port, B2 => n974, ZN => n1179);
   U404 : OAI22_X1 port map( A1 => n902, A2 => n650, B1 => predict_PC_4_2_port,
                           B2 => n2254, ZN => n931);
   U388 : OAI22_X1 port map( A1 => n902, A2 => n640, B1 => predict_PC_4_10_port
                           , B2 => n2254, ZN => n923);
   U392 : OAI22_X1 port map( A1 => n902, A2 => n639, B1 => predict_PC_4_8_port,
                           B2 => n2254, ZN => n925);
   U386 : OAI22_X1 port map( A1 => n902, A2 => n644, B1 => predict_PC_4_11_port
                           , B2 => n2254, ZN => n922);
   U861 : OAI22_X1 port map( A1 => n1151, A2 => target_PC_i(5), B1 => 
                           predict_PC_11_5_port, B2 => n974, ZN => n1177);
   U200 : OAI22_X1 port map( A1 => n800, A2 => target_PC_i(5), B1 => 
                           predict_PC_1_5_port, B2 => n2263, ZN => n826);
   U198 : OAI22_X1 port map( A1 => n800, A2 => target_PC_i(6), B1 => 
                           predict_PC_1_6_port, B2 => n2263, ZN => n825);
   U194 : OAI22_X1 port map( A1 => n800, A2 => n639, B1 => predict_PC_1_8_port,
                           B2 => n2263, ZN => n823);
   U138 : OAI22_X1 port map( A1 => n765, A2 => target_PC_i(3), B1 => 
                           predict_PC_0_3_port, B2 => n2266, ZN => n793);
   U122 : OAI22_X1 port map( A1 => n765, A2 => n644, B1 => predict_PC_0_11_port
                           , B2 => n2266, ZN => n785);
   U340 : OAI22_X1 port map( A1 => n868, A2 => n633, B1 => predict_PC_3_1_port,
                           B2 => n2257, ZN => n898);
   U188 : OAI22_X1 port map( A1 => n800, A2 => n644, B1 => predict_PC_1_11_port
                           , B2 => n2263, ZN => n820);
   U124 : OAI22_X1 port map( A1 => n765, A2 => n640, B1 => predict_PC_0_10_port
                           , B2 => n2266, ZN => n786);
   U204 : OAI22_X1 port map( A1 => n800, A2 => n652, B1 => predict_PC_1_3_port,
                           B2 => n2263, ZN => n828);
   U254 : OAI22_X1 port map( A1 => n834, A2 => n644, B1 => predict_PC_2_11_port
                           , B2 => n2260, ZN => n854);
   U272 : OAI22_X1 port map( A1 => n834, A2 => n650, B1 => predict_PC_2_2_port,
                           B2 => n2260, ZN => n863);
   U274 : OAI22_X1 port map( A1 => n834, A2 => n633, B1 => predict_PC_2_1_port,
                           B2 => n2260, ZN => n864);
   U260 : OAI22_X1 port map( A1 => n834, A2 => n639, B1 => predict_PC_2_8_port,
                           B2 => n2260, ZN => n857);
   U202 : OAI22_X1 port map( A1 => n800, A2 => target_PC_i(4), B1 => 
                           predict_PC_1_4_port, B2 => n2263, ZN => n827);
   U128 : OAI22_X1 port map( A1 => n765, A2 => n639, B1 => predict_PC_0_8_port,
                           B2 => n2266, ZN => n788);
   U140 : OAI22_X1 port map( A1 => n765, A2 => n650, B1 => predict_PC_0_2_port,
                           B2 => n2266, ZN => n794);
   U208 : OAI22_X1 port map( A1 => n800, A2 => n633, B1 => predict_PC_1_1_port,
                           B2 => n2263, ZN => n830);
   U256 : OAI22_X1 port map( A1 => n834, A2 => n640, B1 => predict_PC_2_10_port
                           , B2 => n2260, ZN => n855);
   U268 : OAI22_X1 port map( A1 => n834, A2 => n641, B1 => predict_PC_2_4_port,
                           B2 => n2260, ZN => n861);
   U270 : OAI22_X1 port map( A1 => n834, A2 => n652, B1 => predict_PC_2_3_port,
                           B2 => n2260, ZN => n862);
   U320 : OAI22_X1 port map( A1 => n868, A2 => n644, B1 => predict_PC_3_11_port
                           , B2 => n2257, ZN => n888);
   U206 : OAI22_X1 port map( A1 => n800, A2 => n650, B1 => predict_PC_1_2_port,
                           B2 => n2263, ZN => n829);
   U322 : OAI22_X1 port map( A1 => n868, A2 => n640, B1 => predict_PC_3_10_port
                           , B2 => n2257, ZN => n889);
   U136 : OAI22_X1 port map( A1 => n765, A2 => target_PC_i(4), B1 => 
                           predict_PC_0_4_port, B2 => n2266, ZN => n792);
   U332 : OAI22_X1 port map( A1 => n868, A2 => target_PC_i(5), B1 => 
                           predict_PC_3_5_port, B2 => n2257, ZN => n894);
   U326 : OAI22_X1 port map( A1 => n868, A2 => n639, B1 => predict_PC_3_8_port,
                           B2 => n2257, ZN => n891);
   U132 : OAI22_X1 port map( A1 => n765, A2 => target_PC_i(6), B1 => 
                           predict_PC_0_6_port, B2 => n2266, ZN => n790);
   U266 : OAI22_X1 port map( A1 => n834, A2 => target_PC_i(5), B1 => 
                           predict_PC_2_5_port, B2 => n2260, ZN => n860);
   U334 : OAI22_X1 port map( A1 => n868, A2 => target_PC_i(4), B1 => 
                           predict_PC_3_4_port, B2 => n2257, ZN => n895);
   U190 : OAI22_X1 port map( A1 => n800, A2 => n640, B1 => predict_PC_1_10_port
                           , B2 => n2263, ZN => n821);
   U330 : OAI22_X1 port map( A1 => n868, A2 => target_PC_i(6), B1 => 
                           predict_PC_3_6_port, B2 => n2257, ZN => n893);
   U134 : OAI22_X1 port map( A1 => n765, A2 => target_PC_i(5), B1 => 
                           predict_PC_0_5_port, B2 => n2266, ZN => n791);
   U338 : OAI22_X1 port map( A1 => n868, A2 => n650, B1 => predict_PC_3_2_port,
                           B2 => n2257, ZN => n897);
   U142 : OAI22_X1 port map( A1 => n765, A2 => n633, B1 => predict_PC_0_1_port,
                           B2 => n2266, ZN => n795);
   U336 : OAI22_X1 port map( A1 => n868, A2 => target_PC_i(3), B1 => 
                           predict_PC_3_3_port, B2 => n2257, ZN => n896);
   U264 : OAI22_X1 port map( A1 => n834, A2 => target_PC_i(6), B1 => 
                           predict_PC_2_6_port, B2 => n2260, ZN => n859);
   U1159 : OAI22_X1 port map( A1 => n1284, A2 => n636, B1 => 
                           predict_PC_15_25_port, B2 => n727, ZN => n1350);
   U1145 : OAI22_X1 port map( A1 => n1284, A2 => n649, B1 => 
                           predict_PC_15_26_port, B2 => n727, ZN => n1339);
   U1023 : OAI22_X1 port map( A1 => n1251, A2 => n636, B1 => 
                           predict_PC_14_25_port, B2 => n730, ZN => n1257);
   U888 : OAI22_X1 port map( A1 => n1184, A2 => n636, B1 => 
                           predict_PC_12_25_port, B2 => n737, ZN => n1190);
   U1021 : OAI22_X1 port map( A1 => n1251, A2 => n649, B1 => 
                           predict_PC_14_26_port, B2 => n730, ZN => n1256);
   U955 : OAI22_X1 port map( A1 => n1218, A2 => n636, B1 => 
                           predict_PC_13_25_port, B2 => n733, ZN => n1224);
   U886 : OAI22_X1 port map( A1 => n1184, A2 => n649, B1 => 
                           predict_PC_12_26_port, B2 => n737, ZN => n1189);
   U953 : OAI22_X1 port map( A1 => n1218, A2 => n649, B1 => 
                           predict_PC_13_26_port, B2 => n733, ZN => n1223);
   U554 : OAI22_X1 port map( A1 => n1018, A2 => n649, B1 => 
                           predict_PC_7_26_port, B2 => n988, ZN => n1023);
   U422 : OAI22_X1 port map( A1 => n936, A2 => n649, B1 => predict_PC_5_26_port
                           , B2 => n2253, ZN => n941);
   U821 : OAI22_X1 port map( A1 => n1151, A2 => n636, B1 => 
                           predict_PC_11_25_port, B2 => n976, ZN => n1157);
   U424 : OAI22_X1 port map( A1 => n936, A2 => n636, B1 => predict_PC_5_25_port
                           , B2 => n2253, ZN => n942);
   U687 : OAI22_X1 port map( A1 => n1085, A2 => n649, B1 => 
                           predict_PC_9_26_port, B2 => n982, ZN => n1090);
   U819 : OAI22_X1 port map( A1 => n1151, A2 => n649, B1 => 
                           predict_PC_11_26_port, B2 => n976, ZN => n1156);
   U755 : OAI22_X1 port map( A1 => n1118, A2 => n636, B1 => 
                           predict_PC_10_25_port, B2 => n979, ZN => n1124);
   U556 : OAI22_X1 port map( A1 => n1018, A2 => n636, B1 => 
                           predict_PC_7_25_port, B2 => n988, ZN => n1024);
   U356 : OAI22_X1 port map( A1 => n902, A2 => n649, B1 => predict_PC_4_26_port
                           , B2 => n2256, ZN => n907);
   U623 : OAI22_X1 port map( A1 => n1051, A2 => n636, B1 => 
                           predict_PC_8_25_port, B2 => n985, ZN => n1057);
   U753 : OAI22_X1 port map( A1 => n1118, A2 => n649, B1 => 
                           predict_PC_10_26_port, B2 => n979, ZN => n1123);
   U621 : OAI22_X1 port map( A1 => n1051, A2 => n649, B1 => 
                           predict_PC_8_26_port, B2 => n985, ZN => n1056);
   U488 : OAI22_X1 port map( A1 => n969, A2 => n649, B1 => predict_PC_6_26_port
                           , B2 => n2214, ZN => n990);
   U490 : OAI22_X1 port map( A1 => n969, A2 => n636, B1 => predict_PC_6_25_port
                           , B2 => n2214, ZN => n991);
   U358 : OAI22_X1 port map( A1 => n902, A2 => n636, B1 => predict_PC_4_25_port
                           , B2 => n2256, ZN => n908);
   U689 : OAI22_X1 port map( A1 => n1085, A2 => n636, B1 => 
                           predict_PC_9_25_port, B2 => n982, ZN => n1091);
   U292 : OAI22_X1 port map( A1 => n868, A2 => n636, B1 => predict_PC_3_25_port
                           , B2 => n2259, ZN => n874);
   U158 : OAI22_X1 port map( A1 => n800, A2 => n649, B1 => predict_PC_1_26_port
                           , B2 => n2265, ZN => n805);
   U224 : OAI22_X1 port map( A1 => n834, A2 => n649, B1 => predict_PC_2_26_port
                           , B2 => n2262, ZN => n839);
   U94 : OAI22_X1 port map( A1 => n765, A2 => n636, B1 => predict_PC_0_25_port,
                           B2 => n2268, ZN => n771);
   U290 : OAI22_X1 port map( A1 => n868, A2 => n649, B1 => predict_PC_3_26_port
                           , B2 => n2259, ZN => n873);
   U92 : OAI22_X1 port map( A1 => n765, A2 => n649, B1 => predict_PC_0_26_port,
                           B2 => n2268, ZN => n770);
   U160 : OAI22_X1 port map( A1 => n800, A2 => n636, B1 => predict_PC_1_25_port
                           , B2 => n2265, ZN => n806);
   U226 : OAI22_X1 port map( A1 => n834, A2 => n636, B1 => predict_PC_2_25_port
                           , B2 => n2262, ZN => n840);
   U68 : NAND2_X1 port map( A1 => n2286, A2 => n2288, ZN => n696);
   U67 : AOI22_X1 port map( A1 => n2285, A2 => taken_o_port, B1 => n663, B2 => 
                           n696, ZN => n736);
   U34 : OAI21_X1 port map( B1 => n2285, B2 => n713, A => n1284, ZN => n2096);
   U40 : OAI21_X1 port map( B1 => n2285, B2 => n710, A => n1184, ZN => n2093);
   U38 : OAI21_X1 port map( B1 => n2285, B2 => n711, A => n1218, ZN => n2094);
   U36 : OAI21_X1 port map( B1 => n2285, B2 => n712, A => n1251, ZN => n2095);
   U54 : OAI21_X1 port map( B1 => n2285, B2 => n702, A => n936, ZN => n2086);
   U44 : OAI21_X1 port map( B1 => n2285, B2 => n708, A => n1118, ZN => n2091);
   U48 : OAI21_X1 port map( B1 => n2285, B2 => n706, A => n1051, ZN => n2089);
   U52 : OAI21_X1 port map( B1 => n2285, B2 => n704, A => n969, ZN => n2087);
   U46 : OAI21_X1 port map( B1 => n2285, B2 => n707, A => n1085, ZN => n2090);
   U42 : OAI21_X1 port map( B1 => n2285, B2 => n709, A => n1151, ZN => n2092);
   U50 : OAI21_X1 port map( B1 => n2285, B2 => n705, A => n1018, ZN => n2088);
   U56 : OAI21_X1 port map( B1 => n2285, B2 => n700, A => n902, ZN => n2085);
   U58 : OAI21_X1 port map( B1 => n2285, B2 => n698, A => n868, ZN => n2084);
   U60 : OAI21_X1 port map( B1 => n2285, B2 => n695, A => n834, ZN => n2083);
   U62 : OAI21_X1 port map( B1 => n2285, B2 => n694, A => n800, ZN => n2082);
   U64 : OAI21_X1 port map( B1 => n2285, B2 => n665, A => n765, ZN => n2081);
   U1188 : AOI22_X1 port map( A1 => n2287, A2 => n601, B1 => n678, B2 => n2285,
                           ZN => n1582);
   U1244 : AOI22_X1 port map( A1 => n2287, A2 => n605, B1 => n683, B2 => n2285,
                           ZN => n1574);
   U1216 : AOI22_X1 port map( A1 => n2287, A2 => n603, B1 => n680, B2 => n2285,
                           ZN => n1578);
   U1272 : AOI22_X1 port map( A1 => n2287, A2 => n607, B1 => n685, B2 => n2285,
                           ZN => n1570);
   U1356 : AOI22_X1 port map( A1 => n2287, A2 => n613, B1 => n691, B2 => n2285,
                           ZN => n1558);
   U1412 : AOI22_X1 port map( A1 => n2287, A2 => n617, B1 => n668, B2 => n2285,
                           ZN => n1550);
   U1230 : AOI22_X1 port map( A1 => n2287, A2 => n604, B1 => n681, B2 => n2285,
                           ZN => n1576);
   U1258 : AOI22_X1 port map( A1 => n2287, A2 => n606, B1 => n684, B2 => n2285,
                           ZN => n1572);
   U1342 : AOI22_X1 port map( A1 => n2287, A2 => n612, B1 => n690, B2 => n2285,
                           ZN => n1560);
   U1314 : AOI22_X1 port map( A1 => n2287, A2 => n610, B1 => n688, B2 => n2285,
                           ZN => n1564);
   U1300 : AOI22_X1 port map( A1 => n2287, A2 => n609, B1 => n687, B2 => n2285,
                           ZN => n1566);
   U1202 : AOI22_X1 port map( A1 => n2287, A2 => n602, B1 => n679, B2 => n2285,
                           ZN => n1580);
   U1286 : AOI22_X1 port map( A1 => n2287, A2 => n608, B1 => n686, B2 => n2285,
                           ZN => n1568);
   U1328 : AOI22_X1 port map( A1 => n2287, A2 => n611, B1 => n689, B2 => n2285,
                           ZN => n1562);
   U1454 : AOI22_X1 port map( A1 => n2287, A2 => n620, B1 => n671, B2 => n2285,
                           ZN => n1544);
   U1146 : AOI22_X1 port map( A1 => n2287, A2 => n598, B1 => n675, B2 => n2285,
                           ZN => n1588);
   U1426 : AOI22_X1 port map( A1 => stall_i, A2 => n618, B1 => n669, B2 => 
                           n2285, ZN => n1548);
   U1160 : AOI22_X1 port map( A1 => stall_i, A2 => n599, B1 => n676, B2 => 
                           n2285, ZN => n1586);
   U1482 : AOI22_X1 port map( A1 => stall_i, A2 => n622, B1 => n674, B2 => 
                           n2285, ZN => n1540);
   U1398 : AOI22_X1 port map( A1 => stall_i, A2 => n616, B1 => n667, B2 => 
                           n2285, ZN => n1552);
   U1384 : AOI22_X1 port map( A1 => stall_i, A2 => n615, B1 => n666, B2 => 
                           n2285, ZN => n1554);
   U1370 : AOI22_X1 port map( A1 => stall_i, A2 => n614, B1 => n692, B2 => 
                           n2285, ZN => n1556);
   U1468 : AOI22_X1 port map( A1 => stall_i, A2 => n621, B1 => n672, B2 => 
                           n2285, ZN => n1542);
   U1080 : AOI22_X1 port map( A1 => stall_i, A2 => n593, B1 => n673, B2 => 
                           n2285, ZN => n1598);
   U1174 : AOI22_X1 port map( A1 => stall_i, A2 => n600, B1 => n677, B2 => 
                           n2285, ZN => n1584);
   U1496 : AOI22_X1 port map( A1 => stall_i, A2 => n623, B1 => n682, B2 => 
                           n2285, ZN => n1538);
   U1440 : AOI22_X1 port map( A1 => stall_i, A2 => n619, B1 => n670, B2 => 
                           n2285, ZN => n1546);
   U1513 : AOI22_X1 port map( A1 => stall_i, A2 => n624, B1 => n693, B2 => 
                           n2285, ZN => n1536);
   U33 : OAI22_X1 port map( A1 => n2285, A2 => n660, B1 => n696, B2 => n703, ZN
                           => n2097);
   U32 : OAI22_X1 port map( A1 => n2285, A2 => n662, B1 => n696, B2 => n701, ZN
                           => n2098);
   U31 : OAI22_X1 port map( A1 => n2285, A2 => n661, B1 => n696, B2 => n699, ZN
                           => n2099);
   U30 : OAI22_X1 port map( A1 => n2285, A2 => n664, B1 => n696, B2 => n697, ZN
                           => n2100);
   U941 : NAND2_X1 port map( A1 => n662, A2 => n660, ZN => n797);
   U1512 : NAND2_X1 port map( A1 => n589, A2 => n588, ZN => n900);
   U1008 : NAND2_X1 port map( A1 => n588, A2 => n662, ZN => n832);
   U1076 : NAND2_X1 port map( A1 => n589, A2 => n660, ZN => n866);
   U1547 : NOR2_X1 port map( A1 => n2209, A2 => n2202, ZN => n761);
   U1538 : NAND2_X1 port map( A1 => TAG_i(3), A2 => n699, ZN => n2208);
   U1529 : NAND2_X1 port map( A1 => TAG_i(2), A2 => n697, ZN => n2203);
   U1550 : NAND2_X1 port map( A1 => TAG_i(1), A2 => n703, ZN => n2201);
   U1522 : NAND2_X1 port map( A1 => n699, A2 => n697, ZN => n2199);
   U1543 : NOR2_X1 port map( A1 => n2198, A2 => n2209, ZN => n762);
   U1549 : NOR2_X1 port map( A1 => n2209, A2 => n2201, ZN => n760);
   U1534 : NOR2_X1 port map( A1 => n2201, A2 => n2208, ZN => n758);
   U1537 : NOR2_X1 port map( A1 => n2198, A2 => n2208, ZN => n756);
   U1525 : NOR2_X1 port map( A1 => n2198, A2 => n2203, ZN => n750);
   U1528 : NOR2_X1 port map( A1 => n2201, A2 => n2203, ZN => n748);
   U1544 : NAND2_X1 port map( A1 => n701, A2 => n703, ZN => n2198);
   U1517 : NOR2_X1 port map( A1 => n2198, A2 => n2199, ZN => n747);
   U1601 : NAND3_X1 port map( A1 => n590, A2 => n2286, A3 => n664, ZN => n934);
   U1602 : NAND3_X1 port map( A1 => n591, A2 => n2286, A3 => n661, ZN => n1083)
                           ;
   U1600 : NAND3_X1 port map( A1 => n2286, A2 => n664, A3 => n661, ZN => n798);
   U1607 : NAND3_X1 port map( A1 => n591, A2 => n590, A3 => n2286, ZN => n1216)
                           ;
   U1530 : INV_X1 port map( A => TAG_i(3), ZN => n697);
   U1539 : INV_X1 port map( A => TAG_i(2), ZN => n699);
   U1551 : INV_X1 port map( A => TAG_i(0), ZN => n703);
   U1545 : INV_X1 port map( A => TAG_i(1), ZN => n701);
   U71 : AND4_X1 port map( A1 => n740, A2 => n741, A3 => n742, A4 => n743, ZN 
                           => n739);
   U76 : AND4_X1 port map( A1 => n752, A2 => n753, A3 => n754, A4 => n755, ZN 
                           => n738);
   U1107 : OR2_X1 port map( A1 => n1307, A2 => n1308, ZN => 
                           predicted_next_PC_o_29_port);
   U1133 : OR2_X1 port map( A1 => n1329, A2 => n1330, ZN => 
                           predicted_next_PC_o_27_port);
   U1120 : OR2_X1 port map( A1 => n1318, A2 => n1319, ZN => 
                           predicted_next_PC_o_28_port);
   U1094 : OR2_X1 port map( A1 => n1296, A2 => n1297, ZN => 
                           predicted_next_PC_o_30_port);
   U9 : INV_X1 port map( A => n673, ZN => predicted_next_PC_o_31_port);
   U22 : INV_X1 port map( A => n686, ZN => predicted_next_PC_o_16_port);
   U6 : INV_X1 port map( A => n670, ZN => predicted_next_PC_o_5_port);
   U7 : INV_X1 port map( A => n671, ZN => predicted_next_PC_o_4_port);
   U23 : INV_X1 port map( A => n687, ZN => predicted_next_PC_o_15_port);
   U20 : INV_X1 port map( A => n684, ZN => predicted_next_PC_o_18_port);
   U21 : INV_X1 port map( A => n685, ZN => predicted_next_PC_o_17_port);
   U13 : INV_X1 port map( A => n677, ZN => predicted_next_PC_o_24_port);
   U15 : INV_X1 port map( A => n679, ZN => predicted_next_PC_o_22_port);
   U10 : INV_X1 port map( A => n674, ZN => predicted_next_PC_o_2_port);
   U2 : INV_X1 port map( A => n666, ZN => predicted_next_PC_o_9_port);
   U3 : INV_X1 port map( A => n667, ZN => predicted_next_PC_o_8_port);
   U5 : INV_X1 port map( A => n669, ZN => predicted_next_PC_o_6_port);
   U19 : INV_X1 port map( A => n683, ZN => predicted_next_PC_o_19_port);
   U17 : INV_X1 port map( A => n681, ZN => predicted_next_PC_o_20_port);
   U16 : INV_X1 port map( A => n680, ZN => predicted_next_PC_o_21_port);
   U14 : INV_X1 port map( A => n678, ZN => predicted_next_PC_o_23_port);
   U8 : INV_X1 port map( A => n672, ZN => predicted_next_PC_o_3_port);
   U4 : INV_X1 port map( A => n668, ZN => predicted_next_PC_o_7_port);
   U12 : INV_X1 port map( A => n676, ZN => predicted_next_PC_o_25_port);
   U11 : INV_X1 port map( A => n675, ZN => predicted_next_PC_o_26_port);
   U27 : INV_X1 port map( A => n691, ZN => predicted_next_PC_o_11_port);
   U25 : INV_X1 port map( A => n689, ZN => predicted_next_PC_o_13_port);
   U24 : INV_X1 port map( A => n688, ZN => predicted_next_PC_o_14_port);
   U18 : INV_X1 port map( A => n682, ZN => predicted_next_PC_o_1_port);
   U29 : INV_X1 port map( A => n693, ZN => predicted_next_PC_o_0_port);
   U28 : INV_X1 port map( A => n692, ZN => predicted_next_PC_o_10_port);
   U26 : INV_X1 port map( A => n690, ZN => predicted_next_PC_o_12_port);
   U66 : INV_X1 port map( A => n736, ZN => n2080);
   U1557 : OAI21_X1 port map( B1 => was_taken_i, B2 => n663, A => n592, ZN => 
                           n2212);
   U1340 : INV_X1 port map( A => n1493, ZN => n1561);
   U800 : INV_X1 port map( A => n1147, ZN => n1730);
   U569 : INV_X1 port map( A => n1031, ZN => n1842);
   U429 : INV_X1 port map( A => n945, ZN => n1910);
   U860 : INV_X1 port map( A => n1177, ZN => n1701);
   U992 : INV_X1 port map( A => n1243, ZN => n1638);
   U858 : INV_X1 port map( A => n1176, ZN => n1702);
   U1062 : INV_X1 port map( A => n1277, ZN => n1605);
   U503 : INV_X1 port map( A => n998, ZN => n1874);
   U191 : INV_X1 port map( A => n822, ZN => n2025);
   U804 : INV_X1 port map( A => n1149, ZN => n1728);
   U1000 : INV_X1 port map( A => n1247, ZN => n1634);
   U1060 : INV_X1 port map( A => n1276, ZN => n1606);
   U636 : INV_X1 port map( A => n1064, ZN => n1810);
   U720 : INV_X1 port map( A => n1107, ZN => n1769);
   U197 : INV_X1 port map( A => n825, ZN => n2022);
   U461 : INV_X1 port map( A => n961, ZN => n1894);
   U852 : INV_X1 port map( A => n1173, ZN => n1705);
   U463 : INV_X1 port map( A => n962, ZN => n1893);
   U1072 : INV_X1 port map( A => n1282, ZN => n1600);
   U305 : INV_X1 port map( A => n881, ZN => n1970);
   U455 : INV_X1 port map( A => n958, ZN => n1897);
   U397 : INV_X1 port map( A => n928, ZN => n1925);
   U199 : INV_X1 port map( A => n826, ZN => n2021);
   U449 : INV_X1 port map( A => n955, ZN => n1900);
   U395 : INV_X1 port map( A => n927, ZN => n1926);
   U1054 : INV_X1 port map( A => n1273, ZN => n1609);
   U927 : INV_X1 port map( A => n1210, ZN => n1669);
   U712 : INV_X1 port map( A => n1103, ZN => n1773);
   U1382 : INV_X1 port map( A => n1526, ZN => n1555);
   U994 : INV_X1 port map( A => n1244, ZN => n1637);
   U201 : INV_X1 port map( A => n827, ZN => n2020);
   U836 : INV_X1 port map( A => n1165, ZN => n1713);
   U925 : INV_X1 port map( A => n1209, ZN => n1670);
   U702 : INV_X1 port map( A => n1098, ZN => n1778);
   U437 : INV_X1 port map( A => n949, ZN => n1906);
   U933 : INV_X1 port map( A => n1213, ZN => n1666);
   U323 : INV_X1 port map( A => n890, ZN => n1961);
   U389 : INV_X1 port map( A => n924, ZN => n1929);
   U135 : INV_X1 port map( A => n792, ZN => n2052);
   U333 : INV_X1 port map( A => n895, ZN => n1956);
   U137 : INV_X1 port map( A => n793, ZN => n2051);
   U796 : INV_X1 port map( A => n1145, ZN => n1732);
   U980 : INV_X1 port map( A => n1237, ZN => n1644);
   U595 : INV_X1 port map( A => n1044, ZN => n1829);
   U335 : INV_X1 port map( A => n896, ZN => n1955);
   U660 : INV_X1 port map( A => n1076, ZN => n1798);
   U794 : INV_X1 port map( A => n1144, ZN => n1733);
   U792 : INV_X1 port map( A => n1143, ZN => n1734);
   U1480 : INV_X1 port map( A => n2169, ZN => n1541);
   U768 : INV_X1 port map( A => n1131, ZN => n1746);
   U662 : INV_X1 port map( A => n1077, ZN => n1797);
   U776 : INV_X1 port map( A => n1135, ZN => n1742);
   U173 : INV_X1 port map( A => n813, ZN => n2034);
   U521 : INV_X1 port map( A => n1007, ZN => n1865);
   U1424 : INV_X1 port map( A => n2125, ZN => n1549);
   U601 : INV_X1 port map( A => n1047, ZN => n1826);
   U257 : INV_X1 port map( A => n856, ZN => n1993);
   U529 : INV_X1 port map( A => n1011, ZN => n1861);
   U371 : INV_X1 port map( A => n915, ZN => n1938);
   U263 : INV_X1 port map( A => n859, ZN => n1990);
   U265 : INV_X1 port map( A => n860, ZN => n1989);
   U527 : INV_X1 port map( A => n1010, ZN => n1862);
   U786 : INV_X1 port map( A => n1140, ZN => n1737);
   U331 : INV_X1 port map( A => n894, ZN => n1957);
   U587 : INV_X1 port map( A => n1040, ZN => n1833);
   U732 : INV_X1 port map( A => n1113, ZN => n1763);
   U1508 : INV_X1 port map( A => n2191, ZN => n1537);
   U728 : INV_X1 port map( A => n1111, ZN => n1765);
   U585 : INV_X1 port map( A => n1039, ZN => n1834);
   U919 : INV_X1 port map( A => n1206, ZN => n1673);
   U726 : INV_X1 port map( A => n1110, ZN => n1766);
   U117 : INV_X1 port map( A => n783, ZN => n2061);
   U183 : INV_X1 port map( A => n818, ZN => n2029);
   U125 : INV_X1 port map( A => n787, ZN => n2057);
   U1438 : INV_X1 port map( A => n2136, ZN => n1547);
   U986 : INV_X1 port map( A => n1240, ZN => n1641);
   U730 : INV_X1 port map( A => n1112, ZN => n1764);
   U329 : INV_X1 port map( A => n893, ZN => n1958);
   U654 : INV_X1 port map( A => n1073, ZN => n1801);
   U593 : INV_X1 port map( A => n1043, ZN => n1830);
   U1036 : INV_X1 port map( A => n1264, ZN => n1618);
   U131 : INV_X1 port map( A => n790, ZN => n2054);
   U133 : INV_X1 port map( A => n791, ZN => n2053);
   U840 : INV_X1 port map( A => n1167, ZN => n1711);
   U738 : INV_X1 port map( A => n1116, ZN => n1760);
   U261 : INV_X1 port map( A => n858, ZN => n1991);
   U666 : INV_X1 port map( A => n1079, ZN => n1795);
   U788 : INV_X1 port map( A => n1141, ZN => n1736);
   U784 : INV_X1 port map( A => n1139, ZN => n1738);
   U982 : INV_X1 port map( A => n1238, ZN => n1643);
   U179 : INV_X1 port map( A => n816, ZN => n2031);
   U782 : INV_X1 port map( A => n1138, ZN => n1739);
   U169 : INV_X1 port map( A => n811, ZN => n2036);
   U1032 : INV_X1 port map( A => n1262, ZN => n1620);
   U1200 : INV_X1 port map( A => n1383, ZN => n1581);
   U605 : INV_X1 port map( A => n1049, ZN => n1824);
   U1298 : INV_X1 port map( A => n1460, ZN => n1567);
   U129 : INV_X1 port map( A => n789, ZN => n2055);
   U1038 : INV_X1 port map( A => n1265, ZN => n1617);
   U962 : INV_X1 port map( A => n1228, ZN => n1653);
   U229 : INV_X1 port map( A => n842, ZN => n2007);
   U1034 : INV_X1 port map( A => n1263, ZN => n1619);
   U917 : INV_X1 port map( A => n1205, ZN => n1674);
   U798 : INV_X1 port map( A => n1146, ZN => n1731);
   U915 : INV_X1 port map( A => n1204, ZN => n1675);
   U652 : INV_X1 port map( A => n1072, ZN => n1802);
   U525 : INV_X1 port map( A => n1009, ZN => n1863);
   U828 : INV_X1 port map( A => n1161, ZN => n1717);
   U1270 : INV_X1 port map( A => n1438, ZN => n1571);
   U780 : INV_X1 port map( A => n1137, ZN => n1740);
   U167 : INV_X1 port map( A => n810, ZN => n2037);
   U295 : INV_X1 port map( A => n876, ZN => n1975);
   U692 : INV_X1 port map( A => n1093, ZN => n1783);
   U231 : INV_X1 port map( A => n843, ZN => n2006);
   U656 : INV_X1 port map( A => n1074, ZN => n1800);
   U259 : INV_X1 port map( A => n857, ZN => n1992);
   U341 : INV_X1 port map( A => n899, ZN => n1952);
   U984 : INV_X1 port map( A => n1239, ZN => n1642);
   U267 : INV_X1 port map( A => n861, ZN => n1988);
   U523 : INV_X1 port map( A => n1008, ZN => n1864);
   U139 : INV_X1 port map( A => n794, ZN => n2050);
   U978 : INV_X1 port map( A => n1236, ZN => n1645);
   U964 : INV_X1 port map( A => n1229, ZN => n1652);
   U251 : INV_X1 port map( A => n853, ZN => n1996);
   U513 : INV_X1 port map( A => n1003, ZN => n1869);
   U790 : INV_X1 port map( A => n1142, ZN => n1735);
   U511 : INV_X1 port map( A => n1002, ZN => n1870);
   U772 : INV_X1 port map( A => n1133, ZN => n1744);
   U958 : INV_X1 port map( A => n1226, ZN => n1655);
   U672 : INV_X1 port map( A => n1082, ZN => n1792);
   U175 : INV_X1 port map( A => n814, ZN => n2033);
   U509 : INV_X1 port map( A => n1001, ZN => n1871);
   U770 : INV_X1 port map( A => n1132, ZN => n1745);
   U271 : INV_X1 port map( A => n863, ZN => n1986);
   U247 : INV_X1 port map( A => n851, ZN => n1998);
   U899 : INV_X1 port map( A => n1196, ZN => n1683);
   U1410 : INV_X1 port map( A => n2114, ZN => n1551);
   U515 : INV_X1 port map( A => n1004, ZN => n1868);
   U249 : INV_X1 port map( A => n852, ZN => n1997);
   U970 : INV_X1 port map( A => n1232, ZN => n1649);
   U337 : INV_X1 port map( A => n897, ZN => n1954);
   U909 : INV_X1 port map( A => n1201, ZN => n1678);
   U517 : INV_X1 port map( A => n1005, ZN => n1867);
   U269 : INV_X1 port map( A => n862, ZN => n1987);
   U766 : INV_X1 port map( A => n1130, ZN => n1747);
   U842 : INV_X1 port map( A => n1168, ZN => n1710);
   U824 : INV_X1 port map( A => n1159, ZN => n1719);
   U1284 : INV_X1 port map( A => n1449, ZN => n1569);
   U764 : INV_X1 port map( A => n1129, ZN => n1748);
   U907 : INV_X1 port map( A => n1200, ZN => n1679);
   U762 : INV_X1 port map( A => n1128, ZN => n1749);
   U275 : INV_X1 port map( A => n865, ZN => n1984);
   U599 : INV_X1 port map( A => n1046, ZN => n1827);
   U774 : INV_X1 port map( A => n1134, ZN => n1743);
   U911 : INV_X1 port map( A => n1202, ZN => n1677);
   U968 : INV_X1 port map( A => n1231, ZN => n1650);
   U369 : INV_X1 port map( A => n914, ZN => n1939);
   U531 : INV_X1 port map( A => n1012, ZN => n1860);
   U913 : INV_X1 port map( A => n1203, ZN => n1676);
   U373 : INV_X1 port map( A => n916, ZN => n1937);
   U245 : INV_X1 port map( A => n850, ZN => n1999);
   U760 : INV_X1 port map( A => n1127, ZN => n1750);
   U972 : INV_X1 port map( A => n1233, ZN => n1648);
   U243 : INV_X1 port map( A => n849, ZN => n2000);
   U1026 : INV_X1 port map( A => n1259, ZN => n1623);
   U758 : INV_X1 port map( A => n1126, ZN => n1751);
   U1186 : INV_X1 port map( A => n1372, ZN => n1583);
   U253 : INV_X1 port map( A => n854, ZN => n1995);
   U960 : INV_X1 port map( A => n1227, ZN => n1654);
   U974 : INV_X1 port map( A => n1234, ZN => n1647);
   U519 : INV_X1 port map( A => n1006, ZN => n1866);
   U644 : INV_X1 port map( A => n1068, ZN => n1806);
   U241 : INV_X1 port map( A => n848, ZN => n2001);
   U664 : INV_X1 port map( A => n1078, ZN => n1796);
   U163 : INV_X1 port map( A => n808, ZN => n2039);
   U597 : INV_X1 port map( A => n1045, ZN => n1828);
   U905 : INV_X1 port map( A => n1199, ZN => n1680);
   U255 : INV_X1 port map( A => n855, ZN => n1994);
   U976 : INV_X1 port map( A => n1235, ZN => n1646);
   U177 : INV_X1 port map( A => n815, ZN => n2032);
   U239 : INV_X1 port map( A => n847, ZN => n2002);
   U658 : INV_X1 port map( A => n1075, ZN => n1799);
   U668 : INV_X1 port map( A => n1080, ZN => n1794);
   U1028 : INV_X1 port map( A => n1260, ZN => n1622);
   U143 : INV_X1 port map( A => n796, ZN => n2048);
   U966 : INV_X1 port map( A => n1230, ZN => n1651);
   U237 : INV_X1 port map( A => n846, ZN => n2003);
   U778 : INV_X1 port map( A => n1136, ZN => n1741);
   U642 : INV_X1 port map( A => n1067, ZN => n1807);
   U235 : INV_X1 port map( A => n845, ZN => n2004);
   U171 : INV_X1 port map( A => n812, ZN => n2035);
   U361 : INV_X1 port map( A => n910, ZN => n1943);
   U826 : INV_X1 port map( A => n1160, ZN => n1718);
   U165 : INV_X1 port map( A => n809, ZN => n2038);
   U233 : INV_X1 port map( A => n844, ZN => n2005);
   U1030 : INV_X1 port map( A => n1261, ZN => n1621);
   U533 : INV_X1 port map( A => n1013, ZN => n1859);
   U433 : INV_X1 port map( A => n947, ZN => n1908);
   U710 : INV_X1 port map( A => n1102, ZN => n1774);
   U561 : INV_X1 port map( A => n1027, ZN => n1846);
   U107 : INV_X1 port map( A => n778, ZN => n2066);
   U387 : INV_X1 port map( A => n923, ZN => n1930);
   U694 : INV_X1 port map( A => n1094, ZN => n1782);
   U990 : INV_X1 port map( A => n1242, ZN => n1639);
   U435 : INV_X1 port map( A => n948, ZN => n1907);
   U209 : INV_X1 port map( A => n831, ZN => n2016);
   U937 : INV_X1 port map( A => n1215, ZN => n1664);
   U718 : INV_X1 port map( A => n1106, ZN => n1770);
   U559 : INV_X1 port map( A => n1026, ZN => n1847);
   U363 : INV_X1 port map( A => n911, ZN => n1942);
   U309 : INV_X1 port map( A => n883, ZN => n1968);
   U1228 : INV_X1 port map( A => n1405, ZN => n1577);
   U921 : INV_X1 port map( A => n1207, ZN => n1672);
   U105 : INV_X1 port map( A => n777, ZN => n2067);
   U1050 : INV_X1 port map( A => n1271, ZN => n1611);
   U405 : INV_X1 port map( A => n932, ZN => n1921);
   U439 : INV_X1 port map( A => n950, ZN => n1905);
   U317 : INV_X1 port map( A => n887, ZN => n1964);
   U856 : INV_X1 port map( A => n1175, ZN => n1703);
   U441 : INV_X1 port map( A => n951, ZN => n1904);
   U205 : INV_X1 port map( A => n829, ZN => n2018);
   U499 : INV_X1 port map( A => n996, ZN => n1876);
   U497 : INV_X1 port map( A => n995, ZN => n1877);
   U1396 : INV_X1 port map( A => n2103, ZN => n1553);
   U846 : INV_X1 port map( A => n1170, ZN => n1708);
   U903 : INV_X1 port map( A => n1198, ZN => n1681);
   U1066 : INV_X1 port map( A => n1279, ZN => n1603);
   U716 : INV_X1 port map( A => n1105, ZN => n1771);
   U391 : INV_X1 port map( A => n925, ZN => n1928);
   U495 : INV_X1 port map( A => n994, ZN => n1878);
   U923 : INV_X1 port map( A => n1208, ZN => n1671);
   U187 : INV_X1 port map( A => n820, ZN => n2027);
   U193 : INV_X1 port map( A => n823, ZN => n2024);
   U901 : INV_X1 port map( A => n1197, ZN => n1682);
   U203 : INV_X1 port map( A => n828, ZN => n2019);
   U696 : INV_X1 port map( A => n1095, ZN => n1781);
   U493 : INV_X1 port map( A => n993, ZN => n1879);
   U1052 : INV_X1 port map( A => n1272, ZN => n1610);
   U632 : INV_X1 port map( A => n1062, ZN => n1812);
   U403 : INV_X1 port map( A => n931, ZN => n1922);
   U443 : INV_X1 port map( A => n952, ZN => n1903);
   U103 : INV_X1 port map( A => n776, ZN => n2068);
   U321 : INV_X1 port map( A => n889, ZN => n1962);
   U393 : INV_X1 port map( A => n926, ZN => n1927);
   U848 : INV_X1 port map( A => n1171, ZN => n1707);
   U101 : INV_X1 port map( A => n775, ZN => n2069);
   U996 : INV_X1 port map( A => n1245, ZN => n1636);
   U303 : INV_X1 port map( A => n880, ZN => n1971);
   U630 : INV_X1 port map( A => n1061, ZN => n1813);
   U1058 : INV_X1 port map( A => n1275, ZN => n1607);
   U1068 : INV_X1 port map( A => n1280, ZN => n1602);
   U189 : INV_X1 port map( A => n821, ZN => n2026);
   U99 : INV_X1 port map( A => n774, ZN => n2070);
   U1242 : INV_X1 port map( A => n1416, ZN => n1575);
   U473 : INV_X1 port map( A => n967, ZN => n1888);
   U539 : INV_X1 port map( A => n1016, ZN => n1856);
   U850 : INV_X1 port map( A => n1172, ZN => n1706);
   U97 : INV_X1 port map( A => n773, ZN => n2071);
   U469 : INV_X1 port map( A => n965, ZN => n1890);
   U1452 : INV_X1 port map( A => n2147, ZN => n1545);
   U401 : INV_X1 port map( A => n930, ZN => n1923);
   U399 : INV_X1 port map( A => n929, ZN => n1924);
   U445 : INV_X1 port map( A => n953, ZN => n1902);
   U467 : INV_X1 port map( A => n964, ZN => n1891);
   U1354 : INV_X1 port map( A => n1504, ZN => n1559);
   U1368 : INV_X1 port map( A => n1515, ZN => n1557);
   U1326 : INV_X1 port map( A => n1482, ZN => n1563);
   U638 : INV_X1 port map( A => n1065, ZN => n1809);
   U447 : INV_X1 port map( A => n954, ZN => n1901);
   U465 : INV_X1 port map( A => n963, ZN => n1892);
   U698 : INV_X1 port map( A => n1096, ZN => n1780);
   U714 : INV_X1 port map( A => n1104, ZN => n1772);
   U459 : INV_X1 port map( A => n960, ZN => n1895);
   U998 : INV_X1 port map( A => n1246, ZN => n1635);
   U319 : INV_X1 port map( A => n888, ZN => n1963);
   U307 : INV_X1 port map( A => n882, ZN => n1969);
   U457 : INV_X1 port map( A => n959, ZN => n1896);
   U648 : INV_X1 port map( A => n1070, ZN => n1804);
   U453 : INV_X1 port map( A => n957, ZN => n1898);
   U854 : INV_X1 port map( A => n1174, ZN => n1704);
   U1056 : INV_X1 port map( A => n1274, ZN => n1608);
   U700 : INV_X1 port map( A => n1097, ZN => n1779);
   U195 : INV_X1 port map( A => n824, ZN => n2023);
   U451 : INV_X1 port map( A => n956, ZN => n1899);
   U988 : INV_X1 port map( A => n1241, ZN => n1640);
   U297 : INV_X1 port map( A => n877, ZN => n1974);
   U591 : INV_X1 port map( A => n1042, ZN => n1831);
   U313 : INV_X1 port map( A => n885, ZN => n1966);
   U864 : INV_X1 port map( A => n1179, ZN => n1699);
   U866 : INV_X1 port map( A => n1180, ZN => n1698);
   U706 : INV_X1 port map( A => n1100, ZN => n1776);
   U589 : INV_X1 port map( A => n1041, ZN => n1832);
   U734 : INV_X1 port map( A => n1114, ZN => n1762);
   U127 : INV_X1 port map( A => n788, ZN => n2056);
   U929 : INV_X1 port map( A => n1211, ZN => n1668);
   U646 : INV_X1 port map( A => n1069, ZN => n1805);
   U1256 : INV_X1 port map( A => n1427, ZN => n1573);
   U830 : INV_X1 port map( A => n1162, ZN => n1716);
   U1312 : INV_X1 port map( A => n1471, ZN => n1565);
   U897 : INV_X1 port map( A => n1195, ZN => n1684);
   U535 : INV_X1 port map( A => n1014, ZN => n1858);
   U123 : INV_X1 port map( A => n786, ZN => n2058);
   U626 : INV_X1 port map( A => n1059, ZN => n1815);
   U583 : INV_X1 port map( A => n1038, ZN => n1835);
   U1040 : INV_X1 port map( A => n1266, ZN => n1616);
   U375 : INV_X1 port map( A => n917, ZN => n1936);
   U181 : INV_X1 port map( A => n817, ZN => n2030);
   U895 : INV_X1 port map( A => n1194, ZN => n1685);
   U581 : INV_X1 port map( A => n1037, ZN => n1836);
   U708 : INV_X1 port map( A => n1101, ZN => n1775);
   U862 : INV_X1 port map( A => n1178, ZN => n1700);
   U1004 : INV_X1 port map( A => n1249, ZN => n1632);
   U121 : INV_X1 port map( A => n785, ZN => n2059);
   U579 : INV_X1 port map( A => n1036, ZN => n1837);
   U870 : INV_X1 port map( A => n1182, ZN => n1696);
   U1042 : INV_X1 port map( A => n1267, ZN => n1615);
   U377 : INV_X1 port map( A => n918, ZN => n1935);
   U931 : INV_X1 port map( A => n1212, ZN => n1667);
   U1466 : INV_X1 port map( A => n2158, ZN => n1543);
   U577 : INV_X1 port map( A => n1035, ZN => n1838);
   U119 : INV_X1 port map( A => n784, ZN => n2060);
   U379 : INV_X1 port map( A => n919, ZN => n1934);
   U1044 : INV_X1 port map( A => n1268, ZN => n1614);
   U315 : INV_X1 port map( A => n886, ZN => n1965);
   U365 : INV_X1 port map( A => n912, ZN => n1941);
   U507 : INV_X1 port map( A => n1000, ZN => n1872);
   U381 : INV_X1 port map( A => n920, ZN => n1933);
   U832 : INV_X1 port map( A => n1163, ZN => n1715);
   U1064 : INV_X1 port map( A => n1278, ZN => n1604);
   U1214 : INV_X1 port map( A => n1394, ZN => n1579);
   U575 : INV_X1 port map( A => n1034, ZN => n1839);
   U407 : INV_X1 port map( A => n933, ZN => n1920);
   U650 : INV_X1 port map( A => n1071, ZN => n1803);
   U115 : INV_X1 port map( A => n782, ZN => n2062);
   U571 : INV_X1 port map( A => n1032, ZN => n1841);
   U640 : INV_X1 port map( A => n1066, ZN => n1808);
   U724 : INV_X1 port map( A => n1109, ZN => n1767);
   U383 : INV_X1 port map( A => n921, ZN => n1932);
   U113 : INV_X1 port map( A => n781, ZN => n2063);
   U834 : INV_X1 port map( A => n1164, ZN => n1714);
   U573 : INV_X1 port map( A => n1033, ZN => n1840);
   U722 : INV_X1 port map( A => n1108, ZN => n1768);
   U1046 : INV_X1 port map( A => n1269, ZN => n1613);
   U427 : INV_X1 port map( A => n944, ZN => n1911);
   U501 : INV_X1 port map( A => n997, ZN => n1875);
   U327 : INV_X1 port map( A => n892, ZN => n1959);
   U111 : INV_X1 port map( A => n780, ZN => n2064);
   U844 : INV_X1 port map( A => n1169, ZN => n1709);
   U431 : INV_X1 port map( A => n946, ZN => n1909);
   U385 : INV_X1 port map( A => n922, ZN => n1931);
   U628 : INV_X1 port map( A => n1060, ZN => n1814);
   U893 : INV_X1 port map( A => n1193, ZN => n1686);
   U185 : INV_X1 port map( A => n819, ZN => n2028);
   U299 : INV_X1 port map( A => n878, ZN => n1973);
   U704 : INV_X1 port map( A => n1099, ZN => n1777);
   U311 : INV_X1 port map( A => n884, ZN => n1967);
   U1048 : INV_X1 port map( A => n1270, ZN => n1612);
   U563 : INV_X1 port map( A => n1028, ZN => n1845);
   U301 : INV_X1 port map( A => n879, ZN => n1972);
   U325 : INV_X1 port map( A => n891, ZN => n1960);
   U838 : INV_X1 port map( A => n1166, ZN => n1712);
   U891 : INV_X1 port map( A => n1192, ZN => n1687);
   U367 : INV_X1 port map( A => n913, ZN => n1940);
   U109 : INV_X1 port map( A => n779, ZN => n2065);
   U634 : INV_X1 port map( A => n1063, ZN => n1811);
   U505 : INV_X1 port map( A => n999, ZN => n1873);
   U567 : INV_X1 port map( A => n1030, ZN => n1843);
   U565 : INV_X1 port map( A => n1029, ZN => n1844);
   U802 : INV_X1 port map( A => n1148, ZN => n1729);
   U1494 : INV_X1 port map( A => n2180, ZN => n1539);
   U273 : INV_X1 port map( A => n864, ZN => n1985);
   U471 : INV_X1 port map( A => n966, ZN => n1889);
   U221 : INV_X1 port map( A => n838, ZN => n2011);
   U141 : INV_X1 port map( A => n795, ZN => n2049);
   U537 : INV_X1 port map( A => n1015, ZN => n1857);
   U736 : INV_X1 port map( A => n1115, ZN => n1761);
   U207 : INV_X1 port map( A => n830, ZN => n2017);
   U1002 : INV_X1 port map( A => n1248, ZN => n1633);
   U889 : INV_X1 port map( A => n1191, ZN => n1688);
   U935 : INV_X1 port map( A => n1214, ZN => n1665);
   U1070 : INV_X1 port map( A => n1281, ZN => n1601);
   U603 : INV_X1 port map( A => n1048, ZN => n1825);
   U868 : INV_X1 port map( A => n1181, ZN => n1697);
   U339 : INV_X1 port map( A => n898, ZN => n1953);
   U670 : INV_X1 port map( A => n1081, ZN => n1793);
   U950 : INV_X1 port map( A => n1222, ZN => n1659);
   U952 : INV_X1 port map( A => n1223, ZN => n1658);
   U1018 : INV_X1 port map( A => n1255, ZN => n1627);
   U684 : INV_X1 port map( A => n1089, ZN => n1787);
   U85 : INV_X1 port map( A => n767, ZN => n2077);
   U1131 : INV_X1 port map( A => n1328, ZN => n1591);
   U754 : INV_X1 port map( A => n1124, ZN => n1753);
   U1020 : INV_X1 port map( A => n1256, ZN => n1626);
   U287 : INV_X1 port map( A => n872, ZN => n1979);
   U686 : INV_X1 port map( A => n1090, ZN => n1786);
   U91 : INV_X1 port map( A => n770, ZN => n2074);
   U1022 : INV_X1 port map( A => n1257, ZN => n1625);
   U750 : INV_X1 port map( A => n1122, ZN => n1755);
   U159 : INV_X1 port map( A => n806, ZN => n2041);
   U1144 : INV_X1 port map( A => n1339, ZN => n1589);
   U157 : INV_X1 port map( A => n805, ZN => n2042);
   U155 : INV_X1 port map( A => n804, ZN => n2043);
   U752 : INV_X1 port map( A => n1123, ZN => n1754);
   U289 : INV_X1 port map( A => n873, ZN => n1978);
   U225 : INV_X1 port map( A => n840, ZN => n2009);
   U816 : INV_X1 port map( A => n1155, ZN => n1723);
   U223 : INV_X1 port map( A => n839, ZN => n2010);
   U291 : INV_X1 port map( A => n874, ZN => n1977);
   U89 : INV_X1 port map( A => n769, ZN => n2075);
   U555 : INV_X1 port map( A => n1024, ZN => n1849);
   U885 : INV_X1 port map( A => n1189, ZN => n1690);
   U883 : INV_X1 port map( A => n1188, ZN => n1691);
   U553 : INV_X1 port map( A => n1023, ZN => n1850);
   U551 : INV_X1 port map( A => n1022, ZN => n1851);
   U419 : INV_X1 port map( A => n940, ZN => n1915);
   U421 : INV_X1 port map( A => n941, ZN => n1914);
   U423 : INV_X1 port map( A => n942, ZN => n1913);
   U485 : INV_X1 port map( A => n973, ZN => n1883);
   U487 : INV_X1 port map( A => n990, ZN => n1882);
   U489 : INV_X1 port map( A => n991, ZN => n1881);
   U618 : INV_X1 port map( A => n1055, ZN => n1819);
   U353 : INV_X1 port map( A => n906, ZN => n1947);
   U818 : INV_X1 port map( A => n1156, ZN => n1722);
   U620 : INV_X1 port map( A => n1056, ZN => n1818);
   U820 : INV_X1 port map( A => n1157, ZN => n1721);
   U622 : INV_X1 port map( A => n1057, ZN => n1817);
   U355 : INV_X1 port map( A => n907, ZN => n1946);
   U357 : INV_X1 port map( A => n908, ZN => n1945);
   U359 : INV_X1 port map( A => n909, ZN => n1944);
   U491 : INV_X1 port map( A => n992, ZN => n1880);
   U624 : INV_X1 port map( A => n1058, ZN => n1816);
   U481 : INV_X1 port map( A => n971, ZN => n1885);
   U1105 : INV_X1 port map( A => n1306, ZN => n1595);
   U149 : INV_X1 port map( A => n801, ZN => n2046);
   U217 : INV_X1 port map( A => n836, ZN => n2013);
   U946 : INV_X1 port map( A => n1220, ZN => n1661);
   U479 : INV_X1 port map( A => n970, ZN => n1886);
   U1012 : INV_X1 port map( A => n1252, ZN => n1630);
   U215 : INV_X1 port map( A => n835, ZN => n2014);
   U293 : INV_X1 port map( A => n875, ZN => n1976);
   U690 : INV_X1 port map( A => n1092, ZN => n1784);
   U944 : INV_X1 port map( A => n1219, ZN => n1662);
   U746 : INV_X1 port map( A => n1120, ZN => n1757);
   U1024 : INV_X1 port map( A => n1258, ZN => n1624);
   U93 : INV_X1 port map( A => n771, ZN => n2073);
   U413 : INV_X1 port map( A => n937, ZN => n1918);
   U756 : INV_X1 port map( A => n1125, ZN => n1752);
   U744 : INV_X1 port map( A => n1119, ZN => n1758);
   U283 : INV_X1 port map( A => n870, ZN => n1981);
   U1092 : INV_X1 port map( A => n1295, ZN => n1597);
   U415 : INV_X1 port map( A => n938, ZN => n1917);
   U227 : INV_X1 port map( A => n841, ZN => n2008);
   U822 : INV_X1 port map( A => n1158, ZN => n1720);
   U425 : INV_X1 port map( A => n943, ZN => n1912);
   U557 : INV_X1 port map( A => n1025, ZN => n1848);
   U349 : INV_X1 port map( A => n904, ZN => n1949);
   U151 : INV_X1 port map( A => n802, ZN => n2045);
   U688 : INV_X1 port map( A => n1091, ZN => n1785);
   U678 : INV_X1 port map( A => n1086, ZN => n1790);
   U161 : INV_X1 port map( A => n807, ZN => n2040);
   U1158 : INV_X1 port map( A => n1350, ZN => n1587);
   U281 : INV_X1 port map( A => n869, ZN => n1982);
   U1014 : INV_X1 port map( A => n1253, ZN => n1629);
   U612 : INV_X1 port map( A => n1052, ZN => n1822);
   U956 : INV_X1 port map( A => n1225, ZN => n1656);
   U877 : INV_X1 port map( A => n1185, ZN => n1694);
   U810 : INV_X1 port map( A => n1152, ZN => n1726);
   U95 : INV_X1 port map( A => n772, ZN => n2072);
   U812 : INV_X1 port map( A => n1153, ZN => n1725);
   U610 : INV_X1 port map( A => n1050, ZN => n1823);
   U545 : INV_X1 port map( A => n1019, ZN => n1854);
   U1172 : INV_X1 port map( A => n1361, ZN => n1585);
   U680 : INV_X1 port map( A => n1087, ZN => n1789);
   U347 : INV_X1 port map( A => n903, ZN => n1950);
   U547 : INV_X1 port map( A => n1020, ZN => n1853);
   U887 : INV_X1 port map( A => n1190, ZN => n1689);
   U614 : INV_X1 port map( A => n1053, ZN => n1821);
   U954 : INV_X1 port map( A => n1224, ZN => n1657);
   U879 : INV_X1 port map( A => n1186, ZN => n1693);
   U83 : INV_X1 port map( A => n766, ZN => n2078);
   U814 : INV_X1 port map( A => n1154, ZN => n1724);
   U1016 : INV_X1 port map( A => n1254, ZN => n1628);
   U279 : INV_X1 port map( A => n867, ZN => n1983);
   U345 : INV_X1 port map( A => n901, ZN => n1951);
   U1010 : INV_X1 port map( A => n1250, ZN => n1631);
   U81 : INV_X1 port map( A => n764, ZN => n2079);
   U616 : INV_X1 port map( A => n1054, ZN => n1820);
   U942 : INV_X1 port map( A => n1217, ZN => n1663);
   U682 : INV_X1 port map( A => n1088, ZN => n1788);
   U543 : INV_X1 port map( A => n1017, ZN => n1855);
   U1078 : INV_X1 port map( A => n1283, ZN => n1599);
   U417 : INV_X1 port map( A => n939, ZN => n1916);
   U881 : INV_X1 port map( A => n1187, ZN => n1692);
   U1118 : INV_X1 port map( A => n1317, ZN => n1593);
   U808 : INV_X1 port map( A => n1150, ZN => n1727);
   U748 : INV_X1 port map( A => n1121, ZN => n1756);
   U483 : INV_X1 port map( A => n972, ZN => n1884);
   U411 : INV_X1 port map( A => n935, ZN => n1919);
   U153 : INV_X1 port map( A => n803, ZN => n2044);
   U213 : INV_X1 port map( A => n833, ZN => n2015);
   U351 : INV_X1 port map( A => n905, ZN => n1948);
   U875 : INV_X1 port map( A => n1183, ZN => n1695);
   U742 : INV_X1 port map( A => n1117, ZN => n1759);
   U87 : INV_X1 port map( A => n768, ZN => n2076);
   U948 : INV_X1 port map( A => n1221, ZN => n1660);
   U549 : INV_X1 port map( A => n1021, ZN => n1852);
   U147 : INV_X1 port map( A => n799, ZN => n2047);
   U676 : INV_X1 port map( A => n1084, ZN => n1791);
   U219 : INV_X1 port map( A => n837, ZN => n2012);
   U477 : INV_X1 port map( A => n968, ZN => n1887);
   U285 : INV_X1 port map( A => n871, ZN => n1980);
   U35 : BUF_X1 port map( A => target_PC_i(23), Z => n643);
   U37 : BUF_X1 port map( A => target_PC_i(21), Z => n642);
   U39 : CLKBUF_X1 port map( A => target_PC_i(29), Z => n634);
   U41 : BUF_X1 port map( A => target_PC_i(25), Z => n636);
   U43 : BUF_X1 port map( A => target_PC_i(3), Z => n652);
   U45 : BUF_X1 port map( A => target_PC_i(2), Z => n650);
   U47 : BUF_X1 port map( A => target_PC_i(13), Z => n651);
   U49 : INV_X1 port map( A => stall_i, ZN => n2286);
   U51 : AND2_X1 port map( A1 => n2224, A2 => n8, ZN => n714);
   U53 : BUF_X1 port map( A => target_PC_i(31), Z => n647);
   U55 : AND2_X1 port map( A1 => n9, A2 => n2222, ZN => n717);
   U57 : BUF_X1 port map( A => target_PC_i(24), Z => n635);
   U59 : BUF_X1 port map( A => target_PC_i(27), Z => n653);
   U61 : BUF_X1 port map( A => target_PC_i(1), Z => n633);
   U63 : AND2_X1 port map( A1 => target_PC_i(6), A2 => n618, ZN => n720);
   U65 : BUF_X1 port map( A => target_PC_i(4), Z => n641);
   U69 : BUF_X1 port map( A => target_PC_i(8), Z => n639);
   U70 : BUF_X1 port map( A => target_PC_i(12), Z => n646);
   U82 : BUF_X1 port map( A => target_PC_i(0), Z => n648);
   U84 : INV_X1 port map( A => n765, ZN => n2268);
   U86 : INV_X1 port map( A => n1184, ZN => n734);
   U88 : INV_X1 port map( A => n800, ZN => n2264);
   U90 : INV_X1 port map( A => n868, ZN => n2259);
   U96 : INV_X1 port map( A => n1284, ZN => n726);
   U126 : INV_X1 port map( A => n1018, ZN => n987);
   U130 : INV_X1 port map( A => n1051, ZN => n984);
   U144 : INV_X1 port map( A => n1085, ZN => n982);
   U145 : INV_X1 port map( A => n902, ZN => n2256);
   U146 : INV_X1 port map( A => n902, ZN => n2254);
   U148 : INV_X1 port map( A => n765, ZN => n2266);
   U150 : INV_X1 port map( A => n969, ZN => n2214);
   U152 : INV_X1 port map( A => n834, ZN => n2260);
   U154 : INV_X1 port map( A => n1151, ZN => n976);
   U156 : INV_X1 port map( A => n902, ZN => n2255);
   U162 : INV_X1 port map( A => n969, ZN => n2213);
   U192 : INV_X1 port map( A => n1284, ZN => n727);
   U196 : INV_X1 port map( A => n834, ZN => n2262);
   U210 : INV_X1 port map( A => n868, ZN => n2258);
   U211 : INV_X1 port map( A => n1184, ZN => n735);
   U212 : INV_X1 port map( A => n1118, ZN => n977);
   U214 : INV_X1 port map( A => n1151, ZN => n974);
   U216 : INV_X1 port map( A => n1251, ZN => n728);
   U218 : INV_X1 port map( A => n1218, ZN => n732);
   U220 : INV_X1 port map( A => n1251, ZN => n730);
   U222 : INV_X1 port map( A => n1018, ZN => n988);
   U228 : INV_X1 port map( A => n800, ZN => n2263);
   U258 : INV_X1 port map( A => n765, ZN => n2267);
   U262 : INV_X1 port map( A => n1085, ZN => n980);
   U276 : INV_X1 port map( A => n1051, ZN => n985);
   U277 : INV_X1 port map( A => n1284, ZN => n725);
   U278 : INV_X1 port map( A => n834, ZN => n2261);
   U280 : INV_X1 port map( A => n1085, ZN => n981);
   U282 : INV_X1 port map( A => n1118, ZN => n979);
   U284 : INV_X1 port map( A => n1118, ZN => n978);
   U286 : INV_X1 port map( A => n969, ZN => n989);
   U288 : INV_X1 port map( A => n1184, ZN => n737);
   U294 : INV_X1 port map( A => n936, ZN => n2216);
   U324 : INV_X1 port map( A => n936, ZN => n2215);
   U328 : INV_X1 port map( A => n868, ZN => n2257);
   U342 : INV_X1 port map( A => n936, ZN => n2253);
   U343 : INV_X1 port map( A => n1218, ZN => n733);
   U344 : INV_X1 port map( A => n1251, ZN => n729);
   U346 : INV_X1 port map( A => n1051, ZN => n983);
   U348 : INV_X1 port map( A => n1151, ZN => n975);
   U350 : INV_X1 port map( A => n1018, ZN => n986);
   U352 : INV_X1 port map( A => n800, ZN => n2265);
   U354 : INV_X1 port map( A => n1218, ZN => n731);
   U360 : OR2_X2 port map( A1 => n1216, A2 => n866, ZN => n1251);
   U390 : OR2_X2 port map( A1 => n900, A2 => n1083, ZN => n1151);
   U394 : OR2_X2 port map( A1 => n832, A2 => n934, ZN => n936);
   U408 : OR2_X2 port map( A1 => n866, A2 => n1083, ZN => n1118);
   U409 : OR2_X2 port map( A1 => n866, A2 => n798, ZN => n834);
   U410 : OR2_X2 port map( A1 => n900, A2 => n1216, ZN => n1284);
   U412 : OR2_X2 port map( A1 => n866, A2 => n934, ZN => n969);
   U414 : OR2_X2 port map( A1 => n832, A2 => n1083, ZN => n1085);
   U416 : OR2_X2 port map( A1 => n900, A2 => n798, ZN => n868);
   U418 : OR2_X2 port map( A1 => n1216, A2 => n797, ZN => n1184);
   U420 : OR2_X2 port map( A1 => n797, A2 => n934, ZN => n902);
   U426 : OR2_X2 port map( A1 => n797, A2 => n1083, ZN => n1051);
   U456 : OR2_X2 port map( A1 => n900, A2 => n934, ZN => n1018);
   U460 : OR2_X2 port map( A1 => n1216, A2 => n832, ZN => n1218);
   U474 : OR2_X2 port map( A1 => n832, A2 => n798, ZN => n800);
   U475 : OR2_X2 port map( A1 => n797, A2 => n798, ZN => n765);
   U476 : INV_X2 port map( A => stall_i, ZN => n2285);
   U478 : BUF_X2 port map( A => n762, Z => n2270);
   U480 : BUF_X2 port map( A => n746, Z => n2282);
   U482 : BUF_X2 port map( A => n745, Z => n2283);
   U484 : BUF_X2 port map( A => n744, Z => n2284);
   U486 : BUF_X2 port map( A => n751, Z => n2277);
   U492 : BUF_X2 port map( A => n760, Z => n2272);
   U522 : BUF_X2 port map( A => n749, Z => n2279);
   U526 : BUF_X2 port map( A => n750, Z => n2278);
   U540 : BUF_X2 port map( A => n748, Z => n2280);
   U541 : BUF_X2 port map( A => n763, Z => n2269);
   U542 : BUF_X2 port map( A => n756, Z => n2276);
   U544 : BUF_X2 port map( A => n758, Z => n2274);
   U546 : BUF_X2 port map( A => n757, Z => n2275);
   U548 : BUF_X2 port map( A => n759, Z => n2273);
   U550 : BUF_X2 port map( A => n761, Z => n2271);
   U552 : INV_X1 port map( A => reset, ZN => n2291);
   U558 : INV_X1 port map( A => reset, ZN => n2293);
   U588 : INV_X1 port map( A => reset, ZN => n2310);
   U592 : INV_X1 port map( A => reset, ZN => n2296);
   U606 : INV_X1 port map( A => reset, ZN => n2290);
   U607 : INV_X1 port map( A => reset, ZN => n2302);
   U608 : INV_X1 port map( A => reset, ZN => n2307);
   U609 : INV_X1 port map( A => reset, ZN => n2304);
   U611 : INV_X1 port map( A => reset, ZN => n2289);
   U613 : INV_X1 port map( A => reset, ZN => n2288);
   U615 : INV_X1 port map( A => reset, ZN => n2309);
   U617 : INV_X1 port map( A => reset, ZN => n2297);
   U619 : INV_X1 port map( A => reset, ZN => n2299);
   U625 : INV_X1 port map( A => reset, ZN => n2306);
   U655 : INV_X1 port map( A => reset, ZN => n2295);
   U659 : INV_X1 port map( A => reset, ZN => n2308);
   U673 : INV_X1 port map( A => reset, ZN => n2298);
   U674 : INV_X1 port map( A => reset, ZN => n2294);
   U675 : INV_X1 port map( A => reset, ZN => n2303);
   U677 : INV_X1 port map( A => reset, ZN => n2301);
   U679 : INV_X1 port map( A => reset, ZN => n2300);
   U681 : INV_X1 port map( A => reset, ZN => n2292);
   U683 : INV_X1 port map( A => reset, ZN => n2305);
   U685 : INV_X1 port map( A => reset, ZN => n2311);
   U691 : BUF_X1 port map( A => target_PC_i(14), Z => n630);
   U721 : BUF_X1 port map( A => target_PC_i(19), Z => n645);
   U725 : BUF_X1 port map( A => target_PC_i(17), Z => n631);
   U739 : BUF_X1 port map( A => target_PC_i(22), Z => n632);
   U740 : BUF_X1 port map( A => target_PC_i(16), Z => n637);
   U741 : BUF_X1 port map( A => target_PC_i(20), Z => n638);
   U743 : BUF_X1 port map( A => target_PC_i(26), Z => n649);
   U745 : BUF_X1 port map( A => target_PC_i(10), Z => n640);
   U747 : AND2_X1 port map( A1 => target_PC_i(24), A2 => n600, ZN => n719);
   U749 : AND2_X1 port map( A1 => n7, A2 => n2225, ZN => n715);
   U751 : BUF_X2 port map( A => target_PC_i(11), Z => n644);
   U757 : AND2_X1 port map( A1 => n623, A2 => target_PC_i(1), ZN => n723);
   U787 : AND2_X1 port map( A1 => target_PC_i(31), A2 => n593, ZN => n718);
   U791 : AND4_X1 port map( A1 => n655, A2 => n654, A3 => n656, A4 => n657, ZN 
                           => n2211);
   U805 : AND4_X1 port map( A1 => n2247, A2 => n2246, A3 => n2248, A4 => n2245,
                           ZN => n654);
   U806 : AND4_X1 port map( A1 => n2238, A2 => n2239, A3 => n2237, A4 => n2240,
                           ZN => n655);
   U807 : AND4_X1 port map( A1 => n2232, A2 => n2229, A3 => n2231, A4 => n2230,
                           ZN => n656);
   U809 : AND4_X1 port map( A1 => n2219, A2 => n2218, A3 => n2220, A4 => n2217,
                           ZN => n657);
   U811 : INV_X1 port map( A => n724, ZN => n2210);
   U813 : AND2_X1 port map( A1 => target_PC_i(0), A2 => n624, ZN => n722);
   U815 : INV_X1 port map( A => target_PC_i(29), ZN => n2225);
   U817 : CLKBUF_X1 port map( A => target_PC_i(30), Z => n658);
   U823 : AND2_X1 port map( A1 => n2221, A2 => n6, ZN => n716);
   U853 : INV_X1 port map( A => target_PC_i(27), ZN => n2222);
   U857 : CLKBUF_X1 port map( A => target_PC_i(28), Z => n659);
   U871 : CLKBUF_X1 port map( A => mispredict_o_port, Z => n724);
   U872 : INV_X1 port map( A => target_PC_i(30), ZN => n2221);
   U873 : AND2_X1 port map( A1 => n617, A2 => target_PC_i(7), ZN => n721);
   U874 : INV_X1 port map( A => target_PC_i(28), ZN => n2224);
   U876 : AOI21_X1 port map( B1 => n2211, B2 => n663, A => n2212, ZN => 
                           mispredict_o_port);
   U878 : AOI21_X1 port map( B1 => n738, B2 => n739, A => reset, ZN => 
                           taken_o_port);
   U880 : BUF_X1 port map( A => stall_i, Z => n2287);
   U882 : BUF_X1 port map( A => n747, Z => n2281);
   U884 : AOI221_X1 port map( B1 => target_PC_i(10), B2 => n614, C1 => n613, C2
                           => n644, A => n2249, ZN => n2248);
   U890 : AOI221_X1 port map( B1 => target_PC_i(8), B2 => n616, C1 => 
                           target_PC_i(9), C2 => n615, A => n2250, ZN => n2247)
                           ;
   U920 : AOI221_X1 port map( B1 => target_PC_i(14), B2 => n610, C1 => n609, C2
                           => target_PC_i(15), A => n2251, ZN => n2246);
   U924 : NOR2_X1 port map( A1 => n2200, A2 => n2199, ZN => n746);
   U938 : NOR2_X1 port map( A1 => n2202, A2 => n2199, ZN => n744);
   U939 : NOR2_X1 port map( A1 => n2200, A2 => n2208, ZN => n757);
   U940 : NOR2_X1 port map( A1 => n2200, A2 => n2203, ZN => n751);
   U943 : NOR2_X1 port map( A1 => n2209, A2 => n2200, ZN => n763);
   U945 : NOR2_X1 port map( A1 => n2202, A2 => n2208, ZN => n759);
   U947 : NOR2_X1 port map( A1 => n2202, A2 => n2203, ZN => n749);
   U949 : NOR2_X1 port map( A1 => n2201, A2 => n2199, ZN => n745);
   U951 : OAI22_X1 port map( A1 => target_PC_i(16), A2 => n608, B1 => 
                           target_PC_i(17), B2 => n607, ZN => n2228);
   U957 : OAI22_X1 port map( A1 => target_PC_i(18), A2 => n606, B1 => 
                           target_PC_i(19), B2 => n605, ZN => n2227);
   U987 : OAI22_X1 port map( A1 => n2224, A2 => n8, B1 => n2225, B2 => n7, ZN 
                           => n2226);
   U991 : OAI22_X1 port map( A1 => n2221, A2 => n6, B1 => n2222, B2 => n9, ZN 
                           => n2223);
   U1005 : OAI22_X1 port map( A1 => target_PC_i(22), A2 => n602, B1 => 
                           target_PC_i(23), B2 => n601, ZN => n2233);
   U1006 : OAI22_X1 port map( A1 => target_PC_i(20), A2 => n604, B1 => 
                           target_PC_i(21), B2 => n603, ZN => n2234);
   U1007 : OAI22_X1 port map( A1 => target_PC_i(25), A2 => n599, B1 => 
                           target_PC_i(26), B2 => n598, ZN => n2235);
   U1009 : OAI22_X1 port map( A1 => target_PC_i(31), A2 => n593, B1 => 
                           target_PC_i(24), B2 => n600, ZN => n2236);
   U1011 : OAI22_X1 port map( A1 => target_PC_i(2), A2 => n622, B1 => 
                           target_PC_i(3), B2 => n621, ZN => n2241);
   U1013 : OAI22_X1 port map( A1 => target_PC_i(0), A2 => n624, B1 => 
                           target_PC_i(1), B2 => n623, ZN => n2242);
   U1015 : OAI22_X1 port map( A1 => target_PC_i(6), A2 => n618, B1 => 
                           target_PC_i(7), B2 => n617, ZN => n2243);
   U1017 : OAI22_X1 port map( A1 => target_PC_i(4), A2 => n620, B1 => 
                           target_PC_i(5), B2 => n619, ZN => n2244);
   U1019 : OAI22_X1 port map( A1 => target_PC_i(10), A2 => n614, B1 => 
                           target_PC_i(11), B2 => n613, ZN => n2249);
   U1025 : OAI22_X1 port map( A1 => target_PC_i(8), A2 => n616, B1 => 
                           target_PC_i(9), B2 => n615, ZN => n2250);
   U1055 : OAI22_X1 port map( A1 => target_PC_i(14), A2 => n610, B1 => 
                           target_PC_i(15), B2 => n609, ZN => n2251);
   U1059 : OAI22_X1 port map( A1 => target_PC_i(12), A2 => n612, B1 => 
                           target_PC_i(13), B2 => n611, ZN => n2252);
   U1073 : AOI221_X1 port map( B1 => target_PC_i(16), B2 => n608, C1 => n607, 
                           C2 => target_PC_i(17), A => n2228, ZN => n2217);
   U1074 : AOI221_X1 port map( B1 => target_PC_i(18), B2 => n606, C1 => n605, 
                           C2 => target_PC_i(19), A => n2227, ZN => n2218);
   U1075 : NOR3_X1 port map( A1 => n2226, A2 => n715, A3 => n714, ZN => n2219);
   U1077 : NOR3_X1 port map( A1 => n2223, A2 => n717, A3 => n716, ZN => n2220);
   U1079 : AOI221_X1 port map( B1 => target_PC_i(22), B2 => n602, C1 => 
                           target_PC_i(23), C2 => n601, A => n2233, ZN => n2232
                           );
   U1093 : AOI221_X1 port map( B1 => target_PC_i(20), B2 => n604, C1 => 
                           target_PC_i(21), C2 => n603, A => n2234, ZN => n2231
                           );
   U1106 : AOI221_X1 port map( B1 => target_PC_i(25), B2 => n599, C1 => n598, 
                           C2 => target_PC_i(26), A => n2235, ZN => n2230);
   U1119 : NOR3_X1 port map( A1 => n718, A2 => n719, A3 => n2236, ZN => n2229);
   U1132 : AOI221_X1 port map( B1 => target_PC_i(2), B2 => n622, C1 => n621, C2
                           => target_PC_i(3), A => n2241, ZN => n2240);
   U1173 : NOR3_X1 port map( A1 => n722, A2 => n723, A3 => n2242, ZN => n2239);
   U1383 : NOR3_X1 port map( A1 => n721, A2 => n720, A3 => n2243, ZN => n2238);
   U1411 : AOI221_X1 port map( B1 => target_PC_i(4), B2 => n620, C1 => n619, C2
                           => target_PC_i(5), A => n2244, ZN => n2237);
   U1509 : AOI221_X1 port map( B1 => target_PC_i(12), B2 => n612, C1 => n611, 
                           C2 => target_PC_i(13), A => n2252, ZN => n2245);
   U1510 : OAI22_X1 port map( A1 => n1284, A2 => n647, B1 => 
                           predict_PC_15_31_port, B2 => n727, ZN => n1283);
   U1511 : OAI22_X1 port map( A1 => n1251, A2 => n647, B1 => 
                           predict_PC_14_31_port, B2 => n730, ZN => n1250);
   U1518 : OAI22_X1 port map( A1 => n969, A2 => n647, B1 => 
                           predict_PC_6_31_port, B2 => n2214, ZN => n968);
   U1520 : OAI22_X1 port map( A1 => n1118, A2 => n647, B1 => 
                           predict_PC_10_31_port, B2 => n979, ZN => n1117);
   U1521 : OAI22_X1 port map( A1 => n834, A2 => n647, B1 => 
                           predict_PC_2_31_port, B2 => n2262, ZN => n833);
   U1524 : OAI22_X1 port map( A1 => n765, A2 => n647, B1 => 
                           predict_PC_0_31_port, B2 => n2268, ZN => n764);
   U1527 : OAI22_X1 port map( A1 => n800, A2 => n647, B1 => 
                           predict_PC_1_31_port, B2 => n2265, ZN => n799);
   U1533 : OAI22_X1 port map( A1 => n868, A2 => n647, B1 => 
                           predict_PC_3_31_port, B2 => n2259, ZN => n867);
   U1536 : OAI22_X1 port map( A1 => n936, A2 => n647, B1 => 
                           predict_PC_5_31_port, B2 => n2253, ZN => n935);
   U1541 : OAI22_X1 port map( A1 => n1018, A2 => n647, B1 => 
                           predict_PC_7_31_port, B2 => n988, ZN => n1017);
   U1554 : OAI22_X1 port map( A1 => n1051, A2 => target_PC_i(31), B1 => 
                           predict_PC_8_31_port, B2 => n985, ZN => n1050);
   U1555 : OAI22_X1 port map( A1 => n1085, A2 => n647, B1 => 
                           predict_PC_9_31_port, B2 => n982, ZN => n1084);
   U1556 : OAI22_X1 port map( A1 => n1218, A2 => n647, B1 => 
                           predict_PC_13_31_port, B2 => n733, ZN => n1217);
   U1558 : OAI22_X1 port map( A1 => n1151, A2 => n647, B1 => 
                           predict_PC_11_31_port, B2 => n976, ZN => n1150);
   U1559 : OAI22_X1 port map( A1 => n902, A2 => n647, B1 => 
                           predict_PC_4_31_port, B2 => n2256, ZN => n901);
   U1560 : OAI22_X1 port map( A1 => n1184, A2 => n647, B1 => 
                           predict_PC_12_31_port, B2 => n737, ZN => n1183);
   U1561 : OAI22_X1 port map( A1 => n765, A2 => n648, B1 => predict_PC_0_0_port
                           , B2 => n2266, ZN => n796);
   U1562 : OAI22_X1 port map( A1 => n800, A2 => n648, B1 => predict_PC_1_0_port
                           , B2 => n2263, ZN => n831);
   U1563 : OAI22_X1 port map( A1 => n834, A2 => n648, B1 => predict_PC_2_0_port
                           , B2 => n2260, ZN => n865);
   U1564 : OAI22_X1 port map( A1 => n868, A2 => n648, B1 => predict_PC_3_0_port
                           , B2 => n2257, ZN => n899);
   U1565 : OAI22_X1 port map( A1 => n902, A2 => n648, B1 => predict_PC_4_0_port
                           , B2 => n2254, ZN => n933);
   U1566 : OAI22_X1 port map( A1 => n936, A2 => n648, B1 => predict_PC_5_0_port
                           , B2 => n2215, ZN => n967);
   U1567 : OAI22_X1 port map( A1 => n969, A2 => n648, B1 => predict_PC_6_0_port
                           , B2 => n989, ZN => n1016);
   U1568 : OAI22_X1 port map( A1 => n1018, A2 => n648, B1 => 
                           predict_PC_7_0_port, B2 => n986, ZN => n1049);
   U1569 : OAI22_X1 port map( A1 => n1051, A2 => n648, B1 => 
                           predict_PC_8_0_port, B2 => n983, ZN => n1082);
   U1570 : OAI22_X1 port map( A1 => n1085, A2 => n648, B1 => 
                           predict_PC_9_0_port, B2 => n980, ZN => n1116);
   U1571 : OAI22_X1 port map( A1 => n1118, A2 => target_PC_i(0), B1 => 
                           predict_PC_10_0_port, B2 => n977, ZN => n1149);
   U1572 : OAI22_X1 port map( A1 => n1151, A2 => n648, B1 => 
                           predict_PC_11_0_port, B2 => n974, ZN => n1182);
   U1573 : OAI22_X1 port map( A1 => n1184, A2 => n648, B1 => 
                           predict_PC_12_0_port, B2 => n734, ZN => n1215);
   U1574 : OAI22_X1 port map( A1 => n1218, A2 => n648, B1 => 
                           predict_PC_13_0_port, B2 => n731, ZN => n1249);
   U1575 : OAI22_X1 port map( A1 => n1251, A2 => target_PC_i(0), B1 => 
                           predict_PC_14_0_port, B2 => n728, ZN => n1282);
   U1576 : OAI22_X1 port map( A1 => n1284, A2 => target_PC_i(0), B1 => 
                           predict_PC_15_0_port, B2 => n725, ZN => n2191);
   U1577 : OAI22_X1 port map( A1 => n765, A2 => target_PC_i(9), B1 => 
                           predict_PC_0_9_port, B2 => n2266, ZN => n787);
   U1578 : OAI22_X1 port map( A1 => n1018, A2 => target_PC_i(9), B1 => 
                           predict_PC_7_9_port, B2 => n986, ZN => n1040);
   U1579 : OAI22_X1 port map( A1 => n1251, A2 => target_PC_i(9), B1 => 
                           predict_PC_14_9_port, B2 => n728, ZN => n1273);
   U1580 : OAI22_X1 port map( A1 => n1051, A2 => target_PC_i(9), B1 => 
                           predict_PC_8_9_port, B2 => n983, ZN => n1073);
   U1581 : OAI22_X1 port map( A1 => n1085, A2 => target_PC_i(9), B1 => 
                           predict_PC_9_9_port, B2 => n980, ZN => n1107);
   U1582 : OAI22_X1 port map( A1 => n1118, A2 => target_PC_i(9), B1 => 
                           predict_PC_10_9_port, B2 => n977, ZN => n1140);
   U1583 : OAI22_X1 port map( A1 => n1151, A2 => target_PC_i(9), B1 => 
                           predict_PC_11_9_port, B2 => n974, ZN => n1173);
   U1584 : OAI22_X1 port map( A1 => n1184, A2 => target_PC_i(9), B1 => 
                           predict_PC_12_9_port, B2 => n734, ZN => n1206);
   U1585 : OAI22_X1 port map( A1 => n1218, A2 => target_PC_i(9), B1 => 
                           predict_PC_13_9_port, B2 => n731, ZN => n1240);
   U1586 : OAI22_X1 port map( A1 => n1284, A2 => target_PC_i(9), B1 => 
                           predict_PC_15_9_port, B2 => n725, ZN => n1526);
   U1587 : OAI22_X1 port map( A1 => n969, A2 => target_PC_i(9), B1 => 
                           predict_PC_6_9_port, B2 => n989, ZN => n1007);
   U1588 : OAI22_X1 port map( A1 => n800, A2 => target_PC_i(9), B1 => 
                           predict_PC_1_9_port, B2 => n2263, ZN => n822);
   U1589 : OAI22_X1 port map( A1 => n834, A2 => target_PC_i(9), B1 => 
                           predict_PC_2_9_port, B2 => n2260, ZN => n856);
   U1590 : OAI22_X1 port map( A1 => n868, A2 => target_PC_i(9), B1 => 
                           predict_PC_3_9_port, B2 => n2257, ZN => n890);
   U1591 : OAI22_X1 port map( A1 => n902, A2 => target_PC_i(9), B1 => 
                           predict_PC_4_9_port, B2 => n2254, ZN => n924);
   U1592 : OAI22_X1 port map( A1 => n936, A2 => target_PC_i(9), B1 => 
                           predict_PC_5_9_port, B2 => n2215, ZN => n958);
   U1593 : OAI22_X1 port map( A1 => n1284, A2 => target_PC_i(7), B1 => 
                           predict_PC_15_7_port, B2 => n725, ZN => n2114);
   U1594 : OAI22_X1 port map( A1 => n1251, A2 => target_PC_i(7), B1 => 
                           predict_PC_14_7_port, B2 => n728, ZN => n1275);
   U1595 : OAI22_X1 port map( A1 => n1218, A2 => target_PC_i(7), B1 => 
                           predict_PC_13_7_port, B2 => n731, ZN => n1242);
   U1596 : OAI22_X1 port map( A1 => n1184, A2 => target_PC_i(7), B1 => 
                           predict_PC_12_7_port, B2 => n734, ZN => n1208);
   U1597 : OAI22_X1 port map( A1 => n1151, A2 => target_PC_i(7), B1 => 
                           predict_PC_11_7_port, B2 => n974, ZN => n1175);
   U1598 : OAI22_X1 port map( A1 => n1118, A2 => target_PC_i(7), B1 => 
                           predict_PC_10_7_port, B2 => n977, ZN => n1142);
   U1599 : OAI22_X1 port map( A1 => n1085, A2 => target_PC_i(7), B1 => 
                           predict_PC_9_7_port, B2 => n980, ZN => n1109);
   U1608 : OAI22_X1 port map( A1 => n1051, A2 => target_PC_i(7), B1 => 
                           predict_PC_8_7_port, B2 => n983, ZN => n1075);
   U1609 : OAI22_X1 port map( A1 => n1018, A2 => target_PC_i(7), B1 => 
                           predict_PC_7_7_port, B2 => n986, ZN => n1042);
   U1610 : OAI22_X1 port map( A1 => n969, A2 => target_PC_i(7), B1 => 
                           predict_PC_6_7_port, B2 => n989, ZN => n1009);
   U1611 : OAI22_X1 port map( A1 => n936, A2 => target_PC_i(7), B1 => 
                           predict_PC_5_7_port, B2 => n2215, ZN => n960);
   U1612 : OAI22_X1 port map( A1 => n902, A2 => target_PC_i(7), B1 => 
                           predict_PC_4_7_port, B2 => n2254, ZN => n926);
   U1613 : OAI22_X1 port map( A1 => n868, A2 => target_PC_i(7), B1 => 
                           predict_PC_3_7_port, B2 => n2257, ZN => n892);
   U1614 : OAI22_X1 port map( A1 => n834, A2 => target_PC_i(7), B1 => 
                           predict_PC_2_7_port, B2 => n2260, ZN => n858);
   U1615 : OAI22_X1 port map( A1 => n800, A2 => target_PC_i(7), B1 => 
                           predict_PC_1_7_port, B2 => n2263, ZN => n824);
   U1616 : OAI22_X1 port map( A1 => n765, A2 => target_PC_i(7), B1 => 
                           predict_PC_0_7_port, B2 => n2266, ZN => n789);
   U1617 : OAI22_X1 port map( A1 => n1284, A2 => n635, B1 => 
                           predict_PC_15_24_port, B2 => n727, ZN => n1361);
   U1618 : OAI22_X1 port map( A1 => n1251, A2 => n635, B1 => 
                           predict_PC_14_24_port, B2 => n730, ZN => n1258);
   U1619 : OAI22_X1 port map( A1 => n1218, A2 => n635, B1 => 
                           predict_PC_13_24_port, B2 => n733, ZN => n1225);
   U1620 : OAI22_X1 port map( A1 => n1184, A2 => target_PC_i(24), B1 => 
                           predict_PC_12_24_port, B2 => n737, ZN => n1191);
   U1621 : OAI22_X1 port map( A1 => n1151, A2 => n635, B1 => 
                           predict_PC_11_24_port, B2 => n976, ZN => n1158);
   U1622 : OAI22_X1 port map( A1 => n1118, A2 => n635, B1 => 
                           predict_PC_10_24_port, B2 => n979, ZN => n1125);
   U1623 : OAI22_X1 port map( A1 => n1085, A2 => n635, B1 => 
                           predict_PC_9_24_port, B2 => n982, ZN => n1092);
   U1624 : OAI22_X1 port map( A1 => n1051, A2 => n635, B1 => 
                           predict_PC_8_24_port, B2 => n985, ZN => n1058);
   U1625 : OAI22_X1 port map( A1 => n1018, A2 => n635, B1 => 
                           predict_PC_7_24_port, B2 => n988, ZN => n1025);
   U1626 : OAI22_X1 port map( A1 => n969, A2 => n635, B1 => 
                           predict_PC_6_24_port, B2 => n2214, ZN => n992);
   U1627 : OAI22_X1 port map( A1 => n936, A2 => n635, B1 => 
                           predict_PC_5_24_port, B2 => n2253, ZN => n943);
   U1628 : OAI22_X1 port map( A1 => n902, A2 => n635, B1 => 
                           predict_PC_4_24_port, B2 => n2256, ZN => n909);
   U1629 : OAI22_X1 port map( A1 => n868, A2 => n635, B1 => 
                           predict_PC_3_24_port, B2 => n2259, ZN => n875);
   U1630 : OAI22_X1 port map( A1 => n834, A2 => n635, B1 => 
                           predict_PC_2_24_port, B2 => n2262, ZN => n841);
   U1631 : OAI22_X1 port map( A1 => n800, A2 => n635, B1 => 
                           predict_PC_1_24_port, B2 => n2265, ZN => n807);
   U1632 : OAI22_X1 port map( A1 => n765, A2 => n635, B1 => 
                           predict_PC_0_24_port, B2 => n2268, ZN => n772);
   U1633 : OAI22_X1 port map( A1 => n1284, A2 => n653, B1 => 
                           predict_PC_15_27_port, B2 => n727, ZN => n1328);
   U1634 : OAI22_X1 port map( A1 => n765, A2 => n653, B1 => 
                           predict_PC_0_27_port, B2 => n2268, ZN => n769);
   U1635 : OAI22_X1 port map( A1 => n800, A2 => n653, B1 => 
                           predict_PC_1_27_port, B2 => n2265, ZN => n804);
   U1636 : OAI22_X1 port map( A1 => n1251, A2 => n653, B1 => 
                           predict_PC_14_27_port, B2 => n730, ZN => n1255);
   U1637 : OAI22_X1 port map( A1 => n868, A2 => n653, B1 => 
                           predict_PC_3_27_port, B2 => n2259, ZN => n872);
   U1638 : OAI22_X1 port map( A1 => n1218, A2 => n653, B1 => 
                           predict_PC_13_27_port, B2 => n733, ZN => n1222);
   U1639 : OAI22_X1 port map( A1 => n969, A2 => n653, B1 => 
                           predict_PC_6_27_port, B2 => n2214, ZN => n973);
   U1640 : OAI22_X1 port map( A1 => n936, A2 => n653, B1 => 
                           predict_PC_5_27_port, B2 => n2253, ZN => n940);
   U1641 : OAI22_X1 port map( A1 => n1018, A2 => n653, B1 => 
                           predict_PC_7_27_port, B2 => n988, ZN => n1022);
   U1642 : OAI22_X1 port map( A1 => n902, A2 => n653, B1 => 
                           predict_PC_4_27_port, B2 => n2256, ZN => n906);
   U1643 : OAI22_X1 port map( A1 => n1184, A2 => n653, B1 => 
                           predict_PC_12_27_port, B2 => n737, ZN => n1188);
   U1644 : OAI22_X1 port map( A1 => n834, A2 => target_PC_i(27), B1 => 
                           predict_PC_2_27_port, B2 => n2262, ZN => n838);
   U1645 : OAI22_X1 port map( A1 => n1151, A2 => n653, B1 => 
                           predict_PC_11_27_port, B2 => n976, ZN => n1155);
   U1646 : OAI22_X1 port map( A1 => n1118, A2 => n653, B1 => 
                           predict_PC_10_27_port, B2 => n979, ZN => n1122);
   U1647 : OAI22_X1 port map( A1 => n1085, A2 => n653, B1 => 
                           predict_PC_9_27_port, B2 => n982, ZN => n1089);
   U1648 : OAI22_X1 port map( A1 => n1051, A2 => n653, B1 => 
                           predict_PC_8_27_port, B2 => n985, ZN => n1055);
   U1649 : OAI22_X1 port map( A1 => n1284, A2 => n658, B1 => 
                           predict_PC_15_30_port, B2 => n727, ZN => n1295);
   U1650 : OAI22_X1 port map( A1 => n1184, A2 => n658, B1 => 
                           predict_PC_12_30_port, B2 => n737, ZN => n1185);
   U1651 : OAI22_X1 port map( A1 => n1151, A2 => n658, B1 => 
                           predict_PC_11_30_port, B2 => n976, ZN => n1152);
   U1652 : OAI22_X1 port map( A1 => n800, A2 => n658, B1 => 
                           predict_PC_1_30_port, B2 => n2265, ZN => n801);
   U1653 : OAI22_X1 port map( A1 => n902, A2 => n658, B1 => 
                           predict_PC_4_30_port, B2 => n2256, ZN => n903);
   U1654 : OAI22_X1 port map( A1 => n868, A2 => n658, B1 => 
                           predict_PC_3_30_port, B2 => n2259, ZN => n869);
   U1655 : OAI22_X1 port map( A1 => n834, A2 => n658, B1 => 
                           predict_PC_2_30_port, B2 => n2262, ZN => n835);
   U1656 : OAI22_X1 port map( A1 => n936, A2 => n658, B1 => 
                           predict_PC_5_30_port, B2 => n2253, ZN => n937);
   U1657 : OAI22_X1 port map( A1 => n969, A2 => n658, B1 => 
                           predict_PC_6_30_port, B2 => n2214, ZN => n970);
   U1658 : OAI22_X1 port map( A1 => n1018, A2 => n658, B1 => 
                           predict_PC_7_30_port, B2 => n988, ZN => n1019);
   U1659 : OAI22_X1 port map( A1 => n1118, A2 => n658, B1 => 
                           predict_PC_10_30_port, B2 => n979, ZN => n1119);
   U1660 : OAI22_X1 port map( A1 => n765, A2 => n658, B1 => 
                           predict_PC_0_30_port, B2 => n2268, ZN => n766);
   U1661 : OAI22_X1 port map( A1 => n1085, A2 => n658, B1 => 
                           predict_PC_9_30_port, B2 => n982, ZN => n1086);
   U1662 : OAI22_X1 port map( A1 => n1251, A2 => n658, B1 => 
                           predict_PC_14_30_port, B2 => n730, ZN => n1252);
   U1663 : OAI22_X1 port map( A1 => n1051, A2 => n658, B1 => 
                           predict_PC_8_30_port, B2 => n985, ZN => n1052);
   U1664 : OAI22_X1 port map( A1 => n1218, A2 => n658, B1 => 
                           predict_PC_13_30_port, B2 => n733, ZN => n1219);
   U1665 : OAI22_X1 port map( A1 => n1284, A2 => n659, B1 => 
                           predict_PC_15_28_port, B2 => n727, ZN => n1317);
   U1666 : OAI22_X1 port map( A1 => n1184, A2 => n659, B1 => 
                           predict_PC_12_28_port, B2 => n737, ZN => n1187);
   U1667 : OAI22_X1 port map( A1 => n800, A2 => n659, B1 => 
                           predict_PC_1_28_port, B2 => n2265, ZN => n803);
   U1668 : OAI22_X1 port map( A1 => n1151, A2 => n659, B1 => 
                           predict_PC_11_28_port, B2 => n976, ZN => n1154);
   U1669 : OAI22_X1 port map( A1 => n902, A2 => n659, B1 => 
                           predict_PC_4_28_port, B2 => n2256, ZN => n905);
   U1670 : OAI22_X1 port map( A1 => n868, A2 => n659, B1 => 
                           predict_PC_3_28_port, B2 => n2259, ZN => n871);
   U1671 : OAI22_X1 port map( A1 => n936, A2 => n659, B1 => 
                           predict_PC_5_28_port, B2 => n2253, ZN => n939);
   U1672 : OAI22_X1 port map( A1 => n969, A2 => n659, B1 => 
                           predict_PC_6_28_port, B2 => n2214, ZN => n972);
   U1673 : OAI22_X1 port map( A1 => n1018, A2 => n659, B1 => 
                           predict_PC_7_28_port, B2 => n988, ZN => n1021);
   U1674 : OAI22_X1 port map( A1 => n834, A2 => n659, B1 => 
                           predict_PC_2_28_port, B2 => n2262, ZN => n837);
   U1675 : OAI22_X1 port map( A1 => n1085, A2 => n659, B1 => 
                           predict_PC_9_28_port, B2 => n982, ZN => n1088);
   U1676 : OAI22_X1 port map( A1 => n1118, A2 => n659, B1 => 
                           predict_PC_10_28_port, B2 => n979, ZN => n1121);
   U1677 : OAI22_X1 port map( A1 => n765, A2 => n659, B1 => 
                           predict_PC_0_28_port, B2 => n2268, ZN => n768);
   U1678 : OAI22_X1 port map( A1 => n1251, A2 => n659, B1 => 
                           predict_PC_14_28_port, B2 => n730, ZN => n1254);
   U1679 : OAI22_X1 port map( A1 => n1218, A2 => n659, B1 => 
                           predict_PC_13_28_port, B2 => n733, ZN => n1221);
   U1680 : OAI22_X1 port map( A1 => n1051, A2 => n659, B1 => 
                           predict_PC_8_28_port, B2 => n985, ZN => n1054);
   U1681 : OAI22_X1 port map( A1 => n1284, A2 => n634, B1 => 
                           predict_PC_15_29_port, B2 => n727, ZN => n1306);
   U1682 : OAI22_X1 port map( A1 => n1184, A2 => n634, B1 => 
                           predict_PC_12_29_port, B2 => n737, ZN => n1186);
   U1683 : OAI22_X1 port map( A1 => n800, A2 => n634, B1 => 
                           predict_PC_1_29_port, B2 => n2265, ZN => n802);
   U1684 : OAI22_X1 port map( A1 => n1151, A2 => n634, B1 => 
                           predict_PC_11_29_port, B2 => n976, ZN => n1153);
   U1685 : OAI22_X1 port map( A1 => n902, A2 => n634, B1 => 
                           predict_PC_4_29_port, B2 => n2256, ZN => n904);
   U1686 : OAI22_X1 port map( A1 => n868, A2 => n634, B1 => 
                           predict_PC_3_29_port, B2 => n2259, ZN => n870);
   U1687 : OAI22_X1 port map( A1 => n936, A2 => n634, B1 => 
                           predict_PC_5_29_port, B2 => n2253, ZN => n938);
   U1688 : OAI22_X1 port map( A1 => n969, A2 => n634, B1 => 
                           predict_PC_6_29_port, B2 => n2214, ZN => n971);
   U1689 : OAI22_X1 port map( A1 => n1018, A2 => n634, B1 => 
                           predict_PC_7_29_port, B2 => n988, ZN => n1020);
   U1690 : OAI22_X1 port map( A1 => n834, A2 => n634, B1 => 
                           predict_PC_2_29_port, B2 => n2262, ZN => n836);
   U1691 : OAI22_X1 port map( A1 => n1085, A2 => n634, B1 => 
                           predict_PC_9_29_port, B2 => n982, ZN => n1087);
   U1692 : OAI22_X1 port map( A1 => n1118, A2 => n634, B1 => 
                           predict_PC_10_29_port, B2 => n979, ZN => n1120);
   U1693 : OAI22_X1 port map( A1 => n765, A2 => target_PC_i(29), B1 => 
                           predict_PC_0_29_port, B2 => n2268, ZN => n767);
   U1694 : OAI22_X1 port map( A1 => n1251, A2 => n634, B1 => 
                           predict_PC_14_29_port, B2 => n730, ZN => n1253);
   U1695 : OAI22_X1 port map( A1 => n1218, A2 => n634, B1 => 
                           predict_PC_13_29_port, B2 => n733, ZN => n1220);
   U1696 : OAI22_X1 port map( A1 => n1051, A2 => n634, B1 => 
                           predict_PC_8_29_port, B2 => n985, ZN => n1053);

end SYN_bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity fetch_block is

   port( branch_target_i, sum_addr_i, A_i, NPC4_i : in std_logic_vector (31 
         downto 0);  S_MUX_PC_BUS_i : in std_logic_vector (1 downto 0);  PC_o, 
         PC4_o, PC_BUS_pre_BTB : out std_logic_vector (31 downto 0);  stall_i, 
         take_prediction_i, mispredict_i : in std_logic;  predicted_PC : in 
         std_logic_vector (31 downto 0);  clk, rst : in std_logic);

end fetch_block;

architecture SYN_Struct of fetch_block is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component mux41_1
      port( IN0, IN1, IN2, IN3 : in std_logic_vector (31 downto 0);  CTRL : in 
            std_logic_vector (1 downto 0);  OUT1 : out std_logic_vector (31 
            downto 0));
   end component;
   
   component mux41_0
      port( IN0, IN1, IN2, IN3 : in std_logic_vector (31 downto 0);  CTRL : in 
            std_logic_vector (1 downto 0);  OUT1 : out std_logic_vector (31 
            downto 0));
   end component;
   
   component add4
      port( IN1 : in std_logic_vector (31 downto 0);  OUT1 : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component ff32_en_0
      port( D : in std_logic_vector (31 downto 0);  en, clk, rst : in std_logic
            ;  Q : out std_logic_vector (31 downto 0));
   end component;
   
   signal PC_o_31_port, PC_o_30_port, PC_o_29_port, PC_o_28_port, PC_o_27_port,
      PC_o_26_port, PC_o_25_port, PC_o_24_port, PC_o_23_port, PC_o_22_port, 
      PC_o_21_port, PC_o_20_port, PC_o_19_port, PC_o_18_port, PC_o_17_port, 
      PC_o_16_port, PC_o_15_port, PC_o_14_port, PC_o_13_port, PC_o_12_port, 
      PC_o_11_port, PC_o_10_port, PC_o_9_port, PC_o_8_port, PC_o_7_port, 
      PC_o_6_port, PC_o_5_port, PC_o_4_port, PC_o_3_port, PC_o_2_port, 
      PC_o_1_port, PC_o_0_port, PC4_o_31_port, PC4_o_30_port, PC4_o_29_port, 
      PC4_o_28_port, PC4_o_27_port, PC4_o_26_port, PC4_o_25_port, PC4_o_24_port
      , PC4_o_23_port, PC4_o_22_port, PC4_o_21_port, PC4_o_20_port, 
      PC4_o_19_port, PC4_o_18_port, PC4_o_17_port, PC4_o_16_port, PC4_o_15_port
      , PC4_o_14_port, PC4_o_13_port, PC4_o_12_port, PC4_o_11_port, 
      PC4_o_10_port, PC4_o_9_port, PC4_o_8_port, PC4_o_7_port, PC4_o_6_port, 
      PC4_o_5_port, PC4_o_4_port, PC4_o_3_port, PC4_o_2_port, PC4_o_1_port, 
      PC4_o_0_port, PC_BUS_pre_BTB_31_port, PC_BUS_pre_BTB_30_port, 
      PC_BUS_pre_BTB_29_port, PC_BUS_pre_BTB_28_port, PC_BUS_pre_BTB_27_port, 
      PC_BUS_pre_BTB_26_port, PC_BUS_pre_BTB_25_port, PC_BUS_pre_BTB_24_port, 
      PC_BUS_pre_BTB_23_port, PC_BUS_pre_BTB_22_port, PC_BUS_pre_BTB_21_port, 
      PC_BUS_pre_BTB_19_port, PC_BUS_pre_BTB_18_port, PC_BUS_pre_BTB_17_port, 
      PC_BUS_pre_BTB_15_port, PC_BUS_pre_BTB_14_port, PC_BUS_pre_BTB_13_port, 
      PC_BUS_pre_BTB_12_port, PC_BUS_pre_BTB_11_port, PC_BUS_pre_BTB_10_port, 
      PC_BUS_pre_BTB_9_port, PC_BUS_pre_BTB_7_port, PC_BUS_pre_BTB_6_port, 
      PC_BUS_pre_BTB_5_port, PC_BUS_pre_BTB_4_port, PC_BUS_pre_BTB_3_port, 
      PC_BUS_pre_BTB_2_port, PC_BUS_pre_BTB_1_port, PC_BUS_pre_BTB_0_port, 
      PC_BUS_31_port, PC_BUS_30_port, PC_BUS_29_port, PC_BUS_28_port, 
      PC_BUS_27_port, PC_BUS_26_port, PC_BUS_25_port, PC_BUS_24_port, 
      PC_BUS_23_port, PC_BUS_22_port, PC_BUS_21_port, PC_BUS_20_port, 
      PC_BUS_19_port, PC_BUS_18_port, PC_BUS_17_port, PC_BUS_16_port, 
      PC_BUS_15_port, PC_BUS_14_port, PC_BUS_13_port, PC_BUS_12_port, 
      PC_BUS_11_port, PC_BUS_10_port, PC_BUS_9_port, PC_BUS_8_port, 
      PC_BUS_7_port, PC_BUS_6_port, PC_BUS_5_port, PC_BUS_4_port, PC_BUS_3_port
      , PC_BUS_2_port, PC_BUS_1_port, PC_BUS_0_port, PC_BUS_pre_BTB_16_port, 
      PC_BUS_pre_BTB_20_port, PC_BUS_pre_BTB_8_port, n5 : std_logic;

begin
   PC_o <= ( PC_o_31_port, PC_o_30_port, PC_o_29_port, PC_o_28_port, 
      PC_o_27_port, PC_o_26_port, PC_o_25_port, PC_o_24_port, PC_o_23_port, 
      PC_o_22_port, PC_o_21_port, PC_o_20_port, PC_o_19_port, PC_o_18_port, 
      PC_o_17_port, PC_o_16_port, PC_o_15_port, PC_o_14_port, PC_o_13_port, 
      PC_o_12_port, PC_o_11_port, PC_o_10_port, PC_o_9_port, PC_o_8_port, 
      PC_o_7_port, PC_o_6_port, PC_o_5_port, PC_o_4_port, PC_o_3_port, 
      PC_o_2_port, PC_o_1_port, PC_o_0_port );
   PC4_o <= ( PC4_o_31_port, PC4_o_30_port, PC4_o_29_port, PC4_o_28_port, 
      PC4_o_27_port, PC4_o_26_port, PC4_o_25_port, PC4_o_24_port, PC4_o_23_port
      , PC4_o_22_port, PC4_o_21_port, PC4_o_20_port, PC4_o_19_port, 
      PC4_o_18_port, PC4_o_17_port, PC4_o_16_port, PC4_o_15_port, PC4_o_14_port
      , PC4_o_13_port, PC4_o_12_port, PC4_o_11_port, PC4_o_10_port, 
      PC4_o_9_port, PC4_o_8_port, PC4_o_7_port, PC4_o_6_port, PC4_o_5_port, 
      PC4_o_4_port, PC4_o_3_port, PC4_o_2_port, PC4_o_1_port, PC4_o_0_port );
   PC_BUS_pre_BTB <= ( PC_BUS_pre_BTB_31_port, PC_BUS_pre_BTB_30_port, 
      PC_BUS_pre_BTB_29_port, PC_BUS_pre_BTB_28_port, PC_BUS_pre_BTB_27_port, 
      PC_BUS_pre_BTB_26_port, PC_BUS_pre_BTB_25_port, PC_BUS_pre_BTB_24_port, 
      PC_BUS_pre_BTB_23_port, PC_BUS_pre_BTB_22_port, PC_BUS_pre_BTB_21_port, 
      PC_BUS_pre_BTB_20_port, PC_BUS_pre_BTB_19_port, PC_BUS_pre_BTB_18_port, 
      PC_BUS_pre_BTB_17_port, PC_BUS_pre_BTB_16_port, PC_BUS_pre_BTB_15_port, 
      PC_BUS_pre_BTB_14_port, PC_BUS_pre_BTB_13_port, PC_BUS_pre_BTB_12_port, 
      PC_BUS_pre_BTB_11_port, PC_BUS_pre_BTB_10_port, PC_BUS_pre_BTB_9_port, 
      PC_BUS_pre_BTB_8_port, PC_BUS_pre_BTB_7_port, PC_BUS_pre_BTB_6_port, 
      PC_BUS_pre_BTB_5_port, PC_BUS_pre_BTB_4_port, PC_BUS_pre_BTB_3_port, 
      PC_BUS_pre_BTB_2_port, PC_BUS_pre_BTB_1_port, PC_BUS_pre_BTB_0_port );
   
   PC : ff32_en_0 port map( D(31) => PC_BUS_31_port, D(30) => PC_BUS_30_port, 
                           D(29) => PC_BUS_29_port, D(28) => PC_BUS_28_port, 
                           D(27) => PC_BUS_27_port, D(26) => PC_BUS_26_port, 
                           D(25) => PC_BUS_25_port, D(24) => PC_BUS_24_port, 
                           D(23) => PC_BUS_23_port, D(22) => PC_BUS_22_port, 
                           D(21) => PC_BUS_21_port, D(20) => PC_BUS_20_port, 
                           D(19) => PC_BUS_19_port, D(18) => PC_BUS_18_port, 
                           D(17) => PC_BUS_17_port, D(16) => PC_BUS_16_port, 
                           D(15) => PC_BUS_15_port, D(14) => PC_BUS_14_port, 
                           D(13) => PC_BUS_13_port, D(12) => PC_BUS_12_port, 
                           D(11) => PC_BUS_11_port, D(10) => PC_BUS_10_port, 
                           D(9) => PC_BUS_9_port, D(8) => PC_BUS_8_port, D(7) 
                           => PC_BUS_7_port, D(6) => PC_BUS_6_port, D(5) => 
                           PC_BUS_5_port, D(4) => PC_BUS_4_port, D(3) => 
                           PC_BUS_3_port, D(2) => PC_BUS_2_port, D(1) => 
                           PC_BUS_1_port, D(0) => PC_BUS_0_port, en => n5, clk 
                           => clk, rst => rst, Q(31) => PC_o_31_port, Q(30) => 
                           PC_o_30_port, Q(29) => PC_o_29_port, Q(28) => 
                           PC_o_28_port, Q(27) => PC_o_27_port, Q(26) => 
                           PC_o_26_port, Q(25) => PC_o_25_port, Q(24) => 
                           PC_o_24_port, Q(23) => PC_o_23_port, Q(22) => 
                           PC_o_22_port, Q(21) => PC_o_21_port, Q(20) => 
                           PC_o_20_port, Q(19) => PC_o_19_port, Q(18) => 
                           PC_o_18_port, Q(17) => PC_o_17_port, Q(16) => 
                           PC_o_16_port, Q(15) => PC_o_15_port, Q(14) => 
                           PC_o_14_port, Q(13) => PC_o_13_port, Q(12) => 
                           PC_o_12_port, Q(11) => PC_o_11_port, Q(10) => 
                           PC_o_10_port, Q(9) => PC_o_9_port, Q(8) => 
                           PC_o_8_port, Q(7) => PC_o_7_port, Q(6) => 
                           PC_o_6_port, Q(5) => PC_o_5_port, Q(4) => 
                           PC_o_4_port, Q(3) => PC_o_3_port, Q(2) => 
                           PC_o_2_port, Q(1) => PC_o_1_port, Q(0) => 
                           PC_o_0_port);
   PCADD : add4 port map( IN1(31) => PC_o_31_port, IN1(30) => PC_o_30_port, 
                           IN1(29) => PC_o_29_port, IN1(28) => PC_o_28_port, 
                           IN1(27) => PC_o_27_port, IN1(26) => PC_o_26_port, 
                           IN1(25) => PC_o_25_port, IN1(24) => PC_o_24_port, 
                           IN1(23) => PC_o_23_port, IN1(22) => PC_o_22_port, 
                           IN1(21) => PC_o_21_port, IN1(20) => PC_o_20_port, 
                           IN1(19) => PC_o_19_port, IN1(18) => PC_o_18_port, 
                           IN1(17) => PC_o_17_port, IN1(16) => PC_o_16_port, 
                           IN1(15) => PC_o_15_port, IN1(14) => PC_o_14_port, 
                           IN1(13) => PC_o_13_port, IN1(12) => PC_o_12_port, 
                           IN1(11) => PC_o_11_port, IN1(10) => PC_o_10_port, 
                           IN1(9) => PC_o_9_port, IN1(8) => PC_o_8_port, IN1(7)
                           => PC_o_7_port, IN1(6) => PC_o_6_port, IN1(5) => 
                           PC_o_5_port, IN1(4) => PC_o_4_port, IN1(3) => 
                           PC_o_3_port, IN1(2) => PC_o_2_port, IN1(1) => 
                           PC_o_1_port, IN1(0) => PC_o_0_port, OUT1(31) => 
                           PC4_o_31_port, OUT1(30) => PC4_o_30_port, OUT1(29) 
                           => PC4_o_29_port, OUT1(28) => PC4_o_28_port, 
                           OUT1(27) => PC4_o_27_port, OUT1(26) => PC4_o_26_port
                           , OUT1(25) => PC4_o_25_port, OUT1(24) => 
                           PC4_o_24_port, OUT1(23) => PC4_o_23_port, OUT1(22) 
                           => PC4_o_22_port, OUT1(21) => PC4_o_21_port, 
                           OUT1(20) => PC4_o_20_port, OUT1(19) => PC4_o_19_port
                           , OUT1(18) => PC4_o_18_port, OUT1(17) => 
                           PC4_o_17_port, OUT1(16) => PC4_o_16_port, OUT1(15) 
                           => PC4_o_15_port, OUT1(14) => PC4_o_14_port, 
                           OUT1(13) => PC4_o_13_port, OUT1(12) => PC4_o_12_port
                           , OUT1(11) => PC4_o_11_port, OUT1(10) => 
                           PC4_o_10_port, OUT1(9) => PC4_o_9_port, OUT1(8) => 
                           PC4_o_8_port, OUT1(7) => PC4_o_7_port, OUT1(6) => 
                           PC4_o_6_port, OUT1(5) => PC4_o_5_port, OUT1(4) => 
                           PC4_o_4_port, OUT1(3) => PC4_o_3_port, OUT1(2) => 
                           PC4_o_2_port, OUT1(1) => PC4_o_1_port, OUT1(0) => 
                           PC4_o_0_port);
   MUXTARGET : mux41_0 port map( IN0(31) => NPC4_i(31), IN0(30) => NPC4_i(30), 
                           IN0(29) => NPC4_i(29), IN0(28) => NPC4_i(28), 
                           IN0(27) => NPC4_i(27), IN0(26) => NPC4_i(26), 
                           IN0(25) => NPC4_i(25), IN0(24) => NPC4_i(24), 
                           IN0(23) => NPC4_i(23), IN0(22) => NPC4_i(22), 
                           IN0(21) => NPC4_i(21), IN0(20) => NPC4_i(20), 
                           IN0(19) => NPC4_i(19), IN0(18) => NPC4_i(18), 
                           IN0(17) => NPC4_i(17), IN0(16) => NPC4_i(16), 
                           IN0(15) => NPC4_i(15), IN0(14) => NPC4_i(14), 
                           IN0(13) => NPC4_i(13), IN0(12) => NPC4_i(12), 
                           IN0(11) => NPC4_i(11), IN0(10) => NPC4_i(10), IN0(9)
                           => NPC4_i(9), IN0(8) => NPC4_i(8), IN0(7) => 
                           NPC4_i(7), IN0(6) => NPC4_i(6), IN0(5) => NPC4_i(5),
                           IN0(4) => NPC4_i(4), IN0(3) => NPC4_i(3), IN0(2) => 
                           NPC4_i(2), IN0(1) => NPC4_i(1), IN0(0) => NPC4_i(0),
                           IN1(31) => A_i(31), IN1(30) => A_i(30), IN1(29) => 
                           A_i(29), IN1(28) => A_i(28), IN1(27) => A_i(27), 
                           IN1(26) => A_i(26), IN1(25) => A_i(25), IN1(24) => 
                           A_i(24), IN1(23) => A_i(23), IN1(22) => A_i(22), 
                           IN1(21) => A_i(21), IN1(20) => A_i(20), IN1(19) => 
                           A_i(19), IN1(18) => A_i(18), IN1(17) => A_i(17), 
                           IN1(16) => A_i(16), IN1(15) => A_i(15), IN1(14) => 
                           A_i(14), IN1(13) => A_i(13), IN1(12) => A_i(12), 
                           IN1(11) => A_i(11), IN1(10) => A_i(10), IN1(9) => 
                           A_i(9), IN1(8) => A_i(8), IN1(7) => A_i(7), IN1(6) 
                           => A_i(6), IN1(5) => A_i(5), IN1(4) => A_i(4), 
                           IN1(3) => A_i(3), IN1(2) => A_i(2), IN1(1) => A_i(1)
                           , IN1(0) => A_i(0), IN2(31) => sum_addr_i(31), 
                           IN2(30) => sum_addr_i(30), IN2(29) => sum_addr_i(29)
                           , IN2(28) => sum_addr_i(28), IN2(27) => 
                           sum_addr_i(27), IN2(26) => sum_addr_i(26), IN2(25) 
                           => sum_addr_i(25), IN2(24) => sum_addr_i(24), 
                           IN2(23) => sum_addr_i(23), IN2(22) => sum_addr_i(22)
                           , IN2(21) => sum_addr_i(21), IN2(20) => 
                           sum_addr_i(20), IN2(19) => sum_addr_i(19), IN2(18) 
                           => sum_addr_i(18), IN2(17) => sum_addr_i(17), 
                           IN2(16) => sum_addr_i(16), IN2(15) => sum_addr_i(15)
                           , IN2(14) => sum_addr_i(14), IN2(13) => 
                           sum_addr_i(13), IN2(12) => sum_addr_i(12), IN2(11) 
                           => sum_addr_i(11), IN2(10) => sum_addr_i(10), IN2(9)
                           => sum_addr_i(9), IN2(8) => sum_addr_i(8), IN2(7) =>
                           sum_addr_i(7), IN2(6) => sum_addr_i(6), IN2(5) => 
                           sum_addr_i(5), IN2(4) => sum_addr_i(4), IN2(3) => 
                           sum_addr_i(3), IN2(2) => sum_addr_i(2), IN2(1) => 
                           sum_addr_i(1), IN2(0) => sum_addr_i(0), IN3(31) => 
                           branch_target_i(31), IN3(30) => branch_target_i(30),
                           IN3(29) => branch_target_i(29), IN3(28) => 
                           branch_target_i(28), IN3(27) => branch_target_i(27),
                           IN3(26) => branch_target_i(26), IN3(25) => 
                           branch_target_i(25), IN3(24) => branch_target_i(24),
                           IN3(23) => branch_target_i(23), IN3(22) => 
                           branch_target_i(22), IN3(21) => branch_target_i(21),
                           IN3(20) => branch_target_i(20), IN3(19) => 
                           branch_target_i(19), IN3(18) => branch_target_i(18),
                           IN3(17) => branch_target_i(17), IN3(16) => 
                           branch_target_i(16), IN3(15) => branch_target_i(15),
                           IN3(14) => branch_target_i(14), IN3(13) => 
                           branch_target_i(13), IN3(12) => branch_target_i(12),
                           IN3(11) => branch_target_i(11), IN3(10) => 
                           branch_target_i(10), IN3(9) => branch_target_i(9), 
                           IN3(8) => branch_target_i(8), IN3(7) => 
                           branch_target_i(7), IN3(6) => branch_target_i(6), 
                           IN3(5) => branch_target_i(5), IN3(4) => 
                           branch_target_i(4), IN3(3) => branch_target_i(3), 
                           IN3(2) => branch_target_i(2), IN3(1) => 
                           branch_target_i(1), IN3(0) => branch_target_i(0), 
                           CTRL(1) => S_MUX_PC_BUS_i(1), CTRL(0) => 
                           S_MUX_PC_BUS_i(0), OUT1(31) => 
                           PC_BUS_pre_BTB_31_port, OUT1(30) => 
                           PC_BUS_pre_BTB_30_port, OUT1(29) => 
                           PC_BUS_pre_BTB_29_port, OUT1(28) => 
                           PC_BUS_pre_BTB_28_port, OUT1(27) => 
                           PC_BUS_pre_BTB_27_port, OUT1(26) => 
                           PC_BUS_pre_BTB_26_port, OUT1(25) => 
                           PC_BUS_pre_BTB_25_port, OUT1(24) => 
                           PC_BUS_pre_BTB_24_port, OUT1(23) => 
                           PC_BUS_pre_BTB_23_port, OUT1(22) => 
                           PC_BUS_pre_BTB_22_port, OUT1(21) => 
                           PC_BUS_pre_BTB_21_port, OUT1(20) => 
                           PC_BUS_pre_BTB_20_port, OUT1(19) => 
                           PC_BUS_pre_BTB_19_port, OUT1(18) => 
                           PC_BUS_pre_BTB_18_port, OUT1(17) => 
                           PC_BUS_pre_BTB_17_port, OUT1(16) => 
                           PC_BUS_pre_BTB_16_port, OUT1(15) => 
                           PC_BUS_pre_BTB_15_port, OUT1(14) => 
                           PC_BUS_pre_BTB_14_port, OUT1(13) => 
                           PC_BUS_pre_BTB_13_port, OUT1(12) => 
                           PC_BUS_pre_BTB_12_port, OUT1(11) => 
                           PC_BUS_pre_BTB_11_port, OUT1(10) => 
                           PC_BUS_pre_BTB_10_port, OUT1(9) => 
                           PC_BUS_pre_BTB_9_port, OUT1(8) => 
                           PC_BUS_pre_BTB_8_port, OUT1(7) => 
                           PC_BUS_pre_BTB_7_port, OUT1(6) => 
                           PC_BUS_pre_BTB_6_port, OUT1(5) => 
                           PC_BUS_pre_BTB_5_port, OUT1(4) => 
                           PC_BUS_pre_BTB_4_port, OUT1(3) => 
                           PC_BUS_pre_BTB_3_port, OUT1(2) => 
                           PC_BUS_pre_BTB_2_port, OUT1(1) => 
                           PC_BUS_pre_BTB_1_port, OUT1(0) => 
                           PC_BUS_pre_BTB_0_port);
   MUXPREDICTION : mux41_1 port map( IN0(31) => PC4_o_31_port, IN0(30) => 
                           PC4_o_30_port, IN0(29) => PC4_o_29_port, IN0(28) => 
                           PC4_o_28_port, IN0(27) => PC4_o_27_port, IN0(26) => 
                           PC4_o_26_port, IN0(25) => PC4_o_25_port, IN0(24) => 
                           PC4_o_24_port, IN0(23) => PC4_o_23_port, IN0(22) => 
                           PC4_o_22_port, IN0(21) => PC4_o_21_port, IN0(20) => 
                           PC4_o_20_port, IN0(19) => PC4_o_19_port, IN0(18) => 
                           PC4_o_18_port, IN0(17) => PC4_o_17_port, IN0(16) => 
                           PC4_o_16_port, IN0(15) => PC4_o_15_port, IN0(14) => 
                           PC4_o_14_port, IN0(13) => PC4_o_13_port, IN0(12) => 
                           PC4_o_12_port, IN0(11) => PC4_o_11_port, IN0(10) => 
                           PC4_o_10_port, IN0(9) => PC4_o_9_port, IN0(8) => 
                           PC4_o_8_port, IN0(7) => PC4_o_7_port, IN0(6) => 
                           PC4_o_6_port, IN0(5) => PC4_o_5_port, IN0(4) => 
                           PC4_o_4_port, IN0(3) => PC4_o_3_port, IN0(2) => 
                           PC4_o_2_port, IN0(1) => PC4_o_1_port, IN0(0) => 
                           PC4_o_0_port, IN1(31) => predicted_PC(31), IN1(30) 
                           => predicted_PC(30), IN1(29) => predicted_PC(29), 
                           IN1(28) => predicted_PC(28), IN1(27) => 
                           predicted_PC(27), IN1(26) => predicted_PC(26), 
                           IN1(25) => predicted_PC(25), IN1(24) => 
                           predicted_PC(24), IN1(23) => predicted_PC(23), 
                           IN1(22) => predicted_PC(22), IN1(21) => 
                           predicted_PC(21), IN1(20) => predicted_PC(20), 
                           IN1(19) => predicted_PC(19), IN1(18) => 
                           predicted_PC(18), IN1(17) => predicted_PC(17), 
                           IN1(16) => predicted_PC(16), IN1(15) => 
                           predicted_PC(15), IN1(14) => predicted_PC(14), 
                           IN1(13) => predicted_PC(13), IN1(12) => 
                           predicted_PC(12), IN1(11) => predicted_PC(11), 
                           IN1(10) => predicted_PC(10), IN1(9) => 
                           predicted_PC(9), IN1(8) => predicted_PC(8), IN1(7) 
                           => predicted_PC(7), IN1(6) => predicted_PC(6), 
                           IN1(5) => predicted_PC(5), IN1(4) => predicted_PC(4)
                           , IN1(3) => predicted_PC(3), IN1(2) => 
                           predicted_PC(2), IN1(1) => predicted_PC(1), IN1(0) 
                           => predicted_PC(0), IN2(31) => 
                           PC_BUS_pre_BTB_31_port, IN2(30) => 
                           PC_BUS_pre_BTB_30_port, IN2(29) => 
                           PC_BUS_pre_BTB_29_port, IN2(28) => 
                           PC_BUS_pre_BTB_28_port, IN2(27) => 
                           PC_BUS_pre_BTB_27_port, IN2(26) => 
                           PC_BUS_pre_BTB_26_port, IN2(25) => 
                           PC_BUS_pre_BTB_25_port, IN2(24) => 
                           PC_BUS_pre_BTB_24_port, IN2(23) => 
                           PC_BUS_pre_BTB_23_port, IN2(22) => 
                           PC_BUS_pre_BTB_22_port, IN2(21) => 
                           PC_BUS_pre_BTB_21_port, IN2(20) => 
                           PC_BUS_pre_BTB_20_port, IN2(19) => 
                           PC_BUS_pre_BTB_19_port, IN2(18) => 
                           PC_BUS_pre_BTB_18_port, IN2(17) => 
                           PC_BUS_pre_BTB_17_port, IN2(16) => 
                           PC_BUS_pre_BTB_16_port, IN2(15) => 
                           PC_BUS_pre_BTB_15_port, IN2(14) => 
                           PC_BUS_pre_BTB_14_port, IN2(13) => 
                           PC_BUS_pre_BTB_13_port, IN2(12) => 
                           PC_BUS_pre_BTB_12_port, IN2(11) => 
                           PC_BUS_pre_BTB_11_port, IN2(10) => 
                           PC_BUS_pre_BTB_10_port, IN2(9) => 
                           PC_BUS_pre_BTB_9_port, IN2(8) => 
                           PC_BUS_pre_BTB_8_port, IN2(7) => 
                           PC_BUS_pre_BTB_7_port, IN2(6) => 
                           PC_BUS_pre_BTB_6_port, IN2(5) => 
                           PC_BUS_pre_BTB_5_port, IN2(4) => 
                           PC_BUS_pre_BTB_4_port, IN2(3) => 
                           PC_BUS_pre_BTB_3_port, IN2(2) => 
                           PC_BUS_pre_BTB_2_port, IN2(1) => 
                           PC_BUS_pre_BTB_1_port, IN2(0) => 
                           PC_BUS_pre_BTB_0_port, IN3(31) => 
                           PC_BUS_pre_BTB_31_port, IN3(30) => 
                           PC_BUS_pre_BTB_30_port, IN3(29) => 
                           PC_BUS_pre_BTB_29_port, IN3(28) => 
                           PC_BUS_pre_BTB_28_port, IN3(27) => 
                           PC_BUS_pre_BTB_27_port, IN3(26) => 
                           PC_BUS_pre_BTB_26_port, IN3(25) => 
                           PC_BUS_pre_BTB_25_port, IN3(24) => 
                           PC_BUS_pre_BTB_24_port, IN3(23) => 
                           PC_BUS_pre_BTB_23_port, IN3(22) => 
                           PC_BUS_pre_BTB_22_port, IN3(21) => 
                           PC_BUS_pre_BTB_21_port, IN3(20) => 
                           PC_BUS_pre_BTB_20_port, IN3(19) => 
                           PC_BUS_pre_BTB_19_port, IN3(18) => 
                           PC_BUS_pre_BTB_18_port, IN3(17) => 
                           PC_BUS_pre_BTB_17_port, IN3(16) => 
                           PC_BUS_pre_BTB_16_port, IN3(15) => 
                           PC_BUS_pre_BTB_15_port, IN3(14) => 
                           PC_BUS_pre_BTB_14_port, IN3(13) => 
                           PC_BUS_pre_BTB_13_port, IN3(12) => 
                           PC_BUS_pre_BTB_12_port, IN3(11) => 
                           PC_BUS_pre_BTB_11_port, IN3(10) => 
                           PC_BUS_pre_BTB_10_port, IN3(9) => 
                           PC_BUS_pre_BTB_9_port, IN3(8) => 
                           PC_BUS_pre_BTB_8_port, IN3(7) => 
                           PC_BUS_pre_BTB_7_port, IN3(6) => 
                           PC_BUS_pre_BTB_6_port, IN3(5) => 
                           PC_BUS_pre_BTB_5_port, IN3(4) => 
                           PC_BUS_pre_BTB_4_port, IN3(3) => 
                           PC_BUS_pre_BTB_3_port, IN3(2) => 
                           PC_BUS_pre_BTB_2_port, IN3(1) => 
                           PC_BUS_pre_BTB_1_port, IN3(0) => 
                           PC_BUS_pre_BTB_0_port, CTRL(1) => mispredict_i, 
                           CTRL(0) => take_prediction_i, OUT1(31) => 
                           PC_BUS_31_port, OUT1(30) => PC_BUS_30_port, OUT1(29)
                           => PC_BUS_29_port, OUT1(28) => PC_BUS_28_port, 
                           OUT1(27) => PC_BUS_27_port, OUT1(26) => 
                           PC_BUS_26_port, OUT1(25) => PC_BUS_25_port, OUT1(24)
                           => PC_BUS_24_port, OUT1(23) => PC_BUS_23_port, 
                           OUT1(22) => PC_BUS_22_port, OUT1(21) => 
                           PC_BUS_21_port, OUT1(20) => PC_BUS_20_port, OUT1(19)
                           => PC_BUS_19_port, OUT1(18) => PC_BUS_18_port, 
                           OUT1(17) => PC_BUS_17_port, OUT1(16) => 
                           PC_BUS_16_port, OUT1(15) => PC_BUS_15_port, OUT1(14)
                           => PC_BUS_14_port, OUT1(13) => PC_BUS_13_port, 
                           OUT1(12) => PC_BUS_12_port, OUT1(11) => 
                           PC_BUS_11_port, OUT1(10) => PC_BUS_10_port, OUT1(9) 
                           => PC_BUS_9_port, OUT1(8) => PC_BUS_8_port, OUT1(7) 
                           => PC_BUS_7_port, OUT1(6) => PC_BUS_6_port, OUT1(5) 
                           => PC_BUS_5_port, OUT1(4) => PC_BUS_4_port, OUT1(3) 
                           => PC_BUS_3_port, OUT1(2) => PC_BUS_2_port, OUT1(1) 
                           => PC_BUS_1_port, OUT1(0) => PC_BUS_0_port);
   U1 : INV_X1 port map( A => stall_i, ZN => n5);

end SYN_Struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity top_level is

   port( clock, rst : in std_logic;  IRAM_Addr_o : out std_logic_vector (31 
         downto 0);  IRAM_Dout_i : in std_logic_vector (31 downto 0);  
         DRAM_Enable_o, DRAM_WR_o : out std_logic;  DRAM_Din_o, DRAM_Addr_o : 
         out std_logic_vector (31 downto 0);  DRAM_Dout_i : in std_logic_vector
         (31 downto 0));

end top_level;

architecture SYN_arch of top_level is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component fw_logic
      port( D1_i, rAdec_i, D2_i, D3_i, rA_i, rB_i : in std_logic_vector (4 
            downto 0);  S_mem_W, S_wb_W, S_exe_W : in std_logic;  S_FWAdec, 
            S_FWA, S_FWB : out std_logic_vector (1 downto 0);  S_mem_LOAD_BAR :
            in std_logic);
   end component;
   
   component mem_block
      port( X_i, LOAD_i : in std_logic_vector (31 downto 0);  W_o : out 
            std_logic_vector (31 downto 0);  S_MUX_MEM_i_BAR : in std_logic);
   end component;
   
   component mem_regs
      port( W_i : in std_logic_vector (31 downto 0);  D3_i : in 
            std_logic_vector (4 downto 0);  W_o : out std_logic_vector (31 
            downto 0);  D3_o : out std_logic_vector (4 downto 0);  clk, rst : 
            in std_logic);
   end component;
   
   component execute_block
      port( IMM_i, A_i : in std_logic_vector (31 downto 0);  rB_i, rC_i : in 
            std_logic_vector (4 downto 0);  MUXED_B_i : in std_logic_vector (31
            downto 0);  S_MUX_ALUIN_i : in std_logic;  FW_X_i, FW_W_i : in 
            std_logic_vector (31 downto 0);  S_FW_A_i, S_FW_B_i : in 
            std_logic_vector (1 downto 0);  muxed_dest : out std_logic_vector 
            (4 downto 0);  muxed_B : out std_logic_vector (31 downto 0);  
            S_MUX_DEST_i : in std_logic_vector (1 downto 0);  OP : in 
            std_logic_vector (0 to 4);  ALUW_i : in std_logic_vector (12 downto
            0);  DOUT : out std_logic_vector (31 downto 0);  stall_o : out 
            std_logic;  Clock, Reset : in std_logic);
   end component;
   
   component execute_regs
      port( X_i, S_i : in std_logic_vector (31 downto 0);  D2_i : in 
            std_logic_vector (4 downto 0);  X_o, S_o : out std_logic_vector (31
            downto 0);  D2_o : out std_logic_vector (4 downto 0);  stall_i, clk
            , rst : in std_logic);
   end component;
   
   component decode_regs
      port( A_i, B_i : in std_logic_vector (31 downto 0);  rA_i, rB_i, rC_i : 
            in std_logic_vector (4 downto 0);  IMM_i : in std_logic_vector (31 
            downto 0);  ALUW_i : in std_logic_vector (12 downto 0);  A_o, B_o :
            out std_logic_vector (31 downto 0);  rA_o, rB_o, rC_o : out 
            std_logic_vector (4 downto 0);  IMM_o : out std_logic_vector (31 
            downto 0);  ALUW_o : out std_logic_vector (12 downto 0);  stall_i, 
            clk, rst : in std_logic);
   end component;
   
   component dlx_regfile
      port( Clk, Rst, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, 
            ADD_RD2 : in std_logic_vector (4 downto 0);  DATAIN : in 
            std_logic_vector (31 downto 0);  OUT1, OUT2 : out std_logic_vector 
            (31 downto 0));
   end component;
   
   component 
      dlx_cu_MICROCODE_MEM_SIZE64_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE13
      port( Clk, Rst : in std_logic;  IR_IN : in std_logic_vector (31 downto 0)
            ;  stall_exe_i, mispredict_i : in std_logic;  D1_i, D2_i : in 
            std_logic_vector (4 downto 0);  S1_LATCH_EN, S2_LATCH_EN, 
            S3_LATCH_EN : out std_logic;  S_MUX_PC_BUS : out std_logic_vector 
            (1 downto 0);  S_EXT, S_EXT_SIGN, S_EQ_NEQ : out std_logic;  
            S_MUX_DEST : out std_logic_vector (1 downto 0);  S_MUX_LINK, 
            S_MEM_W_R, S_MEM_EN, S_RF_W_wb, S_RF_W_mem, S_RF_W_exe, S_MUX_ALUIN
            , stall_exe_o, stall_dec_o, stall_fetch_o, stall_btb_o, 
            was_branch_o, was_jmp_o : out std_logic;  ALU_WORD_o : out 
            std_logic_vector (12 downto 0);  ALU_OPCODE : out std_logic_vector 
            (0 to 4);  S_MUX_MEM_BAR : out std_logic);
   end component;
   
   component jump_logic
      port( NPCF_i, IR_i, A_i : in std_logic_vector (31 downto 0);  A_o : out 
            std_logic_vector (31 downto 0);  rA_o, rB_o, rC_o : out 
            std_logic_vector (4 downto 0);  branch_target_o, sum_addr_o, 
            extended_imm : out std_logic_vector (31 downto 0);  taken_o : out 
            std_logic;  FW_X_i, FW_W_i : in std_logic_vector (31 downto 0);  
            S_FW_Adec_i : in std_logic_vector (1 downto 0);  S_EXT_i, 
            S_EXT_SIGN_i, S_MUX_LINK_i, S_EQ_NEQ_i : in std_logic);
   end component;
   
   component fetch_regs
      port( NPCF_i, IR_i : in std_logic_vector (31 downto 0);  NPCF_o, IR_o : 
            out std_logic_vector (31 downto 0);  stall_i, clk, rst : in 
            std_logic);
   end component;
   
   component btb_N_LINES4_SIZE32
      port( clock, reset, stall_i : in std_logic;  TAG_i : in std_logic_vector 
            (3 downto 0);  target_PC_i : in std_logic_vector (31 downto 0);  
            was_taken_i : in std_logic;  predicted_next_PC_o : out 
            std_logic_vector (31 downto 0);  taken_o, mispredict_o : out 
            std_logic);
   end component;
   
   component fetch_block
      port( branch_target_i, sum_addr_i, A_i, NPC4_i : in std_logic_vector (31 
            downto 0);  S_MUX_PC_BUS_i : in std_logic_vector (1 downto 0);  
            PC_o, PC4_o, PC_BUS_pre_BTB : out std_logic_vector (31 downto 0);  
            stall_i, take_prediction_i, mispredict_i : in std_logic;  
            predicted_PC : in std_logic_vector (31 downto 0);  clk, rst : in 
            std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, IRAM_Addr_o_31_port, 
      IRAM_Addr_o_30_port, IRAM_Addr_o_29_port, IRAM_Addr_o_28_port, 
      IRAM_Addr_o_27_port, IRAM_Addr_o_26_port, IRAM_Addr_o_25_port, 
      IRAM_Addr_o_24_port, IRAM_Addr_o_23_port, IRAM_Addr_o_22_port, 
      IRAM_Addr_o_21_port, IRAM_Addr_o_20_port, IRAM_Addr_o_19_port, 
      IRAM_Addr_o_18_port, IRAM_Addr_o_17_port, IRAM_Addr_o_16_port, 
      IRAM_Addr_o_15_port, IRAM_Addr_o_14_port, IRAM_Addr_o_13_port, 
      IRAM_Addr_o_12_port, IRAM_Addr_o_11_port, IRAM_Addr_o_10_port, 
      IRAM_Addr_o_9_port, IRAM_Addr_o_8_port, IRAM_Addr_o_7_port, 
      IRAM_Addr_o_6_port, IRAM_Addr_o_5_port, IRAM_Addr_o_4_port, 
      IRAM_Addr_o_3_port, IRAM_Addr_o_2_port, IRAM_Addr_o_1_port, 
      IRAM_Addr_o_0_port, DRAM_Addr_o_31_port, DRAM_Addr_o_30_port, 
      DRAM_Addr_o_29_port, DRAM_Addr_o_28_port, DRAM_Addr_o_27_port, 
      DRAM_Addr_o_26_port, DRAM_Addr_o_25_port, DRAM_Addr_o_24_port, 
      DRAM_Addr_o_23_port, DRAM_Addr_o_22_port, DRAM_Addr_o_21_port, 
      DRAM_Addr_o_20_port, DRAM_Addr_o_19_port, DRAM_Addr_o_18_port, 
      DRAM_Addr_o_17_port, DRAM_Addr_o_16_port, DRAM_Addr_o_15_port, 
      DRAM_Addr_o_14_port, DRAM_Addr_o_13_port, DRAM_Addr_o_12_port, 
      DRAM_Addr_o_11_port, DRAM_Addr_o_10_port, DRAM_Addr_o_9_port, 
      DRAM_Addr_o_8_port, DRAM_Addr_o_7_port, DRAM_Addr_o_6_port, 
      DRAM_Addr_o_5_port, DRAM_Addr_o_4_port, DRAM_Addr_o_3_port, 
      DRAM_Addr_o_2_port, DRAM_Addr_o_1_port, DRAM_Addr_o_0_port, 
      was_taken_from_jl, was_branch, was_jmp, was_taken, 
      dummy_branch_target_31_port, dummy_branch_target_30_port, 
      dummy_branch_target_29_port, dummy_branch_target_28_port, 
      dummy_branch_target_27_port, dummy_branch_target_26_port, 
      dummy_branch_target_25_port, dummy_branch_target_24_port, 
      dummy_branch_target_23_port, dummy_branch_target_22_port, 
      dummy_branch_target_21_port, dummy_branch_target_20_port, 
      dummy_branch_target_19_port, dummy_branch_target_18_port, 
      dummy_branch_target_17_port, dummy_branch_target_16_port, 
      dummy_branch_target_15_port, dummy_branch_target_14_port, 
      dummy_branch_target_13_port, dummy_branch_target_12_port, 
      dummy_branch_target_11_port, dummy_branch_target_10_port, 
      dummy_branch_target_9_port, dummy_branch_target_8_port, 
      dummy_branch_target_7_port, dummy_branch_target_6_port, 
      dummy_branch_target_5_port, dummy_branch_target_4_port, 
      dummy_branch_target_3_port, dummy_branch_target_2_port, 
      dummy_branch_target_1_port, dummy_branch_target_0_port, 
      dummy_sum_addr_31_port, dummy_sum_addr_30_port, dummy_sum_addr_29_port, 
      dummy_sum_addr_28_port, dummy_sum_addr_27_port, dummy_sum_addr_26_port, 
      dummy_sum_addr_25_port, dummy_sum_addr_24_port, dummy_sum_addr_23_port, 
      dummy_sum_addr_22_port, dummy_sum_addr_21_port, dummy_sum_addr_20_port, 
      dummy_sum_addr_19_port, dummy_sum_addr_18_port, dummy_sum_addr_17_port, 
      dummy_sum_addr_16_port, dummy_sum_addr_15_port, dummy_sum_addr_14_port, 
      dummy_sum_addr_13_port, dummy_sum_addr_12_port, dummy_sum_addr_11_port, 
      dummy_sum_addr_10_port, dummy_sum_addr_9_port, dummy_sum_addr_8_port, 
      dummy_sum_addr_7_port, dummy_sum_addr_6_port, dummy_sum_addr_5_port, 
      dummy_sum_addr_4_port, dummy_sum_addr_3_port, dummy_sum_addr_2_port, 
      dummy_sum_addr_1_port, dummy_sum_addr_0_port, dummy_A_31_port, 
      dummy_A_30_port, dummy_A_29_port, dummy_A_28_port, dummy_A_27_port, 
      dummy_A_26_port, dummy_A_25_port, dummy_A_24_port, dummy_A_23_port, 
      dummy_A_22_port, dummy_A_21_port, dummy_A_20_port, dummy_A_19_port, 
      dummy_A_18_port, dummy_A_17_port, dummy_A_16_port, dummy_A_15_port, 
      dummy_A_14_port, dummy_A_13_port, dummy_A_12_port, dummy_A_11_port, 
      dummy_A_10_port, dummy_A_9_port, dummy_A_8_port, dummy_A_7_port, 
      dummy_A_6_port, dummy_A_5_port, dummy_A_4_port, dummy_A_3_port, 
      dummy_A_2_port, dummy_A_1_port, dummy_A_0_port, NPCF_31_port, 
      NPCF_30_port, NPCF_29_port, NPCF_28_port, NPCF_27_port, NPCF_26_port, 
      NPCF_25_port, NPCF_24_port, NPCF_23_port, NPCF_22_port, NPCF_21_port, 
      NPCF_20_port, NPCF_19_port, NPCF_18_port, NPCF_17_port, NPCF_16_port, 
      NPCF_15_port, NPCF_14_port, NPCF_13_port, NPCF_12_port, NPCF_11_port, 
      NPCF_10_port, NPCF_9_port, NPCF_8_port, NPCF_7_port, NPCF_6_port, 
      NPCF_5_port, NPCF_4_port, NPCF_3_port, NPCF_2_port, NPCF_1_port, 
      NPCF_0_port, dummy_S_MUX_PC_BUS_1_port, dummy_S_MUX_PC_BUS_0_port, 
      PC4_31_port, PC4_30_port, PC4_29_port, PC4_28_port, PC4_27_port, 
      PC4_26_port, PC4_25_port, PC4_24_port, PC4_23_port, PC4_22_port, 
      PC4_21_port, PC4_20_port, PC4_19_port, PC4_18_port, PC4_17_port, 
      PC4_16_port, PC4_15_port, PC4_14_port, PC4_13_port, PC4_12_port, 
      PC4_11_port, PC4_10_port, PC4_9_port, PC4_8_port, PC4_7_port, PC4_6_port,
      PC4_5_port, PC4_4_port, PC4_3_port, PC4_2_port, PC4_1_port, PC4_0_port, 
      TARGET_PC_31_port, TARGET_PC_30_port, TARGET_PC_29_port, 
      TARGET_PC_28_port, TARGET_PC_27_port, TARGET_PC_26_port, 
      TARGET_PC_25_port, TARGET_PC_24_port, TARGET_PC_23_port, 
      TARGET_PC_22_port, TARGET_PC_21_port, TARGET_PC_19_port, 
      TARGET_PC_18_port, TARGET_PC_17_port, TARGET_PC_15_port, 
      TARGET_PC_14_port, TARGET_PC_13_port, TARGET_PC_12_port, 
      TARGET_PC_11_port, TARGET_PC_10_port, TARGET_PC_9_port, TARGET_PC_7_port,
      TARGET_PC_6_port, TARGET_PC_5_port, TARGET_PC_4_port, TARGET_PC_3_port, 
      TARGET_PC_2_port, TARGET_PC_1_port, TARGET_PC_0_port, mispredict, 
      take_prediction, predicted_PC_31_port, predicted_PC_30_port, 
      predicted_PC_29_port, predicted_PC_28_port, predicted_PC_27_port, 
      predicted_PC_26_port, predicted_PC_25_port, predicted_PC_24_port, 
      predicted_PC_23_port, predicted_PC_22_port, predicted_PC_21_port, 
      predicted_PC_20_port, predicted_PC_19_port, predicted_PC_18_port, 
      predicted_PC_17_port, predicted_PC_16_port, predicted_PC_15_port, 
      predicted_PC_14_port, predicted_PC_13_port, predicted_PC_12_port, 
      predicted_PC_11_port, predicted_PC_10_port, predicted_PC_9_port, 
      predicted_PC_8_port, predicted_PC_7_port, predicted_PC_6_port, 
      predicted_PC_5_port, predicted_PC_4_port, predicted_PC_3_port, 
      predicted_PC_2_port, predicted_PC_1_port, predicted_PC_0_port, IR_31_port
      , IR_30_port, IR_29_port, IR_28_port, IR_27_port, IR_26_port, IR_25_port,
      IR_24_port, IR_23_port, IR_22_port, IR_21_port, IR_20_port, IR_19_port, 
      IR_18_port, IR_17_port, IR_16_port, IR_15_port, IR_14_port, IR_13_port, 
      IR_12_port, IR_11_port, IR_10_port, IR_9_port, IR_8_port, IR_7_port, 
      IR_6_port, IR_5_port, IR_4_port, IR_3_port, IR_2_port, IR_1_port, 
      IR_0_port, AtoComp_31_port, AtoComp_30_port, AtoComp_29_port, 
      AtoComp_28_port, AtoComp_27_port, AtoComp_26_port, AtoComp_25_port, 
      AtoComp_24_port, AtoComp_23_port, AtoComp_22_port, AtoComp_21_port, 
      AtoComp_20_port, AtoComp_19_port, AtoComp_18_port, AtoComp_17_port, 
      AtoComp_16_port, AtoComp_15_port, AtoComp_14_port, AtoComp_13_port, 
      AtoComp_12_port, AtoComp_11_port, AtoComp_10_port, AtoComp_9_port, 
      AtoComp_8_port, AtoComp_7_port, AtoComp_6_port, AtoComp_5_port, 
      AtoComp_4_port, AtoComp_3_port, AtoComp_2_port, AtoComp_1_port, 
      AtoComp_0_port, rA2reg_4_port, rA2reg_3_port, rA2reg_2_port, 
      rA2reg_1_port, rA2reg_0_port, rB2reg_4_port, rB2reg_3_port, rB2reg_2_port
      , rB2reg_1_port, rB2reg_0_port, rC2reg_4_port, rC2reg_3_port, 
      rC2reg_2_port, rC2reg_1_port, rC2reg_0_port, help_IMM_31_port, 
      help_IMM_30_port, help_IMM_29_port, help_IMM_28_port, help_IMM_27_port, 
      help_IMM_26_port, help_IMM_25_port, help_IMM_24_port, help_IMM_23_port, 
      help_IMM_22_port, help_IMM_21_port, help_IMM_20_port, help_IMM_19_port, 
      help_IMM_18_port, help_IMM_17_port, help_IMM_16_port, help_IMM_15_port, 
      help_IMM_14_port, help_IMM_13_port, help_IMM_12_port, help_IMM_11_port, 
      help_IMM_10_port, help_IMM_9_port, help_IMM_8_port, help_IMM_7_port, 
      help_IMM_6_port, help_IMM_5_port, help_IMM_4_port, help_IMM_3_port, 
      help_IMM_2_port, help_IMM_1_port, help_IMM_0_port, wb2reg_31_port, 
      wb2reg_30_port, wb2reg_29_port, wb2reg_28_port, wb2reg_27_port, 
      wb2reg_26_port, wb2reg_25_port, wb2reg_24_port, wb2reg_23_port, 
      wb2reg_22_port, wb2reg_21_port, wb2reg_20_port, wb2reg_19_port, 
      wb2reg_18_port, wb2reg_17_port, wb2reg_16_port, wb2reg_15_port, 
      wb2reg_14_port, wb2reg_13_port, wb2reg_12_port, wb2reg_11_port, 
      wb2reg_10_port, wb2reg_9_port, wb2reg_8_port, wb2reg_7_port, 
      wb2reg_6_port, wb2reg_5_port, wb2reg_4_port, wb2reg_3_port, wb2reg_2_port
      , wb2reg_1_port, wb2reg_0_port, dummy_S_FWAdec_1_port, 
      dummy_S_FWAdec_0_port, dummy_S_EXT, dummy_S_EXT_SIGN, dummy_S_MUX_LINK, 
      dummy_S_EQ_NEQ, exe_stall_cu, muxed_dest2exe_4_port, 
      muxed_dest2exe_3_port, muxed_dest2exe_2_port, muxed_dest2exe_1_port, 
      muxed_dest2exe_0_port, D22D3_4_port, D22D3_3_port, D22D3_2_port, 
      D22D3_1_port, D22D3_0_port, dummy_S_MUX_DEST_1_port, 
      dummy_S_MUX_DEST_0_port, dummy_S_MUX_MEM, dummy_S_RF_W_wb, 
      dummy_S_RF_W_mem, dummy_S_MUX_ALUIN, stall_exe, ALUW_dec_12_port, 
      ALUW_dec_11_port, ALUW_dec_10_port, ALUW_dec_9_port, ALUW_dec_8_port, 
      ALUW_dec_7_port, ALUW_dec_6_port, ALUW_dec_5_port, ALUW_dec_4_port, 
      ALUW_dec_3_port, ALUW_dec_2_port, ALUW_dec_1_port, ALUW_dec_0_port, 
      W2wb_31_port, W2wb_30_port, W2wb_29_port, W2wb_28_port, W2wb_27_port, 
      W2wb_26_port, W2wb_25_port, W2wb_24_port, W2wb_23_port, W2wb_22_port, 
      W2wb_21_port, W2wb_20_port, W2wb_19_port, W2wb_18_port, W2wb_17_port, 
      W2wb_16_port, W2wb_15_port, W2wb_14_port, W2wb_13_port, W2wb_12_port, 
      W2wb_11_port, W2wb_10_port, W2wb_9_port, W2wb_8_port, W2wb_7_port, 
      W2wb_6_port, W2wb_5_port, W2wb_4_port, W2wb_3_port, W2wb_2_port, 
      W2wb_1_port, W2wb_0_port, dummy_B_31_port, dummy_B_30_port, 
      dummy_B_29_port, dummy_B_28_port, dummy_B_27_port, dummy_B_26_port, 
      dummy_B_25_port, dummy_B_24_port, dummy_B_23_port, dummy_B_22_port, 
      dummy_B_21_port, dummy_B_20_port, dummy_B_19_port, dummy_B_18_port, 
      dummy_B_17_port, dummy_B_16_port, dummy_B_15_port, dummy_B_14_port, 
      dummy_B_13_port, dummy_B_12_port, dummy_B_11_port, dummy_B_10_port, 
      dummy_B_9_port, dummy_B_8_port, dummy_B_7_port, dummy_B_6_port, 
      dummy_B_5_port, dummy_B_4_port, dummy_B_3_port, dummy_B_2_port, 
      dummy_B_1_port, dummy_B_0_port, A2exe_31_port, A2exe_30_port, 
      A2exe_29_port, A2exe_28_port, A2exe_27_port, A2exe_26_port, A2exe_25_port
      , A2exe_24_port, A2exe_23_port, A2exe_22_port, A2exe_21_port, 
      A2exe_20_port, A2exe_19_port, A2exe_18_port, A2exe_17_port, A2exe_16_port
      , A2exe_15_port, A2exe_14_port, A2exe_13_port, A2exe_12_port, 
      A2exe_11_port, A2exe_10_port, A2exe_9_port, A2exe_8_port, A2exe_7_port, 
      A2exe_6_port, A2exe_5_port, A2exe_4_port, A2exe_3_port, A2exe_2_port, 
      A2exe_1_port, A2exe_0_port, B2exe_31_port, B2exe_30_port, B2exe_29_port, 
      B2exe_28_port, B2exe_27_port, B2exe_26_port, B2exe_25_port, B2exe_24_port
      , B2exe_23_port, B2exe_22_port, B2exe_21_port, B2exe_20_port, 
      B2exe_19_port, B2exe_18_port, B2exe_17_port, B2exe_16_port, B2exe_15_port
      , B2exe_14_port, B2exe_13_port, B2exe_12_port, B2exe_11_port, 
      B2exe_10_port, B2exe_9_port, B2exe_8_port, B2exe_7_port, B2exe_6_port, 
      B2exe_5_port, B2exe_4_port, B2exe_3_port, B2exe_2_port, B2exe_1_port, 
      B2exe_0_port, rA2fw_4_port, rA2fw_3_port, rA2fw_2_port, rA2fw_1_port, 
      rA2fw_0_port, rB2mux_4_port, rB2mux_3_port, rB2mux_2_port, rB2mux_1_port,
      rB2mux_0_port, rC2mux_4_port, rC2mux_3_port, rC2mux_2_port, rC2mux_1_port
      , rC2mux_0_port, IMM2exe_31_port, IMM2exe_30_port, IMM2exe_29_port, 
      IMM2exe_28_port, IMM2exe_27_port, IMM2exe_26_port, IMM2exe_25_port, 
      IMM2exe_24_port, IMM2exe_23_port, IMM2exe_22_port, IMM2exe_21_port, 
      IMM2exe_20_port, IMM2exe_19_port, IMM2exe_18_port, IMM2exe_17_port, 
      IMM2exe_16_port, IMM2exe_15_port, IMM2exe_14_port, IMM2exe_13_port, 
      IMM2exe_12_port, IMM2exe_11_port, IMM2exe_10_port, IMM2exe_9_port, 
      IMM2exe_8_port, IMM2exe_7_port, IMM2exe_6_port, IMM2exe_5_port, 
      IMM2exe_4_port, IMM2exe_3_port, IMM2exe_2_port, IMM2exe_1_port, 
      IMM2exe_0_port, ALUW_12_port, ALUW_11_port, ALUW_10_port, ALUW_9_port, 
      ALUW_8_port, ALUW_7_port, ALUW_6_port, ALUW_5_port, ALUW_4_port, 
      ALUW_3_port, ALUW_2_port, ALUW_1_port, ALUW_0_port, X2mem_31_port, 
      X2mem_30_port, X2mem_29_port, X2mem_28_port, X2mem_27_port, X2mem_26_port
      , X2mem_25_port, X2mem_24_port, X2mem_23_port, X2mem_22_port, 
      X2mem_21_port, X2mem_20_port, X2mem_19_port, X2mem_18_port, X2mem_17_port
      , X2mem_16_port, X2mem_15_port, X2mem_14_port, X2mem_13_port, 
      X2mem_12_port, X2mem_11_port, X2mem_10_port, X2mem_9_port, X2mem_8_port, 
      X2mem_7_port, X2mem_6_port, X2mem_5_port, X2mem_4_port, X2mem_3_port, 
      X2mem_2_port, X2mem_1_port, X2mem_0_port, S2mem_31_port, S2mem_30_port, 
      S2mem_29_port, S2mem_28_port, S2mem_27_port, S2mem_26_port, S2mem_25_port
      , S2mem_24_port, S2mem_23_port, S2mem_22_port, S2mem_21_port, 
      S2mem_20_port, S2mem_19_port, S2mem_18_port, S2mem_17_port, S2mem_16_port
      , S2mem_15_port, S2mem_14_port, S2mem_13_port, S2mem_12_port, 
      S2mem_11_port, S2mem_10_port, S2mem_9_port, S2mem_8_port, S2mem_7_port, 
      S2mem_6_port, S2mem_5_port, S2mem_4_port, S2mem_2_port, S2mem_1_port, 
      dummy_S_FWA2exe_1_port, dummy_S_FWB2exe_1_port, dummy_S_FWB2exe_0_port, 
      D32reg_4_port, D32reg_3_port, D32reg_2_port, D32reg_1_port, D32reg_0_port
      , n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
      n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36
      , n37, n38, n39, n40, n41, n42, n43, n44, net684116, net684117, net684118
      , net684119, net684120, net684121, net684122, net684123, net684124 : 
      std_logic;

begin
   IRAM_Addr_o <= ( IRAM_Addr_o_31_port, IRAM_Addr_o_30_port, 
      IRAM_Addr_o_29_port, IRAM_Addr_o_28_port, IRAM_Addr_o_27_port, 
      IRAM_Addr_o_26_port, IRAM_Addr_o_25_port, IRAM_Addr_o_24_port, 
      IRAM_Addr_o_23_port, IRAM_Addr_o_22_port, IRAM_Addr_o_21_port, 
      IRAM_Addr_o_20_port, IRAM_Addr_o_19_port, IRAM_Addr_o_18_port, 
      IRAM_Addr_o_17_port, IRAM_Addr_o_16_port, IRAM_Addr_o_15_port, 
      IRAM_Addr_o_14_port, IRAM_Addr_o_13_port, IRAM_Addr_o_12_port, 
      IRAM_Addr_o_11_port, IRAM_Addr_o_10_port, IRAM_Addr_o_9_port, 
      IRAM_Addr_o_8_port, IRAM_Addr_o_7_port, IRAM_Addr_o_6_port, 
      IRAM_Addr_o_5_port, IRAM_Addr_o_4_port, IRAM_Addr_o_3_port, 
      IRAM_Addr_o_2_port, IRAM_Addr_o_1_port, IRAM_Addr_o_0_port );
   DRAM_Addr_o <= ( DRAM_Addr_o_31_port, DRAM_Addr_o_30_port, 
      DRAM_Addr_o_29_port, DRAM_Addr_o_28_port, DRAM_Addr_o_27_port, 
      DRAM_Addr_o_26_port, DRAM_Addr_o_25_port, DRAM_Addr_o_24_port, 
      DRAM_Addr_o_23_port, DRAM_Addr_o_22_port, DRAM_Addr_o_21_port, 
      DRAM_Addr_o_20_port, DRAM_Addr_o_19_port, DRAM_Addr_o_18_port, 
      DRAM_Addr_o_17_port, DRAM_Addr_o_16_port, DRAM_Addr_o_15_port, 
      DRAM_Addr_o_14_port, DRAM_Addr_o_13_port, DRAM_Addr_o_12_port, 
      DRAM_Addr_o_11_port, DRAM_Addr_o_10_port, DRAM_Addr_o_9_port, 
      DRAM_Addr_o_8_port, DRAM_Addr_o_7_port, DRAM_Addr_o_6_port, 
      DRAM_Addr_o_5_port, DRAM_Addr_o_4_port, DRAM_Addr_o_3_port, 
      DRAM_Addr_o_2_port, DRAM_Addr_o_1_port, DRAM_Addr_o_0_port );
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   UFETCH_BLOCK : fetch_block port map( branch_target_i(31) => 
                           dummy_branch_target_31_port, branch_target_i(30) => 
                           dummy_branch_target_30_port, branch_target_i(29) => 
                           dummy_branch_target_29_port, branch_target_i(28) => 
                           dummy_branch_target_28_port, branch_target_i(27) => 
                           dummy_branch_target_27_port, branch_target_i(26) => 
                           dummy_branch_target_26_port, branch_target_i(25) => 
                           dummy_branch_target_25_port, branch_target_i(24) => 
                           dummy_branch_target_24_port, branch_target_i(23) => 
                           dummy_branch_target_23_port, branch_target_i(22) => 
                           dummy_branch_target_22_port, branch_target_i(21) => 
                           dummy_branch_target_21_port, branch_target_i(20) => 
                           dummy_branch_target_20_port, branch_target_i(19) => 
                           dummy_branch_target_19_port, branch_target_i(18) => 
                           dummy_branch_target_18_port, branch_target_i(17) => 
                           dummy_branch_target_17_port, branch_target_i(16) => 
                           dummy_branch_target_16_port, branch_target_i(15) => 
                           dummy_branch_target_15_port, branch_target_i(14) => 
                           dummy_branch_target_14_port, branch_target_i(13) => 
                           dummy_branch_target_13_port, branch_target_i(12) => 
                           dummy_branch_target_12_port, branch_target_i(11) => 
                           dummy_branch_target_11_port, branch_target_i(10) => 
                           dummy_branch_target_10_port, branch_target_i(9) => 
                           dummy_branch_target_9_port, branch_target_i(8) => 
                           dummy_branch_target_8_port, branch_target_i(7) => 
                           dummy_branch_target_7_port, branch_target_i(6) => 
                           dummy_branch_target_6_port, branch_target_i(5) => 
                           dummy_branch_target_5_port, branch_target_i(4) => 
                           dummy_branch_target_4_port, branch_target_i(3) => 
                           dummy_branch_target_3_port, branch_target_i(2) => 
                           dummy_branch_target_2_port, branch_target_i(1) => 
                           dummy_branch_target_1_port, branch_target_i(0) => 
                           dummy_branch_target_0_port, sum_addr_i(31) => 
                           dummy_sum_addr_31_port, sum_addr_i(30) => 
                           dummy_sum_addr_30_port, sum_addr_i(29) => 
                           dummy_sum_addr_29_port, sum_addr_i(28) => 
                           dummy_sum_addr_28_port, sum_addr_i(27) => 
                           dummy_sum_addr_27_port, sum_addr_i(26) => 
                           dummy_sum_addr_26_port, sum_addr_i(25) => 
                           dummy_sum_addr_25_port, sum_addr_i(24) => 
                           dummy_sum_addr_24_port, sum_addr_i(23) => 
                           dummy_sum_addr_23_port, sum_addr_i(22) => 
                           dummy_sum_addr_22_port, sum_addr_i(21) => 
                           dummy_sum_addr_21_port, sum_addr_i(20) => 
                           dummy_sum_addr_20_port, sum_addr_i(19) => 
                           dummy_sum_addr_19_port, sum_addr_i(18) => 
                           dummy_sum_addr_18_port, sum_addr_i(17) => 
                           dummy_sum_addr_17_port, sum_addr_i(16) => 
                           dummy_sum_addr_16_port, sum_addr_i(15) => 
                           dummy_sum_addr_15_port, sum_addr_i(14) => 
                           dummy_sum_addr_14_port, sum_addr_i(13) => 
                           dummy_sum_addr_13_port, sum_addr_i(12) => 
                           dummy_sum_addr_12_port, sum_addr_i(11) => 
                           dummy_sum_addr_11_port, sum_addr_i(10) => 
                           dummy_sum_addr_10_port, sum_addr_i(9) => 
                           dummy_sum_addr_9_port, sum_addr_i(8) => 
                           dummy_sum_addr_8_port, sum_addr_i(7) => 
                           dummy_sum_addr_7_port, sum_addr_i(6) => 
                           dummy_sum_addr_6_port, sum_addr_i(5) => 
                           dummy_sum_addr_5_port, sum_addr_i(4) => 
                           dummy_sum_addr_4_port, sum_addr_i(3) => 
                           dummy_sum_addr_3_port, sum_addr_i(2) => 
                           dummy_sum_addr_2_port, sum_addr_i(1) => 
                           dummy_sum_addr_1_port, sum_addr_i(0) => 
                           dummy_sum_addr_0_port, A_i(31) => dummy_A_31_port, 
                           A_i(30) => dummy_A_30_port, A_i(29) => 
                           dummy_A_29_port, A_i(28) => dummy_A_28_port, A_i(27)
                           => dummy_A_27_port, A_i(26) => dummy_A_26_port, 
                           A_i(25) => dummy_A_25_port, A_i(24) => 
                           dummy_A_24_port, A_i(23) => dummy_A_23_port, A_i(22)
                           => dummy_A_22_port, A_i(21) => dummy_A_21_port, 
                           A_i(20) => dummy_A_20_port, A_i(19) => 
                           dummy_A_19_port, A_i(18) => dummy_A_18_port, A_i(17)
                           => dummy_A_17_port, A_i(16) => dummy_A_16_port, 
                           A_i(15) => dummy_A_15_port, A_i(14) => 
                           dummy_A_14_port, A_i(13) => dummy_A_13_port, A_i(12)
                           => dummy_A_12_port, A_i(11) => dummy_A_11_port, 
                           A_i(10) => dummy_A_10_port, A_i(9) => dummy_A_9_port
                           , A_i(8) => dummy_A_8_port, A_i(7) => dummy_A_7_port
                           , A_i(6) => dummy_A_6_port, A_i(5) => dummy_A_5_port
                           , A_i(4) => dummy_A_4_port, A_i(3) => dummy_A_3_port
                           , A_i(2) => dummy_A_2_port, A_i(1) => dummy_A_1_port
                           , A_i(0) => dummy_A_0_port, NPC4_i(31) => 
                           NPCF_31_port, NPC4_i(30) => NPCF_30_port, NPC4_i(29)
                           => NPCF_29_port, NPC4_i(28) => NPCF_28_port, 
                           NPC4_i(27) => NPCF_27_port, NPC4_i(26) => 
                           NPCF_26_port, NPC4_i(25) => NPCF_25_port, NPC4_i(24)
                           => NPCF_24_port, NPC4_i(23) => NPCF_23_port, 
                           NPC4_i(22) => NPCF_22_port, NPC4_i(21) => 
                           NPCF_21_port, NPC4_i(20) => NPCF_20_port, NPC4_i(19)
                           => NPCF_19_port, NPC4_i(18) => NPCF_18_port, 
                           NPC4_i(17) => NPCF_17_port, NPC4_i(16) => 
                           NPCF_16_port, NPC4_i(15) => NPCF_15_port, NPC4_i(14)
                           => NPCF_14_port, NPC4_i(13) => NPCF_13_port, 
                           NPC4_i(12) => NPCF_12_port, NPC4_i(11) => 
                           NPCF_11_port, NPC4_i(10) => NPCF_10_port, NPC4_i(9) 
                           => NPCF_9_port, NPC4_i(8) => NPCF_8_port, NPC4_i(7) 
                           => NPCF_7_port, NPC4_i(6) => NPCF_6_port, NPC4_i(5) 
                           => NPCF_5_port, NPC4_i(4) => NPCF_4_port, NPC4_i(3) 
                           => NPCF_3_port, NPC4_i(2) => NPCF_2_port, NPC4_i(1) 
                           => NPCF_1_port, NPC4_i(0) => NPCF_0_port, 
                           S_MUX_PC_BUS_i(1) => dummy_S_MUX_PC_BUS_1_port, 
                           S_MUX_PC_BUS_i(0) => dummy_S_MUX_PC_BUS_0_port, 
                           PC_o(31) => IRAM_Addr_o_31_port, PC_o(30) => 
                           IRAM_Addr_o_30_port, PC_o(29) => IRAM_Addr_o_29_port
                           , PC_o(28) => IRAM_Addr_o_28_port, PC_o(27) => 
                           IRAM_Addr_o_27_port, PC_o(26) => IRAM_Addr_o_26_port
                           , PC_o(25) => IRAM_Addr_o_25_port, PC_o(24) => 
                           IRAM_Addr_o_24_port, PC_o(23) => IRAM_Addr_o_23_port
                           , PC_o(22) => IRAM_Addr_o_22_port, PC_o(21) => 
                           IRAM_Addr_o_21_port, PC_o(20) => IRAM_Addr_o_20_port
                           , PC_o(19) => IRAM_Addr_o_19_port, PC_o(18) => 
                           IRAM_Addr_o_18_port, PC_o(17) => IRAM_Addr_o_17_port
                           , PC_o(16) => IRAM_Addr_o_16_port, PC_o(15) => 
                           IRAM_Addr_o_15_port, PC_o(14) => IRAM_Addr_o_14_port
                           , PC_o(13) => IRAM_Addr_o_13_port, PC_o(12) => 
                           IRAM_Addr_o_12_port, PC_o(11) => IRAM_Addr_o_11_port
                           , PC_o(10) => IRAM_Addr_o_10_port, PC_o(9) => 
                           IRAM_Addr_o_9_port, PC_o(8) => IRAM_Addr_o_8_port, 
                           PC_o(7) => IRAM_Addr_o_7_port, PC_o(6) => 
                           IRAM_Addr_o_6_port, PC_o(5) => IRAM_Addr_o_5_port, 
                           PC_o(4) => IRAM_Addr_o_4_port, PC_o(3) => 
                           IRAM_Addr_o_3_port, PC_o(2) => IRAM_Addr_o_2_port, 
                           PC_o(1) => IRAM_Addr_o_1_port, PC_o(0) => 
                           IRAM_Addr_o_0_port, PC4_o(31) => PC4_31_port, 
                           PC4_o(30) => PC4_30_port, PC4_o(29) => PC4_29_port, 
                           PC4_o(28) => PC4_28_port, PC4_o(27) => PC4_27_port, 
                           PC4_o(26) => PC4_26_port, PC4_o(25) => PC4_25_port, 
                           PC4_o(24) => PC4_24_port, PC4_o(23) => PC4_23_port, 
                           PC4_o(22) => PC4_22_port, PC4_o(21) => PC4_21_port, 
                           PC4_o(20) => PC4_20_port, PC4_o(19) => PC4_19_port, 
                           PC4_o(18) => PC4_18_port, PC4_o(17) => PC4_17_port, 
                           PC4_o(16) => PC4_16_port, PC4_o(15) => PC4_15_port, 
                           PC4_o(14) => PC4_14_port, PC4_o(13) => PC4_13_port, 
                           PC4_o(12) => PC4_12_port, PC4_o(11) => PC4_11_port, 
                           PC4_o(10) => PC4_10_port, PC4_o(9) => PC4_9_port, 
                           PC4_o(8) => PC4_8_port, PC4_o(7) => PC4_7_port, 
                           PC4_o(6) => PC4_6_port, PC4_o(5) => PC4_5_port, 
                           PC4_o(4) => PC4_4_port, PC4_o(3) => PC4_3_port, 
                           PC4_o(2) => PC4_2_port, PC4_o(1) => PC4_1_port, 
                           PC4_o(0) => PC4_0_port, PC_BUS_pre_BTB(31) => 
                           TARGET_PC_31_port, PC_BUS_pre_BTB(30) => 
                           TARGET_PC_30_port, PC_BUS_pre_BTB(29) => 
                           TARGET_PC_29_port, PC_BUS_pre_BTB(28) => 
                           TARGET_PC_28_port, PC_BUS_pre_BTB(27) => 
                           TARGET_PC_27_port, PC_BUS_pre_BTB(26) => 
                           TARGET_PC_26_port, PC_BUS_pre_BTB(25) => 
                           TARGET_PC_25_port, PC_BUS_pre_BTB(24) => 
                           TARGET_PC_24_port, PC_BUS_pre_BTB(23) => 
                           TARGET_PC_23_port, PC_BUS_pre_BTB(22) => 
                           TARGET_PC_22_port, PC_BUS_pre_BTB(21) => 
                           TARGET_PC_21_port, PC_BUS_pre_BTB(20) => n15, 
                           PC_BUS_pre_BTB(19) => TARGET_PC_19_port, 
                           PC_BUS_pre_BTB(18) => TARGET_PC_18_port, 
                           PC_BUS_pre_BTB(17) => TARGET_PC_17_port, 
                           PC_BUS_pre_BTB(16) => n14, PC_BUS_pre_BTB(15) => 
                           TARGET_PC_15_port, PC_BUS_pre_BTB(14) => 
                           TARGET_PC_14_port, PC_BUS_pre_BTB(13) => 
                           TARGET_PC_13_port, PC_BUS_pre_BTB(12) => 
                           TARGET_PC_12_port, PC_BUS_pre_BTB(11) => 
                           TARGET_PC_11_port, PC_BUS_pre_BTB(10) => 
                           TARGET_PC_10_port, PC_BUS_pre_BTB(9) => 
                           TARGET_PC_9_port, PC_BUS_pre_BTB(8) => n16, 
                           PC_BUS_pre_BTB(7) => TARGET_PC_7_port, 
                           PC_BUS_pre_BTB(6) => TARGET_PC_6_port, 
                           PC_BUS_pre_BTB(5) => TARGET_PC_5_port, 
                           PC_BUS_pre_BTB(4) => TARGET_PC_4_port, 
                           PC_BUS_pre_BTB(3) => TARGET_PC_3_port, 
                           PC_BUS_pre_BTB(2) => TARGET_PC_2_port, 
                           PC_BUS_pre_BTB(1) => TARGET_PC_1_port, 
                           PC_BUS_pre_BTB(0) => TARGET_PC_0_port, stall_i => 
                           n11, take_prediction_i => take_prediction, 
                           mispredict_i => mispredict, predicted_PC(31) => 
                           predicted_PC_31_port, predicted_PC(30) => 
                           predicted_PC_30_port, predicted_PC(29) => 
                           predicted_PC_29_port, predicted_PC(28) => 
                           predicted_PC_28_port, predicted_PC(27) => 
                           predicted_PC_27_port, predicted_PC(26) => 
                           predicted_PC_26_port, predicted_PC(25) => 
                           predicted_PC_25_port, predicted_PC(24) => 
                           predicted_PC_24_port, predicted_PC(23) => 
                           predicted_PC_23_port, predicted_PC(22) => 
                           predicted_PC_22_port, predicted_PC(21) => 
                           predicted_PC_21_port, predicted_PC(20) => 
                           predicted_PC_20_port, predicted_PC(19) => 
                           predicted_PC_19_port, predicted_PC(18) => 
                           predicted_PC_18_port, predicted_PC(17) => 
                           predicted_PC_17_port, predicted_PC(16) => 
                           predicted_PC_16_port, predicted_PC(15) => 
                           predicted_PC_15_port, predicted_PC(14) => 
                           predicted_PC_14_port, predicted_PC(13) => 
                           predicted_PC_13_port, predicted_PC(12) => 
                           predicted_PC_12_port, predicted_PC(11) => 
                           predicted_PC_11_port, predicted_PC(10) => 
                           predicted_PC_10_port, predicted_PC(9) => 
                           predicted_PC_9_port, predicted_PC(8) => 
                           predicted_PC_8_port, predicted_PC(7) => 
                           predicted_PC_7_port, predicted_PC(6) => 
                           predicted_PC_6_port, predicted_PC(5) => 
                           predicted_PC_5_port, predicted_PC(4) => 
                           predicted_PC_4_port, predicted_PC(3) => 
                           predicted_PC_3_port, predicted_PC(2) => 
                           predicted_PC_2_port, predicted_PC(1) => 
                           predicted_PC_1_port, predicted_PC(0) => 
                           predicted_PC_0_port, clk => clock, rst => rst);
   UBTB : btb_N_LINES4_SIZE32 port map( clock => clock, reset => rst, stall_i 
                           => n10, TAG_i(3) => IRAM_Addr_o_5_port, TAG_i(2) => 
                           IRAM_Addr_o_4_port, TAG_i(1) => IRAM_Addr_o_3_port, 
                           TAG_i(0) => IRAM_Addr_o_2_port, target_PC_i(31) => 
                           TARGET_PC_31_port, target_PC_i(30) => 
                           TARGET_PC_30_port, target_PC_i(29) => 
                           TARGET_PC_29_port, target_PC_i(28) => 
                           TARGET_PC_28_port, target_PC_i(27) => 
                           TARGET_PC_27_port, target_PC_i(26) => 
                           TARGET_PC_26_port, target_PC_i(25) => 
                           TARGET_PC_25_port, target_PC_i(24) => 
                           TARGET_PC_24_port, target_PC_i(23) => 
                           TARGET_PC_23_port, target_PC_i(22) => 
                           TARGET_PC_22_port, target_PC_i(21) => 
                           TARGET_PC_21_port, target_PC_i(20) => n15, 
                           target_PC_i(19) => TARGET_PC_19_port, 
                           target_PC_i(18) => TARGET_PC_18_port, 
                           target_PC_i(17) => TARGET_PC_17_port, 
                           target_PC_i(16) => n14, target_PC_i(15) => 
                           TARGET_PC_15_port, target_PC_i(14) => 
                           TARGET_PC_14_port, target_PC_i(13) => 
                           TARGET_PC_13_port, target_PC_i(12) => 
                           TARGET_PC_12_port, target_PC_i(11) => 
                           TARGET_PC_11_port, target_PC_i(10) => 
                           TARGET_PC_10_port, target_PC_i(9) => 
                           TARGET_PC_9_port, target_PC_i(8) => n16, 
                           target_PC_i(7) => TARGET_PC_7_port, target_PC_i(6) 
                           => TARGET_PC_6_port, target_PC_i(5) => 
                           TARGET_PC_5_port, target_PC_i(4) => TARGET_PC_4_port
                           , target_PC_i(3) => TARGET_PC_3_port, target_PC_i(2)
                           => TARGET_PC_2_port, target_PC_i(1) => 
                           TARGET_PC_1_port, target_PC_i(0) => TARGET_PC_0_port
                           , was_taken_i => was_taken, predicted_next_PC_o(31) 
                           => predicted_PC_31_port, predicted_next_PC_o(30) => 
                           predicted_PC_30_port, predicted_next_PC_o(29) => 
                           predicted_PC_29_port, predicted_next_PC_o(28) => 
                           predicted_PC_28_port, predicted_next_PC_o(27) => 
                           predicted_PC_27_port, predicted_next_PC_o(26) => 
                           predicted_PC_26_port, predicted_next_PC_o(25) => 
                           predicted_PC_25_port, predicted_next_PC_o(24) => 
                           predicted_PC_24_port, predicted_next_PC_o(23) => 
                           predicted_PC_23_port, predicted_next_PC_o(22) => 
                           predicted_PC_22_port, predicted_next_PC_o(21) => 
                           predicted_PC_21_port, predicted_next_PC_o(20) => 
                           predicted_PC_20_port, predicted_next_PC_o(19) => 
                           predicted_PC_19_port, predicted_next_PC_o(18) => 
                           predicted_PC_18_port, predicted_next_PC_o(17) => 
                           predicted_PC_17_port, predicted_next_PC_o(16) => 
                           predicted_PC_16_port, predicted_next_PC_o(15) => 
                           predicted_PC_15_port, predicted_next_PC_o(14) => 
                           predicted_PC_14_port, predicted_next_PC_o(13) => 
                           predicted_PC_13_port, predicted_next_PC_o(12) => 
                           predicted_PC_12_port, predicted_next_PC_o(11) => 
                           predicted_PC_11_port, predicted_next_PC_o(10) => 
                           predicted_PC_10_port, predicted_next_PC_o(9) => 
                           predicted_PC_9_port, predicted_next_PC_o(8) => 
                           predicted_PC_8_port, predicted_next_PC_o(7) => 
                           predicted_PC_7_port, predicted_next_PC_o(6) => 
                           predicted_PC_6_port, predicted_next_PC_o(5) => 
                           predicted_PC_5_port, predicted_next_PC_o(4) => 
                           predicted_PC_4_port, predicted_next_PC_o(3) => 
                           predicted_PC_3_port, predicted_next_PC_o(2) => 
                           predicted_PC_2_port, predicted_next_PC_o(1) => 
                           predicted_PC_1_port, predicted_next_PC_o(0) => 
                           predicted_PC_0_port, taken_o => take_prediction, 
                           mispredict_o => mispredict);
   UFEETCH_REGS : fetch_regs port map( NPCF_i(31) => PC4_31_port, NPCF_i(30) =>
                           PC4_30_port, NPCF_i(29) => PC4_29_port, NPCF_i(28) 
                           => PC4_28_port, NPCF_i(27) => PC4_27_port, 
                           NPCF_i(26) => PC4_26_port, NPCF_i(25) => PC4_25_port
                           , NPCF_i(24) => PC4_24_port, NPCF_i(23) => 
                           PC4_23_port, NPCF_i(22) => PC4_22_port, NPCF_i(21) 
                           => PC4_21_port, NPCF_i(20) => PC4_20_port, 
                           NPCF_i(19) => PC4_19_port, NPCF_i(18) => PC4_18_port
                           , NPCF_i(17) => PC4_17_port, NPCF_i(16) => 
                           PC4_16_port, NPCF_i(15) => PC4_15_port, NPCF_i(14) 
                           => PC4_14_port, NPCF_i(13) => PC4_13_port, 
                           NPCF_i(12) => PC4_12_port, NPCF_i(11) => PC4_11_port
                           , NPCF_i(10) => PC4_10_port, NPCF_i(9) => PC4_9_port
                           , NPCF_i(8) => PC4_8_port, NPCF_i(7) => PC4_7_port, 
                           NPCF_i(6) => PC4_6_port, NPCF_i(5) => PC4_5_port, 
                           NPCF_i(4) => PC4_4_port, NPCF_i(3) => PC4_3_port, 
                           NPCF_i(2) => PC4_2_port, NPCF_i(1) => PC4_1_port, 
                           NPCF_i(0) => PC4_0_port, IR_i(31) => IRAM_Dout_i(31)
                           , IR_i(30) => IRAM_Dout_i(30), IR_i(29) => 
                           IRAM_Dout_i(29), IR_i(28) => IRAM_Dout_i(28), 
                           IR_i(27) => IRAM_Dout_i(27), IR_i(26) => 
                           IRAM_Dout_i(26), IR_i(25) => IRAM_Dout_i(25), 
                           IR_i(24) => IRAM_Dout_i(24), IR_i(23) => 
                           IRAM_Dout_i(23), IR_i(22) => IRAM_Dout_i(22), 
                           IR_i(21) => IRAM_Dout_i(21), IR_i(20) => 
                           IRAM_Dout_i(20), IR_i(19) => IRAM_Dout_i(19), 
                           IR_i(18) => IRAM_Dout_i(18), IR_i(17) => 
                           IRAM_Dout_i(17), IR_i(16) => IRAM_Dout_i(16), 
                           IR_i(15) => IRAM_Dout_i(15), IR_i(14) => 
                           IRAM_Dout_i(14), IR_i(13) => IRAM_Dout_i(13), 
                           IR_i(12) => IRAM_Dout_i(12), IR_i(11) => 
                           IRAM_Dout_i(11), IR_i(10) => IRAM_Dout_i(10), 
                           IR_i(9) => IRAM_Dout_i(9), IR_i(8) => IRAM_Dout_i(8)
                           , IR_i(7) => IRAM_Dout_i(7), IR_i(6) => 
                           IRAM_Dout_i(6), IR_i(5) => IRAM_Dout_i(5), IR_i(4) 
                           => IRAM_Dout_i(4), IR_i(3) => IRAM_Dout_i(3), 
                           IR_i(2) => IRAM_Dout_i(2), IR_i(1) => IRAM_Dout_i(1)
                           , IR_i(0) => IRAM_Dout_i(0), NPCF_o(31) => 
                           NPCF_31_port, NPCF_o(30) => NPCF_30_port, NPCF_o(29)
                           => NPCF_29_port, NPCF_o(28) => NPCF_28_port, 
                           NPCF_o(27) => NPCF_27_port, NPCF_o(26) => 
                           NPCF_26_port, NPCF_o(25) => NPCF_25_port, NPCF_o(24)
                           => NPCF_24_port, NPCF_o(23) => NPCF_23_port, 
                           NPCF_o(22) => NPCF_22_port, NPCF_o(21) => 
                           NPCF_21_port, NPCF_o(20) => NPCF_20_port, NPCF_o(19)
                           => NPCF_19_port, NPCF_o(18) => NPCF_18_port, 
                           NPCF_o(17) => NPCF_17_port, NPCF_o(16) => 
                           NPCF_16_port, NPCF_o(15) => NPCF_15_port, NPCF_o(14)
                           => NPCF_14_port, NPCF_o(13) => NPCF_13_port, 
                           NPCF_o(12) => NPCF_12_port, NPCF_o(11) => 
                           NPCF_11_port, NPCF_o(10) => NPCF_10_port, NPCF_o(9) 
                           => NPCF_9_port, NPCF_o(8) => NPCF_8_port, NPCF_o(7) 
                           => NPCF_7_port, NPCF_o(6) => NPCF_6_port, NPCF_o(5) 
                           => NPCF_5_port, NPCF_o(4) => NPCF_4_port, NPCF_o(3) 
                           => NPCF_3_port, NPCF_o(2) => NPCF_2_port, NPCF_o(1) 
                           => NPCF_1_port, NPCF_o(0) => NPCF_0_port, IR_o(31) 
                           => IR_31_port, IR_o(30) => IR_30_port, IR_o(29) => 
                           IR_29_port, IR_o(28) => IR_28_port, IR_o(27) => 
                           IR_27_port, IR_o(26) => IR_26_port, IR_o(25) => 
                           IR_25_port, IR_o(24) => IR_24_port, IR_o(23) => 
                           IR_23_port, IR_o(22) => IR_22_port, IR_o(21) => 
                           IR_21_port, IR_o(20) => IR_20_port, IR_o(19) => 
                           IR_19_port, IR_o(18) => IR_18_port, IR_o(17) => 
                           IR_17_port, IR_o(16) => IR_16_port, IR_o(15) => 
                           IR_15_port, IR_o(14) => IR_14_port, IR_o(13) => 
                           IR_13_port, IR_o(12) => IR_12_port, IR_o(11) => 
                           IR_11_port, IR_o(10) => IR_10_port, IR_o(9) => 
                           IR_9_port, IR_o(8) => IR_8_port, IR_o(7) => 
                           IR_7_port, IR_o(6) => IR_6_port, IR_o(5) => 
                           IR_5_port, IR_o(4) => IR_4_port, IR_o(3) => 
                           IR_3_port, IR_o(2) => IR_2_port, IR_o(1) => 
                           IR_1_port, IR_o(0) => IR_0_port, stall_i => n12, clk
                           => clock, rst => rst);
   UJUMP_LOGIC : jump_logic port map( NPCF_i(31) => NPCF_31_port, NPCF_i(30) =>
                           NPCF_30_port, NPCF_i(29) => NPCF_29_port, NPCF_i(28)
                           => NPCF_28_port, NPCF_i(27) => NPCF_27_port, 
                           NPCF_i(26) => NPCF_26_port, NPCF_i(25) => 
                           NPCF_25_port, NPCF_i(24) => NPCF_24_port, NPCF_i(23)
                           => NPCF_23_port, NPCF_i(22) => NPCF_22_port, 
                           NPCF_i(21) => NPCF_21_port, NPCF_i(20) => 
                           NPCF_20_port, NPCF_i(19) => NPCF_19_port, NPCF_i(18)
                           => NPCF_18_port, NPCF_i(17) => NPCF_17_port, 
                           NPCF_i(16) => NPCF_16_port, NPCF_i(15) => 
                           NPCF_15_port, NPCF_i(14) => NPCF_14_port, NPCF_i(13)
                           => NPCF_13_port, NPCF_i(12) => NPCF_12_port, 
                           NPCF_i(11) => NPCF_11_port, NPCF_i(10) => 
                           NPCF_10_port, NPCF_i(9) => NPCF_9_port, NPCF_i(8) =>
                           NPCF_8_port, NPCF_i(7) => NPCF_7_port, NPCF_i(6) => 
                           NPCF_6_port, NPCF_i(5) => NPCF_5_port, NPCF_i(4) => 
                           NPCF_4_port, NPCF_i(3) => NPCF_3_port, NPCF_i(2) => 
                           NPCF_2_port, NPCF_i(1) => NPCF_1_port, NPCF_i(0) => 
                           NPCF_0_port, IR_i(31) => n23, IR_i(30) => n24, 
                           IR_i(29) => n25, IR_i(28) => n26, IR_i(27) => n27, 
                           IR_i(26) => n28, IR_i(25) => IR_25_port, IR_i(24) =>
                           IR_24_port, IR_i(23) => IR_23_port, IR_i(22) => 
                           IR_22_port, IR_i(21) => IR_21_port, IR_i(20) => 
                           IR_20_port, IR_i(19) => IR_19_port, IR_i(18) => 
                           IR_18_port, IR_i(17) => IR_17_port, IR_i(16) => 
                           IR_16_port, IR_i(15) => IR_15_port, IR_i(14) => 
                           IR_14_port, IR_i(13) => IR_13_port, IR_i(12) => 
                           IR_12_port, IR_i(11) => IR_11_port, IR_i(10) => 
                           IR_10_port, IR_i(9) => IR_9_port, IR_i(8) => 
                           IR_8_port, IR_i(7) => IR_7_port, IR_i(6) => 
                           IR_6_port, IR_i(5) => IR_5_port, IR_i(4) => 
                           IR_4_port, IR_i(3) => IR_3_port, IR_i(2) => 
                           IR_2_port, IR_i(1) => IR_1_port, IR_i(0) => 
                           IR_0_port, A_i(31) => AtoComp_31_port, A_i(30) => 
                           AtoComp_30_port, A_i(29) => AtoComp_29_port, A_i(28)
                           => AtoComp_28_port, A_i(27) => AtoComp_27_port, 
                           A_i(26) => AtoComp_26_port, A_i(25) => 
                           AtoComp_25_port, A_i(24) => AtoComp_24_port, A_i(23)
                           => AtoComp_23_port, A_i(22) => AtoComp_22_port, 
                           A_i(21) => AtoComp_21_port, A_i(20) => 
                           AtoComp_20_port, A_i(19) => AtoComp_19_port, A_i(18)
                           => AtoComp_18_port, A_i(17) => AtoComp_17_port, 
                           A_i(16) => AtoComp_16_port, A_i(15) => 
                           AtoComp_15_port, A_i(14) => AtoComp_14_port, A_i(13)
                           => AtoComp_13_port, A_i(12) => AtoComp_12_port, 
                           A_i(11) => AtoComp_11_port, A_i(10) => 
                           AtoComp_10_port, A_i(9) => AtoComp_9_port, A_i(8) =>
                           AtoComp_8_port, A_i(7) => AtoComp_7_port, A_i(6) => 
                           AtoComp_6_port, A_i(5) => AtoComp_5_port, A_i(4) => 
                           AtoComp_4_port, A_i(3) => AtoComp_3_port, A_i(2) => 
                           AtoComp_2_port, A_i(1) => AtoComp_1_port, A_i(0) => 
                           AtoComp_0_port, A_o(31) => dummy_A_31_port, A_o(30) 
                           => dummy_A_30_port, A_o(29) => dummy_A_29_port, 
                           A_o(28) => dummy_A_28_port, A_o(27) => 
                           dummy_A_27_port, A_o(26) => dummy_A_26_port, A_o(25)
                           => dummy_A_25_port, A_o(24) => dummy_A_24_port, 
                           A_o(23) => dummy_A_23_port, A_o(22) => 
                           dummy_A_22_port, A_o(21) => dummy_A_21_port, A_o(20)
                           => dummy_A_20_port, A_o(19) => dummy_A_19_port, 
                           A_o(18) => dummy_A_18_port, A_o(17) => 
                           dummy_A_17_port, A_o(16) => dummy_A_16_port, A_o(15)
                           => dummy_A_15_port, A_o(14) => dummy_A_14_port, 
                           A_o(13) => dummy_A_13_port, A_o(12) => 
                           dummy_A_12_port, A_o(11) => dummy_A_11_port, A_o(10)
                           => dummy_A_10_port, A_o(9) => dummy_A_9_port, A_o(8)
                           => dummy_A_8_port, A_o(7) => dummy_A_7_port, A_o(6) 
                           => dummy_A_6_port, A_o(5) => dummy_A_5_port, A_o(4) 
                           => dummy_A_4_port, A_o(3) => dummy_A_3_port, A_o(2) 
                           => dummy_A_2_port, A_o(1) => dummy_A_1_port, A_o(0) 
                           => dummy_A_0_port, rA_o(4) => rA2reg_4_port, rA_o(3)
                           => rA2reg_3_port, rA_o(2) => rA2reg_2_port, rA_o(1) 
                           => rA2reg_1_port, rA_o(0) => rA2reg_0_port, rB_o(4) 
                           => rB2reg_4_port, rB_o(3) => rB2reg_3_port, rB_o(2) 
                           => rB2reg_2_port, rB_o(1) => rB2reg_1_port, rB_o(0) 
                           => rB2reg_0_port, rC_o(4) => rC2reg_4_port, rC_o(3) 
                           => rC2reg_3_port, rC_o(2) => rC2reg_2_port, rC_o(1) 
                           => rC2reg_1_port, rC_o(0) => rC2reg_0_port, 
                           branch_target_o(31) => dummy_branch_target_31_port, 
                           branch_target_o(30) => dummy_branch_target_30_port, 
                           branch_target_o(29) => dummy_branch_target_29_port, 
                           branch_target_o(28) => dummy_branch_target_28_port, 
                           branch_target_o(27) => dummy_branch_target_27_port, 
                           branch_target_o(26) => dummy_branch_target_26_port, 
                           branch_target_o(25) => dummy_branch_target_25_port, 
                           branch_target_o(24) => dummy_branch_target_24_port, 
                           branch_target_o(23) => dummy_branch_target_23_port, 
                           branch_target_o(22) => dummy_branch_target_22_port, 
                           branch_target_o(21) => dummy_branch_target_21_port, 
                           branch_target_o(20) => dummy_branch_target_20_port, 
                           branch_target_o(19) => dummy_branch_target_19_port, 
                           branch_target_o(18) => dummy_branch_target_18_port, 
                           branch_target_o(17) => dummy_branch_target_17_port, 
                           branch_target_o(16) => dummy_branch_target_16_port, 
                           branch_target_o(15) => dummy_branch_target_15_port, 
                           branch_target_o(14) => dummy_branch_target_14_port, 
                           branch_target_o(13) => dummy_branch_target_13_port, 
                           branch_target_o(12) => dummy_branch_target_12_port, 
                           branch_target_o(11) => dummy_branch_target_11_port, 
                           branch_target_o(10) => dummy_branch_target_10_port, 
                           branch_target_o(9) => dummy_branch_target_9_port, 
                           branch_target_o(8) => dummy_branch_target_8_port, 
                           branch_target_o(7) => dummy_branch_target_7_port, 
                           branch_target_o(6) => dummy_branch_target_6_port, 
                           branch_target_o(5) => dummy_branch_target_5_port, 
                           branch_target_o(4) => dummy_branch_target_4_port, 
                           branch_target_o(3) => dummy_branch_target_3_port, 
                           branch_target_o(2) => dummy_branch_target_2_port, 
                           branch_target_o(1) => dummy_branch_target_1_port, 
                           branch_target_o(0) => dummy_branch_target_0_port, 
                           sum_addr_o(31) => dummy_sum_addr_31_port, 
                           sum_addr_o(30) => dummy_sum_addr_30_port, 
                           sum_addr_o(29) => dummy_sum_addr_29_port, 
                           sum_addr_o(28) => dummy_sum_addr_28_port, 
                           sum_addr_o(27) => dummy_sum_addr_27_port, 
                           sum_addr_o(26) => dummy_sum_addr_26_port, 
                           sum_addr_o(25) => dummy_sum_addr_25_port, 
                           sum_addr_o(24) => dummy_sum_addr_24_port, 
                           sum_addr_o(23) => dummy_sum_addr_23_port, 
                           sum_addr_o(22) => dummy_sum_addr_22_port, 
                           sum_addr_o(21) => dummy_sum_addr_21_port, 
                           sum_addr_o(20) => dummy_sum_addr_20_port, 
                           sum_addr_o(19) => dummy_sum_addr_19_port, 
                           sum_addr_o(18) => dummy_sum_addr_18_port, 
                           sum_addr_o(17) => dummy_sum_addr_17_port, 
                           sum_addr_o(16) => dummy_sum_addr_16_port, 
                           sum_addr_o(15) => dummy_sum_addr_15_port, 
                           sum_addr_o(14) => dummy_sum_addr_14_port, 
                           sum_addr_o(13) => dummy_sum_addr_13_port, 
                           sum_addr_o(12) => dummy_sum_addr_12_port, 
                           sum_addr_o(11) => dummy_sum_addr_11_port, 
                           sum_addr_o(10) => dummy_sum_addr_10_port, 
                           sum_addr_o(9) => dummy_sum_addr_9_port, 
                           sum_addr_o(8) => dummy_sum_addr_8_port, 
                           sum_addr_o(7) => dummy_sum_addr_7_port, 
                           sum_addr_o(6) => dummy_sum_addr_6_port, 
                           sum_addr_o(5) => dummy_sum_addr_5_port, 
                           sum_addr_o(4) => dummy_sum_addr_4_port, 
                           sum_addr_o(3) => dummy_sum_addr_3_port, 
                           sum_addr_o(2) => dummy_sum_addr_2_port, 
                           sum_addr_o(1) => dummy_sum_addr_1_port, 
                           sum_addr_o(0) => dummy_sum_addr_0_port, 
                           extended_imm(31) => help_IMM_31_port, 
                           extended_imm(30) => help_IMM_30_port, 
                           extended_imm(29) => help_IMM_29_port, 
                           extended_imm(28) => help_IMM_28_port, 
                           extended_imm(27) => help_IMM_27_port, 
                           extended_imm(26) => help_IMM_26_port, 
                           extended_imm(25) => help_IMM_25_port, 
                           extended_imm(24) => help_IMM_24_port, 
                           extended_imm(23) => help_IMM_23_port, 
                           extended_imm(22) => help_IMM_22_port, 
                           extended_imm(21) => help_IMM_21_port, 
                           extended_imm(20) => help_IMM_20_port, 
                           extended_imm(19) => help_IMM_19_port, 
                           extended_imm(18) => help_IMM_18_port, 
                           extended_imm(17) => help_IMM_17_port, 
                           extended_imm(16) => help_IMM_16_port, 
                           extended_imm(15) => help_IMM_15_port, 
                           extended_imm(14) => help_IMM_14_port, 
                           extended_imm(13) => help_IMM_13_port, 
                           extended_imm(12) => help_IMM_12_port, 
                           extended_imm(11) => help_IMM_11_port, 
                           extended_imm(10) => help_IMM_10_port, 
                           extended_imm(9) => help_IMM_9_port, extended_imm(8) 
                           => help_IMM_8_port, extended_imm(7) => 
                           help_IMM_7_port, extended_imm(6) => help_IMM_6_port,
                           extended_imm(5) => help_IMM_5_port, extended_imm(4) 
                           => help_IMM_4_port, extended_imm(3) => 
                           help_IMM_3_port, extended_imm(2) => help_IMM_2_port,
                           extended_imm(1) => help_IMM_1_port, extended_imm(0) 
                           => help_IMM_0_port, taken_o => was_taken_from_jl, 
                           FW_X_i(31) => DRAM_Addr_o_31_port, FW_X_i(30) => 
                           DRAM_Addr_o_30_port, FW_X_i(29) => 
                           DRAM_Addr_o_29_port, FW_X_i(28) => 
                           DRAM_Addr_o_28_port, FW_X_i(27) => 
                           DRAM_Addr_o_27_port, FW_X_i(26) => 
                           DRAM_Addr_o_26_port, FW_X_i(25) => 
                           DRAM_Addr_o_25_port, FW_X_i(24) => 
                           DRAM_Addr_o_24_port, FW_X_i(23) => 
                           DRAM_Addr_o_23_port, FW_X_i(22) => 
                           DRAM_Addr_o_22_port, FW_X_i(21) => 
                           DRAM_Addr_o_21_port, FW_X_i(20) => 
                           DRAM_Addr_o_20_port, FW_X_i(19) => 
                           DRAM_Addr_o_19_port, FW_X_i(18) => 
                           DRAM_Addr_o_18_port, FW_X_i(17) => 
                           DRAM_Addr_o_17_port, FW_X_i(16) => 
                           DRAM_Addr_o_16_port, FW_X_i(15) => 
                           DRAM_Addr_o_15_port, FW_X_i(14) => 
                           DRAM_Addr_o_14_port, FW_X_i(13) => 
                           DRAM_Addr_o_13_port, FW_X_i(12) => 
                           DRAM_Addr_o_12_port, FW_X_i(11) => 
                           DRAM_Addr_o_11_port, FW_X_i(10) => 
                           DRAM_Addr_o_10_port, FW_X_i(9) => DRAM_Addr_o_9_port
                           , FW_X_i(8) => DRAM_Addr_o_8_port, FW_X_i(7) => 
                           DRAM_Addr_o_7_port, FW_X_i(6) => DRAM_Addr_o_6_port,
                           FW_X_i(5) => DRAM_Addr_o_5_port, FW_X_i(4) => 
                           DRAM_Addr_o_4_port, FW_X_i(3) => DRAM_Addr_o_3_port,
                           FW_X_i(2) => DRAM_Addr_o_2_port, FW_X_i(1) => 
                           DRAM_Addr_o_1_port, FW_X_i(0) => DRAM_Addr_o_0_port,
                           FW_W_i(31) => wb2reg_31_port, FW_W_i(30) => 
                           wb2reg_30_port, FW_W_i(29) => wb2reg_29_port, 
                           FW_W_i(28) => wb2reg_28_port, FW_W_i(27) => 
                           wb2reg_27_port, FW_W_i(26) => wb2reg_26_port, 
                           FW_W_i(25) => wb2reg_25_port, FW_W_i(24) => 
                           wb2reg_24_port, FW_W_i(23) => wb2reg_23_port, 
                           FW_W_i(22) => wb2reg_22_port, FW_W_i(21) => 
                           wb2reg_21_port, FW_W_i(20) => wb2reg_20_port, 
                           FW_W_i(19) => wb2reg_19_port, FW_W_i(18) => 
                           wb2reg_18_port, FW_W_i(17) => wb2reg_17_port, 
                           FW_W_i(16) => wb2reg_16_port, FW_W_i(15) => 
                           wb2reg_15_port, FW_W_i(14) => wb2reg_14_port, 
                           FW_W_i(13) => wb2reg_13_port, FW_W_i(12) => 
                           wb2reg_12_port, FW_W_i(11) => wb2reg_11_port, 
                           FW_W_i(10) => wb2reg_10_port, FW_W_i(9) => 
                           wb2reg_9_port, FW_W_i(8) => wb2reg_8_port, FW_W_i(7)
                           => wb2reg_7_port, FW_W_i(6) => wb2reg_6_port, 
                           FW_W_i(5) => wb2reg_5_port, FW_W_i(4) => 
                           wb2reg_4_port, FW_W_i(3) => wb2reg_3_port, FW_W_i(2)
                           => wb2reg_2_port, FW_W_i(1) => wb2reg_1_port, 
                           FW_W_i(0) => wb2reg_0_port, S_FW_Adec_i(1) => 
                           dummy_S_FWAdec_1_port, S_FW_Adec_i(0) => 
                           dummy_S_FWAdec_0_port, S_EXT_i => dummy_S_EXT, 
                           S_EXT_SIGN_i => dummy_S_EXT_SIGN, S_MUX_LINK_i => 
                           dummy_S_MUX_LINK, S_EQ_NEQ_i => dummy_S_EQ_NEQ);
   UCU : 
                           dlx_cu_MICROCODE_MEM_SIZE64_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE13 
                           port map( Clk => clock, Rst => rst, IR_IN(31) => 
                           IR_31_port, IR_IN(30) => IR_30_port, IR_IN(29) => 
                           IR_29_port, IR_IN(28) => IR_28_port, IR_IN(27) => 
                           IR_27_port, IR_IN(26) => IR_26_port, IR_IN(25) => 
                           IR_25_port, IR_IN(24) => IR_24_port, IR_IN(23) => 
                           IR_23_port, IR_IN(22) => IR_22_port, IR_IN(21) => 
                           IR_21_port, IR_IN(20) => IR_20_port, IR_IN(19) => 
                           IR_19_port, IR_IN(18) => IR_18_port, IR_IN(17) => 
                           IR_17_port, IR_IN(16) => IR_16_port, IR_IN(15) => 
                           n29, IR_IN(14) => n30, IR_IN(13) => n31, IR_IN(12) 
                           => n32, IR_IN(11) => n33, IR_IN(10) => IR_10_port, 
                           IR_IN(9) => IR_9_port, IR_IN(8) => IR_8_port, 
                           IR_IN(7) => IR_7_port, IR_IN(6) => IR_6_port, 
                           IR_IN(5) => IR_5_port, IR_IN(4) => IR_4_port, 
                           IR_IN(3) => IR_3_port, IR_IN(2) => IR_2_port, 
                           IR_IN(1) => IR_1_port, IR_IN(0) => IR_0_port, 
                           stall_exe_i => exe_stall_cu, mispredict_i => n21, 
                           D1_i(4) => muxed_dest2exe_4_port, D1_i(3) => 
                           muxed_dest2exe_3_port, D1_i(2) => 
                           muxed_dest2exe_2_port, D1_i(1) => 
                           muxed_dest2exe_1_port, D1_i(0) => 
                           muxed_dest2exe_0_port, D2_i(4) => D22D3_4_port, 
                           D2_i(3) => n19, D2_i(2) => n20, D2_i(1) => n17, 
                           D2_i(0) => n18, S1_LATCH_EN => net684116, 
                           S2_LATCH_EN => net684117, S3_LATCH_EN => net684118, 
                           S_MUX_PC_BUS(1) => dummy_S_MUX_PC_BUS_1_port, 
                           S_MUX_PC_BUS(0) => dummy_S_MUX_PC_BUS_0_port, S_EXT 
                           => dummy_S_EXT, S_EXT_SIGN => dummy_S_EXT_SIGN, 
                           S_EQ_NEQ => dummy_S_EQ_NEQ, S_MUX_DEST(1) => 
                           dummy_S_MUX_DEST_1_port, S_MUX_DEST(0) => 
                           dummy_S_MUX_DEST_0_port, S_MUX_LINK => 
                           dummy_S_MUX_LINK, S_MEM_W_R => DRAM_WR_o, S_MEM_EN 
                           => DRAM_Enable_o, S_RF_W_wb => dummy_S_RF_W_wb, 
                           S_RF_W_mem => dummy_S_RF_W_mem, S_RF_W_exe => 
                           net684119, S_MUX_ALUIN => dummy_S_MUX_ALUIN, 
                           stall_exe_o => stall_exe, stall_dec_o => n12, 
                           stall_fetch_o => n11, stall_btb_o => n10, 
                           was_branch_o => was_branch, was_jmp_o => was_jmp, 
                           ALU_WORD_o(12) => ALUW_dec_12_port, ALU_WORD_o(11) 
                           => ALUW_dec_11_port, ALU_WORD_o(10) => 
                           ALUW_dec_10_port, ALU_WORD_o(9) => ALUW_dec_9_port, 
                           ALU_WORD_o(8) => ALUW_dec_8_port, ALU_WORD_o(7) => 
                           ALUW_dec_7_port, ALU_WORD_o(6) => ALUW_dec_6_port, 
                           ALU_WORD_o(5) => ALUW_dec_5_port, ALU_WORD_o(4) => 
                           ALUW_dec_4_port, ALU_WORD_o(3) => ALUW_dec_3_port, 
                           ALU_WORD_o(2) => ALUW_dec_2_port, ALU_WORD_o(1) => 
                           ALUW_dec_1_port, ALU_WORD_o(0) => ALUW_dec_0_port, 
                           ALU_OPCODE(0) => net684120, ALU_OPCODE(1) => 
                           net684121, ALU_OPCODE(2) => net684122, ALU_OPCODE(3)
                           => net684123, ALU_OPCODE(4) => net684124, 
                           S_MUX_MEM_BAR => dummy_S_MUX_MEM);
   RF : dlx_regfile port map( Clk => clock, Rst => rst, ENABLE => n22, RD1 => 
                           X_Logic1_port, RD2 => X_Logic1_port, WR => 
                           dummy_S_RF_W_mem, ADD_WR(4) => D22D3_4_port, 
                           ADD_WR(3) => n19, ADD_WR(2) => n20, ADD_WR(1) => n17
                           , ADD_WR(0) => n18, ADD_RD1(4) => IRAM_Dout_i(25), 
                           ADD_RD1(3) => IRAM_Dout_i(24), ADD_RD1(2) => 
                           IRAM_Dout_i(23), ADD_RD1(1) => IRAM_Dout_i(22), 
                           ADD_RD1(0) => IRAM_Dout_i(21), ADD_RD2(4) => 
                           IRAM_Dout_i(20), ADD_RD2(3) => IRAM_Dout_i(19), 
                           ADD_RD2(2) => IRAM_Dout_i(18), ADD_RD2(1) => 
                           IRAM_Dout_i(17), ADD_RD2(0) => IRAM_Dout_i(16), 
                           DATAIN(31) => W2wb_31_port, DATAIN(30) => 
                           W2wb_30_port, DATAIN(29) => W2wb_29_port, DATAIN(28)
                           => W2wb_28_port, DATAIN(27) => W2wb_27_port, 
                           DATAIN(26) => W2wb_26_port, DATAIN(25) => 
                           W2wb_25_port, DATAIN(24) => W2wb_24_port, DATAIN(23)
                           => W2wb_23_port, DATAIN(22) => W2wb_22_port, 
                           DATAIN(21) => W2wb_21_port, DATAIN(20) => 
                           W2wb_20_port, DATAIN(19) => W2wb_19_port, DATAIN(18)
                           => W2wb_18_port, DATAIN(17) => W2wb_17_port, 
                           DATAIN(16) => W2wb_16_port, DATAIN(15) => 
                           W2wb_15_port, DATAIN(14) => W2wb_14_port, DATAIN(13)
                           => W2wb_13_port, DATAIN(12) => W2wb_12_port, 
                           DATAIN(11) => W2wb_11_port, DATAIN(10) => 
                           W2wb_10_port, DATAIN(9) => W2wb_9_port, DATAIN(8) =>
                           W2wb_8_port, DATAIN(7) => W2wb_7_port, DATAIN(6) => 
                           W2wb_6_port, DATAIN(5) => W2wb_5_port, DATAIN(4) => 
                           W2wb_4_port, DATAIN(3) => W2wb_3_port, DATAIN(2) => 
                           W2wb_2_port, DATAIN(1) => W2wb_1_port, DATAIN(0) => 
                           W2wb_0_port, OUT1(31) => AtoComp_31_port, OUT1(30) 
                           => AtoComp_30_port, OUT1(29) => AtoComp_29_port, 
                           OUT1(28) => AtoComp_28_port, OUT1(27) => 
                           AtoComp_27_port, OUT1(26) => AtoComp_26_port, 
                           OUT1(25) => AtoComp_25_port, OUT1(24) => 
                           AtoComp_24_port, OUT1(23) => AtoComp_23_port, 
                           OUT1(22) => AtoComp_22_port, OUT1(21) => 
                           AtoComp_21_port, OUT1(20) => AtoComp_20_port, 
                           OUT1(19) => AtoComp_19_port, OUT1(18) => 
                           AtoComp_18_port, OUT1(17) => AtoComp_17_port, 
                           OUT1(16) => AtoComp_16_port, OUT1(15) => 
                           AtoComp_15_port, OUT1(14) => AtoComp_14_port, 
                           OUT1(13) => AtoComp_13_port, OUT1(12) => 
                           AtoComp_12_port, OUT1(11) => AtoComp_11_port, 
                           OUT1(10) => AtoComp_10_port, OUT1(9) => 
                           AtoComp_9_port, OUT1(8) => AtoComp_8_port, OUT1(7) 
                           => AtoComp_7_port, OUT1(6) => AtoComp_6_port, 
                           OUT1(5) => AtoComp_5_port, OUT1(4) => AtoComp_4_port
                           , OUT1(3) => AtoComp_3_port, OUT1(2) => 
                           AtoComp_2_port, OUT1(1) => AtoComp_1_port, OUT1(0) 
                           => AtoComp_0_port, OUT2(31) => dummy_B_31_port, 
                           OUT2(30) => dummy_B_30_port, OUT2(29) => 
                           dummy_B_29_port, OUT2(28) => dummy_B_28_port, 
                           OUT2(27) => dummy_B_27_port, OUT2(26) => 
                           dummy_B_26_port, OUT2(25) => dummy_B_25_port, 
                           OUT2(24) => dummy_B_24_port, OUT2(23) => 
                           dummy_B_23_port, OUT2(22) => dummy_B_22_port, 
                           OUT2(21) => dummy_B_21_port, OUT2(20) => 
                           dummy_B_20_port, OUT2(19) => dummy_B_19_port, 
                           OUT2(18) => dummy_B_18_port, OUT2(17) => 
                           dummy_B_17_port, OUT2(16) => dummy_B_16_port, 
                           OUT2(15) => dummy_B_15_port, OUT2(14) => 
                           dummy_B_14_port, OUT2(13) => dummy_B_13_port, 
                           OUT2(12) => dummy_B_12_port, OUT2(11) => 
                           dummy_B_11_port, OUT2(10) => dummy_B_10_port, 
                           OUT2(9) => dummy_B_9_port, OUT2(8) => dummy_B_8_port
                           , OUT2(7) => dummy_B_7_port, OUT2(6) => 
                           dummy_B_6_port, OUT2(5) => dummy_B_5_port, OUT2(4) 
                           => dummy_B_4_port, OUT2(3) => dummy_B_3_port, 
                           OUT2(2) => dummy_B_2_port, OUT2(1) => dummy_B_1_port
                           , OUT2(0) => dummy_B_0_port);
   UDECODE_REGS : decode_regs port map( A_i(31) => AtoComp_31_port, A_i(30) => 
                           AtoComp_30_port, A_i(29) => AtoComp_29_port, A_i(28)
                           => AtoComp_28_port, A_i(27) => AtoComp_27_port, 
                           A_i(26) => AtoComp_26_port, A_i(25) => 
                           AtoComp_25_port, A_i(24) => AtoComp_24_port, A_i(23)
                           => AtoComp_23_port, A_i(22) => AtoComp_22_port, 
                           A_i(21) => AtoComp_21_port, A_i(20) => 
                           AtoComp_20_port, A_i(19) => AtoComp_19_port, A_i(18)
                           => AtoComp_18_port, A_i(17) => AtoComp_17_port, 
                           A_i(16) => AtoComp_16_port, A_i(15) => 
                           AtoComp_15_port, A_i(14) => AtoComp_14_port, A_i(13)
                           => AtoComp_13_port, A_i(12) => AtoComp_12_port, 
                           A_i(11) => AtoComp_11_port, A_i(10) => 
                           AtoComp_10_port, A_i(9) => AtoComp_9_port, A_i(8) =>
                           AtoComp_8_port, A_i(7) => AtoComp_7_port, A_i(6) => 
                           AtoComp_6_port, A_i(5) => AtoComp_5_port, A_i(4) => 
                           AtoComp_4_port, A_i(3) => AtoComp_3_port, A_i(2) => 
                           AtoComp_2_port, A_i(1) => AtoComp_1_port, A_i(0) => 
                           AtoComp_0_port, B_i(31) => dummy_B_31_port, B_i(30) 
                           => dummy_B_30_port, B_i(29) => dummy_B_29_port, 
                           B_i(28) => dummy_B_28_port, B_i(27) => 
                           dummy_B_27_port, B_i(26) => dummy_B_26_port, B_i(25)
                           => dummy_B_25_port, B_i(24) => dummy_B_24_port, 
                           B_i(23) => dummy_B_23_port, B_i(22) => 
                           dummy_B_22_port, B_i(21) => dummy_B_21_port, B_i(20)
                           => dummy_B_20_port, B_i(19) => dummy_B_19_port, 
                           B_i(18) => dummy_B_18_port, B_i(17) => 
                           dummy_B_17_port, B_i(16) => dummy_B_16_port, B_i(15)
                           => dummy_B_15_port, B_i(14) => dummy_B_14_port, 
                           B_i(13) => dummy_B_13_port, B_i(12) => 
                           dummy_B_12_port, B_i(11) => dummy_B_11_port, B_i(10)
                           => dummy_B_10_port, B_i(9) => dummy_B_9_port, B_i(8)
                           => dummy_B_8_port, B_i(7) => dummy_B_7_port, B_i(6) 
                           => dummy_B_6_port, B_i(5) => dummy_B_5_port, B_i(4) 
                           => dummy_B_4_port, B_i(3) => dummy_B_3_port, B_i(2) 
                           => dummy_B_2_port, B_i(1) => dummy_B_1_port, B_i(0) 
                           => dummy_B_0_port, rA_i(4) => rA2reg_4_port, rA_i(3)
                           => rA2reg_3_port, rA_i(2) => rA2reg_2_port, rA_i(1) 
                           => rA2reg_1_port, rA_i(0) => rA2reg_0_port, rB_i(4) 
                           => rB2reg_4_port, rB_i(3) => rB2reg_3_port, rB_i(2) 
                           => rB2reg_2_port, rB_i(1) => rB2reg_1_port, rB_i(0) 
                           => rB2reg_0_port, rC_i(4) => rC2reg_4_port, rC_i(3) 
                           => rC2reg_3_port, rC_i(2) => rC2reg_2_port, rC_i(1) 
                           => rC2reg_1_port, rC_i(0) => rC2reg_0_port, 
                           IMM_i(31) => help_IMM_31_port, IMM_i(30) => 
                           help_IMM_30_port, IMM_i(29) => help_IMM_29_port, 
                           IMM_i(28) => help_IMM_28_port, IMM_i(27) => 
                           help_IMM_27_port, IMM_i(26) => help_IMM_26_port, 
                           IMM_i(25) => help_IMM_25_port, IMM_i(24) => 
                           help_IMM_24_port, IMM_i(23) => help_IMM_23_port, 
                           IMM_i(22) => help_IMM_22_port, IMM_i(21) => 
                           help_IMM_21_port, IMM_i(20) => help_IMM_20_port, 
                           IMM_i(19) => help_IMM_19_port, IMM_i(18) => 
                           help_IMM_18_port, IMM_i(17) => help_IMM_17_port, 
                           IMM_i(16) => help_IMM_16_port, IMM_i(15) => 
                           help_IMM_15_port, IMM_i(14) => help_IMM_14_port, 
                           IMM_i(13) => help_IMM_13_port, IMM_i(12) => 
                           help_IMM_12_port, IMM_i(11) => help_IMM_11_port, 
                           IMM_i(10) => help_IMM_10_port, IMM_i(9) => 
                           help_IMM_9_port, IMM_i(8) => help_IMM_8_port, 
                           IMM_i(7) => help_IMM_7_port, IMM_i(6) => 
                           help_IMM_6_port, IMM_i(5) => help_IMM_5_port, 
                           IMM_i(4) => help_IMM_4_port, IMM_i(3) => 
                           help_IMM_3_port, IMM_i(2) => help_IMM_2_port, 
                           IMM_i(1) => help_IMM_1_port, IMM_i(0) => 
                           help_IMM_0_port, ALUW_i(12) => ALUW_dec_12_port, 
                           ALUW_i(11) => ALUW_dec_11_port, ALUW_i(10) => 
                           ALUW_dec_10_port, ALUW_i(9) => ALUW_dec_9_port, 
                           ALUW_i(8) => ALUW_dec_8_port, ALUW_i(7) => 
                           ALUW_dec_7_port, ALUW_i(6) => ALUW_dec_6_port, 
                           ALUW_i(5) => ALUW_dec_5_port, ALUW_i(4) => 
                           ALUW_dec_4_port, ALUW_i(3) => ALUW_dec_3_port, 
                           ALUW_i(2) => ALUW_dec_2_port, ALUW_i(1) => 
                           ALUW_dec_1_port, ALUW_i(0) => ALUW_dec_0_port, 
                           A_o(31) => A2exe_31_port, A_o(30) => A2exe_30_port, 
                           A_o(29) => A2exe_29_port, A_o(28) => A2exe_28_port, 
                           A_o(27) => A2exe_27_port, A_o(26) => A2exe_26_port, 
                           A_o(25) => A2exe_25_port, A_o(24) => A2exe_24_port, 
                           A_o(23) => A2exe_23_port, A_o(22) => A2exe_22_port, 
                           A_o(21) => A2exe_21_port, A_o(20) => A2exe_20_port, 
                           A_o(19) => A2exe_19_port, A_o(18) => A2exe_18_port, 
                           A_o(17) => A2exe_17_port, A_o(16) => A2exe_16_port, 
                           A_o(15) => A2exe_15_port, A_o(14) => A2exe_14_port, 
                           A_o(13) => A2exe_13_port, A_o(12) => A2exe_12_port, 
                           A_o(11) => A2exe_11_port, A_o(10) => A2exe_10_port, 
                           A_o(9) => A2exe_9_port, A_o(8) => A2exe_8_port, 
                           A_o(7) => A2exe_7_port, A_o(6) => A2exe_6_port, 
                           A_o(5) => A2exe_5_port, A_o(4) => A2exe_4_port, 
                           A_o(3) => A2exe_3_port, A_o(2) => A2exe_2_port, 
                           A_o(1) => A2exe_1_port, A_o(0) => A2exe_0_port, 
                           B_o(31) => B2exe_31_port, B_o(30) => B2exe_30_port, 
                           B_o(29) => B2exe_29_port, B_o(28) => B2exe_28_port, 
                           B_o(27) => B2exe_27_port, B_o(26) => B2exe_26_port, 
                           B_o(25) => B2exe_25_port, B_o(24) => B2exe_24_port, 
                           B_o(23) => B2exe_23_port, B_o(22) => B2exe_22_port, 
                           B_o(21) => B2exe_21_port, B_o(20) => B2exe_20_port, 
                           B_o(19) => B2exe_19_port, B_o(18) => B2exe_18_port, 
                           B_o(17) => B2exe_17_port, B_o(16) => B2exe_16_port, 
                           B_o(15) => B2exe_15_port, B_o(14) => B2exe_14_port, 
                           B_o(13) => B2exe_13_port, B_o(12) => B2exe_12_port, 
                           B_o(11) => B2exe_11_port, B_o(10) => B2exe_10_port, 
                           B_o(9) => B2exe_9_port, B_o(8) => B2exe_8_port, 
                           B_o(7) => B2exe_7_port, B_o(6) => B2exe_6_port, 
                           B_o(5) => B2exe_5_port, B_o(4) => B2exe_4_port, 
                           B_o(3) => B2exe_3_port, B_o(2) => B2exe_2_port, 
                           B_o(1) => B2exe_1_port, B_o(0) => B2exe_0_port, 
                           rA_o(4) => rA2fw_4_port, rA_o(3) => rA2fw_3_port, 
                           rA_o(2) => rA2fw_2_port, rA_o(1) => rA2fw_1_port, 
                           rA_o(0) => rA2fw_0_port, rB_o(4) => rB2mux_4_port, 
                           rB_o(3) => rB2mux_3_port, rB_o(2) => rB2mux_2_port, 
                           rB_o(1) => rB2mux_1_port, rB_o(0) => rB2mux_0_port, 
                           rC_o(4) => rC2mux_4_port, rC_o(3) => rC2mux_3_port, 
                           rC_o(2) => rC2mux_2_port, rC_o(1) => rC2mux_1_port, 
                           rC_o(0) => rC2mux_0_port, IMM_o(31) => 
                           IMM2exe_31_port, IMM_o(30) => IMM2exe_30_port, 
                           IMM_o(29) => IMM2exe_29_port, IMM_o(28) => 
                           IMM2exe_28_port, IMM_o(27) => IMM2exe_27_port, 
                           IMM_o(26) => IMM2exe_26_port, IMM_o(25) => 
                           IMM2exe_25_port, IMM_o(24) => IMM2exe_24_port, 
                           IMM_o(23) => IMM2exe_23_port, IMM_o(22) => 
                           IMM2exe_22_port, IMM_o(21) => IMM2exe_21_port, 
                           IMM_o(20) => IMM2exe_20_port, IMM_o(19) => 
                           IMM2exe_19_port, IMM_o(18) => IMM2exe_18_port, 
                           IMM_o(17) => IMM2exe_17_port, IMM_o(16) => 
                           IMM2exe_16_port, IMM_o(15) => IMM2exe_15_port, 
                           IMM_o(14) => IMM2exe_14_port, IMM_o(13) => 
                           IMM2exe_13_port, IMM_o(12) => IMM2exe_12_port, 
                           IMM_o(11) => IMM2exe_11_port, IMM_o(10) => 
                           IMM2exe_10_port, IMM_o(9) => IMM2exe_9_port, 
                           IMM_o(8) => IMM2exe_8_port, IMM_o(7) => 
                           IMM2exe_7_port, IMM_o(6) => IMM2exe_6_port, IMM_o(5)
                           => IMM2exe_5_port, IMM_o(4) => IMM2exe_4_port, 
                           IMM_o(3) => IMM2exe_3_port, IMM_o(2) => 
                           IMM2exe_2_port, IMM_o(1) => IMM2exe_1_port, IMM_o(0)
                           => IMM2exe_0_port, ALUW_o(12) => ALUW_12_port, 
                           ALUW_o(11) => ALUW_11_port, ALUW_o(10) => 
                           ALUW_10_port, ALUW_o(9) => ALUW_9_port, ALUW_o(8) =>
                           ALUW_8_port, ALUW_o(7) => ALUW_7_port, ALUW_o(6) => 
                           ALUW_6_port, ALUW_o(5) => ALUW_5_port, ALUW_o(4) => 
                           ALUW_4_port, ALUW_o(3) => ALUW_3_port, ALUW_o(2) => 
                           ALUW_2_port, ALUW_o(1) => ALUW_1_port, ALUW_o(0) => 
                           ALUW_0_port, stall_i => stall_exe, clk => clock, rst
                           => rst);
   UEXECUTE_REGS : execute_regs port map( X_i(31) => X2mem_31_port, X_i(30) => 
                           X2mem_30_port, X_i(29) => X2mem_29_port, X_i(28) => 
                           X2mem_28_port, X_i(27) => X2mem_27_port, X_i(26) => 
                           X2mem_26_port, X_i(25) => X2mem_25_port, X_i(24) => 
                           X2mem_24_port, X_i(23) => X2mem_23_port, X_i(22) => 
                           X2mem_22_port, X_i(21) => X2mem_21_port, X_i(20) => 
                           X2mem_20_port, X_i(19) => X2mem_19_port, X_i(18) => 
                           X2mem_18_port, X_i(17) => X2mem_17_port, X_i(16) => 
                           X2mem_16_port, X_i(15) => X2mem_15_port, X_i(14) => 
                           X2mem_14_port, X_i(13) => X2mem_13_port, X_i(12) => 
                           X2mem_12_port, X_i(11) => X2mem_11_port, X_i(10) => 
                           X2mem_10_port, X_i(9) => X2mem_9_port, X_i(8) => 
                           X2mem_8_port, X_i(7) => X2mem_7_port, X_i(6) => 
                           X2mem_6_port, X_i(5) => X2mem_5_port, X_i(4) => 
                           X2mem_4_port, X_i(3) => X2mem_3_port, X_i(2) => 
                           X2mem_2_port, X_i(1) => X2mem_1_port, X_i(0) => 
                           X2mem_0_port, S_i(31) => S2mem_31_port, S_i(30) => 
                           S2mem_30_port, S_i(29) => S2mem_29_port, S_i(28) => 
                           S2mem_28_port, S_i(27) => S2mem_27_port, S_i(26) => 
                           S2mem_26_port, S_i(25) => S2mem_25_port, S_i(24) => 
                           S2mem_24_port, S_i(23) => S2mem_23_port, S_i(22) => 
                           S2mem_22_port, S_i(21) => S2mem_21_port, S_i(20) => 
                           S2mem_20_port, S_i(19) => S2mem_19_port, S_i(18) => 
                           S2mem_18_port, S_i(17) => S2mem_17_port, S_i(16) => 
                           S2mem_16_port, S_i(15) => S2mem_15_port, S_i(14) => 
                           S2mem_14_port, S_i(13) => S2mem_13_port, S_i(12) => 
                           S2mem_12_port, S_i(11) => S2mem_11_port, S_i(10) => 
                           S2mem_10_port, S_i(9) => S2mem_9_port, S_i(8) => 
                           S2mem_8_port, S_i(7) => S2mem_7_port, S_i(6) => 
                           S2mem_6_port, S_i(5) => S2mem_5_port, S_i(4) => 
                           S2mem_4_port, S_i(3) => n9, S_i(2) => S2mem_2_port, 
                           S_i(1) => S2mem_1_port, S_i(0) => n8, D2_i(4) => 
                           muxed_dest2exe_4_port, D2_i(3) => 
                           muxed_dest2exe_3_port, D2_i(2) => 
                           muxed_dest2exe_2_port, D2_i(1) => 
                           muxed_dest2exe_1_port, D2_i(0) => 
                           muxed_dest2exe_0_port, X_o(31) => 
                           DRAM_Addr_o_31_port, X_o(30) => DRAM_Addr_o_30_port,
                           X_o(29) => DRAM_Addr_o_29_port, X_o(28) => 
                           DRAM_Addr_o_28_port, X_o(27) => DRAM_Addr_o_27_port,
                           X_o(26) => DRAM_Addr_o_26_port, X_o(25) => 
                           DRAM_Addr_o_25_port, X_o(24) => DRAM_Addr_o_24_port,
                           X_o(23) => DRAM_Addr_o_23_port, X_o(22) => 
                           DRAM_Addr_o_22_port, X_o(21) => DRAM_Addr_o_21_port,
                           X_o(20) => DRAM_Addr_o_20_port, X_o(19) => 
                           DRAM_Addr_o_19_port, X_o(18) => DRAM_Addr_o_18_port,
                           X_o(17) => DRAM_Addr_o_17_port, X_o(16) => 
                           DRAM_Addr_o_16_port, X_o(15) => DRAM_Addr_o_15_port,
                           X_o(14) => DRAM_Addr_o_14_port, X_o(13) => 
                           DRAM_Addr_o_13_port, X_o(12) => DRAM_Addr_o_12_port,
                           X_o(11) => DRAM_Addr_o_11_port, X_o(10) => 
                           DRAM_Addr_o_10_port, X_o(9) => DRAM_Addr_o_9_port, 
                           X_o(8) => DRAM_Addr_o_8_port, X_o(7) => 
                           DRAM_Addr_o_7_port, X_o(6) => DRAM_Addr_o_6_port, 
                           X_o(5) => DRAM_Addr_o_5_port, X_o(4) => 
                           DRAM_Addr_o_4_port, X_o(3) => DRAM_Addr_o_3_port, 
                           X_o(2) => DRAM_Addr_o_2_port, X_o(1) => 
                           DRAM_Addr_o_1_port, X_o(0) => DRAM_Addr_o_0_port, 
                           S_o(31) => DRAM_Din_o(31), S_o(30) => DRAM_Din_o(30)
                           , S_o(29) => DRAM_Din_o(29), S_o(28) => 
                           DRAM_Din_o(28), S_o(27) => DRAM_Din_o(27), S_o(26) 
                           => DRAM_Din_o(26), S_o(25) => DRAM_Din_o(25), 
                           S_o(24) => DRAM_Din_o(24), S_o(23) => DRAM_Din_o(23)
                           , S_o(22) => DRAM_Din_o(22), S_o(21) => 
                           DRAM_Din_o(21), S_o(20) => DRAM_Din_o(20), S_o(19) 
                           => DRAM_Din_o(19), S_o(18) => DRAM_Din_o(18), 
                           S_o(17) => DRAM_Din_o(17), S_o(16) => DRAM_Din_o(16)
                           , S_o(15) => DRAM_Din_o(15), S_o(14) => 
                           DRAM_Din_o(14), S_o(13) => DRAM_Din_o(13), S_o(12) 
                           => DRAM_Din_o(12), S_o(11) => DRAM_Din_o(11), 
                           S_o(10) => DRAM_Din_o(10), S_o(9) => DRAM_Din_o(9), 
                           S_o(8) => DRAM_Din_o(8), S_o(7) => DRAM_Din_o(7), 
                           S_o(6) => DRAM_Din_o(6), S_o(5) => DRAM_Din_o(5), 
                           S_o(4) => DRAM_Din_o(4), S_o(3) => DRAM_Din_o(3), 
                           S_o(2) => DRAM_Din_o(2), S_o(1) => DRAM_Din_o(1), 
                           S_o(0) => DRAM_Din_o(0), D2_o(4) => D22D3_4_port, 
                           D2_o(3) => D22D3_3_port, D2_o(2) => D22D3_2_port, 
                           D2_o(1) => D22D3_1_port, D2_o(0) => D22D3_0_port, 
                           stall_i => X_Logic0_port, clk => clock, rst => rst);
   UEXECUTE_BLOCK : execute_block port map( IMM_i(31) => IMM2exe_31_port, 
                           IMM_i(30) => IMM2exe_30_port, IMM_i(29) => 
                           IMM2exe_29_port, IMM_i(28) => IMM2exe_28_port, 
                           IMM_i(27) => IMM2exe_27_port, IMM_i(26) => 
                           IMM2exe_26_port, IMM_i(25) => IMM2exe_25_port, 
                           IMM_i(24) => IMM2exe_24_port, IMM_i(23) => 
                           IMM2exe_23_port, IMM_i(22) => IMM2exe_22_port, 
                           IMM_i(21) => IMM2exe_21_port, IMM_i(20) => 
                           IMM2exe_20_port, IMM_i(19) => IMM2exe_19_port, 
                           IMM_i(18) => IMM2exe_18_port, IMM_i(17) => 
                           IMM2exe_17_port, IMM_i(16) => IMM2exe_16_port, 
                           IMM_i(15) => IMM2exe_15_port, IMM_i(14) => 
                           IMM2exe_14_port, IMM_i(13) => IMM2exe_13_port, 
                           IMM_i(12) => IMM2exe_12_port, IMM_i(11) => 
                           IMM2exe_11_port, IMM_i(10) => IMM2exe_10_port, 
                           IMM_i(9) => IMM2exe_9_port, IMM_i(8) => 
                           IMM2exe_8_port, IMM_i(7) => IMM2exe_7_port, IMM_i(6)
                           => IMM2exe_6_port, IMM_i(5) => IMM2exe_5_port, 
                           IMM_i(4) => IMM2exe_4_port, IMM_i(3) => 
                           IMM2exe_3_port, IMM_i(2) => IMM2exe_2_port, IMM_i(1)
                           => IMM2exe_1_port, IMM_i(0) => IMM2exe_0_port, 
                           A_i(31) => A2exe_31_port, A_i(30) => A2exe_30_port, 
                           A_i(29) => A2exe_29_port, A_i(28) => A2exe_28_port, 
                           A_i(27) => A2exe_27_port, A_i(26) => A2exe_26_port, 
                           A_i(25) => A2exe_25_port, A_i(24) => A2exe_24_port, 
                           A_i(23) => A2exe_23_port, A_i(22) => A2exe_22_port, 
                           A_i(21) => A2exe_21_port, A_i(20) => A2exe_20_port, 
                           A_i(19) => A2exe_19_port, A_i(18) => A2exe_18_port, 
                           A_i(17) => A2exe_17_port, A_i(16) => A2exe_16_port, 
                           A_i(15) => A2exe_15_port, A_i(14) => A2exe_14_port, 
                           A_i(13) => A2exe_13_port, A_i(12) => A2exe_12_port, 
                           A_i(11) => A2exe_11_port, A_i(10) => A2exe_10_port, 
                           A_i(9) => A2exe_9_port, A_i(8) => A2exe_8_port, 
                           A_i(7) => A2exe_7_port, A_i(6) => A2exe_6_port, 
                           A_i(5) => A2exe_5_port, A_i(4) => A2exe_4_port, 
                           A_i(3) => A2exe_3_port, A_i(2) => A2exe_2_port, 
                           A_i(1) => A2exe_1_port, A_i(0) => A2exe_0_port, 
                           rB_i(4) => rB2mux_4_port, rB_i(3) => rB2mux_3_port, 
                           rB_i(2) => rB2mux_2_port, rB_i(1) => rB2mux_1_port, 
                           rB_i(0) => rB2mux_0_port, rC_i(4) => rC2mux_4_port, 
                           rC_i(3) => rC2mux_3_port, rC_i(2) => rC2mux_2_port, 
                           rC_i(1) => rC2mux_1_port, rC_i(0) => rC2mux_0_port, 
                           MUXED_B_i(31) => B2exe_31_port, MUXED_B_i(30) => 
                           B2exe_30_port, MUXED_B_i(29) => B2exe_29_port, 
                           MUXED_B_i(28) => B2exe_28_port, MUXED_B_i(27) => 
                           B2exe_27_port, MUXED_B_i(26) => B2exe_26_port, 
                           MUXED_B_i(25) => B2exe_25_port, MUXED_B_i(24) => 
                           B2exe_24_port, MUXED_B_i(23) => B2exe_23_port, 
                           MUXED_B_i(22) => B2exe_22_port, MUXED_B_i(21) => 
                           B2exe_21_port, MUXED_B_i(20) => B2exe_20_port, 
                           MUXED_B_i(19) => B2exe_19_port, MUXED_B_i(18) => 
                           B2exe_18_port, MUXED_B_i(17) => B2exe_17_port, 
                           MUXED_B_i(16) => B2exe_16_port, MUXED_B_i(15) => 
                           B2exe_15_port, MUXED_B_i(14) => B2exe_14_port, 
                           MUXED_B_i(13) => B2exe_13_port, MUXED_B_i(12) => 
                           B2exe_12_port, MUXED_B_i(11) => B2exe_11_port, 
                           MUXED_B_i(10) => B2exe_10_port, MUXED_B_i(9) => 
                           B2exe_9_port, MUXED_B_i(8) => B2exe_8_port, 
                           MUXED_B_i(7) => B2exe_7_port, MUXED_B_i(6) => 
                           B2exe_6_port, MUXED_B_i(5) => B2exe_5_port, 
                           MUXED_B_i(4) => B2exe_4_port, MUXED_B_i(3) => 
                           B2exe_3_port, MUXED_B_i(2) => B2exe_2_port, 
                           MUXED_B_i(1) => B2exe_1_port, MUXED_B_i(0) => 
                           B2exe_0_port, S_MUX_ALUIN_i => dummy_S_MUX_ALUIN, 
                           FW_X_i(31) => DRAM_Addr_o_31_port, FW_X_i(30) => 
                           DRAM_Addr_o_30_port, FW_X_i(29) => 
                           DRAM_Addr_o_29_port, FW_X_i(28) => 
                           DRAM_Addr_o_28_port, FW_X_i(27) => 
                           DRAM_Addr_o_27_port, FW_X_i(26) => 
                           DRAM_Addr_o_26_port, FW_X_i(25) => 
                           DRAM_Addr_o_25_port, FW_X_i(24) => 
                           DRAM_Addr_o_24_port, FW_X_i(23) => 
                           DRAM_Addr_o_23_port, FW_X_i(22) => 
                           DRAM_Addr_o_22_port, FW_X_i(21) => 
                           DRAM_Addr_o_21_port, FW_X_i(20) => 
                           DRAM_Addr_o_20_port, FW_X_i(19) => 
                           DRAM_Addr_o_19_port, FW_X_i(18) => 
                           DRAM_Addr_o_18_port, FW_X_i(17) => 
                           DRAM_Addr_o_17_port, FW_X_i(16) => 
                           DRAM_Addr_o_16_port, FW_X_i(15) => 
                           DRAM_Addr_o_15_port, FW_X_i(14) => 
                           DRAM_Addr_o_14_port, FW_X_i(13) => 
                           DRAM_Addr_o_13_port, FW_X_i(12) => 
                           DRAM_Addr_o_12_port, FW_X_i(11) => 
                           DRAM_Addr_o_11_port, FW_X_i(10) => 
                           DRAM_Addr_o_10_port, FW_X_i(9) => DRAM_Addr_o_9_port
                           , FW_X_i(8) => DRAM_Addr_o_8_port, FW_X_i(7) => 
                           DRAM_Addr_o_7_port, FW_X_i(6) => DRAM_Addr_o_6_port,
                           FW_X_i(5) => DRAM_Addr_o_5_port, FW_X_i(4) => 
                           DRAM_Addr_o_4_port, FW_X_i(3) => DRAM_Addr_o_3_port,
                           FW_X_i(2) => DRAM_Addr_o_2_port, FW_X_i(1) => 
                           DRAM_Addr_o_1_port, FW_X_i(0) => DRAM_Addr_o_0_port,
                           FW_W_i(31) => wb2reg_31_port, FW_W_i(30) => 
                           wb2reg_30_port, FW_W_i(29) => wb2reg_29_port, 
                           FW_W_i(28) => wb2reg_28_port, FW_W_i(27) => 
                           wb2reg_27_port, FW_W_i(26) => wb2reg_26_port, 
                           FW_W_i(25) => wb2reg_25_port, FW_W_i(24) => 
                           wb2reg_24_port, FW_W_i(23) => wb2reg_23_port, 
                           FW_W_i(22) => wb2reg_22_port, FW_W_i(21) => 
                           wb2reg_21_port, FW_W_i(20) => wb2reg_20_port, 
                           FW_W_i(19) => wb2reg_19_port, FW_W_i(18) => 
                           wb2reg_18_port, FW_W_i(17) => wb2reg_17_port, 
                           FW_W_i(16) => wb2reg_16_port, FW_W_i(15) => 
                           wb2reg_15_port, FW_W_i(14) => wb2reg_14_port, 
                           FW_W_i(13) => wb2reg_13_port, FW_W_i(12) => 
                           wb2reg_12_port, FW_W_i(11) => wb2reg_11_port, 
                           FW_W_i(10) => wb2reg_10_port, FW_W_i(9) => 
                           wb2reg_9_port, FW_W_i(8) => wb2reg_8_port, FW_W_i(7)
                           => wb2reg_7_port, FW_W_i(6) => wb2reg_6_port, 
                           FW_W_i(5) => wb2reg_5_port, FW_W_i(4) => 
                           wb2reg_4_port, FW_W_i(3) => wb2reg_3_port, FW_W_i(2)
                           => wb2reg_2_port, FW_W_i(1) => wb2reg_1_port, 
                           FW_W_i(0) => wb2reg_0_port, S_FW_A_i(1) => 
                           dummy_S_FWA2exe_1_port, S_FW_A_i(0) => n13, 
                           S_FW_B_i(1) => dummy_S_FWB2exe_1_port, S_FW_B_i(0) 
                           => dummy_S_FWB2exe_0_port, muxed_dest(4) => 
                           muxed_dest2exe_4_port, muxed_dest(3) => 
                           muxed_dest2exe_3_port, muxed_dest(2) => 
                           muxed_dest2exe_2_port, muxed_dest(1) => 
                           muxed_dest2exe_1_port, muxed_dest(0) => 
                           muxed_dest2exe_0_port, muxed_B(31) => S2mem_31_port,
                           muxed_B(30) => S2mem_30_port, muxed_B(29) => 
                           S2mem_29_port, muxed_B(28) => S2mem_28_port, 
                           muxed_B(27) => S2mem_27_port, muxed_B(26) => 
                           S2mem_26_port, muxed_B(25) => S2mem_25_port, 
                           muxed_B(24) => S2mem_24_port, muxed_B(23) => 
                           S2mem_23_port, muxed_B(22) => S2mem_22_port, 
                           muxed_B(21) => S2mem_21_port, muxed_B(20) => 
                           S2mem_20_port, muxed_B(19) => S2mem_19_port, 
                           muxed_B(18) => S2mem_18_port, muxed_B(17) => 
                           S2mem_17_port, muxed_B(16) => S2mem_16_port, 
                           muxed_B(15) => S2mem_15_port, muxed_B(14) => 
                           S2mem_14_port, muxed_B(13) => S2mem_13_port, 
                           muxed_B(12) => S2mem_12_port, muxed_B(11) => 
                           S2mem_11_port, muxed_B(10) => S2mem_10_port, 
                           muxed_B(9) => S2mem_9_port, muxed_B(8) => 
                           S2mem_8_port, muxed_B(7) => S2mem_7_port, muxed_B(6)
                           => S2mem_6_port, muxed_B(5) => S2mem_5_port, 
                           muxed_B(4) => S2mem_4_port, muxed_B(3) => n9, 
                           muxed_B(2) => S2mem_2_port, muxed_B(1) => 
                           S2mem_1_port, muxed_B(0) => n8, S_MUX_DEST_i(1) => 
                           dummy_S_MUX_DEST_1_port, S_MUX_DEST_i(0) => 
                           dummy_S_MUX_DEST_0_port, OP(0) => n34, OP(1) => n35,
                           OP(2) => n36, OP(3) => n37, OP(4) => n38, ALUW_i(12)
                           => ALUW_12_port, ALUW_i(11) => ALUW_11_port, 
                           ALUW_i(10) => ALUW_10_port, ALUW_i(9) => ALUW_9_port
                           , ALUW_i(8) => ALUW_8_port, ALUW_i(7) => ALUW_7_port
                           , ALUW_i(6) => ALUW_6_port, ALUW_i(5) => ALUW_5_port
                           , ALUW_i(4) => ALUW_4_port, ALUW_i(3) => ALUW_3_port
                           , ALUW_i(2) => ALUW_2_port, ALUW_i(1) => ALUW_1_port
                           , ALUW_i(0) => ALUW_0_port, DOUT(31) => 
                           X2mem_31_port, DOUT(30) => X2mem_30_port, DOUT(29) 
                           => X2mem_29_port, DOUT(28) => X2mem_28_port, 
                           DOUT(27) => X2mem_27_port, DOUT(26) => X2mem_26_port
                           , DOUT(25) => X2mem_25_port, DOUT(24) => 
                           X2mem_24_port, DOUT(23) => X2mem_23_port, DOUT(22) 
                           => X2mem_22_port, DOUT(21) => X2mem_21_port, 
                           DOUT(20) => X2mem_20_port, DOUT(19) => X2mem_19_port
                           , DOUT(18) => X2mem_18_port, DOUT(17) => 
                           X2mem_17_port, DOUT(16) => X2mem_16_port, DOUT(15) 
                           => X2mem_15_port, DOUT(14) => X2mem_14_port, 
                           DOUT(13) => X2mem_13_port, DOUT(12) => X2mem_12_port
                           , DOUT(11) => X2mem_11_port, DOUT(10) => 
                           X2mem_10_port, DOUT(9) => X2mem_9_port, DOUT(8) => 
                           X2mem_8_port, DOUT(7) => X2mem_7_port, DOUT(6) => 
                           X2mem_6_port, DOUT(5) => X2mem_5_port, DOUT(4) => 
                           X2mem_4_port, DOUT(3) => X2mem_3_port, DOUT(2) => 
                           X2mem_2_port, DOUT(1) => X2mem_1_port, DOUT(0) => 
                           X2mem_0_port, stall_o => exe_stall_cu, Clock => 
                           clock, Reset => rst);
   UMEM_REGS : mem_regs port map( W_i(31) => W2wb_31_port, W_i(30) => 
                           W2wb_30_port, W_i(29) => W2wb_29_port, W_i(28) => 
                           W2wb_28_port, W_i(27) => W2wb_27_port, W_i(26) => 
                           W2wb_26_port, W_i(25) => W2wb_25_port, W_i(24) => 
                           W2wb_24_port, W_i(23) => W2wb_23_port, W_i(22) => 
                           W2wb_22_port, W_i(21) => W2wb_21_port, W_i(20) => 
                           W2wb_20_port, W_i(19) => W2wb_19_port, W_i(18) => 
                           W2wb_18_port, W_i(17) => W2wb_17_port, W_i(16) => 
                           W2wb_16_port, W_i(15) => W2wb_15_port, W_i(14) => 
                           W2wb_14_port, W_i(13) => W2wb_13_port, W_i(12) => 
                           W2wb_12_port, W_i(11) => W2wb_11_port, W_i(10) => 
                           W2wb_10_port, W_i(9) => W2wb_9_port, W_i(8) => 
                           W2wb_8_port, W_i(7) => W2wb_7_port, W_i(6) => 
                           W2wb_6_port, W_i(5) => W2wb_5_port, W_i(4) => 
                           W2wb_4_port, W_i(3) => W2wb_3_port, W_i(2) => 
                           W2wb_2_port, W_i(1) => W2wb_1_port, W_i(0) => 
                           W2wb_0_port, D3_i(4) => D22D3_4_port, D3_i(3) => n19
                           , D3_i(2) => n20, D3_i(1) => n17, D3_i(0) => n18, 
                           W_o(31) => wb2reg_31_port, W_o(30) => wb2reg_30_port
                           , W_o(29) => wb2reg_29_port, W_o(28) => 
                           wb2reg_28_port, W_o(27) => wb2reg_27_port, W_o(26) 
                           => wb2reg_26_port, W_o(25) => wb2reg_25_port, 
                           W_o(24) => wb2reg_24_port, W_o(23) => wb2reg_23_port
                           , W_o(22) => wb2reg_22_port, W_o(21) => 
                           wb2reg_21_port, W_o(20) => wb2reg_20_port, W_o(19) 
                           => wb2reg_19_port, W_o(18) => wb2reg_18_port, 
                           W_o(17) => wb2reg_17_port, W_o(16) => wb2reg_16_port
                           , W_o(15) => wb2reg_15_port, W_o(14) => 
                           wb2reg_14_port, W_o(13) => wb2reg_13_port, W_o(12) 
                           => wb2reg_12_port, W_o(11) => wb2reg_11_port, 
                           W_o(10) => wb2reg_10_port, W_o(9) => wb2reg_9_port, 
                           W_o(8) => wb2reg_8_port, W_o(7) => wb2reg_7_port, 
                           W_o(6) => wb2reg_6_port, W_o(5) => wb2reg_5_port, 
                           W_o(4) => wb2reg_4_port, W_o(3) => wb2reg_3_port, 
                           W_o(2) => wb2reg_2_port, W_o(1) => wb2reg_1_port, 
                           W_o(0) => wb2reg_0_port, D3_o(4) => D32reg_4_port, 
                           D3_o(3) => D32reg_3_port, D3_o(2) => D32reg_2_port, 
                           D3_o(1) => D32reg_1_port, D3_o(0) => D32reg_0_port, 
                           clk => clock, rst => rst);
   UMEM_BLOCK : mem_block port map( X_i(31) => DRAM_Addr_o_31_port, X_i(30) => 
                           DRAM_Addr_o_30_port, X_i(29) => DRAM_Addr_o_29_port,
                           X_i(28) => DRAM_Addr_o_28_port, X_i(27) => 
                           DRAM_Addr_o_27_port, X_i(26) => DRAM_Addr_o_26_port,
                           X_i(25) => DRAM_Addr_o_25_port, X_i(24) => 
                           DRAM_Addr_o_24_port, X_i(23) => DRAM_Addr_o_23_port,
                           X_i(22) => DRAM_Addr_o_22_port, X_i(21) => 
                           DRAM_Addr_o_21_port, X_i(20) => DRAM_Addr_o_20_port,
                           X_i(19) => DRAM_Addr_o_19_port, X_i(18) => 
                           DRAM_Addr_o_18_port, X_i(17) => DRAM_Addr_o_17_port,
                           X_i(16) => DRAM_Addr_o_16_port, X_i(15) => 
                           DRAM_Addr_o_15_port, X_i(14) => DRAM_Addr_o_14_port,
                           X_i(13) => DRAM_Addr_o_13_port, X_i(12) => 
                           DRAM_Addr_o_12_port, X_i(11) => DRAM_Addr_o_11_port,
                           X_i(10) => DRAM_Addr_o_10_port, X_i(9) => 
                           DRAM_Addr_o_9_port, X_i(8) => DRAM_Addr_o_8_port, 
                           X_i(7) => DRAM_Addr_o_7_port, X_i(6) => 
                           DRAM_Addr_o_6_port, X_i(5) => DRAM_Addr_o_5_port, 
                           X_i(4) => DRAM_Addr_o_4_port, X_i(3) => 
                           DRAM_Addr_o_3_port, X_i(2) => DRAM_Addr_o_2_port, 
                           X_i(1) => DRAM_Addr_o_1_port, X_i(0) => 
                           DRAM_Addr_o_0_port, LOAD_i(31) => DRAM_Dout_i(31), 
                           LOAD_i(30) => DRAM_Dout_i(30), LOAD_i(29) => 
                           DRAM_Dout_i(29), LOAD_i(28) => DRAM_Dout_i(28), 
                           LOAD_i(27) => DRAM_Dout_i(27), LOAD_i(26) => 
                           DRAM_Dout_i(26), LOAD_i(25) => DRAM_Dout_i(25), 
                           LOAD_i(24) => DRAM_Dout_i(24), LOAD_i(23) => 
                           DRAM_Dout_i(23), LOAD_i(22) => DRAM_Dout_i(22), 
                           LOAD_i(21) => DRAM_Dout_i(21), LOAD_i(20) => 
                           DRAM_Dout_i(20), LOAD_i(19) => DRAM_Dout_i(19), 
                           LOAD_i(18) => DRAM_Dout_i(18), LOAD_i(17) => 
                           DRAM_Dout_i(17), LOAD_i(16) => DRAM_Dout_i(16), 
                           LOAD_i(15) => DRAM_Dout_i(15), LOAD_i(14) => 
                           DRAM_Dout_i(14), LOAD_i(13) => DRAM_Dout_i(13), 
                           LOAD_i(12) => DRAM_Dout_i(12), LOAD_i(11) => 
                           DRAM_Dout_i(11), LOAD_i(10) => DRAM_Dout_i(10), 
                           LOAD_i(9) => DRAM_Dout_i(9), LOAD_i(8) => 
                           DRAM_Dout_i(8), LOAD_i(7) => DRAM_Dout_i(7), 
                           LOAD_i(6) => DRAM_Dout_i(6), LOAD_i(5) => 
                           DRAM_Dout_i(5), LOAD_i(4) => DRAM_Dout_i(4), 
                           LOAD_i(3) => DRAM_Dout_i(3), LOAD_i(2) => 
                           DRAM_Dout_i(2), LOAD_i(1) => DRAM_Dout_i(1), 
                           LOAD_i(0) => DRAM_Dout_i(0), W_o(31) => W2wb_31_port
                           , W_o(30) => W2wb_30_port, W_o(29) => W2wb_29_port, 
                           W_o(28) => W2wb_28_port, W_o(27) => W2wb_27_port, 
                           W_o(26) => W2wb_26_port, W_o(25) => W2wb_25_port, 
                           W_o(24) => W2wb_24_port, W_o(23) => W2wb_23_port, 
                           W_o(22) => W2wb_22_port, W_o(21) => W2wb_21_port, 
                           W_o(20) => W2wb_20_port, W_o(19) => W2wb_19_port, 
                           W_o(18) => W2wb_18_port, W_o(17) => W2wb_17_port, 
                           W_o(16) => W2wb_16_port, W_o(15) => W2wb_15_port, 
                           W_o(14) => W2wb_14_port, W_o(13) => W2wb_13_port, 
                           W_o(12) => W2wb_12_port, W_o(11) => W2wb_11_port, 
                           W_o(10) => W2wb_10_port, W_o(9) => W2wb_9_port, 
                           W_o(8) => W2wb_8_port, W_o(7) => W2wb_7_port, W_o(6)
                           => W2wb_6_port, W_o(5) => W2wb_5_port, W_o(4) => 
                           W2wb_4_port, W_o(3) => W2wb_3_port, W_o(2) => 
                           W2wb_2_port, W_o(1) => W2wb_1_port, W_o(0) => 
                           W2wb_0_port, S_MUX_MEM_i_BAR => dummy_S_MUX_MEM);
   UFW_LOGIC : fw_logic port map( D1_i(4) => n39, D1_i(3) => n40, D1_i(2) => 
                           n41, D1_i(1) => n42, D1_i(0) => n43, rAdec_i(4) => 
                           IR_25_port, rAdec_i(3) => IR_24_port, rAdec_i(2) => 
                           IR_23_port, rAdec_i(1) => IR_22_port, rAdec_i(0) => 
                           IR_21_port, D2_i(4) => D22D3_4_port, D2_i(3) => 
                           D22D3_3_port, D2_i(2) => D22D3_2_port, D2_i(1) => 
                           D22D3_1_port, D2_i(0) => D22D3_0_port, D3_i(4) => 
                           D32reg_4_port, D3_i(3) => D32reg_3_port, D3_i(2) => 
                           D32reg_2_port, D3_i(1) => D32reg_1_port, D3_i(0) => 
                           D32reg_0_port, rA_i(4) => rA2fw_4_port, rA_i(3) => 
                           rA2fw_3_port, rA_i(2) => rA2fw_2_port, rA_i(1) => 
                           rA2fw_1_port, rA_i(0) => rA2fw_0_port, rB_i(4) => 
                           rB2mux_4_port, rB_i(3) => rB2mux_3_port, rB_i(2) => 
                           rB2mux_2_port, rB_i(1) => rB2mux_1_port, rB_i(0) => 
                           rB2mux_0_port, S_mem_W => dummy_S_RF_W_mem, S_wb_W 
                           => dummy_S_RF_W_wb, S_exe_W => n44, S_FWAdec(1) => 
                           dummy_S_FWAdec_1_port, S_FWAdec(0) => 
                           dummy_S_FWAdec_0_port, S_FWA(1) => 
                           dummy_S_FWA2exe_1_port, S_FWA(0) => n13, S_FWB(1) =>
                           dummy_S_FWB2exe_1_port, S_FWB(0) => 
                           dummy_S_FWB2exe_0_port, S_mem_LOAD_BAR => 
                           dummy_S_MUX_MEM);
   U9 : INV_X2 port map( A => n7, ZN => was_taken);
   U10 : AOI21_X1 port map( B1 => was_taken_from_jl, B2 => was_branch, A => 
                           was_jmp, ZN => n7);
   U11 : INV_X1 port map( A => n12, ZN => n22);
   U12 : BUF_X1 port map( A => D22D3_0_port, Z => n18);
   U13 : CLKBUF_X1 port map( A => mispredict, Z => n21);
   U14 : BUF_X1 port map( A => D22D3_1_port, Z => n17);
   U15 : BUF_X1 port map( A => D22D3_3_port, Z => n19);
   U16 : BUF_X1 port map( A => D22D3_2_port, Z => n20);
   n23 <= '0';
   n24 <= '0';
   n25 <= '0';
   n26 <= '0';
   n27 <= '0';
   n28 <= '0';
   n29 <= '0';
   n30 <= '0';
   n31 <= '0';
   n32 <= '0';
   n33 <= '0';
   n34 <= '0';
   n35 <= '0';
   n36 <= '0';
   n37 <= '0';
   n38 <= '0';
   n39 <= '0';
   n40 <= '0';
   n41 <= '0';
   n42 <= '0';
   n43 <= '0';
   n44 <= '0';

end SYN_arch;
