
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_top_level is

-- define attributes
attribute ENUM_ENCODING : STRING;

-- define any necessary types
type aluOp is (NOP, SLLS, SRLS, SRAS, ADDS, ADDUS, SUBS, SUBUS, ANDS, ORS, 
   XORS, SEQS, SNES, SLTS, SGTS, SLES, SGES, MOVI2SS, MOVS2IS, MOVFS, MOVDS, 
   MOVFP2IS, MOVI2FP, MOVI2TS, MOVT2IS, SLTUS, SGTUS, SLEUS, SGEUS, MULTU, 
   MULTS);
attribute ENUM_ENCODING of aluOp : type is 
   "00000 00001 00010 00011 00100 00101 00110 00111 01000 01001 01010 01011 01100 01101 01110 01111 10000 10001 10010 10011 10100 10101 10110 10111 11000 11001 11010 11011 11100 11101 11110";
type UNSIGNED is array (INTEGER range <>) of std_logic;
   
   -- Declarations for conversion functions.
   function std_logic_vector_to_aluOp(arg : in std_logic_vector( 1 to 5 )) 
               return aluOp;
   function aluOp_to_std_logic_vector(arg : in aluOp) return std_logic_vector;

end CONV_PACK_top_level;

package body CONV_PACK_top_level is
   
   -- std_logic_vector to enum type function
   function std_logic_vector_to_aluOp(arg : in std_logic_vector( 1 to 5 )) 
   return aluOp is
   -- synopsys built_in SYN_FEED_THRU;
   begin
      case arg is
         when "00000" => return NOP;
         when "00001" => return SLLS;
         when "00010" => return SRLS;
         when "00011" => return SRAS;
         when "00100" => return ADDS;
         when "00101" => return ADDUS;
         when "00110" => return SUBS;
         when "00111" => return SUBUS;
         when "01000" => return ANDS;
         when "01001" => return ORS;
         when "01010" => return XORS;
         when "01011" => return SEQS;
         when "01100" => return SNES;
         when "01101" => return SLTS;
         when "01110" => return SGTS;
         when "01111" => return SLES;
         when "10000" => return SGES;
         when "10001" => return MOVI2SS;
         when "10010" => return MOVS2IS;
         when "10011" => return MOVFS;
         when "10100" => return MOVDS;
         when "10101" => return MOVFP2IS;
         when "10110" => return MOVI2FP;
         when "10111" => return MOVI2TS;
         when "11000" => return MOVT2IS;
         when "11001" => return SLTUS;
         when "11010" => return SGTUS;
         when "11011" => return SLEUS;
         when "11100" => return SGEUS;
         when "11101" => return MULTU;
         when "11110" => return MULTS;
         when others => assert FALSE -- this should not happen.
               report "un-convertible value"
               severity warning;
               return NOP;
      end case;
   end;
   
   -- enum type to std_logic_vector function
   function aluOp_to_std_logic_vector(arg : in aluOp) return std_logic_vector 
   is
   -- synopsys built_in SYN_FEED_THRU;
   begin
      case arg is
         when NOP => return "00000";
         when SLLS => return "00001";
         when SRLS => return "00010";
         when SRAS => return "00011";
         when ADDS => return "00100";
         when ADDUS => return "00101";
         when SUBS => return "00110";
         when SUBUS => return "00111";
         when ANDS => return "01000";
         when ORS => return "01001";
         when XORS => return "01010";
         when SEQS => return "01011";
         when SNES => return "01100";
         when SLTS => return "01101";
         when SGTS => return "01110";
         when SLES => return "01111";
         when SGES => return "10000";
         when MOVI2SS => return "10001";
         when MOVS2IS => return "10010";
         when MOVFS => return "10011";
         when MOVDS => return "10100";
         when MOVFP2IS => return "10101";
         when MOVI2FP => return "10110";
         when MOVI2TS => return "10111";
         when MOVT2IS => return "11000";
         when SLTUS => return "11001";
         when SGTUS => return "11010";
         when SLEUS => return "11011";
         when SGEUS => return "11100";
         when MULTU => return "11101";
         when MULTS => return "11110";
         when others => assert FALSE -- this should not happen.
               report "un-convertible value"
               severity warning;
               return "00000";
      end case;
   end;

end CONV_PACK_top_level;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_16 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_16;

architecture SYN_USE_DEFA_ARCH_NAME of 
   SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_16 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net3615 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net3615);
   main_gate : AND2_X1 port map( A1 => net3615, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_15 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_15;

architecture SYN_USE_DEFA_ARCH_NAME of 
   SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_15 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net3615 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net3615);
   main_gate : AND2_X1 port map( A1 => net3615, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_14 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_14;

architecture SYN_USE_DEFA_ARCH_NAME of 
   SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_14 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net3615 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net3615);
   main_gate : AND2_X1 port map( A1 => net3615, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_13 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_13;

architecture SYN_USE_DEFA_ARCH_NAME of 
   SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_13 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net3615 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net3615);
   main_gate : AND2_X1 port map( A1 => net3615, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_12 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_12;

architecture SYN_USE_DEFA_ARCH_NAME of 
   SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_12 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net3615 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net3615);
   main_gate : AND2_X1 port map( A1 => net3615, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_11 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_11;

architecture SYN_USE_DEFA_ARCH_NAME of 
   SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_11 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net3615 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net3615);
   main_gate : AND2_X1 port map( A1 => net3615, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_10 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_10;

architecture SYN_USE_DEFA_ARCH_NAME of 
   SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_10 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net3615 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net3615);
   main_gate : AND2_X1 port map( A1 => net3615, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_9 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_9;

architecture SYN_USE_DEFA_ARCH_NAME of 
   SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_9 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net3615 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net3615);
   main_gate : AND2_X1 port map( A1 => net3615, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_8 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_8;

architecture SYN_USE_DEFA_ARCH_NAME of 
   SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_8 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net3615 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net3615);
   main_gate : AND2_X1 port map( A1 => net3615, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_7 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_7;

architecture SYN_USE_DEFA_ARCH_NAME of 
   SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_7 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net3615 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net3615);
   main_gate : AND2_X1 port map( A1 => net3615, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_6 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_6;

architecture SYN_USE_DEFA_ARCH_NAME of 
   SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_6 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net3615 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net3615);
   main_gate : AND2_X1 port map( A1 => net3615, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_5 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_5;

architecture SYN_USE_DEFA_ARCH_NAME of 
   SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_5 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net3615 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net3615);
   main_gate : AND2_X1 port map( A1 => net3615, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_4 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_4;

architecture SYN_USE_DEFA_ARCH_NAME of 
   SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_4 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net3615 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net3615);
   main_gate : AND2_X1 port map( A1 => net3615, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_3 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_3;

architecture SYN_USE_DEFA_ARCH_NAME of 
   SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_3 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net3615 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net3615);
   main_gate : AND2_X1 port map( A1 => net3615, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_2 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_2;

architecture SYN_USE_DEFA_ARCH_NAME of 
   SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_2 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net3615 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net3615);
   main_gate : AND2_X1 port map( A1 => net3615, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_1 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_1;

architecture SYN_USE_DEFA_ARCH_NAME of 
   SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_1 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net3615 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net3615);
   main_gate : AND2_X1 port map( A1 => net3615, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_ff32_en_1 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_ff32_en_1;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_ff32_en_1 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net3600 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net3600);
   main_gate : AND2_X1 port map( A1 => net3600, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_dlx_regfile_33 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_dlx_regfile_33;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_dlx_regfile_33 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net3385 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net3385);
   main_gate : AND2_X1 port map( A1 => net3385, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_dlx_regfile_32 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_dlx_regfile_32;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_dlx_regfile_32 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net3385 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net3385);
   main_gate : AND2_X1 port map( A1 => net3385, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_dlx_regfile_31 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_dlx_regfile_31;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_dlx_regfile_31 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net3385 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net3385);
   main_gate : AND2_X1 port map( A1 => net3385, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_dlx_regfile_30 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_dlx_regfile_30;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_dlx_regfile_30 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net3385 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net3385);
   main_gate : AND2_X1 port map( A1 => net3385, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_dlx_regfile_29 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_dlx_regfile_29;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_dlx_regfile_29 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net3385 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net3385);
   main_gate : AND2_X1 port map( A1 => net3385, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_dlx_regfile_28 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_dlx_regfile_28;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_dlx_regfile_28 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net3385 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net3385);
   main_gate : AND2_X1 port map( A1 => net3385, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_dlx_regfile_27 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_dlx_regfile_27;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_dlx_regfile_27 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net3385 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net3385);
   main_gate : AND2_X1 port map( A1 => net3385, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_dlx_regfile_26 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_dlx_regfile_26;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_dlx_regfile_26 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net3385 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net3385);
   main_gate : AND2_X1 port map( A1 => net3385, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_dlx_regfile_25 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_dlx_regfile_25;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_dlx_regfile_25 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net3385 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net3385);
   main_gate : AND2_X1 port map( A1 => net3385, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_dlx_regfile_24 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_dlx_regfile_24;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_dlx_regfile_24 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net3385 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net3385);
   main_gate : AND2_X1 port map( A1 => net3385, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_dlx_regfile_23 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_dlx_regfile_23;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_dlx_regfile_23 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net3385 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net3385);
   main_gate : AND2_X1 port map( A1 => net3385, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_dlx_regfile_22 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_dlx_regfile_22;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_dlx_regfile_22 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net3385 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net3385);
   main_gate : AND2_X1 port map( A1 => net3385, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_dlx_regfile_21 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_dlx_regfile_21;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_dlx_regfile_21 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net3385 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net3385);
   main_gate : AND2_X1 port map( A1 => net3385, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_dlx_regfile_20 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_dlx_regfile_20;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_dlx_regfile_20 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net3385 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net3385);
   main_gate : AND2_X1 port map( A1 => net3385, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_dlx_regfile_19 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_dlx_regfile_19;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_dlx_regfile_19 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net3385 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net3385);
   main_gate : AND2_X1 port map( A1 => net3385, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_dlx_regfile_18 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_dlx_regfile_18;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_dlx_regfile_18 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net3385 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net3385);
   main_gate : AND2_X1 port map( A1 => net3385, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_dlx_regfile_17 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_dlx_regfile_17;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_dlx_regfile_17 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net3385 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net3385);
   main_gate : AND2_X1 port map( A1 => net3385, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_dlx_regfile_16 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_dlx_regfile_16;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_dlx_regfile_16 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net3385 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net3385);
   main_gate : AND2_X1 port map( A1 => net3385, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_dlx_regfile_15 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_dlx_regfile_15;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_dlx_regfile_15 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net3385 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net3385);
   main_gate : AND2_X1 port map( A1 => net3385, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_dlx_regfile_14 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_dlx_regfile_14;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_dlx_regfile_14 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net3385 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net3385);
   main_gate : AND2_X1 port map( A1 => net3385, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_dlx_regfile_13 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_dlx_regfile_13;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_dlx_regfile_13 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net3385 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net3385);
   main_gate : AND2_X1 port map( A1 => net3385, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_dlx_regfile_12 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_dlx_regfile_12;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_dlx_regfile_12 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net3385 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net3385);
   main_gate : AND2_X1 port map( A1 => net3385, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_dlx_regfile_11 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_dlx_regfile_11;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_dlx_regfile_11 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net3385 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net3385);
   main_gate : AND2_X1 port map( A1 => net3385, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_dlx_regfile_10 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_dlx_regfile_10;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_dlx_regfile_10 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net3385 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net3385);
   main_gate : AND2_X1 port map( A1 => net3385, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_dlx_regfile_9 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_dlx_regfile_9;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_dlx_regfile_9 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net3385 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net3385);
   main_gate : AND2_X1 port map( A1 => net3385, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_dlx_regfile_8 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_dlx_regfile_8;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_dlx_regfile_8 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net3385 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net3385);
   main_gate : AND2_X1 port map( A1 => net3385, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_dlx_regfile_7 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_dlx_regfile_7;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_dlx_regfile_7 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net3385 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net3385);
   main_gate : AND2_X1 port map( A1 => net3385, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_dlx_regfile_6 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_dlx_regfile_6;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_dlx_regfile_6 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net3385 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net3385);
   main_gate : AND2_X1 port map( A1 => net3385, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_dlx_regfile_5 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_dlx_regfile_5;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_dlx_regfile_5 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net3385 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net3385);
   main_gate : AND2_X1 port map( A1 => net3385, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_dlx_regfile_4 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_dlx_regfile_4;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_dlx_regfile_4 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net3385 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net3385);
   main_gate : AND2_X1 port map( A1 => net3385, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_dlx_regfile_3 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_dlx_regfile_3;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_dlx_regfile_3 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net3385 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net3385);
   main_gate : AND2_X1 port map( A1 => net3385, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_dlx_regfile_2 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_dlx_regfile_2;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_dlx_regfile_2 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net3385 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net3385);
   main_gate : AND2_X1 port map( A1 => net3385, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_dlx_regfile_1 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_dlx_regfile_1;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_dlx_regfile_1 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net3385 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net3385);
   main_gate : AND2_X1 port map( A1 => net3385, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_ff32_en_SIZE5_3 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_ff32_en_SIZE5_3;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_ff32_en_SIZE5_3 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net3355 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net3355);
   main_gate : AND2_X1 port map( A1 => net3355, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_ff32_en_SIZE5_2 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_ff32_en_SIZE5_2;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_ff32_en_SIZE5_2 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net3355 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net3355);
   main_gate : AND2_X1 port map( A1 => net3355, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_ff32_en_SIZE32_5 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_ff32_en_SIZE32_5;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_ff32_en_SIZE32_5 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net3340 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net3340);
   main_gate : AND2_X1 port map( A1 => net3340, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_ff32_en_SIZE32_4 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_ff32_en_SIZE32_4;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_ff32_en_SIZE32_4 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net3340 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net3340);
   main_gate : AND2_X1 port map( A1 => net3340, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_ff32_en_SIZE32_1 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_ff32_en_SIZE32_1;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_ff32_en_SIZE32_1 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net3340 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net3340);
   main_gate : AND2_X1 port map( A1 => net3340, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_127 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_127;

architecture SYN_BEHAVIORAL of FA_127 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U1 : XNOR2_X1 port map( A => n6, B => B, ZN => S);
   U5 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => B, A2 => Ci, ZN => n4);
   U3 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_126 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_126;

architecture SYN_BEHAVIORAL of FA_126 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U5 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => B, A2 => Ci, ZN => n4);
   U3 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U1 : XNOR2_X1 port map( A => n6, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_125 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_125;

architecture SYN_BEHAVIORAL of FA_125 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n2);
   U1 : XNOR2_X1 port map( A => n2, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_120 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_120;

architecture SYN_BEHAVIORAL of FA_120 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => S);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_119 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_119;

architecture SYN_BEHAVIORAL of FA_119 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U5 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => B, A2 => Ci, ZN => n4);
   U3 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U1 : XNOR2_X1 port map( A => n6, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_118 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_118;

architecture SYN_BEHAVIORAL of FA_118 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U5 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => B, A2 => Ci, ZN => n4);
   U3 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U1 : XNOR2_X1 port map( A => n6, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_117 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_117;

architecture SYN_BEHAVIORAL of FA_117 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n2);
   U1 : XNOR2_X1 port map( A => n2, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_116 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_116;

architecture SYN_BEHAVIORAL of FA_116 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => A, A2 => B, ZN => Co);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_115 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_115;

architecture SYN_BEHAVIORAL of FA_115 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U5 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => B, A2 => Ci, ZN => n4);
   U3 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U1 : XNOR2_X1 port map( A => n6, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_114 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_114;

architecture SYN_BEHAVIORAL of FA_114 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U5 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => B, A2 => Ci, ZN => n4);
   U3 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U1 : XNOR2_X1 port map( A => n6, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_113 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_113;

architecture SYN_BEHAVIORAL of FA_113 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n2);
   U1 : XNOR2_X1 port map( A => n2, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_112 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_112;

architecture SYN_BEHAVIORAL of FA_112 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => S);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_111 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_111;

architecture SYN_BEHAVIORAL of FA_111 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U5 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => B, A2 => Ci, ZN => n4);
   U3 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U1 : XNOR2_X1 port map( A => n6, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_110 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_110;

architecture SYN_BEHAVIORAL of FA_110 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U5 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => B, A2 => Ci, ZN => n4);
   U3 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U1 : XNOR2_X1 port map( A => n6, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_109 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_109;

architecture SYN_BEHAVIORAL of FA_109 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n2);
   U1 : XNOR2_X1 port map( A => n2, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_108 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_108;

architecture SYN_BEHAVIORAL of FA_108 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => A, A2 => B, ZN => Co);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_107 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_107;

architecture SYN_BEHAVIORAL of FA_107 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U5 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => B, A2 => Ci, ZN => n4);
   U3 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U1 : XNOR2_X1 port map( A => n6, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_106 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_106;

architecture SYN_BEHAVIORAL of FA_106 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U5 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => B, A2 => Ci, ZN => n4);
   U3 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U1 : XNOR2_X1 port map( A => n6, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_105 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_105;

architecture SYN_BEHAVIORAL of FA_105 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n2);
   U1 : XNOR2_X1 port map( A => n2, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_104 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_104;

architecture SYN_BEHAVIORAL of FA_104 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => S);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_103 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_103;

architecture SYN_BEHAVIORAL of FA_103 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U5 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => B, A2 => Ci, ZN => n4);
   U3 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U1 : XNOR2_X1 port map( A => n6, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_102 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_102;

architecture SYN_BEHAVIORAL of FA_102 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U5 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => B, A2 => Ci, ZN => n4);
   U3 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U1 : XNOR2_X1 port map( A => n6, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_101 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_101;

architecture SYN_BEHAVIORAL of FA_101 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n2);
   U1 : XNOR2_X1 port map( A => n2, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_100 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_100;

architecture SYN_BEHAVIORAL of FA_100 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => A, A2 => B, ZN => Co);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_99 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_99;

architecture SYN_BEHAVIORAL of FA_99 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U5 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => B, A2 => Ci, ZN => n4);
   U3 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U1 : XNOR2_X1 port map( A => n6, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_98 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_98;

architecture SYN_BEHAVIORAL of FA_98 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U5 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => B, A2 => Ci, ZN => n4);
   U3 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U1 : XNOR2_X1 port map( A => n6, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_97 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_97;

architecture SYN_BEHAVIORAL of FA_97 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n2);
   U1 : XNOR2_X1 port map( A => n2, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_96 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_96;

architecture SYN_BEHAVIORAL of FA_96 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => S);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_95 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_95;

architecture SYN_BEHAVIORAL of FA_95 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U1 : XNOR2_X1 port map( A => n6, B => B, ZN => S);
   U4 : NAND2_X1 port map( A1 => B, A2 => Ci, ZN => n4);
   U5 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_94 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_94;

architecture SYN_BEHAVIORAL of FA_94 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U1 : XNOR2_X1 port map( A => n6, B => B, ZN => S);
   U4 : NAND2_X1 port map( A1 => B, A2 => Ci, ZN => n4);
   U5 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_93 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_93;

architecture SYN_BEHAVIORAL of FA_93 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n1);
   U2 : XOR2_X1 port map( A => Ci, B => n1, Z => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_92 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_92;

architecture SYN_BEHAVIORAL of FA_92 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => A, A2 => B, ZN => Co);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_91 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_91;

architecture SYN_BEHAVIORAL of FA_91 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U1 : XNOR2_X1 port map( A => n6, B => B, ZN => S);
   U4 : NAND2_X1 port map( A1 => B, A2 => Ci, ZN => n4);
   U5 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_90 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_90;

architecture SYN_BEHAVIORAL of FA_90 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U1 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U3 : XNOR2_X1 port map( A => n6, B => B, ZN => S);
   U4 : NAND2_X1 port map( A1 => B, A2 => Ci, ZN => n4);
   U5 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_89 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_89;

architecture SYN_BEHAVIORAL of FA_89 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n1);
   U2 : XOR2_X1 port map( A => Ci, B => n1, Z => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_88 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_88;

architecture SYN_BEHAVIORAL of FA_88 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => S);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_87 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_87;

architecture SYN_BEHAVIORAL of FA_87 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U1 : NAND2_X1 port map( A1 => B, A2 => Ci, ZN => n5);
   U3 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n4);
   U4 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U5 : XNOR2_X1 port map( A => n6, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_86 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_86;

architecture SYN_BEHAVIORAL of FA_86 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => Ci, ZN => n5);
   U2 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n4);
   U3 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U4 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U5 : XNOR2_X1 port map( A => n6, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_85 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_85;

architecture SYN_BEHAVIORAL of FA_85 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => Ci, ZN => n2);
   U2 : XNOR2_X1 port map( A => n2, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_84 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_84;

architecture SYN_BEHAVIORAL of FA_84 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => A, A2 => B, ZN => Co);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_83 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_83;

architecture SYN_BEHAVIORAL of FA_83 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U1 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U3 : XNOR2_X1 port map( A => n6, B => B, ZN => S);
   U4 : NAND2_X1 port map( A1 => B, A2 => Ci, ZN => n4);
   U5 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_82 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_82;

architecture SYN_BEHAVIORAL of FA_82 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U1 : XNOR2_X1 port map( A => n6, B => B, ZN => S);
   U3 : NAND2_X1 port map( A1 => B, A2 => Ci, ZN => n4);
   U4 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U5 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_81 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_81;

architecture SYN_BEHAVIORAL of FA_81 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n2, B => B, ZN => S);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_80 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_80;

architecture SYN_BEHAVIORAL of FA_80 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n3);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => Co);
   U3 : XNOR2_X1 port map( A => n3, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_79 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_79;

architecture SYN_BEHAVIORAL of FA_79 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U1 : XNOR2_X1 port map( A => n6, B => B, ZN => S);
   U4 : NAND2_X1 port map( A1 => B, A2 => Ci, ZN => n4);
   U5 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_78 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_78;

architecture SYN_BEHAVIORAL of FA_78 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U1 : XNOR2_X1 port map( A => n6, B => B, ZN => S);
   U3 : NAND2_X1 port map( A1 => B, A2 => Ci, ZN => n4);
   U4 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n5);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_77 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_77;

architecture SYN_BEHAVIORAL of FA_77 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n2, B => B, ZN => S);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_76 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_76;

architecture SYN_BEHAVIORAL of FA_76 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => A, A2 => B, ZN => Co);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_75 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_75;

architecture SYN_BEHAVIORAL of FA_75 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U1 : XNOR2_X1 port map( A => n6, B => B, ZN => S);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U4 : NAND2_X1 port map( A1 => B, A2 => Ci, ZN => n4);
   U5 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_74 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_74;

architecture SYN_BEHAVIORAL of FA_74 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U1 : XNOR2_X1 port map( A => n6, B => B, ZN => S);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U4 : NAND2_X1 port map( A1 => B, A2 => Ci, ZN => n4);
   U5 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_73 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_73;

architecture SYN_BEHAVIORAL of FA_73 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n2);
   U1 : XNOR2_X1 port map( A => n2, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_72 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_72;

architecture SYN_BEHAVIORAL of FA_72 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => S);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_71 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_71;

architecture SYN_BEHAVIORAL of FA_71 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U3 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U1 : XNOR2_X1 port map( A => n6, B => B, ZN => S);
   U4 : NAND2_X1 port map( A1 => B, A2 => Ci, ZN => n4);
   U5 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_70 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_70;

architecture SYN_BEHAVIORAL of FA_70 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n4 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n4);
   U1 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n2);
   U3 : NAND2_X1 port map( A1 => n2, A2 => n3, ZN => Co);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => B, ZN => n3);
   U5 : XNOR2_X1 port map( A => n4, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_69 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_69;

architecture SYN_BEHAVIORAL of FA_69 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal net48795 : std_logic;

begin
   
   U1 : FA_X1 port map( A => B, B => A, CI => Ci, CO => net48795, S => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_68 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_68;

architecture SYN_BEHAVIORAL of FA_68 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => A, A2 => B, ZN => Co);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_67 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_67;

architecture SYN_BEHAVIORAL of FA_67 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n4 : std_logic;

begin
   
   U1 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n2);
   U2 : NAND2_X1 port map( A1 => n2, A2 => n3, ZN => Co);
   U3 : NAND2_X1 port map( A1 => Ci, A2 => B, ZN => n3);
   U4 : XNOR2_X1 port map( A => n4, B => B, ZN => S);
   U5 : XNOR2_X1 port map( A => A, B => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_66 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_66;

architecture SYN_BEHAVIORAL of FA_66 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n4 : std_logic;

begin
   
   U1 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n2);
   U2 : NAND2_X1 port map( A1 => n2, A2 => n3, ZN => Co);
   U3 : NAND2_X1 port map( A1 => Ci, A2 => B, ZN => n3);
   U4 : XNOR2_X1 port map( A => n4, B => B, ZN => S);
   U5 : XNOR2_X1 port map( A => Ci, B => A, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_65 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_65;

architecture SYN_BEHAVIORAL of FA_65 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => Ci, ZN => n2);
   U2 : XNOR2_X1 port map( A => n2, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_64 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_64;

architecture SYN_BEHAVIORAL of FA_64 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => S);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_63 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_63;

architecture SYN_BEHAVIORAL of FA_63 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U3 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U1 : XNOR2_X1 port map( A => n6, B => B, ZN => S);
   U4 : NAND2_X1 port map( A1 => B, A2 => Ci, ZN => n4);
   U5 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_62 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_62;

architecture SYN_BEHAVIORAL of FA_62 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U1 : XNOR2_X1 port map( A => n6, B => B, ZN => S);
   U4 : NAND2_X1 port map( A1 => B, A2 => Ci, ZN => n4);
   U5 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_61 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_61;

architecture SYN_BEHAVIORAL of FA_61 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n2);
   U1 : XNOR2_X1 port map( A => n2, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_60 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_60;

architecture SYN_BEHAVIORAL of FA_60 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => A, A2 => B, ZN => Co);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_59 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_59;

architecture SYN_BEHAVIORAL of FA_59 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U3 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U1 : XNOR2_X1 port map( A => n6, B => B, ZN => S);
   U4 : NAND2_X1 port map( A1 => B, A2 => Ci, ZN => n4);
   U5 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_58 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_58;

architecture SYN_BEHAVIORAL of FA_58 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U1 : XNOR2_X1 port map( A => n6, B => B, ZN => S);
   U4 : NAND2_X1 port map( A1 => B, A2 => Ci, ZN => n4);
   U5 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_57 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_57;

architecture SYN_BEHAVIORAL of FA_57 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n2);
   U1 : XNOR2_X1 port map( A => n2, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_56 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_56;

architecture SYN_BEHAVIORAL of FA_56 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => S);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_55 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_55;

architecture SYN_BEHAVIORAL of FA_55 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U1 : NAND2_X1 port map( A1 => B, A2 => Ci, ZN => n4);
   U4 : XNOR2_X1 port map( A => n6, B => B, ZN => S);
   U5 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_54 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_54;

architecture SYN_BEHAVIORAL of FA_54 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U3 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U1 : XNOR2_X1 port map( A => n6, B => B, ZN => S);
   U4 : NAND2_X1 port map( A1 => B, A2 => Ci, ZN => n4);
   U5 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_53 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_53;

architecture SYN_BEHAVIORAL of FA_53 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n2);
   U1 : XNOR2_X1 port map( A => n2, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_52 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_52;

architecture SYN_BEHAVIORAL of FA_52 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => S);
   U2 : OR2_X1 port map( A1 => A, A2 => B, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_51 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_51;

architecture SYN_BEHAVIORAL of FA_51 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U1 : NAND2_X1 port map( A1 => B, A2 => Ci, ZN => n4);
   U4 : XNOR2_X1 port map( A => n6, B => B, ZN => S);
   U5 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_50 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_50;

architecture SYN_BEHAVIORAL of FA_50 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U3 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U1 : XNOR2_X1 port map( A => n6, B => B, ZN => S);
   U4 : NAND2_X1 port map( A1 => B, A2 => Ci, ZN => n4);
   U5 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_49 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_49;

architecture SYN_BEHAVIORAL of FA_49 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n2);
   U1 : XNOR2_X1 port map( A => n2, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_48 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_48;

architecture SYN_BEHAVIORAL of FA_48 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => S);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_47 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_47;

architecture SYN_BEHAVIORAL of FA_47 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U1 : XNOR2_X1 port map( A => n6, B => B, ZN => S);
   U4 : NAND2_X1 port map( A1 => B, A2 => Ci, ZN => n4);
   U5 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_46 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_46;

architecture SYN_BEHAVIORAL of FA_46 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U1 : XNOR2_X1 port map( A => n6, B => B, ZN => S);
   U4 : NAND2_X1 port map( A1 => B, A2 => Ci, ZN => n4);
   U5 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_45 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_45;

architecture SYN_BEHAVIORAL of FA_45 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal net48794 : std_logic;

begin
   
   U1 : FA_X1 port map( A => B, B => A, CI => Ci, CO => net48794, S => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_44 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_44;

architecture SYN_BEHAVIORAL of FA_44 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => S);
   U2 : OR2_X1 port map( A1 => A, A2 => B, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_43 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_43;

architecture SYN_BEHAVIORAL of FA_43 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U1 : XNOR2_X1 port map( A => n6, B => B, ZN => S);
   U4 : NAND2_X1 port map( A1 => B, A2 => Ci, ZN => n4);
   U5 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_42 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_42;

architecture SYN_BEHAVIORAL of FA_42 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U1 : XNOR2_X1 port map( A => n6, B => B, ZN => S);
   U4 : NAND2_X1 port map( A1 => B, A2 => Ci, ZN => n4);
   U5 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_41 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_41;

architecture SYN_BEHAVIORAL of FA_41 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U2 : XOR2_X1 port map( A => B, B => n2, Z => n1);
   U3 : XNOR2_X1 port map( A => Ci, B => n1, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_40 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_40;

architecture SYN_BEHAVIORAL of FA_40 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Co);
   U2 : INV_X1 port map( A => A, ZN => n3);
   U3 : XNOR2_X1 port map( A => n3, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_39 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_39;

architecture SYN_BEHAVIORAL of FA_39 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U1 : XNOR2_X1 port map( A => n6, B => B, ZN => S);
   U4 : NAND2_X1 port map( A1 => B, A2 => Ci, ZN => n4);
   U5 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_38 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_38;

architecture SYN_BEHAVIORAL of FA_38 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U3 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U1 : XNOR2_X1 port map( A => n6, B => B, ZN => S);
   U4 : NAND2_X1 port map( A1 => B, A2 => Ci, ZN => n4);
   U5 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_37 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_37;

architecture SYN_BEHAVIORAL of FA_37 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n2);
   U1 : XNOR2_X1 port map( A => n2, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_36 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_36;

architecture SYN_BEHAVIORAL of FA_36 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => A, A2 => B, ZN => Co);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_35 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_35;

architecture SYN_BEHAVIORAL of FA_35 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U1 : XNOR2_X1 port map( A => n6, B => B, ZN => S);
   U4 : NAND2_X1 port map( A1 => B, A2 => Ci, ZN => n4);
   U5 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_34 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_34;

architecture SYN_BEHAVIORAL of FA_34 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U3 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U1 : XNOR2_X1 port map( A => n6, B => B, ZN => S);
   U4 : NAND2_X1 port map( A1 => B, A2 => Ci, ZN => n4);
   U5 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_33 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_33;

architecture SYN_BEHAVIORAL of FA_33 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n2);
   U1 : XNOR2_X1 port map( A => n2, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_32 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_32;

architecture SYN_BEHAVIORAL of FA_32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n3, B => B, ZN => S);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => Co);
   U3 : INV_X1 port map( A => A, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_31 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_31;

architecture SYN_BEHAVIORAL of FA_31 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U1 : XNOR2_X1 port map( A => n6, B => B, ZN => S);
   U4 : NAND2_X1 port map( A1 => B, A2 => Ci, ZN => n4);
   U5 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_30 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_30;

architecture SYN_BEHAVIORAL of FA_30 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U3 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U1 : XNOR2_X1 port map( A => n6, B => B, ZN => S);
   U4 : NAND2_X1 port map( A1 => B, A2 => Ci, ZN => n4);
   U5 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_29 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_29;

architecture SYN_BEHAVIORAL of FA_29 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n1);
   U2 : XNOR2_X1 port map( A => Ci, B => n1, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_28 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_28;

architecture SYN_BEHAVIORAL of FA_28 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => S);
   U2 : OR2_X1 port map( A1 => A, A2 => B, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_27 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_27;

architecture SYN_BEHAVIORAL of FA_27 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U1 : XNOR2_X1 port map( A => n6, B => B, ZN => S);
   U4 : NAND2_X1 port map( A1 => B, A2 => Ci, ZN => n4);
   U5 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_26 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_26;

architecture SYN_BEHAVIORAL of FA_26 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U3 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U1 : XNOR2_X1 port map( A => n6, B => B, ZN => S);
   U4 : NAND2_X1 port map( A1 => B, A2 => Ci, ZN => n4);
   U5 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_25 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_25;

architecture SYN_BEHAVIORAL of FA_25 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n1);
   U2 : XNOR2_X1 port map( A => Ci, B => n1, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_24 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_24;

architecture SYN_BEHAVIORAL of FA_24 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n3);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => Co);
   U3 : XNOR2_X1 port map( A => n3, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_23 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_23;

architecture SYN_BEHAVIORAL of FA_23 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U1 : XNOR2_X1 port map( A => n6, B => B, ZN => S);
   U4 : NAND2_X1 port map( A1 => B, A2 => Ci, ZN => n4);
   U5 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_22 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_22;

architecture SYN_BEHAVIORAL of FA_22 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U1 : XNOR2_X1 port map( A => n6, B => B, ZN => S);
   U4 : NAND2_X1 port map( A1 => B, A2 => Ci, ZN => n4);
   U5 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_21 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_21;

architecture SYN_BEHAVIORAL of FA_21 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n2);
   U1 : XNOR2_X1 port map( A => n2, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_20 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_20;

architecture SYN_BEHAVIORAL of FA_20 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => A, A2 => B, ZN => Co);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_19 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_19;

architecture SYN_BEHAVIORAL of FA_19 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U1 : XNOR2_X1 port map( A => n6, B => B, ZN => S);
   U4 : NAND2_X1 port map( A1 => B, A2 => Ci, ZN => n4);
   U5 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_18 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_18;

architecture SYN_BEHAVIORAL of FA_18 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U1 : XNOR2_X1 port map( A => n6, B => B, ZN => S);
   U4 : NAND2_X1 port map( A1 => B, A2 => Ci, ZN => n4);
   U5 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_17 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_17;

architecture SYN_BEHAVIORAL of FA_17 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n2);
   U1 : XNOR2_X1 port map( A => n2, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_16 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_16;

architecture SYN_BEHAVIORAL of FA_16 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => S);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_15 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_15;

architecture SYN_BEHAVIORAL of FA_15 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U3 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U1 : XNOR2_X1 port map( A => n6, B => B, ZN => S);
   U4 : NAND2_X1 port map( A1 => B, A2 => Ci, ZN => n4);
   U5 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_14 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_14;

architecture SYN_BEHAVIORAL of FA_14 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U1 : XNOR2_X1 port map( A => n6, B => B, ZN => S);
   U4 : NAND2_X1 port map( A1 => B, A2 => Ci, ZN => n4);
   U5 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_13 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_13;

architecture SYN_BEHAVIORAL of FA_13 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n2);
   U1 : XNOR2_X1 port map( A => n2, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_12 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_12;

architecture SYN_BEHAVIORAL of FA_12 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => A, A2 => B, ZN => Co);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_11 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_11;

architecture SYN_BEHAVIORAL of FA_11 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U3 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U1 : XNOR2_X1 port map( A => n6, B => B, ZN => S);
   U4 : NAND2_X1 port map( A1 => B, A2 => Ci, ZN => n4);
   U5 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_10 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_10;

architecture SYN_BEHAVIORAL of FA_10 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U1 : XNOR2_X1 port map( A => n6, B => B, ZN => S);
   U4 : NAND2_X1 port map( A1 => B, A2 => Ci, ZN => n4);
   U5 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_9 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_9;

architecture SYN_BEHAVIORAL of FA_9 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n2);
   U1 : XNOR2_X1 port map( A => n2, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_8 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_8;

architecture SYN_BEHAVIORAL of FA_8 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n3, B => B, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n3);
   U3 : AND2_X1 port map( A1 => B, A2 => A, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_7 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_7;

architecture SYN_BEHAVIORAL of FA_7 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U1 : XNOR2_X1 port map( A => n6, B => B, ZN => S);
   U3 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => B, A2 => Ci, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_6 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_6;

architecture SYN_BEHAVIORAL of FA_6 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U5 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n5);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U1 : XNOR2_X1 port map( A => n6, B => B, ZN => S);
   U3 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U4 : NAND2_X1 port map( A1 => B, A2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_5 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_5;

architecture SYN_BEHAVIORAL of FA_5 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => Ci, ZN => n2);
   U2 : XNOR2_X1 port map( A => n2, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_4 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_4;

architecture SYN_BEHAVIORAL of FA_4 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => S);
   U2 : OR2_X1 port map( A1 => A, A2 => B, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_3 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_3;

architecture SYN_BEHAVIORAL of FA_3 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U1 : XNOR2_X1 port map( A => n6, B => B, ZN => S);
   U4 : NAND2_X1 port map( A1 => B, A2 => Ci, ZN => n4);
   U5 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_2 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_2;

architecture SYN_BEHAVIORAL of FA_2 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U5 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => B, A2 => Ci, ZN => n4);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U1 : XNOR2_X1 port map( A => n6, B => B, ZN => S);
   U3 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_1 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1;

architecture SYN_BEHAVIORAL of FA_1 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n2);
   U1 : XNOR2_X1 port map( A => n2, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity mux21_SIZE4_15 is

   port( IN0, IN1 : in std_logic_vector (3 downto 0);  CTRL : in std_logic;  
         OUT1 : out std_logic_vector (3 downto 0));

end mux21_SIZE4_15;

architecture SYN_Bhe of mux21_SIZE4_15 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => IN0(3), B => IN1(3), S => CTRL, Z => OUT1(3));
   U2 : MUX2_X1 port map( A => IN0(2), B => IN1(2), S => CTRL, Z => OUT1(2));
   U3 : MUX2_X1 port map( A => IN0(1), B => IN1(1), S => CTRL, Z => OUT1(1));
   U4 : MUX2_X1 port map( A => IN0(0), B => IN1(0), S => CTRL, Z => OUT1(0));

end SYN_Bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity mux21_SIZE4_14 is

   port( IN0, IN1 : in std_logic_vector (3 downto 0);  CTRL : in std_logic;  
         OUT1 : out std_logic_vector (3 downto 0));

end mux21_SIZE4_14;

architecture SYN_Bhe of mux21_SIZE4_14 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => IN0(3), B => IN1(3), S => CTRL, Z => OUT1(3));
   U2 : MUX2_X1 port map( A => IN0(2), B => IN1(2), S => CTRL, Z => OUT1(2));
   U3 : MUX2_X1 port map( A => IN0(1), B => IN1(1), S => CTRL, Z => OUT1(1));
   U4 : MUX2_X1 port map( A => IN0(0), B => IN1(0), S => CTRL, Z => OUT1(0));

end SYN_Bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity mux21_SIZE4_13 is

   port( IN0, IN1 : in std_logic_vector (3 downto 0);  CTRL : in std_logic;  
         OUT1 : out std_logic_vector (3 downto 0));

end mux21_SIZE4_13;

architecture SYN_Bhe of mux21_SIZE4_13 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => IN0(3), B => IN1(3), S => CTRL, Z => OUT1(3));
   U2 : MUX2_X1 port map( A => IN0(2), B => IN1(2), S => CTRL, Z => OUT1(2));
   U3 : MUX2_X1 port map( A => IN0(1), B => IN1(1), S => CTRL, Z => OUT1(1));
   U4 : MUX2_X1 port map( A => IN0(0), B => IN1(0), S => CTRL, Z => OUT1(0));

end SYN_Bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity mux21_SIZE4_12 is

   port( IN0, IN1 : in std_logic_vector (3 downto 0);  CTRL : in std_logic;  
         OUT1 : out std_logic_vector (3 downto 0));

end mux21_SIZE4_12;

architecture SYN_Bhe of mux21_SIZE4_12 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : MUX2_X1 port map( A => IN0(2), B => IN1(2), S => CTRL, Z => OUT1(2));
   U3 : MUX2_X1 port map( A => IN0(1), B => IN1(1), S => CTRL, Z => OUT1(1));
   U1 : MUX2_X1 port map( A => IN0(3), B => IN1(3), S => CTRL, Z => OUT1(3));
   U4 : MUX2_X1 port map( A => IN0(0), B => IN1(0), S => CTRL, Z => OUT1(0));

end SYN_Bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity mux21_SIZE4_11 is

   port( IN0, IN1 : in std_logic_vector (3 downto 0);  CTRL : in std_logic;  
         OUT1 : out std_logic_vector (3 downto 0));

end mux21_SIZE4_11;

architecture SYN_Bhe of mux21_SIZE4_11 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : MUX2_X1 port map( A => IN0(2), B => IN1(2), S => CTRL, Z => OUT1(2));
   U3 : MUX2_X1 port map( A => IN0(1), B => IN1(1), S => CTRL, Z => OUT1(1));
   U1 : MUX2_X1 port map( A => IN0(0), B => IN1(0), S => CTRL, Z => OUT1(0));
   U4 : MUX2_X1 port map( A => IN0(3), B => IN1(3), S => CTRL, Z => OUT1(3));

end SYN_Bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity mux21_SIZE4_10 is

   port( IN0, IN1 : in std_logic_vector (3 downto 0);  CTRL : in std_logic;  
         OUT1 : out std_logic_vector (3 downto 0));

end mux21_SIZE4_10;

architecture SYN_Bhe of mux21_SIZE4_10 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : MUX2_X1 port map( A => IN0(2), B => IN1(2), S => CTRL, Z => OUT1(2));
   U3 : MUX2_X1 port map( A => IN0(1), B => IN1(1), S => CTRL, Z => OUT1(1));
   U4 : MUX2_X1 port map( A => IN0(0), B => IN1(0), S => CTRL, Z => OUT1(0));
   U1 : MUX2_X1 port map( A => IN0(3), B => IN1(3), S => CTRL, Z => OUT1(3));

end SYN_Bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity mux21_SIZE4_9 is

   port( IN0, IN1 : in std_logic_vector (3 downto 0);  CTRL : in std_logic;  
         OUT1 : out std_logic_vector (3 downto 0));

end mux21_SIZE4_9;

architecture SYN_Bhe of mux21_SIZE4_9 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U3 : MUX2_X1 port map( A => IN0(1), B => IN1(1), S => CTRL, Z => OUT1(1));
   U1 : MUX2_X1 port map( A => IN0(3), B => IN1(3), S => CTRL, Z => OUT1(3));
   U2 : MUX2_X1 port map( A => IN0(0), B => IN1(0), S => CTRL, Z => OUT1(0));
   U4 : MUX2_X1 port map( A => IN0(2), B => IN1(2), S => CTRL, Z => OUT1(2));

end SYN_Bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity mux21_SIZE4_8 is

   port( IN0, IN1 : in std_logic_vector (3 downto 0);  CTRL : in std_logic;  
         OUT1 : out std_logic_vector (3 downto 0));

end mux21_SIZE4_8;

architecture SYN_Bhe of mux21_SIZE4_8 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => IN0(3), B => IN1(3), S => CTRL, Z => OUT1(3));
   U2 : MUX2_X1 port map( A => IN0(2), B => IN1(2), S => CTRL, Z => OUT1(2));
   U3 : MUX2_X1 port map( A => IN0(1), B => IN1(1), S => CTRL, Z => OUT1(1));
   U4 : MUX2_X1 port map( A => IN0(0), B => IN1(0), S => CTRL, Z => OUT1(0));

end SYN_Bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity mux21_SIZE4_7 is

   port( IN0, IN1 : in std_logic_vector (3 downto 0);  CTRL : in std_logic;  
         OUT1 : out std_logic_vector (3 downto 0));

end mux21_SIZE4_7;

architecture SYN_Bhe of mux21_SIZE4_7 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => IN0(3), B => IN1(3), S => CTRL, Z => OUT1(3));
   U3 : MUX2_X1 port map( A => IN0(1), B => IN1(1), S => CTRL, Z => OUT1(1));
   U2 : MUX2_X1 port map( A => IN0(0), B => IN1(0), S => CTRL, Z => OUT1(0));
   U4 : MUX2_X1 port map( A => IN0(2), B => IN1(2), S => CTRL, Z => OUT1(2));

end SYN_Bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity mux21_SIZE4_6 is

   port( IN0, IN1 : in std_logic_vector (3 downto 0);  CTRL : in std_logic;  
         OUT1 : out std_logic_vector (3 downto 0));

end mux21_SIZE4_6;

architecture SYN_Bhe of mux21_SIZE4_6 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : MUX2_X1 port map( A => IN0(2), B => IN1(2), S => CTRL, Z => OUT1(2));
   U3 : MUX2_X1 port map( A => IN0(1), B => IN1(1), S => CTRL, Z => OUT1(1));
   U1 : MUX2_X1 port map( A => IN0(0), B => IN1(0), S => CTRL, Z => OUT1(0));
   U4 : MUX2_X1 port map( A => IN0(3), B => IN1(3), S => CTRL, Z => OUT1(3));

end SYN_Bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity mux21_SIZE4_5 is

   port( IN0, IN1 : in std_logic_vector (3 downto 0);  CTRL : in std_logic;  
         OUT1 : out std_logic_vector (3 downto 0));

end mux21_SIZE4_5;

architecture SYN_Bhe of mux21_SIZE4_5 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => IN0(3), B => IN1(3), S => CTRL, Z => OUT1(3));
   U2 : MUX2_X1 port map( A => IN0(2), B => IN1(2), S => CTRL, Z => OUT1(2));
   U3 : MUX2_X1 port map( A => IN0(1), B => IN1(1), S => CTRL, Z => OUT1(1));
   U4 : MUX2_X1 port map( A => IN0(0), B => IN1(0), S => CTRL, Z => OUT1(0));

end SYN_Bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity mux21_SIZE4_4 is

   port( IN0, IN1 : in std_logic_vector (3 downto 0);  CTRL : in std_logic;  
         OUT1 : out std_logic_vector (3 downto 0));

end mux21_SIZE4_4;

architecture SYN_Bhe of mux21_SIZE4_4 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : MUX2_X1 port map( A => IN0(2), B => IN1(2), S => CTRL, Z => OUT1(2));
   U4 : MUX2_X1 port map( A => IN0(0), B => IN1(0), S => CTRL, Z => OUT1(0));
   U1 : MUX2_X1 port map( A => IN0(3), B => IN1(3), S => CTRL, Z => OUT1(3));
   U3 : MUX2_X1 port map( A => IN0(1), B => IN1(1), S => CTRL, Z => OUT1(1));

end SYN_Bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity mux21_SIZE4_3 is

   port( IN0, IN1 : in std_logic_vector (3 downto 0);  CTRL : in std_logic;  
         OUT1 : out std_logic_vector (3 downto 0));

end mux21_SIZE4_3;

architecture SYN_Bhe of mux21_SIZE4_3 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => IN0(0), B => IN1(0), S => CTRL, Z => OUT1(0));
   U2 : MUX2_X1 port map( A => IN0(3), B => IN1(3), S => CTRL, Z => OUT1(3));
   U3 : MUX2_X1 port map( A => IN0(1), B => IN1(1), S => CTRL, Z => OUT1(1));
   U4 : MUX2_X1 port map( A => IN0(2), B => IN1(2), S => CTRL, Z => OUT1(2));

end SYN_Bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity mux21_SIZE4_2 is

   port( IN0, IN1 : in std_logic_vector (3 downto 0);  CTRL : in std_logic;  
         OUT1 : out std_logic_vector (3 downto 0));

end mux21_SIZE4_2;

architecture SYN_Bhe of mux21_SIZE4_2 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => IN0(3), B => IN1(3), S => CTRL, Z => OUT1(3));
   U2 : MUX2_X1 port map( A => IN0(2), B => IN1(2), S => CTRL, Z => OUT1(2));
   U3 : MUX2_X1 port map( A => IN0(1), B => IN1(1), S => CTRL, Z => OUT1(1));
   U4 : MUX2_X1 port map( A => IN0(0), B => IN1(0), S => CTRL, Z => OUT1(0));

end SYN_Bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity mux21_SIZE4_1 is

   port( IN0, IN1 : in std_logic_vector (3 downto 0);  CTRL : in std_logic;  
         OUT1 : out std_logic_vector (3 downto 0));

end mux21_SIZE4_1;

architecture SYN_Bhe of mux21_SIZE4_1 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : MUX2_X1 port map( A => IN0(2), B => IN1(2), S => CTRL, Z => OUT1(2));
   U4 : MUX2_X1 port map( A => IN0(0), B => IN1(0), S => CTRL, Z => OUT1(0));
   U1 : MUX2_X1 port map( A => IN0(1), B => IN1(1), S => CTRL, Z => OUT1(1));
   U3 : MUX2_X1 port map( A => IN0(3), B => IN1(3), S => CTRL, Z => OUT1(3));

end SYN_Bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity RCA_N4_30 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_30;

architecture SYN_STRUCTURAL of RCA_N4_30 is

   component FA_117
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_118
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_119
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_120
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal n1, CTMP_3_port, CTMP_2_port, CTMP_1_port, net48793 : std_logic;

begin
   
   FAI_1 : FA_120 port map( A => A(0), B => B(0), Ci => n1, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_119 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_118 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_117 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => net48793);
   n1 <= '0';

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity RCA_N4_29 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_29;

architecture SYN_STRUCTURAL of RCA_N4_29 is

   component FA_113
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_114
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_115
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_116
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal n1, CTMP_3_port, CTMP_2_port, CTMP_1_port, net48792 : std_logic;

begin
   
   FAI_1 : FA_116 port map( A => A(0), B => B(0), Ci => n1, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_115 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_114 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_113 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => net48792);
   n1 <= '1';

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity RCA_N4_28 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_28;

architecture SYN_STRUCTURAL of RCA_N4_28 is

   component FA_109
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_110
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_111
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_112
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal n1, CTMP_3_port, CTMP_2_port, CTMP_1_port, net48791 : std_logic;

begin
   
   FAI_1 : FA_112 port map( A => A(0), B => B(0), Ci => n1, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_111 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_110 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_109 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => net48791);
   n1 <= '0';

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity RCA_N4_27 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_27;

architecture SYN_STRUCTURAL of RCA_N4_27 is

   component FA_105
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_106
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_107
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_108
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal n1, CTMP_3_port, CTMP_2_port, CTMP_1_port, net48790 : std_logic;

begin
   
   FAI_1 : FA_108 port map( A => A(0), B => B(0), Ci => n1, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_107 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_106 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_105 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => net48790);
   n1 <= '1';

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity RCA_N4_26 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_26;

architecture SYN_STRUCTURAL of RCA_N4_26 is

   component FA_101
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_102
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_103
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_104
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal n1, CTMP_3_port, CTMP_2_port, CTMP_1_port, net48789 : std_logic;

begin
   
   FAI_1 : FA_104 port map( A => A(0), B => B(0), Ci => n1, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_103 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_102 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_101 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => net48789);
   n1 <= '0';

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity RCA_N4_25 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_25;

architecture SYN_STRUCTURAL of RCA_N4_25 is

   component FA_97
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_98
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_99
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_100
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal n1, CTMP_3_port, CTMP_2_port, CTMP_1_port, net48788 : std_logic;

begin
   
   FAI_1 : FA_100 port map( A => A(0), B => B(0), Ci => n1, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_99 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_98 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_97 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => net48788);
   n1 <= '1';

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity RCA_N4_24 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_24;

architecture SYN_STRUCTURAL of RCA_N4_24 is

   component FA_93
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_94
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_95
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_96
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal n1, CTMP_3_port, CTMP_2_port, CTMP_1_port, net48787 : std_logic;

begin
   
   FAI_1 : FA_96 port map( A => A(0), B => B(0), Ci => n1, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_95 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_94 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_93 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => net48787);
   n1 <= '0';

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity RCA_N4_23 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_23;

architecture SYN_STRUCTURAL of RCA_N4_23 is

   component FA_89
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_90
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_91
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_92
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal n1, CTMP_3_port, CTMP_2_port, CTMP_1_port, net48786 : std_logic;

begin
   
   FAI_1 : FA_92 port map( A => A(0), B => B(0), Ci => n1, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_91 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_90 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_89 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => net48786);
   n1 <= '1';

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity RCA_N4_22 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_22;

architecture SYN_STRUCTURAL of RCA_N4_22 is

   component FA_85
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_86
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_87
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_88
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal n1, CTMP_3_port, CTMP_2_port, CTMP_1_port, net48785 : std_logic;

begin
   
   FAI_1 : FA_88 port map( A => A(0), B => B(0), Ci => n1, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_87 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_86 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_85 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => net48785);
   n1 <= '0';

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity RCA_N4_21 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_21;

architecture SYN_STRUCTURAL of RCA_N4_21 is

   component FA_81
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_82
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_83
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_84
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal n1, CTMP_3_port, CTMP_2_port, CTMP_1_port, net48784 : std_logic;

begin
   
   FAI_1 : FA_84 port map( A => A(0), B => B(0), Ci => n1, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_83 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_82 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_81 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => net48784);
   n1 <= '1';

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity RCA_N4_20 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_20;

architecture SYN_STRUCTURAL of RCA_N4_20 is

   component FA_77
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_78
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_79
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_80
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal n1, CTMP_3_port, CTMP_2_port, CTMP_1_port, net48783 : std_logic;

begin
   
   FAI_1 : FA_80 port map( A => A(0), B => B(0), Ci => n1, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_79 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_78 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_77 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => net48783);
   n1 <= '0';

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity RCA_N4_19 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_19;

architecture SYN_STRUCTURAL of RCA_N4_19 is

   component FA_73
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_74
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_75
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_76
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal n1, CTMP_3_port, CTMP_2_port, CTMP_1_port, net48782 : std_logic;

begin
   
   FAI_1 : FA_76 port map( A => A(0), B => B(0), Ci => n1, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_75 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_74 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_73 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => net48782);
   n1 <= '1';

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity RCA_N4_18 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_18;

architecture SYN_STRUCTURAL of RCA_N4_18 is

   component FA_69
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_70
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_71
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_72
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal n1, CTMP_3_port, CTMP_2_port, CTMP_1_port, net48781 : std_logic;

begin
   
   FAI_1 : FA_72 port map( A => A(0), B => B(0), Ci => n1, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_71 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_70 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_69 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => net48781);
   n1 <= '0';

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity RCA_N4_17 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_17;

architecture SYN_STRUCTURAL of RCA_N4_17 is

   component FA_65
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_66
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_67
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_68
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal n1, CTMP_3_port, CTMP_2_port, CTMP_1_port, net48780 : std_logic;

begin
   
   FAI_1 : FA_68 port map( A => A(0), B => B(0), Ci => n1, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_67 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_66 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_65 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => net48780);
   n1 <= '1';

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity RCA_N4_16 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_16;

architecture SYN_STRUCTURAL of RCA_N4_16 is

   component FA_61
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_62
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_63
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_64
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal n1, CTMP_3_port, CTMP_2_port, CTMP_1_port, net48779 : std_logic;

begin
   
   FAI_1 : FA_64 port map( A => A(0), B => B(0), Ci => n1, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_63 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_62 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_61 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => net48779);
   n1 <= '0';

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity RCA_N4_15 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_15;

architecture SYN_STRUCTURAL of RCA_N4_15 is

   component FA_57
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_58
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_59
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_60
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal n1, CTMP_3_port, CTMP_2_port, CTMP_1_port, net48778 : std_logic;

begin
   
   FAI_1 : FA_60 port map( A => A(0), B => B(0), Ci => n1, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_59 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_58 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_57 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => net48778);
   n1 <= '1';

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity RCA_N4_14 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_14;

architecture SYN_STRUCTURAL of RCA_N4_14 is

   component FA_53
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_54
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_55
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_56
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal n1, CTMP_3_port, CTMP_2_port, CTMP_1_port, net48777 : std_logic;

begin
   
   FAI_1 : FA_56 port map( A => A(0), B => B(0), Ci => n1, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_55 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_54 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_53 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => net48777);
   n1 <= '0';

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity RCA_N4_13 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_13;

architecture SYN_STRUCTURAL of RCA_N4_13 is

   component FA_49
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_50
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_51
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_52
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal n1, CTMP_3_port, CTMP_2_port, CTMP_1_port, net48776 : std_logic;

begin
   
   FAI_1 : FA_52 port map( A => A(0), B => B(0), Ci => n1, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_51 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_50 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_49 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => net48776);
   n1 <= '1';

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity RCA_N4_12 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_12;

architecture SYN_STRUCTURAL of RCA_N4_12 is

   component FA_45
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_46
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_47
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_48
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal n1, CTMP_3_port, CTMP_2_port, CTMP_1_port, net48775 : std_logic;

begin
   
   FAI_1 : FA_48 port map( A => A(0), B => B(0), Ci => n1, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_47 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_46 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_45 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => net48775);
   n1 <= '0';

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity RCA_N4_11 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_11;

architecture SYN_STRUCTURAL of RCA_N4_11 is

   component FA_41
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_42
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_43
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_44
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal n1, CTMP_3_port, CTMP_2_port, CTMP_1_port, net48774 : std_logic;

begin
   
   FAI_1 : FA_44 port map( A => A(0), B => B(0), Ci => n1, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_43 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_42 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_41 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => net48774);
   n1 <= '1';

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity RCA_N4_10 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_10;

architecture SYN_STRUCTURAL of RCA_N4_10 is

   component FA_37
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_38
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_39
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_40
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal n1, CTMP_3_port, CTMP_2_port, CTMP_1_port, net48773 : std_logic;

begin
   
   FAI_1 : FA_40 port map( A => A(0), B => B(0), Ci => n1, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_39 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_38 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_37 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => net48773);
   n1 <= '0';

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity RCA_N4_9 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_9;

architecture SYN_STRUCTURAL of RCA_N4_9 is

   component FA_33
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_34
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_35
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_36
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal n1, CTMP_3_port, CTMP_2_port, CTMP_1_port, net48772 : std_logic;

begin
   
   FAI_1 : FA_36 port map( A => A(0), B => B(0), Ci => n1, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_35 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_34 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_33 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => net48772);
   n1 <= '1';

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity RCA_N4_8 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_8;

architecture SYN_STRUCTURAL of RCA_N4_8 is

   component FA_29
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_30
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_31
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_32
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal n1, CTMP_3_port, CTMP_2_port, CTMP_1_port, net48771 : std_logic;

begin
   
   FAI_1 : FA_32 port map( A => A(0), B => B(0), Ci => n1, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_31 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_30 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_29 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => net48771);
   n1 <= '0';

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity RCA_N4_7 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_7;

architecture SYN_STRUCTURAL of RCA_N4_7 is

   component FA_25
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_26
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_27
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_28
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal n1, CTMP_3_port, CTMP_2_port, CTMP_1_port, net48770 : std_logic;

begin
   
   FAI_1 : FA_28 port map( A => A(0), B => B(0), Ci => n1, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_27 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_26 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_25 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => net48770);
   n1 <= '1';

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity RCA_N4_6 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_6;

architecture SYN_STRUCTURAL of RCA_N4_6 is

   component FA_21
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_22
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_23
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_24
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal n1, CTMP_3_port, CTMP_2_port, CTMP_1_port, net48769 : std_logic;

begin
   
   FAI_1 : FA_24 port map( A => A(0), B => B(0), Ci => n1, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_23 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_22 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_21 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => net48769);
   n1 <= '0';

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity RCA_N4_5 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_5;

architecture SYN_STRUCTURAL of RCA_N4_5 is

   component FA_17
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_18
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_19
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_20
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal n1, CTMP_3_port, CTMP_2_port, CTMP_1_port, net48768 : std_logic;

begin
   
   FAI_1 : FA_20 port map( A => A(0), B => B(0), Ci => n1, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_19 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_18 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_17 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => net48768);
   n1 <= '1';

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity RCA_N4_4 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_4;

architecture SYN_STRUCTURAL of RCA_N4_4 is

   component FA_13
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_14
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_15
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_16
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal n1, CTMP_3_port, CTMP_2_port, CTMP_1_port, net48767 : std_logic;

begin
   
   FAI_1 : FA_16 port map( A => A(0), B => B(0), Ci => n1, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_15 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_14 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_13 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => net48767);
   n1 <= '0';

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity RCA_N4_3 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_3;

architecture SYN_STRUCTURAL of RCA_N4_3 is

   component FA_9
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_10
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_11
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_12
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal n1, CTMP_3_port, CTMP_2_port, CTMP_1_port, net48766 : std_logic;

begin
   
   FAI_1 : FA_12 port map( A => A(0), B => B(0), Ci => n1, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_11 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_10 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_9 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => net48766);
   n1 <= '1';

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity RCA_N4_2 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_2;

architecture SYN_STRUCTURAL of RCA_N4_2 is

   component FA_5
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_6
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_7
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_8
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal n1, CTMP_3_port, CTMP_2_port, CTMP_1_port, net48765 : std_logic;

begin
   
   FAI_1 : FA_8 port map( A => A(0), B => B(0), Ci => n1, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_7 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_6 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_5 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => net48765);
   n1 <= '0';

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity RCA_N4_1 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_1;

architecture SYN_STRUCTURAL of RCA_N4_1 is

   component FA_1
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_2
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_3
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_4
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal n1, CTMP_3_port, CTMP_2_port, CTMP_1_port, net48764 : std_logic;

begin
   
   FAI_1 : FA_4 port map( A => A(0), B => B(0), Ci => n1, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_3 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_2 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_1 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => net48764);
   n1 <= '1';

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity shift_N9_2 is

   port( Clock, ALOAD : in std_logic;  D : in std_logic_vector (8 downto 0);  
         SO : out std_logic);

end shift_N9_2;

architecture SYN_archi of shift_N9_2 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component SDFF_X1
      port( D, SI, SE, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal tmp_8_port, tmp_7_port, tmp_6_port, tmp_5_port, tmp_4_port, 
      tmp_3_port, tmp_2_port, tmp_1_port, N11, n1, n10, n11_port, n12, n13, n14
      , n15, n16, n17 : std_logic;

begin
   
   tmp_reg_8_inst : DFF_X1 port map( D => N11, CK => Clock, Q => tmp_8_port, QN
                           => n1);
   tmp_reg_7_inst : SDFF_X1 port map( D => tmp_8_port, SI => D(7), SE => ALOAD,
                           CK => Clock, Q => tmp_7_port, QN => n10);
   tmp_reg_6_inst : SDFF_X1 port map( D => tmp_7_port, SI => D(6), SE => ALOAD,
                           CK => Clock, Q => tmp_6_port, QN => n11_port);
   tmp_reg_5_inst : SDFF_X1 port map( D => tmp_6_port, SI => D(5), SE => ALOAD,
                           CK => Clock, Q => tmp_5_port, QN => n12);
   tmp_reg_4_inst : SDFF_X1 port map( D => tmp_5_port, SI => D(4), SE => ALOAD,
                           CK => Clock, Q => tmp_4_port, QN => n13);
   tmp_reg_3_inst : SDFF_X1 port map( D => tmp_4_port, SI => D(3), SE => ALOAD,
                           CK => Clock, Q => tmp_3_port, QN => n14);
   tmp_reg_2_inst : SDFF_X1 port map( D => tmp_3_port, SI => D(2), SE => ALOAD,
                           CK => Clock, Q => tmp_2_port, QN => n15);
   tmp_reg_1_inst : SDFF_X1 port map( D => tmp_2_port, SI => D(1), SE => ALOAD,
                           CK => Clock, Q => tmp_1_port, QN => n16);
   tmp_reg_0_inst : SDFF_X1 port map( D => tmp_1_port, SI => D(0), SE => ALOAD,
                           CK => Clock, Q => SO, QN => n17);
   U3 : AND2_X1 port map( A1 => ALOAD, A2 => D(8), ZN => N11);

end SYN_archi;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity shift_N9_1 is

   port( Clock, ALOAD : in std_logic;  D : in std_logic_vector (8 downto 0);  
         SO : out std_logic);

end shift_N9_1;

architecture SYN_archi of shift_N9_1 is

   component SDFF_X2
      port( D, SI, SE, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component SDFF_X1
      port( D, SI, SE, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal tmp_8_port, tmp_7_port, tmp_6_port, tmp_5_port, tmp_4_port, 
      tmp_3_port, tmp_2_port, tmp_1_port, N11, n1, n2, n10, n11_port, n12, n13,
      n14, n15, n16 : std_logic;

begin
   
   tmp_reg_8_inst : DFF_X1 port map( D => N11, CK => Clock, Q => tmp_8_port, QN
                           => n2);
   tmp_reg_7_inst : SDFF_X1 port map( D => tmp_8_port, SI => D(7), SE => ALOAD,
                           CK => Clock, Q => tmp_7_port, QN => n10);
   tmp_reg_6_inst : SDFF_X1 port map( D => tmp_7_port, SI => D(6), SE => ALOAD,
                           CK => Clock, Q => tmp_6_port, QN => n11_port);
   tmp_reg_5_inst : SDFF_X1 port map( D => tmp_6_port, SI => D(5), SE => ALOAD,
                           CK => Clock, Q => tmp_5_port, QN => n12);
   tmp_reg_4_inst : SDFF_X1 port map( D => tmp_5_port, SI => D(4), SE => ALOAD,
                           CK => Clock, Q => tmp_4_port, QN => n13);
   tmp_reg_3_inst : SDFF_X1 port map( D => tmp_4_port, SI => D(3), SE => ALOAD,
                           CK => Clock, Q => tmp_3_port, QN => n14);
   tmp_reg_2_inst : SDFF_X1 port map( D => tmp_3_port, SI => D(2), SE => ALOAD,
                           CK => Clock, Q => tmp_2_port, QN => n15);
   tmp_reg_1_inst : SDFF_X1 port map( D => tmp_2_port, SI => D(1), SE => ALOAD,
                           CK => Clock, Q => tmp_1_port, QN => n16);
   U3 : AND2_X1 port map( A1 => ALOAD, A2 => D(8), ZN => N11);
   tmp_reg_0_inst : SDFF_X2 port map( D => tmp_1_port, SI => D(0), SE => ALOAD,
                           CK => Clock, Q => SO, QN => n1);

end SYN_archi;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity booth_encoder_8 is

   port( B_in : in std_logic_vector (2 downto 0);  A_out : out std_logic_vector
         (2 downto 0));

end booth_encoder_8;

architecture SYN_bhe of booth_encoder_8 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI33_X1
      port( A1, A2, A3, B1, B2, B3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n6, n7, n8, n9 : std_logic;

begin
   
   U6 : OAI33_X1 port map( A1 => B_in(0), A2 => B_in(1), A3 => n6, B1 => n9, B2
                           => n8, B3 => B_in(2), ZN => A_out(0));
   U4 : NAND2_X1 port map( A1 => B_in(2), A2 => n9, ZN => n7);
   U9 : INV_X1 port map( A => B_in(2), ZN => n6);
   U3 : INV_X1 port map( A => B_in(1), ZN => n8);
   U5 : INV_X1 port map( A => B_in(0), ZN => n9);
   U7 : OAI221_X1 port map( B1 => B_in(1), B2 => n9, C1 => n8, C2 => B_in(2), A
                           => n7, ZN => A_out(2));
   U8 : AOI21_X1 port map( B1 => B_in(0), B2 => B_in(1), A => n6, ZN => 
                           A_out(1));

end SYN_bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity booth_encoder_7 is

   port( B_in : in std_logic_vector (2 downto 0);  A_out : out std_logic_vector
         (2 downto 0));

end booth_encoder_7;

architecture SYN_bhe of booth_encoder_7 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI33_X1
      port( A1, A2, A3, B1, B2, B3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n6, n7, n8, n9 : std_logic;

begin
   
   U6 : OAI33_X1 port map( A1 => B_in(0), A2 => B_in(1), A3 => n6, B1 => n9, B2
                           => n8, B3 => B_in(2), ZN => A_out(0));
   U5 : AOI21_X1 port map( B1 => B_in(0), B2 => B_in(1), A => n6, ZN => 
                           A_out(1));
   U8 : INV_X1 port map( A => B_in(0), ZN => n9);
   U7 : INV_X1 port map( A => B_in(1), ZN => n8);
   U3 : INV_X1 port map( A => B_in(2), ZN => n6);
   U4 : OAI221_X1 port map( B1 => B_in(1), B2 => n9, C1 => n8, C2 => B_in(2), A
                           => n7, ZN => A_out(2));
   U9 : NAND2_X1 port map( A1 => B_in(2), A2 => n9, ZN => n7);

end SYN_bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity booth_encoder_6 is

   port( B_in : in std_logic_vector (2 downto 0);  A_out : out std_logic_vector
         (2 downto 0));

end booth_encoder_6;

architecture SYN_bhe of booth_encoder_6 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI33_X1
      port( A1, A2, A3, B1, B2, B3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n5, n6, n7 : std_logic;

begin
   
   U6 : OAI33_X1 port map( A1 => B_in(0), A2 => B_in(1), A3 => n1, B1 => n7, B2
                           => n6, B3 => B_in(2), ZN => A_out(0));
   U3 : INV_X1 port map( A => B_in(2), ZN => n1);
   U4 : INV_X1 port map( A => B_in(1), ZN => n6);
   U5 : INV_X1 port map( A => B_in(0), ZN => n7);
   U7 : NAND2_X1 port map( A1 => B_in(2), A2 => n7, ZN => n5);
   U8 : OAI221_X1 port map( B1 => B_in(1), B2 => n7, C1 => n6, C2 => B_in(2), A
                           => n5, ZN => A_out(2));
   U9 : AOI21_X1 port map( B1 => B_in(0), B2 => B_in(1), A => n1, ZN => 
                           A_out(1));

end SYN_bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity booth_encoder_5 is

   port( B_in : in std_logic_vector (2 downto 0);  A_out : out std_logic_vector
         (2 downto 0));

end booth_encoder_5;

architecture SYN_bhe of booth_encoder_5 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI33_X1
      port( A1, A2, A3, B1, B2, B3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n5, n6, n7 : std_logic;

begin
   
   U6 : OAI33_X1 port map( A1 => B_in(0), A2 => B_in(1), A3 => n1, B1 => n7, B2
                           => n6, B3 => B_in(2), ZN => A_out(0));
   U7 : INV_X1 port map( A => B_in(1), ZN => n6);
   U3 : INV_X1 port map( A => B_in(2), ZN => n1);
   U4 : INV_X1 port map( A => B_in(0), ZN => n7);
   U5 : AOI21_X1 port map( B1 => B_in(0), B2 => B_in(1), A => n1, ZN => 
                           A_out(1));
   U8 : OAI221_X1 port map( B1 => B_in(1), B2 => n7, C1 => n6, C2 => B_in(2), A
                           => n5, ZN => A_out(2));
   U9 : NAND2_X1 port map( A1 => B_in(2), A2 => n7, ZN => n5);

end SYN_bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity booth_encoder_4 is

   port( B_in : in std_logic_vector (2 downto 0);  A_out : out std_logic_vector
         (2 downto 0));

end booth_encoder_4;

architecture SYN_bhe of booth_encoder_4 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI33_X1
      port( A1, A2, A3, B1, B2, B3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n5, n6, n7 : std_logic;

begin
   
   U6 : OAI33_X1 port map( A1 => B_in(0), A2 => B_in(1), A3 => n1, B1 => n7, B2
                           => n6, B3 => B_in(2), ZN => A_out(0));
   U3 : INV_X1 port map( A => B_in(2), ZN => n1);
   U4 : INV_X1 port map( A => B_in(1), ZN => n6);
   U5 : INV_X1 port map( A => B_in(0), ZN => n7);
   U7 : OAI221_X1 port map( B1 => B_in(1), B2 => n7, C1 => n6, C2 => B_in(2), A
                           => n5, ZN => A_out(2));
   U8 : NAND2_X1 port map( A1 => B_in(2), A2 => n7, ZN => n5);
   U9 : AOI21_X1 port map( B1 => B_in(0), B2 => B_in(1), A => n1, ZN => 
                           A_out(1));

end SYN_bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity booth_encoder_3 is

   port( B_in : in std_logic_vector (2 downto 0);  A_out : out std_logic_vector
         (2 downto 0));

end booth_encoder_3;

architecture SYN_bhe of booth_encoder_3 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI33_X1
      port( A1, A2, A3, B1, B2, B3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n5, n6, n7 : std_logic;

begin
   
   U6 : OAI33_X1 port map( A1 => B_in(0), A2 => B_in(1), A3 => n1, B1 => n7, B2
                           => n6, B3 => B_in(2), ZN => A_out(0));
   U3 : INV_X1 port map( A => B_in(2), ZN => n1);
   U4 : INV_X1 port map( A => B_in(1), ZN => n6);
   U5 : INV_X1 port map( A => B_in(0), ZN => n7);
   U7 : AOI21_X1 port map( B1 => B_in(0), B2 => B_in(1), A => n1, ZN => 
                           A_out(1));
   U8 : OAI221_X1 port map( B1 => B_in(1), B2 => n7, C1 => n6, C2 => B_in(2), A
                           => n5, ZN => A_out(2));
   U9 : NAND2_X1 port map( A1 => B_in(2), A2 => n7, ZN => n5);

end SYN_bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity booth_encoder_2 is

   port( B_in : in std_logic_vector (2 downto 0);  A_out : out std_logic_vector
         (2 downto 0));

end booth_encoder_2;

architecture SYN_bhe of booth_encoder_2 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI33_X1
      port( A1, A2, A3, B1, B2, B3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n5, n6, n7 : std_logic;

begin
   
   U6 : OAI33_X1 port map( A1 => B_in(0), A2 => B_in(1), A3 => n1, B1 => n7, B2
                           => n6, B3 => B_in(2), ZN => A_out(0));
   U7 : INV_X1 port map( A => B_in(1), ZN => n6);
   U3 : INV_X1 port map( A => B_in(0), ZN => n7);
   U4 : INV_X1 port map( A => B_in(2), ZN => n1);
   U5 : NAND2_X1 port map( A1 => B_in(2), A2 => n7, ZN => n5);
   U8 : OAI221_X1 port map( B1 => B_in(1), B2 => n7, C1 => n6, C2 => B_in(2), A
                           => n5, ZN => A_out(2));
   U9 : AOI21_X1 port map( B1 => B_in(0), B2 => B_in(1), A => n1, ZN => 
                           A_out(1));

end SYN_bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity booth_encoder_1 is

   port( B_in : in std_logic_vector (2 downto 0);  A_out : out std_logic_vector
         (2 downto 0));

end booth_encoder_1;

architecture SYN_bhe of booth_encoder_1 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI33_X1
      port( A1, A2, A3, B1, B2, B3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4, n5 : std_logic;

begin
   
   U6 : OAI33_X1 port map( A1 => B_in(0), A2 => B_in(1), A3 => n4, B1 => n5, B2
                           => n4, B3 => B_in(2), ZN => A_out(0));
   U4 : NAND2_X1 port map( A1 => B_in(2), A2 => n5, ZN => n1);
   U3 : OAI221_X1 port map( B1 => B_in(1), B2 => n5, C1 => n4, C2 => B_in(2), A
                           => n1, ZN => A_out(2));
   U5 : INV_X1 port map( A => B_in(0), ZN => n5);
   U7 : INV_X1 port map( A => B_in(1), ZN => n4);
   U8 : AOI21_X1 port map( B1 => B_in(0), B2 => B_in(1), A => n4, ZN => 
                           A_out(1));

end SYN_bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity carry_sel_gen_N4_15 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end carry_sel_gen_N4_15;

architecture SYN_STRUCTURAL of carry_sel_gen_N4_15 is

   component mux21_SIZE4_15
      port( IN0, IN1 : in std_logic_vector (3 downto 0);  CTRL : in std_logic; 
            OUT1 : out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_N4_29
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_30
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, nocarry_sum_to_mux_3_port, 
      nocarry_sum_to_mux_2_port, nocarry_sum_to_mux_1_port, 
      nocarry_sum_to_mux_0_port, carry_sum_to_mux_3_port, 
      carry_sum_to_mux_2_port, carry_sum_to_mux_1_port, carry_sum_to_mux_0_port
      , net48762, net48763 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   rca_nocarry : RCA_N4_30 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           nocarry_sum_to_mux_3_port, S(2) => 
                           nocarry_sum_to_mux_2_port, S(1) => 
                           nocarry_sum_to_mux_1_port, S(0) => 
                           nocarry_sum_to_mux_0_port, Co => net48763);
   rca_carry : RCA_N4_29 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           carry_sum_to_mux_3_port, S(2) => 
                           carry_sum_to_mux_2_port, S(1) => 
                           carry_sum_to_mux_1_port, S(0) => 
                           carry_sum_to_mux_0_port, Co => net48762);
   outmux : mux21_SIZE4_15 port map( IN0(3) => nocarry_sum_to_mux_3_port, 
                           IN0(2) => nocarry_sum_to_mux_2_port, IN0(1) => 
                           nocarry_sum_to_mux_1_port, IN0(0) => 
                           nocarry_sum_to_mux_0_port, IN1(3) => 
                           carry_sum_to_mux_3_port, IN1(2) => 
                           carry_sum_to_mux_2_port, IN1(1) => 
                           carry_sum_to_mux_1_port, IN1(0) => 
                           carry_sum_to_mux_0_port, CTRL => Ci, OUT1(3) => S(3)
                           , OUT1(2) => S(2), OUT1(1) => S(1), OUT1(0) => S(0))
                           ;

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity carry_sel_gen_N4_14 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end carry_sel_gen_N4_14;

architecture SYN_STRUCTURAL of carry_sel_gen_N4_14 is

   component mux21_SIZE4_14
      port( IN0, IN1 : in std_logic_vector (3 downto 0);  CTRL : in std_logic; 
            OUT1 : out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_N4_27
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_28
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, nocarry_sum_to_mux_3_port, 
      nocarry_sum_to_mux_2_port, nocarry_sum_to_mux_1_port, 
      nocarry_sum_to_mux_0_port, carry_sum_to_mux_3_port, 
      carry_sum_to_mux_2_port, carry_sum_to_mux_1_port, carry_sum_to_mux_0_port
      , net48760, net48761 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   rca_nocarry : RCA_N4_28 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           nocarry_sum_to_mux_3_port, S(2) => 
                           nocarry_sum_to_mux_2_port, S(1) => 
                           nocarry_sum_to_mux_1_port, S(0) => 
                           nocarry_sum_to_mux_0_port, Co => net48761);
   rca_carry : RCA_N4_27 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           carry_sum_to_mux_3_port, S(2) => 
                           carry_sum_to_mux_2_port, S(1) => 
                           carry_sum_to_mux_1_port, S(0) => 
                           carry_sum_to_mux_0_port, Co => net48760);
   outmux : mux21_SIZE4_14 port map( IN0(3) => nocarry_sum_to_mux_3_port, 
                           IN0(2) => nocarry_sum_to_mux_2_port, IN0(1) => 
                           nocarry_sum_to_mux_1_port, IN0(0) => 
                           nocarry_sum_to_mux_0_port, IN1(3) => 
                           carry_sum_to_mux_3_port, IN1(2) => 
                           carry_sum_to_mux_2_port, IN1(1) => 
                           carry_sum_to_mux_1_port, IN1(0) => 
                           carry_sum_to_mux_0_port, CTRL => Ci, OUT1(3) => S(3)
                           , OUT1(2) => S(2), OUT1(1) => S(1), OUT1(0) => S(0))
                           ;

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity carry_sel_gen_N4_13 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end carry_sel_gen_N4_13;

architecture SYN_STRUCTURAL of carry_sel_gen_N4_13 is

   component mux21_SIZE4_13
      port( IN0, IN1 : in std_logic_vector (3 downto 0);  CTRL : in std_logic; 
            OUT1 : out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_N4_25
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_26
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, nocarry_sum_to_mux_3_port, 
      nocarry_sum_to_mux_2_port, nocarry_sum_to_mux_1_port, 
      nocarry_sum_to_mux_0_port, carry_sum_to_mux_3_port, 
      carry_sum_to_mux_2_port, carry_sum_to_mux_1_port, carry_sum_to_mux_0_port
      , net48758, net48759 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   rca_nocarry : RCA_N4_26 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           nocarry_sum_to_mux_3_port, S(2) => 
                           nocarry_sum_to_mux_2_port, S(1) => 
                           nocarry_sum_to_mux_1_port, S(0) => 
                           nocarry_sum_to_mux_0_port, Co => net48759);
   rca_carry : RCA_N4_25 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           carry_sum_to_mux_3_port, S(2) => 
                           carry_sum_to_mux_2_port, S(1) => 
                           carry_sum_to_mux_1_port, S(0) => 
                           carry_sum_to_mux_0_port, Co => net48758);
   outmux : mux21_SIZE4_13 port map( IN0(3) => nocarry_sum_to_mux_3_port, 
                           IN0(2) => nocarry_sum_to_mux_2_port, IN0(1) => 
                           nocarry_sum_to_mux_1_port, IN0(0) => 
                           nocarry_sum_to_mux_0_port, IN1(3) => 
                           carry_sum_to_mux_3_port, IN1(2) => 
                           carry_sum_to_mux_2_port, IN1(1) => 
                           carry_sum_to_mux_1_port, IN1(0) => 
                           carry_sum_to_mux_0_port, CTRL => Ci, OUT1(3) => S(3)
                           , OUT1(2) => S(2), OUT1(1) => S(1), OUT1(0) => S(0))
                           ;

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity carry_sel_gen_N4_12 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end carry_sel_gen_N4_12;

architecture SYN_STRUCTURAL of carry_sel_gen_N4_12 is

   component mux21_SIZE4_12
      port( IN0, IN1 : in std_logic_vector (3 downto 0);  CTRL : in std_logic; 
            OUT1 : out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_N4_23
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_24
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, nocarry_sum_to_mux_3_port, 
      nocarry_sum_to_mux_2_port, nocarry_sum_to_mux_1_port, 
      nocarry_sum_to_mux_0_port, carry_sum_to_mux_3_port, 
      carry_sum_to_mux_2_port, carry_sum_to_mux_1_port, carry_sum_to_mux_0_port
      , net48756, net48757 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   rca_nocarry : RCA_N4_24 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           nocarry_sum_to_mux_3_port, S(2) => 
                           nocarry_sum_to_mux_2_port, S(1) => 
                           nocarry_sum_to_mux_1_port, S(0) => 
                           nocarry_sum_to_mux_0_port, Co => net48757);
   rca_carry : RCA_N4_23 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           carry_sum_to_mux_3_port, S(2) => 
                           carry_sum_to_mux_2_port, S(1) => 
                           carry_sum_to_mux_1_port, S(0) => 
                           carry_sum_to_mux_0_port, Co => net48756);
   outmux : mux21_SIZE4_12 port map( IN0(3) => nocarry_sum_to_mux_3_port, 
                           IN0(2) => nocarry_sum_to_mux_2_port, IN0(1) => 
                           nocarry_sum_to_mux_1_port, IN0(0) => 
                           nocarry_sum_to_mux_0_port, IN1(3) => 
                           carry_sum_to_mux_3_port, IN1(2) => 
                           carry_sum_to_mux_2_port, IN1(1) => 
                           carry_sum_to_mux_1_port, IN1(0) => 
                           carry_sum_to_mux_0_port, CTRL => Ci, OUT1(3) => S(3)
                           , OUT1(2) => S(2), OUT1(1) => S(1), OUT1(0) => S(0))
                           ;

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity carry_sel_gen_N4_11 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end carry_sel_gen_N4_11;

architecture SYN_STRUCTURAL of carry_sel_gen_N4_11 is

   component mux21_SIZE4_11
      port( IN0, IN1 : in std_logic_vector (3 downto 0);  CTRL : in std_logic; 
            OUT1 : out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_N4_21
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_22
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, nocarry_sum_to_mux_3_port, 
      nocarry_sum_to_mux_2_port, nocarry_sum_to_mux_1_port, 
      nocarry_sum_to_mux_0_port, carry_sum_to_mux_3_port, 
      carry_sum_to_mux_2_port, carry_sum_to_mux_1_port, carry_sum_to_mux_0_port
      , net48754, net48755 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   rca_nocarry : RCA_N4_22 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           nocarry_sum_to_mux_3_port, S(2) => 
                           nocarry_sum_to_mux_2_port, S(1) => 
                           nocarry_sum_to_mux_1_port, S(0) => 
                           nocarry_sum_to_mux_0_port, Co => net48755);
   rca_carry : RCA_N4_21 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           carry_sum_to_mux_3_port, S(2) => 
                           carry_sum_to_mux_2_port, S(1) => 
                           carry_sum_to_mux_1_port, S(0) => 
                           carry_sum_to_mux_0_port, Co => net48754);
   outmux : mux21_SIZE4_11 port map( IN0(3) => nocarry_sum_to_mux_3_port, 
                           IN0(2) => nocarry_sum_to_mux_2_port, IN0(1) => 
                           nocarry_sum_to_mux_1_port, IN0(0) => 
                           nocarry_sum_to_mux_0_port, IN1(3) => 
                           carry_sum_to_mux_3_port, IN1(2) => 
                           carry_sum_to_mux_2_port, IN1(1) => 
                           carry_sum_to_mux_1_port, IN1(0) => 
                           carry_sum_to_mux_0_port, CTRL => Ci, OUT1(3) => S(3)
                           , OUT1(2) => S(2), OUT1(1) => S(1), OUT1(0) => S(0))
                           ;

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity carry_sel_gen_N4_10 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end carry_sel_gen_N4_10;

architecture SYN_STRUCTURAL of carry_sel_gen_N4_10 is

   component mux21_SIZE4_10
      port( IN0, IN1 : in std_logic_vector (3 downto 0);  CTRL : in std_logic; 
            OUT1 : out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_N4_19
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_20
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, nocarry_sum_to_mux_3_port, 
      nocarry_sum_to_mux_2_port, nocarry_sum_to_mux_1_port, 
      nocarry_sum_to_mux_0_port, carry_sum_to_mux_3_port, 
      carry_sum_to_mux_2_port, carry_sum_to_mux_1_port, carry_sum_to_mux_0_port
      , net48752, net48753 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   rca_nocarry : RCA_N4_20 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           nocarry_sum_to_mux_3_port, S(2) => 
                           nocarry_sum_to_mux_2_port, S(1) => 
                           nocarry_sum_to_mux_1_port, S(0) => 
                           nocarry_sum_to_mux_0_port, Co => net48753);
   rca_carry : RCA_N4_19 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           carry_sum_to_mux_3_port, S(2) => 
                           carry_sum_to_mux_2_port, S(1) => 
                           carry_sum_to_mux_1_port, S(0) => 
                           carry_sum_to_mux_0_port, Co => net48752);
   outmux : mux21_SIZE4_10 port map( IN0(3) => nocarry_sum_to_mux_3_port, 
                           IN0(2) => nocarry_sum_to_mux_2_port, IN0(1) => 
                           nocarry_sum_to_mux_1_port, IN0(0) => 
                           nocarry_sum_to_mux_0_port, IN1(3) => 
                           carry_sum_to_mux_3_port, IN1(2) => 
                           carry_sum_to_mux_2_port, IN1(1) => 
                           carry_sum_to_mux_1_port, IN1(0) => 
                           carry_sum_to_mux_0_port, CTRL => Ci, OUT1(3) => S(3)
                           , OUT1(2) => S(2), OUT1(1) => S(1), OUT1(0) => S(0))
                           ;

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity carry_sel_gen_N4_9 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end carry_sel_gen_N4_9;

architecture SYN_STRUCTURAL of carry_sel_gen_N4_9 is

   component mux21_SIZE4_9
      port( IN0, IN1 : in std_logic_vector (3 downto 0);  CTRL : in std_logic; 
            OUT1 : out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_N4_17
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_18
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, nocarry_sum_to_mux_3_port, 
      nocarry_sum_to_mux_2_port, nocarry_sum_to_mux_1_port, 
      nocarry_sum_to_mux_0_port, carry_sum_to_mux_3_port, 
      carry_sum_to_mux_2_port, carry_sum_to_mux_1_port, carry_sum_to_mux_0_port
      , net48750, net48751 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   rca_nocarry : RCA_N4_18 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           nocarry_sum_to_mux_3_port, S(2) => 
                           nocarry_sum_to_mux_2_port, S(1) => 
                           nocarry_sum_to_mux_1_port, S(0) => 
                           nocarry_sum_to_mux_0_port, Co => net48751);
   rca_carry : RCA_N4_17 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           carry_sum_to_mux_3_port, S(2) => 
                           carry_sum_to_mux_2_port, S(1) => 
                           carry_sum_to_mux_1_port, S(0) => 
                           carry_sum_to_mux_0_port, Co => net48750);
   outmux : mux21_SIZE4_9 port map( IN0(3) => nocarry_sum_to_mux_3_port, IN0(2)
                           => nocarry_sum_to_mux_2_port, IN0(1) => 
                           nocarry_sum_to_mux_1_port, IN0(0) => 
                           nocarry_sum_to_mux_0_port, IN1(3) => 
                           carry_sum_to_mux_3_port, IN1(2) => 
                           carry_sum_to_mux_2_port, IN1(1) => 
                           carry_sum_to_mux_1_port, IN1(0) => 
                           carry_sum_to_mux_0_port, CTRL => Ci, OUT1(3) => S(3)
                           , OUT1(2) => S(2), OUT1(1) => S(1), OUT1(0) => S(0))
                           ;

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity carry_sel_gen_N4_8 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end carry_sel_gen_N4_8;

architecture SYN_STRUCTURAL of carry_sel_gen_N4_8 is

   component mux21_SIZE4_8
      port( IN0, IN1 : in std_logic_vector (3 downto 0);  CTRL : in std_logic; 
            OUT1 : out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_N4_15
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_16
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, nocarry_sum_to_mux_3_port, 
      nocarry_sum_to_mux_2_port, nocarry_sum_to_mux_1_port, 
      nocarry_sum_to_mux_0_port, carry_sum_to_mux_3_port, 
      carry_sum_to_mux_2_port, carry_sum_to_mux_1_port, carry_sum_to_mux_0_port
      , net48748, net48749 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   rca_nocarry : RCA_N4_16 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           nocarry_sum_to_mux_3_port, S(2) => 
                           nocarry_sum_to_mux_2_port, S(1) => 
                           nocarry_sum_to_mux_1_port, S(0) => 
                           nocarry_sum_to_mux_0_port, Co => net48749);
   rca_carry : RCA_N4_15 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           carry_sum_to_mux_3_port, S(2) => 
                           carry_sum_to_mux_2_port, S(1) => 
                           carry_sum_to_mux_1_port, S(0) => 
                           carry_sum_to_mux_0_port, Co => net48748);
   outmux : mux21_SIZE4_8 port map( IN0(3) => nocarry_sum_to_mux_3_port, IN0(2)
                           => nocarry_sum_to_mux_2_port, IN0(1) => 
                           nocarry_sum_to_mux_1_port, IN0(0) => 
                           nocarry_sum_to_mux_0_port, IN1(3) => 
                           carry_sum_to_mux_3_port, IN1(2) => 
                           carry_sum_to_mux_2_port, IN1(1) => 
                           carry_sum_to_mux_1_port, IN1(0) => 
                           carry_sum_to_mux_0_port, CTRL => Ci, OUT1(3) => S(3)
                           , OUT1(2) => S(2), OUT1(1) => S(1), OUT1(0) => S(0))
                           ;

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity carry_sel_gen_N4_7 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end carry_sel_gen_N4_7;

architecture SYN_STRUCTURAL of carry_sel_gen_N4_7 is

   component mux21_SIZE4_7
      port( IN0, IN1 : in std_logic_vector (3 downto 0);  CTRL : in std_logic; 
            OUT1 : out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_N4_13
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_14
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, nocarry_sum_to_mux_3_port, 
      nocarry_sum_to_mux_2_port, nocarry_sum_to_mux_1_port, 
      nocarry_sum_to_mux_0_port, carry_sum_to_mux_3_port, 
      carry_sum_to_mux_2_port, carry_sum_to_mux_1_port, carry_sum_to_mux_0_port
      , net48746, net48747 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   rca_nocarry : RCA_N4_14 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           nocarry_sum_to_mux_3_port, S(2) => 
                           nocarry_sum_to_mux_2_port, S(1) => 
                           nocarry_sum_to_mux_1_port, S(0) => 
                           nocarry_sum_to_mux_0_port, Co => net48747);
   rca_carry : RCA_N4_13 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           carry_sum_to_mux_3_port, S(2) => 
                           carry_sum_to_mux_2_port, S(1) => 
                           carry_sum_to_mux_1_port, S(0) => 
                           carry_sum_to_mux_0_port, Co => net48746);
   outmux : mux21_SIZE4_7 port map( IN0(3) => nocarry_sum_to_mux_3_port, IN0(2)
                           => nocarry_sum_to_mux_2_port, IN0(1) => 
                           nocarry_sum_to_mux_1_port, IN0(0) => 
                           nocarry_sum_to_mux_0_port, IN1(3) => 
                           carry_sum_to_mux_3_port, IN1(2) => 
                           carry_sum_to_mux_2_port, IN1(1) => 
                           carry_sum_to_mux_1_port, IN1(0) => 
                           carry_sum_to_mux_0_port, CTRL => Ci, OUT1(3) => S(3)
                           , OUT1(2) => S(2), OUT1(1) => S(1), OUT1(0) => S(0))
                           ;

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity carry_sel_gen_N4_6 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end carry_sel_gen_N4_6;

architecture SYN_STRUCTURAL of carry_sel_gen_N4_6 is

   component mux21_SIZE4_6
      port( IN0, IN1 : in std_logic_vector (3 downto 0);  CTRL : in std_logic; 
            OUT1 : out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_N4_11
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_12
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, nocarry_sum_to_mux_3_port, 
      nocarry_sum_to_mux_2_port, nocarry_sum_to_mux_1_port, 
      nocarry_sum_to_mux_0_port, carry_sum_to_mux_3_port, 
      carry_sum_to_mux_2_port, carry_sum_to_mux_1_port, carry_sum_to_mux_0_port
      , net48744, net48745 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   rca_nocarry : RCA_N4_12 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           nocarry_sum_to_mux_3_port, S(2) => 
                           nocarry_sum_to_mux_2_port, S(1) => 
                           nocarry_sum_to_mux_1_port, S(0) => 
                           nocarry_sum_to_mux_0_port, Co => net48745);
   rca_carry : RCA_N4_11 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           carry_sum_to_mux_3_port, S(2) => 
                           carry_sum_to_mux_2_port, S(1) => 
                           carry_sum_to_mux_1_port, S(0) => 
                           carry_sum_to_mux_0_port, Co => net48744);
   outmux : mux21_SIZE4_6 port map( IN0(3) => nocarry_sum_to_mux_3_port, IN0(2)
                           => nocarry_sum_to_mux_2_port, IN0(1) => 
                           nocarry_sum_to_mux_1_port, IN0(0) => 
                           nocarry_sum_to_mux_0_port, IN1(3) => 
                           carry_sum_to_mux_3_port, IN1(2) => 
                           carry_sum_to_mux_2_port, IN1(1) => 
                           carry_sum_to_mux_1_port, IN1(0) => 
                           carry_sum_to_mux_0_port, CTRL => Ci, OUT1(3) => S(3)
                           , OUT1(2) => S(2), OUT1(1) => S(1), OUT1(0) => S(0))
                           ;

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity carry_sel_gen_N4_5 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end carry_sel_gen_N4_5;

architecture SYN_STRUCTURAL of carry_sel_gen_N4_5 is

   component mux21_SIZE4_5
      port( IN0, IN1 : in std_logic_vector (3 downto 0);  CTRL : in std_logic; 
            OUT1 : out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_N4_9
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_10
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, nocarry_sum_to_mux_3_port, 
      nocarry_sum_to_mux_2_port, nocarry_sum_to_mux_1_port, 
      nocarry_sum_to_mux_0_port, carry_sum_to_mux_3_port, 
      carry_sum_to_mux_2_port, carry_sum_to_mux_1_port, carry_sum_to_mux_0_port
      , net48742, net48743 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   rca_nocarry : RCA_N4_10 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           nocarry_sum_to_mux_3_port, S(2) => 
                           nocarry_sum_to_mux_2_port, S(1) => 
                           nocarry_sum_to_mux_1_port, S(0) => 
                           nocarry_sum_to_mux_0_port, Co => net48743);
   rca_carry : RCA_N4_9 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           carry_sum_to_mux_3_port, S(2) => 
                           carry_sum_to_mux_2_port, S(1) => 
                           carry_sum_to_mux_1_port, S(0) => 
                           carry_sum_to_mux_0_port, Co => net48742);
   outmux : mux21_SIZE4_5 port map( IN0(3) => nocarry_sum_to_mux_3_port, IN0(2)
                           => nocarry_sum_to_mux_2_port, IN0(1) => 
                           nocarry_sum_to_mux_1_port, IN0(0) => 
                           nocarry_sum_to_mux_0_port, IN1(3) => 
                           carry_sum_to_mux_3_port, IN1(2) => 
                           carry_sum_to_mux_2_port, IN1(1) => 
                           carry_sum_to_mux_1_port, IN1(0) => 
                           carry_sum_to_mux_0_port, CTRL => Ci, OUT1(3) => S(3)
                           , OUT1(2) => S(2), OUT1(1) => S(1), OUT1(0) => S(0))
                           ;

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity carry_sel_gen_N4_4 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end carry_sel_gen_N4_4;

architecture SYN_STRUCTURAL of carry_sel_gen_N4_4 is

   component mux21_SIZE4_4
      port( IN0, IN1 : in std_logic_vector (3 downto 0);  CTRL : in std_logic; 
            OUT1 : out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_N4_7
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_8
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, nocarry_sum_to_mux_3_port, 
      nocarry_sum_to_mux_2_port, nocarry_sum_to_mux_1_port, 
      nocarry_sum_to_mux_0_port, carry_sum_to_mux_3_port, 
      carry_sum_to_mux_2_port, carry_sum_to_mux_1_port, carry_sum_to_mux_0_port
      , net48740, net48741 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   rca_nocarry : RCA_N4_8 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           nocarry_sum_to_mux_3_port, S(2) => 
                           nocarry_sum_to_mux_2_port, S(1) => 
                           nocarry_sum_to_mux_1_port, S(0) => 
                           nocarry_sum_to_mux_0_port, Co => net48741);
   rca_carry : RCA_N4_7 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           carry_sum_to_mux_3_port, S(2) => 
                           carry_sum_to_mux_2_port, S(1) => 
                           carry_sum_to_mux_1_port, S(0) => 
                           carry_sum_to_mux_0_port, Co => net48740);
   outmux : mux21_SIZE4_4 port map( IN0(3) => nocarry_sum_to_mux_3_port, IN0(2)
                           => nocarry_sum_to_mux_2_port, IN0(1) => 
                           nocarry_sum_to_mux_1_port, IN0(0) => 
                           nocarry_sum_to_mux_0_port, IN1(3) => 
                           carry_sum_to_mux_3_port, IN1(2) => 
                           carry_sum_to_mux_2_port, IN1(1) => 
                           carry_sum_to_mux_1_port, IN1(0) => 
                           carry_sum_to_mux_0_port, CTRL => Ci, OUT1(3) => S(3)
                           , OUT1(2) => S(2), OUT1(1) => S(1), OUT1(0) => S(0))
                           ;

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity carry_sel_gen_N4_3 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end carry_sel_gen_N4_3;

architecture SYN_STRUCTURAL of carry_sel_gen_N4_3 is

   component mux21_SIZE4_3
      port( IN0, IN1 : in std_logic_vector (3 downto 0);  CTRL : in std_logic; 
            OUT1 : out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_N4_5
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_6
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, nocarry_sum_to_mux_3_port, 
      nocarry_sum_to_mux_2_port, nocarry_sum_to_mux_1_port, 
      nocarry_sum_to_mux_0_port, carry_sum_to_mux_3_port, 
      carry_sum_to_mux_2_port, carry_sum_to_mux_1_port, carry_sum_to_mux_0_port
      , net48738, net48739 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   rca_nocarry : RCA_N4_6 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           nocarry_sum_to_mux_3_port, S(2) => 
                           nocarry_sum_to_mux_2_port, S(1) => 
                           nocarry_sum_to_mux_1_port, S(0) => 
                           nocarry_sum_to_mux_0_port, Co => net48739);
   rca_carry : RCA_N4_5 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           carry_sum_to_mux_3_port, S(2) => 
                           carry_sum_to_mux_2_port, S(1) => 
                           carry_sum_to_mux_1_port, S(0) => 
                           carry_sum_to_mux_0_port, Co => net48738);
   outmux : mux21_SIZE4_3 port map( IN0(3) => nocarry_sum_to_mux_3_port, IN0(2)
                           => nocarry_sum_to_mux_2_port, IN0(1) => 
                           nocarry_sum_to_mux_1_port, IN0(0) => 
                           nocarry_sum_to_mux_0_port, IN1(3) => 
                           carry_sum_to_mux_3_port, IN1(2) => 
                           carry_sum_to_mux_2_port, IN1(1) => 
                           carry_sum_to_mux_1_port, IN1(0) => 
                           carry_sum_to_mux_0_port, CTRL => Ci, OUT1(3) => S(3)
                           , OUT1(2) => S(2), OUT1(1) => S(1), OUT1(0) => S(0))
                           ;

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity carry_sel_gen_N4_2 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end carry_sel_gen_N4_2;

architecture SYN_STRUCTURAL of carry_sel_gen_N4_2 is

   component mux21_SIZE4_2
      port( IN0, IN1 : in std_logic_vector (3 downto 0);  CTRL : in std_logic; 
            OUT1 : out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_N4_3
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_4
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, nocarry_sum_to_mux_3_port, 
      nocarry_sum_to_mux_2_port, nocarry_sum_to_mux_1_port, 
      nocarry_sum_to_mux_0_port, carry_sum_to_mux_3_port, 
      carry_sum_to_mux_2_port, carry_sum_to_mux_1_port, carry_sum_to_mux_0_port
      , net48736, net48737 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   rca_nocarry : RCA_N4_4 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           nocarry_sum_to_mux_3_port, S(2) => 
                           nocarry_sum_to_mux_2_port, S(1) => 
                           nocarry_sum_to_mux_1_port, S(0) => 
                           nocarry_sum_to_mux_0_port, Co => net48737);
   rca_carry : RCA_N4_3 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           carry_sum_to_mux_3_port, S(2) => 
                           carry_sum_to_mux_2_port, S(1) => 
                           carry_sum_to_mux_1_port, S(0) => 
                           carry_sum_to_mux_0_port, Co => net48736);
   outmux : mux21_SIZE4_2 port map( IN0(3) => nocarry_sum_to_mux_3_port, IN0(2)
                           => nocarry_sum_to_mux_2_port, IN0(1) => 
                           nocarry_sum_to_mux_1_port, IN0(0) => 
                           nocarry_sum_to_mux_0_port, IN1(3) => 
                           carry_sum_to_mux_3_port, IN1(2) => 
                           carry_sum_to_mux_2_port, IN1(1) => 
                           carry_sum_to_mux_1_port, IN1(0) => 
                           carry_sum_to_mux_0_port, CTRL => Ci, OUT1(3) => S(3)
                           , OUT1(2) => S(2), OUT1(1) => S(1), OUT1(0) => S(0))
                           ;

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity carry_sel_gen_N4_1 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end carry_sel_gen_N4_1;

architecture SYN_STRUCTURAL of carry_sel_gen_N4_1 is

   component mux21_SIZE4_1
      port( IN0, IN1 : in std_logic_vector (3 downto 0);  CTRL : in std_logic; 
            OUT1 : out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_N4_1
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_2
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, nocarry_sum_to_mux_3_port, 
      nocarry_sum_to_mux_2_port, nocarry_sum_to_mux_1_port, 
      nocarry_sum_to_mux_0_port, carry_sum_to_mux_3_port, 
      carry_sum_to_mux_2_port, carry_sum_to_mux_1_port, carry_sum_to_mux_0_port
      , net48734, net48735 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   rca_nocarry : RCA_N4_2 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           nocarry_sum_to_mux_3_port, S(2) => 
                           nocarry_sum_to_mux_2_port, S(1) => 
                           nocarry_sum_to_mux_1_port, S(0) => 
                           nocarry_sum_to_mux_0_port, Co => net48735);
   rca_carry : RCA_N4_1 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           carry_sum_to_mux_3_port, S(2) => 
                           carry_sum_to_mux_2_port, S(1) => 
                           carry_sum_to_mux_1_port, S(0) => 
                           carry_sum_to_mux_0_port, Co => net48734);
   outmux : mux21_SIZE4_1 port map( IN0(3) => nocarry_sum_to_mux_3_port, IN0(2)
                           => nocarry_sum_to_mux_2_port, IN0(1) => 
                           nocarry_sum_to_mux_1_port, IN0(0) => 
                           nocarry_sum_to_mux_0_port, IN1(3) => 
                           carry_sum_to_mux_3_port, IN1(2) => 
                           carry_sum_to_mux_2_port, IN1(1) => 
                           carry_sum_to_mux_1_port, IN1(0) => 
                           carry_sum_to_mux_0_port, CTRL => Ci, OUT1(3) => S(3)
                           , OUT1(2) => S(2), OUT1(1) => S(1), OUT1(0) => S(0))
                           ;

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_53 is

   port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic);

end pg_53;

architecture SYN_beh of pg_53 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U3 : AOI21_X1 port map( B1 => g_prec, B2 => p, A => g, ZN => n1);
   U1 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);
   U2 : INV_X1 port map( A => n1, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_52 is

   port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic);

end pg_52;

architecture SYN_beh of pg_52 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U3 : AOI21_X1 port map( B1 => g_prec, B2 => p, A => g, ZN => n1);
   U1 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);
   U2 : INV_X1 port map( A => n1, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_51 is

   port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic);

end pg_51;

architecture SYN_beh of pg_51 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U3 : AOI21_X1 port map( B1 => g_prec, B2 => p, A => g, ZN => n1);
   U1 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);
   U2 : INV_X1 port map( A => n1, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_50 is

   port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic);

end pg_50;

architecture SYN_beh of pg_50 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U3 : AOI21_X1 port map( B1 => g_prec, B2 => p, A => g, ZN => n1);
   U1 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);
   U2 : INV_X1 port map( A => n1, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_49 is

   port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic);

end pg_49;

architecture SYN_beh of pg_49 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U3 : AOI21_X1 port map( B1 => g_prec, B2 => p, A => g, ZN => n1);
   U1 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);
   U2 : INV_X1 port map( A => n1, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_48 is

   port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic);

end pg_48;

architecture SYN_beh of pg_48 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U3 : AOI21_X1 port map( B1 => g_prec, B2 => p, A => g, ZN => n1);
   U1 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);
   U2 : INV_X1 port map( A => n1, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_47 is

   port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic);

end pg_47;

architecture SYN_beh of pg_47 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);
   U2 : INV_X1 port map( A => g, ZN => n2);
   U3 : NAND2_X1 port map( A1 => p, A2 => g_prec, ZN => n1);
   U4 : NAND2_X1 port map( A1 => n1, A2 => n2, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_46 is

   port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic);

end pg_46;

architecture SYN_beh of pg_46 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => g, ZN => n2);
   U2 : AND2_X1 port map( A1 => p_prec, A2 => p, ZN => p_out);
   U3 : NAND2_X1 port map( A1 => g_prec, A2 => p, ZN => n1);
   U4 : NAND2_X1 port map( A1 => n1, A2 => n2, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_45 is

   port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic);

end pg_45;

architecture SYN_beh of pg_45 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => g, ZN => n2);
   U2 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);
   U3 : NAND2_X1 port map( A1 => p, A2 => g_prec, ZN => n1);
   U4 : NAND2_X1 port map( A1 => n1, A2 => n2, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_44 is

   port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic);

end pg_44;

architecture SYN_beh of pg_44 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => p, B2 => g_prec, A => g, ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => g_out);
   U3 : AND2_X1 port map( A1 => p_prec, A2 => p, ZN => p_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_43 is

   port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic);

end pg_43;

architecture SYN_beh of pg_43 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);
   U2 : AOI21_X1 port map( B1 => g_prec, B2 => p, A => g, ZN => n1);
   U3 : INV_X1 port map( A => n1, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_42 is

   port( g, p, g_prec, p_prec : in std_logic;  p_out, g_out_BAR : out std_logic
         );

end pg_42;

architecture SYN_beh of pg_42 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);
   U2 : AOI21_X1 port map( B1 => p, B2 => g_prec, A => g, ZN => g_out_BAR);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_39 is

   port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic);

end pg_39;

architecture SYN_beh of pg_39 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U3 : AOI21_X1 port map( B1 => g_prec, B2 => p, A => g, ZN => n1);
   U1 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);
   U2 : INV_X1 port map( A => n1, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_38 is

   port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic);

end pg_38;

architecture SYN_beh of pg_38 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U3 : AOI21_X1 port map( B1 => g_prec, B2 => p, A => g, ZN => n1);
   U1 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);
   U2 : INV_X1 port map( A => n1, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_37 is

   port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic);

end pg_37;

architecture SYN_beh of pg_37 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U3 : AOI21_X1 port map( B1 => g_prec, B2 => p, A => g, ZN => n1);
   U1 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);
   U2 : INV_X1 port map( A => n1, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_36 is

   port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic);

end pg_36;

architecture SYN_beh of pg_36 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);
   U2 : INV_X1 port map( A => g, ZN => n2);
   U3 : NAND2_X1 port map( A1 => n1, A2 => n2, ZN => g_out);
   U4 : NAND2_X1 port map( A1 => g_prec, A2 => p, ZN => n1);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_35 is

   port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic);

end pg_35;

architecture SYN_beh of pg_35 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);
   U2 : INV_X1 port map( A => g, ZN => n2);
   U3 : NAND2_X1 port map( A1 => n1, A2 => n2, ZN => g_out);
   U4 : NAND2_X1 port map( A1 => g_prec, A2 => p, ZN => n1);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_34 is

   port( p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic;  
         g_BAR : in std_logic);

end pg_34;

architecture SYN_beh of pg_34 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);
   U2 : NAND2_X1 port map( A1 => g_prec, A2 => p, ZN => n1);
   U3 : NAND2_X1 port map( A1 => n1, A2 => g_BAR, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_32 is

   port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic);

end pg_32;

architecture SYN_beh of pg_32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U3 : AOI21_X1 port map( B1 => g_prec, B2 => p, A => g, ZN => n1);
   U1 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);
   U2 : INV_X1 port map( A => n1, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_31 is

   port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic);

end pg_31;

architecture SYN_beh of pg_31 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);
   U2 : INV_X1 port map( A => n1, ZN => g_out);
   U3 : AOI21_X1 port map( B1 => g_prec, B2 => p, A => g, ZN => n1);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_29 is

   port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic);

end pg_29;

architecture SYN_beh of pg_29 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);
   U2 : INV_X1 port map( A => g, ZN => n2);
   U3 : NAND2_X1 port map( A1 => n1, A2 => n2, ZN => g_out);
   U4 : NAND2_X1 port map( A1 => g_prec, A2 => p, ZN => n1);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_27 is

   port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic);

end pg_27;

architecture SYN_beh of pg_27 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => g, ZN => n2);
   U2 : AND2_X1 port map( A1 => p_prec, A2 => p, ZN => p_out);
   U3 : NAND2_X1 port map( A1 => p, A2 => g_prec, ZN => n1);
   U4 : NAND2_X1 port map( A1 => n1, A2 => n2, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_26 is

   port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic);

end pg_26;

architecture SYN_beh of pg_26 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => g_prec, B2 => p, A => g, ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => g_out);
   U3 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_25 is

   port( g, p, g_prec, p_prec : in std_logic;  p_out, g_out_BAR : out std_logic
         );

end pg_25;

architecture SYN_beh of pg_25 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p_prec, A2 => p, ZN => p_out);
   U2 : AOI21_X1 port map( B1 => p, B2 => g_prec, A => g, ZN => g_out_BAR);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_24 is

   port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic);

end pg_24;

architecture SYN_beh of pg_24 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => g_prec, B2 => p, A => g, ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => g_out);
   U3 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_23 is

   port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic);

end pg_23;

architecture SYN_beh of pg_23 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => g, ZN => n2);
   U2 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);
   U3 : NAND2_X1 port map( A1 => p, A2 => g_prec, ZN => n1);
   U4 : NAND2_X1 port map( A1 => n1, A2 => n2, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_22 is

   port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic);

end pg_22;

architecture SYN_beh of pg_22 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => g_out);
   U2 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);
   U3 : AOI21_X1 port map( B1 => p, B2 => g_prec, A => g, ZN => n1);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_21 is

   port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic);

end pg_21;

architecture SYN_beh of pg_21 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => g_out);
   U2 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);
   U3 : AOI21_X1 port map( B1 => p, B2 => g_prec, A => g, ZN => n1);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_20 is

   port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic);

end pg_20;

architecture SYN_beh of pg_20 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);
   U2 : INV_X1 port map( A => n1, ZN => g_out);
   U3 : AOI21_X1 port map( B1 => g_prec, B2 => p, A => g, ZN => n1);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_19 is

   port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic);

end pg_19;

architecture SYN_beh of pg_19 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => g_out);
   U2 : AND2_X1 port map( A1 => p_prec, A2 => p, ZN => p_out);
   U3 : AOI21_X1 port map( B1 => p, B2 => g_prec, A => g, ZN => n1);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_18 is

   port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic);

end pg_18;

architecture SYN_beh of pg_18 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => g_out);
   U2 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);
   U3 : AOI21_X1 port map( B1 => p, B2 => g_prec, A => g, ZN => n3);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_17 is

   port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic);

end pg_17;

architecture SYN_beh of pg_17 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => g_out);
   U2 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);
   U3 : AOI21_X1 port map( B1 => p, B2 => g_prec, A => g, ZN => n1);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_16 is

   port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic);

end pg_16;

architecture SYN_beh of pg_16 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U2 : INV_X1 port map( A => n1, ZN => g_out);
   U1 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);
   U3 : AOI21_X1 port map( B1 => g_prec, B2 => p, A => g, ZN => n1);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_15 is

   port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic);

end pg_15;

architecture SYN_beh of pg_15 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U2 : INV_X1 port map( A => n1, ZN => g_out);
   U1 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);
   U3 : AOI21_X1 port map( B1 => g_prec, B2 => p, A => g, ZN => n1);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_14 is

   port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic);

end pg_14;

architecture SYN_beh of pg_14 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U3 : AOI21_X1 port map( B1 => g_prec, B2 => p, A => g, ZN => n1);
   U1 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);
   U2 : INV_X1 port map( A => n1, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_13 is

   port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic);

end pg_13;

architecture SYN_beh of pg_13 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U3 : AOI21_X1 port map( B1 => g_prec, B2 => p, A => g, ZN => n1);
   U1 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);
   U2 : INV_X1 port map( A => n1, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_12 is

   port( p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic;  
         g_BAR : in std_logic);

end pg_12;

architecture SYN_beh of pg_12 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);
   U2 : NAND2_X1 port map( A1 => g_prec, A2 => p, ZN => n1);
   U3 : NAND2_X1 port map( A1 => n1, A2 => g_BAR, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_11 is

   port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic);

end pg_11;

architecture SYN_beh of pg_11 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => g_out);
   U2 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);
   U3 : AOI21_X1 port map( B1 => g_prec, B2 => p, A => g, ZN => n1);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_10 is

   port( g, p, g_prec, p_prec : in std_logic;  p_out, g_out_BAR : out std_logic
         );

end pg_10;

architecture SYN_beh of pg_10 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);
   U2 : AOI21_X1 port map( B1 => g_prec, B2 => p, A => g, ZN => g_out_BAR);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_9 is

   port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic);

end pg_9;

architecture SYN_beh of pg_9 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);
   U2 : INV_X1 port map( A => n1, ZN => g_out);
   U3 : AOI21_X1 port map( B1 => p, B2 => g_prec, A => g, ZN => n1);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_8 is

   port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic);

end pg_8;

architecture SYN_beh of pg_8 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => g_out);
   U2 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);
   U3 : AOI21_X1 port map( B1 => p, B2 => g_prec, A => g, ZN => n1);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_7 is

   port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic);

end pg_7;

architecture SYN_beh of pg_7 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U3 : AOI21_X1 port map( B1 => g_prec, B2 => p, A => g, ZN => n1);
   U1 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);
   U2 : INV_X1 port map( A => n1, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_6 is

   port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic);

end pg_6;

architecture SYN_beh of pg_6 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U3 : AOI21_X1 port map( B1 => g_prec, B2 => p, A => g, ZN => n1);
   U1 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);
   U2 : INV_X1 port map( A => n1, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_5 is

   port( p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic;  
         g_BAR : in std_logic);

end pg_5;

architecture SYN_beh of pg_5 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);
   U2 : NAND2_X1 port map( A1 => g_prec, A2 => p, ZN => n1);
   U3 : NAND2_X1 port map( A1 => n1, A2 => g_BAR, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_4 is

   port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic);

end pg_4;

architecture SYN_beh of pg_4 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);
   U2 : INV_X1 port map( A => n1, ZN => g_out);
   U3 : AOI21_X1 port map( B1 => g_prec, B2 => p, A => g, ZN => n1);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_3 is

   port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic);

end pg_3;

architecture SYN_beh of pg_3 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);
   U2 : INV_X1 port map( A => n1, ZN => g_out);
   U3 : AOI21_X1 port map( B1 => g_prec, B2 => p, A => g, ZN => n1);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_2 is

   port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic);

end pg_2;

architecture SYN_beh of pg_2 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);
   U2 : INV_X1 port map( A => n1, ZN => g_out);
   U3 : AOI21_X1 port map( B1 => g_prec, B2 => p, A => g, ZN => n1);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_1 is

   port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic);

end pg_1;

architecture SYN_beh of pg_1 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);
   U2 : INV_X1 port map( A => n1, ZN => g_out);
   U3 : AOI21_X1 port map( B1 => g_prec, B2 => p, A => g, ZN => n1);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity g_19 is

   port( g, p, g_prec : in std_logic;  g_out : out std_logic);

end g_19;

architecture SYN_beh of g_19 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U2 : AOI21_X1 port map( B1 => p, B2 => g_prec, A => g, ZN => n1);
   U1 : INV_X1 port map( A => n1, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity g_18 is

   port( g, p, g_prec : in std_logic;  g_out : out std_logic);

end g_18;

architecture SYN_beh of g_18 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U2 : AOI21_X1 port map( B1 => p, B2 => g_prec, A => g, ZN => n1);
   U1 : INV_X1 port map( A => n1, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity g_17 is

   port( g, p, g_prec : in std_logic;  g_out : out std_logic);

end g_17;

architecture SYN_beh of g_17 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U2 : AOI21_X1 port map( B1 => p, B2 => g_prec, A => g, ZN => n1);
   U1 : INV_X1 port map( A => n1, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity g_16 is

   port( g, p, g_prec : in std_logic;  g_out : out std_logic);

end g_16;

architecture SYN_beh of g_16 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U2 : AOI21_X1 port map( B1 => p, B2 => g_prec, A => g, ZN => n1);
   U1 : INV_X1 port map( A => n1, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity g_15 is

   port( g, p, g_prec : in std_logic;  g_out : out std_logic);

end g_15;

architecture SYN_beh of g_15 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U2 : AOI21_X1 port map( B1 => p, B2 => g_prec, A => g, ZN => n1);
   U1 : INV_X1 port map( A => n1, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity g_14 is

   port( g, p, g_prec : in std_logic;  g_out : out std_logic);

end g_14;

architecture SYN_beh of g_14 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => g_out);
   U2 : AOI21_X1 port map( B1 => p, B2 => g_prec, A => g, ZN => n1);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity g_13 is

   port( g, p, g_prec : in std_logic;  g_out : out std_logic);

end g_13;

architecture SYN_beh of g_13 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => g_out);
   U2 : AOI21_X1 port map( B1 => p, B2 => g_prec, A => g, ZN => n1);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity g_12 is

   port( g, p, g_prec : in std_logic;  g_out : out std_logic);

end g_12;

architecture SYN_beh of g_12 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : OR2_X2 port map( A1 => g, A2 => n1, ZN => g_out);
   U2 : AND2_X1 port map( A1 => p, A2 => g_prec, ZN => n1);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity g_10 is

   port( g, p, g_prec : in std_logic;  g_out : out std_logic);

end g_10;

architecture SYN_beh of g_10 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => g, ZN => n3);
   U2 : NAND2_X1 port map( A1 => n2, A2 => n3, ZN => g_out);
   U3 : NAND2_X1 port map( A1 => p, A2 => g_prec, ZN => n2);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity g_9 is

   port( g, p, g_prec : in std_logic;  g_out : out std_logic);

end g_9;

architecture SYN_beh of g_9 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => g, ZN => n2);
   U2 : NAND2_X1 port map( A1 => n1, A2 => n2, ZN => g_out);
   U3 : NAND2_X1 port map( A1 => g_prec, A2 => p, ZN => n1);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity g_8 is

   port( g, p, g_prec : in std_logic;  g_out : out std_logic);

end g_8;

architecture SYN_beh of g_8 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => g_out);
   U2 : AOI21_X1 port map( B1 => g_prec, B2 => p, A => g, ZN => n1);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity g_7 is

   port( g, p, g_prec : in std_logic;  g_out : out std_logic);

end g_7;

architecture SYN_beh of g_7 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => g_out);
   U2 : INV_X1 port map( A => g, ZN => n1);
   U3 : NAND2_X1 port map( A1 => g_prec, A2 => p, ZN => n2);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity g_6 is

   port( g, p, g_prec : in std_logic;  g_out : out std_logic);

end g_6;

architecture SYN_beh of g_6 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => g_prec, B2 => p, A => g, ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity g_5 is

   port( g, p, g_prec : in std_logic;  g_out : out std_logic);

end g_5;

architecture SYN_beh of g_5 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => g_out);
   U2 : AOI21_X1 port map( B1 => g_prec, B2 => p, A => g, ZN => n1);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity g_4 is

   port( g, p, g_prec : in std_logic;  g_out : out std_logic);

end g_4;

architecture SYN_beh of g_4 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n1, A2 => n2, ZN => g_out);
   U2 : INV_X1 port map( A => g, ZN => n2);
   U3 : NAND2_X1 port map( A1 => g_prec, A2 => p, ZN => n1);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity g_3 is

   port( g, p, g_prec : in std_logic;  g_out : out std_logic);

end g_3;

architecture SYN_beh of g_3 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => g_out);
   U2 : AOI21_X1 port map( B1 => p, B2 => g_prec, A => g, ZN => n1);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity g_2 is

   port( g, p, g_prec : in std_logic;  g_out : out std_logic);

end g_2;

architecture SYN_beh of g_2 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => g_out);
   U2 : AOI21_X1 port map( B1 => g_prec, B2 => p, A => g, ZN => n1);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity g_1 is

   port( g, p, g_prec : in std_logic;  g_out_BAR : out std_logic);

end g_1;

architecture SYN_beh of g_1 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AOI21_X1 port map( B1 => p, B2 => g_prec, A => g, ZN => g_out_BAR);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_63 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_63;

architecture SYN_beh of pg_net_63 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_62 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_62;

architecture SYN_beh of pg_net_62 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_61 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_61;

architecture SYN_beh of pg_net_61 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_60 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_60;

architecture SYN_beh of pg_net_60 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_59 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_59;

architecture SYN_beh of pg_net_59 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_58 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_58;

architecture SYN_beh of pg_net_58 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_57 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_57;

architecture SYN_beh of pg_net_57 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_56 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_56;

architecture SYN_beh of pg_net_56 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_55 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_55;

architecture SYN_beh of pg_net_55 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_54 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_54;

architecture SYN_beh of pg_net_54 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_53 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_53;

architecture SYN_beh of pg_net_53 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_52 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_52;

architecture SYN_beh of pg_net_52 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_51 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_51;

architecture SYN_beh of pg_net_51 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_50 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_50;

architecture SYN_beh of pg_net_50 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_49 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_49;

architecture SYN_beh of pg_net_49 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_48 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_48;

architecture SYN_beh of pg_net_48 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);
   U2 : INV_X1 port map( A => a, ZN => n1);
   U3 : XNOR2_X1 port map( A => b, B => n1, ZN => p_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_47 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_47;

architecture SYN_beh of pg_net_47 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);
   U2 : INV_X1 port map( A => a, ZN => n1);
   U3 : XNOR2_X1 port map( A => b, B => n1, ZN => p_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_46 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_46;

architecture SYN_beh of pg_net_46 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_45 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_45;

architecture SYN_beh of pg_net_45 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_44 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_44;

architecture SYN_beh of pg_net_44 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U2 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_43 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_43;

architecture SYN_beh of pg_net_43 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);
   U2 : INV_X1 port map( A => a, ZN => n1);
   U3 : XNOR2_X1 port map( A => b, B => n1, ZN => p_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_42 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_42;

architecture SYN_beh of pg_net_42 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);
   U2 : INV_X1 port map( A => a, ZN => n1);
   U3 : XNOR2_X1 port map( A => b, B => n1, ZN => p_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_41 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_41;

architecture SYN_beh of pg_net_41 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => a, A2 => b, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_40 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_40;

architecture SYN_beh of pg_net_40 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_39 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_39;

architecture SYN_beh of pg_net_39 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_38 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_38;

architecture SYN_beh of pg_net_38 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_33 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_33;

architecture SYN_beh of pg_net_33 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_32 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_32;

architecture SYN_beh of pg_net_32 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n4, n5 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);
   U2 : INV_X1 port map( A => b, ZN => n2);
   U3 : INV_X1 port map( A => a, ZN => n3);
   U4 : NAND2_X1 port map( A1 => n2, A2 => a, ZN => n5);
   U5 : NAND2_X1 port map( A1 => b, A2 => n3, ZN => n4);
   U6 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => p_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_31 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_31;

architecture SYN_beh of pg_net_31 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_30 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_30;

architecture SYN_beh of pg_net_30 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_29 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_29;

architecture SYN_beh of pg_net_29 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_28 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_28;

architecture SYN_beh of pg_net_28 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);
   U2 : XOR2_X1 port map( A => a, B => b, Z => p_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_27 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_27;

architecture SYN_beh of pg_net_27 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);
   U2 : INV_X1 port map( A => a, ZN => n1);
   U3 : XNOR2_X1 port map( A => b, B => n1, ZN => p_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_26 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_26;

architecture SYN_beh of pg_net_26 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_25 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_25;

architecture SYN_beh of pg_net_25 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => a, A2 => b, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_24 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_24;

architecture SYN_beh of pg_net_24 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_23 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_23;

architecture SYN_beh of pg_net_23 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_22 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_22;

architecture SYN_beh of pg_net_22 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_21 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_21;

architecture SYN_beh of pg_net_21 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_20 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_20;

architecture SYN_beh of pg_net_20 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_19 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_19;

architecture SYN_beh of pg_net_19 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_18 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_18;

architecture SYN_beh of pg_net_18 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_17 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_17;

architecture SYN_beh of pg_net_17 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_16 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_16;

architecture SYN_beh of pg_net_16 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_15 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_15;

architecture SYN_beh of pg_net_15 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_14 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_14;

architecture SYN_beh of pg_net_14 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_13 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_13;

architecture SYN_beh of pg_net_13 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_12 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_12;

architecture SYN_beh of pg_net_12 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_11 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_11;

architecture SYN_beh of pg_net_11 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_10 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_10;

architecture SYN_beh of pg_net_10 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_9 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_9;

architecture SYN_beh of pg_net_9 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_8 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_8;

architecture SYN_beh of pg_net_8 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_7 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_7;

architecture SYN_beh of pg_net_7 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_6 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_6;

architecture SYN_beh of pg_net_6 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_5 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_5;

architecture SYN_beh of pg_net_5 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_4 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_4;

architecture SYN_beh of pg_net_4 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_3 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_3;

architecture SYN_beh of pg_net_3 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_2 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_2;

architecture SYN_beh of pg_net_2 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_1 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_1;

architecture SYN_beh of pg_net_1 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : CLKBUF_X1 port map( A => b, Z => n1);
   U3 : AND2_X1 port map( A1 => n1, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity sum_gen_N32_1 is

   port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic_vector 
         (8 downto 0);  S : out std_logic_vector (31 downto 0));

end sum_gen_N32_1;

architecture SYN_STRUCTURAL of sum_gen_N32_1 is

   component carry_sel_gen_N4_1
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component carry_sel_gen_N4_2
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component carry_sel_gen_N4_3
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component carry_sel_gen_N4_4
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component carry_sel_gen_N4_5
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component carry_sel_gen_N4_6
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component carry_sel_gen_N4_7
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component carry_sel_gen_N4_8
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal net3145, net3146, net3147, net3148, net3149, net3150, net3151, 
      net3152 : std_logic;

begin
   
   csel_N_0 : carry_sel_gen_N4_8 port map( A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), Ci => Cin(0), S(3) => S(3), 
                           S(2) => S(2), S(1) => S(1), S(0) => S(0), Co => 
                           net3152);
   csel_N_1 : carry_sel_gen_N4_7 port map( A(3) => A(7), A(2) => A(6), A(1) => 
                           A(5), A(0) => A(4), B(3) => B(7), B(2) => B(6), B(1)
                           => B(5), B(0) => B(4), Ci => Cin(1), S(3) => S(7), 
                           S(2) => S(6), S(1) => S(5), S(0) => S(4), Co => 
                           net3151);
   csel_N_2 : carry_sel_gen_N4_6 port map( A(3) => A(11), A(2) => A(10), A(1) 
                           => A(9), A(0) => A(8), B(3) => B(11), B(2) => B(10),
                           B(1) => B(9), B(0) => B(8), Ci => Cin(2), S(3) => 
                           S(11), S(2) => S(10), S(1) => S(9), S(0) => S(8), Co
                           => net3150);
   csel_N_3 : carry_sel_gen_N4_5 port map( A(3) => A(15), A(2) => A(14), A(1) 
                           => A(13), A(0) => A(12), B(3) => B(15), B(2) => 
                           B(14), B(1) => B(13), B(0) => B(12), Ci => Cin(3), 
                           S(3) => S(15), S(2) => S(14), S(1) => S(13), S(0) =>
                           S(12), Co => net3149);
   csel_N_4 : carry_sel_gen_N4_4 port map( A(3) => A(19), A(2) => A(18), A(1) 
                           => A(17), A(0) => A(16), B(3) => B(19), B(2) => 
                           B(18), B(1) => B(17), B(0) => B(16), Ci => Cin(4), 
                           S(3) => S(19), S(2) => S(18), S(1) => S(17), S(0) =>
                           S(16), Co => net3148);
   csel_N_5 : carry_sel_gen_N4_3 port map( A(3) => A(23), A(2) => A(22), A(1) 
                           => A(21), A(0) => A(20), B(3) => B(23), B(2) => 
                           B(22), B(1) => B(21), B(0) => B(20), Ci => Cin(5), 
                           S(3) => S(23), S(2) => S(22), S(1) => S(21), S(0) =>
                           S(20), Co => net3147);
   csel_N_6 : carry_sel_gen_N4_2 port map( A(3) => A(27), A(2) => A(26), A(1) 
                           => A(25), A(0) => A(24), B(3) => B(27), B(2) => 
                           B(26), B(1) => B(25), B(0) => B(24), Ci => Cin(6), 
                           S(3) => S(27), S(2) => S(26), S(1) => S(25), S(0) =>
                           S(24), Co => net3146);
   csel_N_7 : carry_sel_gen_N4_1 port map( A(3) => A(31), A(2) => A(30), A(1) 
                           => A(29), A(0) => A(28), B(3) => B(31), B(2) => 
                           B(30), B(1) => B(29), B(0) => B(28), Ci => Cin(7), 
                           S(3) => S(31), S(2) => S(30), S(1) => S(29), S(0) =>
                           S(28), Co => net3145);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity carry_tree_N32_logN5_1 is

   port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  
         Cout_7_BAR, Cout_6_port, Cout_5_port, Cout_4_port, Cout_3_port, 
         Cout_2_port, Cout_1_port, Cout_0_port : out std_logic);

end carry_tree_N32_logN5_1;

architecture SYN_arch of carry_tree_N32_logN5_1 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component pg_1
      port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic
            );
   end component;
   
   component pg_2
      port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic
            );
   end component;
   
   component pg_3
      port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic
            );
   end component;
   
   component pg_4
      port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic
            );
   end component;
   
   component pg_5
      port( p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic;  
            g_BAR : in std_logic);
   end component;
   
   component g_1
      port( g, p, g_prec : in std_logic;  g_out_BAR : out std_logic);
   end component;
   
   component g_2
      port( g, p, g_prec : in std_logic;  g_out : out std_logic);
   end component;
   
   component g_3
      port( g, p, g_prec : in std_logic;  g_out : out std_logic);
   end component;
   
   component g_4
      port( g, p, g_prec : in std_logic;  g_out : out std_logic);
   end component;
   
   component g_5
      port( g, p, g_prec : in std_logic;  g_out : out std_logic);
   end component;
   
   component g_6
      port( g, p, g_prec : in std_logic;  g_out : out std_logic);
   end component;
   
   component g_7
      port( g, p, g_prec : in std_logic;  g_out : out std_logic);
   end component;
   
   component pg_6
      port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic
            );
   end component;
   
   component pg_7
      port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic
            );
   end component;
   
   component pg_8
      port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic
            );
   end component;
   
   component pg_9
      port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic
            );
   end component;
   
   component pg_10
      port( g, p, g_prec, p_prec : in std_logic;  p_out, g_out_BAR : out 
            std_logic);
   end component;
   
   component pg_11
      port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic
            );
   end component;
   
   component pg_12
      port( p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic;  
            g_BAR : in std_logic);
   end component;
   
   component g_8
      port( g, p, g_prec : in std_logic;  g_out : out std_logic);
   end component;
   
   component pg_13
      port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic
            );
   end component;
   
   component pg_14
      port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic
            );
   end component;
   
   component pg_15
      port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic
            );
   end component;
   
   component pg_16
      port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic
            );
   end component;
   
   component pg_17
      port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic
            );
   end component;
   
   component pg_18
      port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic
            );
   end component;
   
   component pg_19
      port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic
            );
   end component;
   
   component pg_20
      port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic
            );
   end component;
   
   component pg_21
      port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic
            );
   end component;
   
   component pg_22
      port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic
            );
   end component;
   
   component pg_23
      port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic
            );
   end component;
   
   component pg_24
      port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic
            );
   end component;
   
   component pg_25
      port( g, p, g_prec, p_prec : in std_logic;  p_out, g_out_BAR : out 
            std_logic);
   end component;
   
   component pg_26
      port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic
            );
   end component;
   
   component pg_27
      port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic
            );
   end component;
   
   component g_9
      port( g, p, g_prec : in std_logic;  g_out : out std_logic);
   end component;
   
   component g_10
      port( g, p, g_prec : in std_logic;  g_out : out std_logic);
   end component;
   
   component pg_net_1
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_2
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_3
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_4
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_5
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_6
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_7
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_8
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_9
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_10
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_11
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_12
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_13
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_14
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_15
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_16
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_17
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_18
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_19
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_20
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_21
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_22
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_23
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_24
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_25
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_26
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_27
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_28
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_29
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_30
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_31
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_32
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   signal n7, n8, Cout_0_port2, p_net_31_port, p_net_30_port, p_net_29_port, 
      p_net_28_port, p_net_27_port, p_net_26_port, p_net_25_port, p_net_24_port
      , p_net_23_port, p_net_22_port, p_net_20_port, p_net_19_port, 
      p_net_18_port, p_net_17_port, p_net_16_port, p_net_15_port, p_net_14_port
      , p_net_13_port, p_net_12_port, p_net_11_port, p_net_10_port, 
      p_net_9_port, p_net_8_port, p_net_7_port, p_net_6_port, p_net_5_port, 
      p_net_4_port, p_net_3_port, p_net_2_port, p_net_1_port, g_net_31_port, 
      g_net_30_port, g_net_29_port, g_net_28_port, g_net_27_port, g_net_26_port
      , g_net_25_port, g_net_24_port, g_net_23_port, g_net_22_port, 
      g_net_21_port, g_net_20_port, g_net_19_port, g_net_18_port, g_net_17_port
      , g_net_16_port, g_net_15_port, g_net_14_port, g_net_13_port, 
      g_net_12_port, g_net_11_port, g_net_10_port, g_net_9_port, g_net_8_port, 
      g_net_7_port, g_net_6_port, g_net_5_port, g_net_4_port, g_net_3_port, 
      g_net_2_port, g_net_1_port, g_net_0_port, magic_pro_1_port, 
      magic_pro_0_port, pg_1_15_1_port, pg_1_15_0_port, pg_1_14_1_port, 
      pg_1_14_0_port, pg_1_13_1_port, pg_1_13_0_port, pg_1_12_1_port, 
      pg_1_12_0_port, pg_1_11_1_port, pg_1_11_0_port, pg_1_10_1_port, 
      pg_1_10_0_port, pg_1_9_1_port, pg_1_9_0_port, pg_1_8_1_port, 
      pg_1_8_0_port, pg_1_7_1_port, pg_1_7_0_port, pg_1_6_1_port, pg_1_6_0_port
      , pg_1_5_1_port, pg_1_5_0_port, pg_1_4_1_port, pg_1_4_0_port, 
      pg_1_3_1_port, pg_1_3_0_port, pg_1_2_1_port, pg_1_2_0_port, pg_1_1_1_port
      , pg_1_1_0_port, pg_1_0_0_port, pg_n_4_7_1_port, pg_n_4_7_0_port, 
      pg_n_4_6_1_port, pg_n_4_6_0_port, pg_n_3_7_1_port, pg_n_3_7_0_port, 
      pg_n_3_5_1_port, pg_n_3_5_0_port, pg_n_3_3_1_port, pg_n_3_3_0_port, 
      pg_n_2_7_1_port, pg_n_2_7_0_port, pg_n_2_6_1_port, pg_n_2_6_0_port, 
      pg_n_2_5_1_port, pg_n_2_5_0_port, pg_n_2_4_1_port, pg_n_2_4_0_port, 
      pg_n_2_3_1_port, pg_n_2_3_0_port, pg_n_2_2_1_port, pg_n_2_2_0_port, 
      pg_n_2_1_1_port, pg_n_2_1_0_port, n1, n4, Cout_1_port2, Cout_3_port2 : 
      std_logic;

begin
   Cout_3_port <= Cout_3_port2;
   Cout_1_port <= Cout_1_port2;
   Cout_0_port <= Cout_0_port2;
   
   pg_net_x_1 : pg_net_32 port map( a => A(1), b => B(1), g_out => g_net_1_port
                           , p_out => p_net_1_port);
   pg_net_x_2 : pg_net_31 port map( a => A(2), b => B(2), g_out => g_net_2_port
                           , p_out => p_net_2_port);
   pg_net_x_3 : pg_net_30 port map( a => A(3), b => B(3), g_out => g_net_3_port
                           , p_out => p_net_3_port);
   pg_net_x_4 : pg_net_29 port map( a => A(4), b => B(4), g_out => g_net_4_port
                           , p_out => p_net_4_port);
   pg_net_x_5 : pg_net_28 port map( a => A(5), b => B(5), g_out => g_net_5_port
                           , p_out => p_net_5_port);
   pg_net_x_6 : pg_net_27 port map( a => A(6), b => B(6), g_out => g_net_6_port
                           , p_out => p_net_6_port);
   pg_net_x_7 : pg_net_26 port map( a => A(7), b => B(7), g_out => g_net_7_port
                           , p_out => p_net_7_port);
   pg_net_x_8 : pg_net_25 port map( a => A(8), b => B(8), g_out => g_net_8_port
                           , p_out => p_net_8_port);
   pg_net_x_9 : pg_net_24 port map( a => A(9), b => B(9), g_out => g_net_9_port
                           , p_out => p_net_9_port);
   pg_net_x_10 : pg_net_23 port map( a => A(10), b => B(10), g_out => 
                           g_net_10_port, p_out => p_net_10_port);
   pg_net_x_11 : pg_net_22 port map( a => A(11), b => B(11), g_out => 
                           g_net_11_port, p_out => p_net_11_port);
   pg_net_x_12 : pg_net_21 port map( a => A(12), b => B(12), g_out => 
                           g_net_12_port, p_out => p_net_12_port);
   pg_net_x_13 : pg_net_20 port map( a => A(13), b => B(13), g_out => 
                           g_net_13_port, p_out => p_net_13_port);
   pg_net_x_14 : pg_net_19 port map( a => A(14), b => B(14), g_out => 
                           g_net_14_port, p_out => p_net_14_port);
   pg_net_x_15 : pg_net_18 port map( a => A(15), b => B(15), g_out => 
                           g_net_15_port, p_out => p_net_15_port);
   pg_net_x_16 : pg_net_17 port map( a => A(16), b => B(16), g_out => 
                           g_net_16_port, p_out => p_net_16_port);
   pg_net_x_17 : pg_net_16 port map( a => A(17), b => B(17), g_out => 
                           g_net_17_port, p_out => p_net_17_port);
   pg_net_x_18 : pg_net_15 port map( a => A(18), b => B(18), g_out => 
                           g_net_18_port, p_out => p_net_18_port);
   pg_net_x_19 : pg_net_14 port map( a => A(19), b => B(19), g_out => 
                           g_net_19_port, p_out => p_net_19_port);
   pg_net_x_20 : pg_net_13 port map( a => A(20), b => B(20), g_out => 
                           g_net_20_port, p_out => p_net_20_port);
   pg_net_x_21 : pg_net_12 port map( a => A(21), b => B(21), g_out => 
                           g_net_21_port, p_out => n1);
   pg_net_x_22 : pg_net_11 port map( a => A(22), b => B(22), g_out => 
                           g_net_22_port, p_out => p_net_22_port);
   pg_net_x_23 : pg_net_10 port map( a => A(23), b => B(23), g_out => 
                           g_net_23_port, p_out => p_net_23_port);
   pg_net_x_24 : pg_net_9 port map( a => A(24), b => B(24), g_out => 
                           g_net_24_port, p_out => p_net_24_port);
   pg_net_x_25 : pg_net_8 port map( a => A(25), b => B(25), g_out => 
                           g_net_25_port, p_out => p_net_25_port);
   pg_net_x_26 : pg_net_7 port map( a => A(26), b => B(26), g_out => 
                           g_net_26_port, p_out => p_net_26_port);
   pg_net_x_27 : pg_net_6 port map( a => A(27), b => B(27), g_out => 
                           g_net_27_port, p_out => p_net_27_port);
   pg_net_x_28 : pg_net_5 port map( a => A(28), b => B(28), g_out => 
                           g_net_28_port, p_out => p_net_28_port);
   pg_net_x_29 : pg_net_4 port map( a => A(29), b => B(29), g_out => 
                           g_net_29_port, p_out => p_net_29_port);
   pg_net_x_30 : pg_net_3 port map( a => A(30), b => B(30), g_out => 
                           g_net_30_port, p_out => p_net_30_port);
   pg_net_x_31 : pg_net_2 port map( a => A(31), b => B(31), g_out => 
                           g_net_31_port, p_out => p_net_31_port);
   pg_net_0_MAGIC : pg_net_1 port map( a => A(0), b => B(0), g_out => 
                           magic_pro_0_port, p_out => magic_pro_1_port);
   xG_0_0_MAGIC : g_10 port map( g => magic_pro_0_port, p => magic_pro_1_port, 
                           g_prec => Cin, g_out => g_net_0_port);
   xG_1_0 : g_9 port map( g => g_net_1_port, p => p_net_1_port, g_prec => 
                           g_net_0_port, g_out => pg_1_0_0_port);
   xPG_1_1 : pg_27 port map( g => g_net_3_port, p => p_net_3_port, g_prec => 
                           g_net_2_port, p_prec => p_net_2_port, g_out => 
                           pg_1_1_0_port, p_out => pg_1_1_1_port);
   xPG_1_2 : pg_26 port map( g => g_net_5_port, p => p_net_5_port, g_prec => 
                           g_net_4_port, p_prec => p_net_4_port, g_out => 
                           pg_1_2_0_port, p_out => pg_1_2_1_port);
   xPG_1_3 : pg_25 port map( g => g_net_7_port, p => p_net_7_port, g_prec => 
                           g_net_6_port, p_prec => p_net_6_port, p_out => 
                           pg_1_3_1_port, g_out_BAR => pg_1_3_0_port);
   xPG_1_4 : pg_24 port map( g => g_net_9_port, p => p_net_9_port, g_prec => 
                           g_net_8_port, p_prec => p_net_8_port, g_out => 
                           pg_1_4_0_port, p_out => pg_1_4_1_port);
   xPG_1_5 : pg_23 port map( g => g_net_11_port, p => p_net_11_port, g_prec => 
                           g_net_10_port, p_prec => p_net_10_port, g_out => 
                           pg_1_5_0_port, p_out => pg_1_5_1_port);
   xPG_1_6 : pg_22 port map( g => g_net_13_port, p => p_net_13_port, g_prec => 
                           g_net_12_port, p_prec => p_net_12_port, g_out => 
                           pg_1_6_0_port, p_out => pg_1_6_1_port);
   xPG_1_7 : pg_21 port map( g => g_net_15_port, p => p_net_15_port, g_prec => 
                           g_net_14_port, p_prec => p_net_14_port, g_out => 
                           pg_1_7_0_port, p_out => pg_1_7_1_port);
   xPG_1_8 : pg_20 port map( g => g_net_17_port, p => p_net_17_port, g_prec => 
                           g_net_16_port, p_prec => p_net_16_port, g_out => 
                           pg_1_8_0_port, p_out => pg_1_8_1_port);
   xPG_1_9 : pg_19 port map( g => g_net_19_port, p => p_net_19_port, g_prec => 
                           g_net_18_port, p_prec => p_net_18_port, g_out => 
                           pg_1_9_0_port, p_out => pg_1_9_1_port);
   xPG_1_10 : pg_18 port map( g => g_net_21_port, p => n1, g_prec => 
                           g_net_20_port, p_prec => p_net_20_port, g_out => 
                           pg_1_10_0_port, p_out => pg_1_10_1_port);
   xPG_1_11 : pg_17 port map( g => g_net_23_port, p => p_net_23_port, g_prec =>
                           g_net_22_port, p_prec => p_net_22_port, g_out => 
                           pg_1_11_0_port, p_out => pg_1_11_1_port);
   xPG_1_12 : pg_16 port map( g => g_net_25_port, p => p_net_25_port, g_prec =>
                           g_net_24_port, p_prec => p_net_24_port, g_out => 
                           pg_1_12_0_port, p_out => pg_1_12_1_port);
   xPG_1_13 : pg_15 port map( g => g_net_27_port, p => p_net_27_port, g_prec =>
                           g_net_26_port, p_prec => p_net_26_port, g_out => 
                           pg_1_13_0_port, p_out => pg_1_13_1_port);
   xPG_1_14 : pg_14 port map( g => g_net_29_port, p => p_net_29_port, g_prec =>
                           g_net_28_port, p_prec => p_net_28_port, g_out => 
                           pg_1_14_0_port, p_out => pg_1_14_1_port);
   xPG_1_15 : pg_13 port map( g => g_net_31_port, p => p_net_31_port, g_prec =>
                           g_net_30_port, p_prec => p_net_30_port, g_out => 
                           pg_1_15_0_port, p_out => pg_1_15_1_port);
   xG_2_0 : g_8 port map( g => pg_1_1_0_port, p => pg_1_1_1_port, g_prec => 
                           pg_1_0_0_port, g_out => Cout_0_port2);
   xPG_2_1 : pg_12 port map( p => pg_1_3_1_port, g_prec => pg_1_2_0_port, 
                           p_prec => pg_1_2_1_port, g_out => pg_n_2_1_0_port, 
                           p_out => pg_n_2_1_1_port, g_BAR => pg_1_3_0_port);
   xPG_2_2 : pg_11 port map( g => pg_1_5_0_port, p => pg_1_5_1_port, g_prec => 
                           pg_1_4_0_port, p_prec => pg_1_4_1_port, g_out => 
                           pg_n_2_2_0_port, p_out => pg_n_2_2_1_port);
   xPG_2_3 : pg_10 port map( g => pg_1_7_0_port, p => pg_1_7_1_port, g_prec => 
                           pg_1_6_0_port, p_prec => pg_1_6_1_port, p_out => 
                           pg_n_2_3_1_port, g_out_BAR => pg_n_2_3_0_port);
   xPG_2_4 : pg_9 port map( g => pg_1_9_0_port, p => pg_1_9_1_port, g_prec => 
                           pg_1_8_0_port, p_prec => pg_1_8_1_port, g_out => 
                           pg_n_2_4_0_port, p_out => pg_n_2_4_1_port);
   xPG_2_5 : pg_8 port map( g => pg_1_11_0_port, p => pg_1_11_1_port, g_prec =>
                           pg_1_10_0_port, p_prec => pg_1_10_1_port, g_out => 
                           pg_n_2_5_0_port, p_out => pg_n_2_5_1_port);
   xPG_2_6 : pg_7 port map( g => pg_1_13_0_port, p => pg_1_13_1_port, g_prec =>
                           pg_1_12_0_port, p_prec => pg_1_12_1_port, g_out => 
                           pg_n_2_6_0_port, p_out => pg_n_2_6_1_port);
   xPG_2_7 : pg_6 port map( g => pg_1_15_0_port, p => pg_1_15_1_port, g_prec =>
                           pg_1_14_0_port, p_prec => pg_1_14_1_port, g_out => 
                           pg_n_2_7_0_port, p_out => pg_n_2_7_1_port);
   xG_3_1 : g_7 port map( g => pg_n_2_1_0_port, p => pg_n_2_1_1_port, g_prec =>
                           Cout_0_port2, g_out => n8);
   xG_4_2 : g_6 port map( g => pg_n_2_2_0_port, p => pg_n_2_2_1_port, g_prec =>
                           Cout_1_port2, g_out => Cout_2_port);
   xG_4_3 : g_5 port map( g => pg_n_3_3_0_port, p => pg_n_3_3_1_port, g_prec =>
                           n8, g_out => n7);
   xG_5_4 : g_4 port map( g => pg_n_2_4_0_port, p => pg_n_2_4_1_port, g_prec =>
                           n7, g_out => Cout_4_port);
   xG_5_5 : g_3 port map( g => n4, p => pg_n_3_5_1_port, g_prec => n7, g_out =>
                           Cout_5_port);
   xG_5_6 : g_2 port map( g => pg_n_4_6_0_port, p => pg_n_4_6_1_port, g_prec =>
                           n7, g_out => Cout_6_port);
   xG_5_7 : g_1 port map( g => pg_n_4_7_0_port, p => pg_n_4_7_1_port, g_prec =>
                           Cout_3_port2, g_out_BAR => Cout_7_BAR);
   xPG_3_3 : pg_5 port map( p => pg_n_2_3_1_port, g_prec => pg_n_2_2_0_port, 
                           p_prec => pg_n_2_2_1_port, g_out => pg_n_3_3_0_port,
                           p_out => pg_n_3_3_1_port, g_BAR => pg_n_2_3_0_port);
   xPG_3_5 : pg_4 port map( g => pg_n_2_5_0_port, p => pg_n_2_5_1_port, g_prec 
                           => pg_n_2_4_0_port, p_prec => pg_n_2_4_1_port, g_out
                           => pg_n_3_5_0_port, p_out => pg_n_3_5_1_port);
   xPG_3_7 : pg_3 port map( g => pg_n_2_7_0_port, p => pg_n_2_7_1_port, g_prec 
                           => pg_n_2_6_0_port, p_prec => pg_n_2_6_1_port, g_out
                           => pg_n_3_7_0_port, p_out => pg_n_3_7_1_port);
   xPG_4_6 : pg_2 port map( g => pg_n_2_6_0_port, p => pg_n_2_6_1_port, g_prec 
                           => pg_n_3_5_0_port, p_prec => pg_n_3_5_1_port, g_out
                           => pg_n_4_6_0_port, p_out => pg_n_4_6_1_port);
   xPG_4_7 : pg_1 port map( g => pg_n_3_7_0_port, p => pg_n_3_7_1_port, g_prec 
                           => n4, p_prec => pg_n_3_5_1_port, g_out => 
                           pg_n_4_7_0_port, p_out => pg_n_4_7_1_port);
   U1 : CLKBUF_X2 port map( A => n8, Z => Cout_1_port2);
   U2 : BUF_X1 port map( A => n7, Z => Cout_3_port2);
   U3 : CLKBUF_X1 port map( A => pg_n_3_5_0_port, Z => n4);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity xor_gen_N32_1 is

   port( A : in std_logic_vector (31 downto 0);  B : in std_logic;  S : out 
         std_logic_vector (31 downto 0));

end xor_gen_N32_1;

architecture SYN_bhe of xor_gen_N32_1 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X2
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n4, n5 : std_logic;

begin
   
   U8 : XOR2_X1 port map( A => B, B => A(31), Z => S(31));
   U9 : XOR2_X1 port map( A => B, B => A(30), Z => S(30));
   U11 : XOR2_X1 port map( A => B, B => A(29), Z => S(29));
   U13 : XOR2_X1 port map( A => B, B => A(27), Z => S(27));
   U14 : XOR2_X1 port map( A => B, B => A(26), Z => S(26));
   U16 : XOR2_X1 port map( A => B, B => A(24), Z => S(24));
   U20 : XOR2_X1 port map( A => B, B => A(20), Z => S(20));
   U22 : XOR2_X1 port map( A => B, B => A(19), Z => S(19));
   U25 : XOR2_X1 port map( A => B, B => A(16), Z => S(16));
   U26 : XOR2_X1 port map( A => B, B => A(15), Z => S(15));
   U30 : XOR2_X1 port map( A => B, B => A(11), Z => S(11));
   U32 : XOR2_X1 port map( A => B, B => A(0), Z => S(0));
   U1 : MUX2_X1 port map( A => B, B => n2, S => A(23), Z => S(23));
   U2 : XOR2_X1 port map( A => B, B => A(5), Z => S(5));
   U3 : MUX2_X1 port map( A => B, B => n2, S => A(10), Z => S(10));
   U4 : MUX2_X1 port map( A => B, B => n2, S => A(6), Z => S(6));
   U5 : XNOR2_X1 port map( A => A(3), B => n2, ZN => S(3));
   U6 : XOR2_X1 port map( A => B, B => A(13), Z => S(13));
   U7 : MUX2_X1 port map( A => B, B => n2, S => A(7), Z => S(7));
   U10 : XOR2_X2 port map( A => A(2), B => B, Z => S(2));
   U12 : XOR2_X2 port map( A => A(1), B => B, Z => S(1));
   U15 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => S(21));
   U17 : INV_X1 port map( A => A(21), ZN => n3);
   U18 : XOR2_X1 port map( A => A(8), B => B, Z => S(8));
   U19 : XOR2_X1 port map( A => B, B => A(4), Z => S(4));
   U21 : INV_X1 port map( A => B, ZN => n2);
   U23 : XOR2_X1 port map( A => B, B => A(12), Z => S(12));
   U24 : XOR2_X1 port map( A => B, B => A(18), Z => S(18));
   U27 : XOR2_X1 port map( A => B, B => A(25), Z => S(25));
   U28 : XOR2_X1 port map( A => B, B => A(28), Z => S(28));
   U29 : XOR2_X1 port map( A => B, B => A(22), Z => S(22));
   U31 : XOR2_X1 port map( A => B, B => A(17), Z => S(17));
   U33 : XOR2_X1 port map( A => B, B => A(14), Z => S(14));
   U34 : XOR2_X1 port map( A => B, B => A(9), Z => S(9));
   U35 : NAND2_X1 port map( A1 => B, A2 => n3, ZN => n4);
   U36 : NAND2_X1 port map( A1 => n2, A2 => A(21), ZN => n5);

end SYN_bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity ff32_en_SIZE5_3 is

   port( D : in std_logic_vector (4 downto 0);  en, clk, rst : in std_logic;  Q
         : out std_logic_vector (4 downto 0));

end ff32_en_SIZE5_3;

architecture SYN_behavioral of ff32_en_SIZE5_3 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_ff32_en_SIZE5_3
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   signal net3361, n1, n4, n5, n7, n8, n9 : std_logic;

begin
   
   Q_reg_4_inst : DFFR_X1 port map( D => D(4), CK => net3361, RN => n5, Q => 
                           Q(4), QN => n7);
   Q_reg_2_inst : DFFR_X1 port map( D => D(2), CK => net3361, RN => n5, Q => 
                           Q(2), QN => n8);
   Q_reg_1_inst : DFFR_X1 port map( D => D(1), CK => net3361, RN => n5, Q => 
                           Q(1), QN => n9);
   clk_gate_Q_reg : SNPS_CLOCK_GATE_HIGH_ff32_en_SIZE5_3 port map( CLK => clk, 
                           EN => en, ENCLK => net3361);
   Q_reg_3_inst : DFFR_X1 port map( D => D(3), CK => net3361, RN => n5, Q => 
                           Q(3), QN => n4);
   Q_reg_0_inst : DFFR_X1 port map( D => D(0), CK => net3361, RN => n5, Q => 
                           Q(0), QN => n1);
   U2 : INV_X1 port map( A => rst, ZN => n5);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity ff32_en_SIZE5_2 is

   port( D : in std_logic_vector (4 downto 0);  en, clk, rst : in std_logic;  Q
         : out std_logic_vector (4 downto 0));

end ff32_en_SIZE5_2;

architecture SYN_behavioral of ff32_en_SIZE5_2 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_ff32_en_SIZE5_2
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal net3361, n5, n7, n8, n9, n10, n11 : std_logic;

begin
   
   Q_reg_4_inst : DFFR_X1 port map( D => D(4), CK => net3361, RN => n5, Q => 
                           Q(4), QN => n7);
   Q_reg_3_inst : DFFR_X1 port map( D => D(3), CK => net3361, RN => n5, Q => 
                           Q(3), QN => n8);
   Q_reg_2_inst : DFFR_X1 port map( D => D(2), CK => net3361, RN => n5, Q => 
                           Q(2), QN => n9);
   Q_reg_1_inst : DFFR_X1 port map( D => D(1), CK => net3361, RN => n5, Q => 
                           Q(1), QN => n10);
   Q_reg_0_inst : DFFR_X1 port map( D => D(0), CK => net3361, RN => n5, Q => 
                           Q(0), QN => n11);
   clk_gate_Q_reg : SNPS_CLOCK_GATE_HIGH_ff32_en_SIZE5_2 port map( CLK => clk, 
                           EN => en, ENCLK => net3361);
   U2 : INV_X1 port map( A => rst, ZN => n5);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity ff32_en_SIZE5_1 is

   port( D : in std_logic_vector (4 downto 0);  en, clk, rst : in std_logic;  Q
         : out std_logic_vector (4 downto 0));

end ff32_en_SIZE5_1;

architecture SYN_behavioral of ff32_en_SIZE5_1 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6, n7, net48733 : std_logic;

begin
   
   Q_reg_3_inst : DFFR_X1 port map( D => D(3), CK => clk, RN => n6, Q => Q(3), 
                           QN => n7);
   Q_reg_1_inst : DFFR_X1 port map( D => D(1), CK => clk, RN => n6, Q => Q(1), 
                           QN => n5);
   Q_reg_2_inst : DFFR_X1 port map( D => D(2), CK => clk, RN => n6, Q => Q(2), 
                           QN => net48733);
   Q_reg_0_inst : DFFR_X1 port map( D => D(0), CK => clk, RN => n6, Q => Q(0), 
                           QN => n2);
   Q_reg_4_inst : DFFR_X1 port map( D => D(4), CK => clk, RN => n6, Q => Q(4), 
                           QN => n1);
   U2 : INV_X1 port map( A => rst, ZN => n6);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity ff32_en_SIZE32_5 is

   port( D : in std_logic_vector (31 downto 0);  en, clk, rst : in std_logic;  
         Q : out std_logic_vector (31 downto 0));

end ff32_en_SIZE32_5;

architecture SYN_behavioral of ff32_en_SIZE32_5 is

   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_ff32_en_SIZE32_5
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal net3346, n32, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, 
      n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59
      , n60, n61, n62, n63, n64, n65 : std_logic;

begin
   
   Q_reg_31_inst : DFFR_X1 port map( D => D(31), CK => net3346, RN => n32, Q =>
                           Q(31), QN => n34);
   Q_reg_30_inst : DFFR_X1 port map( D => D(30), CK => net3346, RN => n32, Q =>
                           Q(30), QN => n35);
   Q_reg_29_inst : DFFR_X1 port map( D => D(29), CK => net3346, RN => n32, Q =>
                           Q(29), QN => n36);
   Q_reg_28_inst : DFFR_X1 port map( D => D(28), CK => net3346, RN => n32, Q =>
                           Q(28), QN => n37);
   Q_reg_27_inst : DFFR_X1 port map( D => D(27), CK => net3346, RN => n32, Q =>
                           Q(27), QN => n38);
   Q_reg_26_inst : DFFR_X1 port map( D => D(26), CK => net3346, RN => n32, Q =>
                           Q(26), QN => n39);
   Q_reg_25_inst : DFFR_X1 port map( D => D(25), CK => net3346, RN => n32, Q =>
                           Q(25), QN => n40);
   Q_reg_24_inst : DFFR_X1 port map( D => D(24), CK => net3346, RN => n32, Q =>
                           Q(24), QN => n41);
   Q_reg_23_inst : DFFR_X1 port map( D => D(23), CK => net3346, RN => n32, Q =>
                           Q(23), QN => n42);
   Q_reg_22_inst : DFFR_X1 port map( D => D(22), CK => net3346, RN => n32, Q =>
                           Q(22), QN => n43);
   Q_reg_21_inst : DFFR_X1 port map( D => D(21), CK => net3346, RN => n32, Q =>
                           Q(21), QN => n44);
   Q_reg_20_inst : DFFR_X1 port map( D => D(20), CK => net3346, RN => n32, Q =>
                           Q(20), QN => n45);
   Q_reg_19_inst : DFFR_X1 port map( D => D(19), CK => net3346, RN => n32, Q =>
                           Q(19), QN => n46);
   Q_reg_18_inst : DFFR_X1 port map( D => D(18), CK => net3346, RN => n32, Q =>
                           Q(18), QN => n47);
   Q_reg_17_inst : DFFR_X1 port map( D => D(17), CK => net3346, RN => n32, Q =>
                           Q(17), QN => n48);
   Q_reg_16_inst : DFFR_X1 port map( D => D(16), CK => net3346, RN => n32, Q =>
                           Q(16), QN => n49);
   Q_reg_15_inst : DFFR_X1 port map( D => D(15), CK => net3346, RN => n32, Q =>
                           Q(15), QN => n50);
   Q_reg_14_inst : DFFR_X1 port map( D => D(14), CK => net3346, RN => n32, Q =>
                           Q(14), QN => n51);
   Q_reg_13_inst : DFFR_X1 port map( D => D(13), CK => net3346, RN => n32, Q =>
                           Q(13), QN => n52);
   Q_reg_12_inst : DFFR_X1 port map( D => D(12), CK => net3346, RN => n32, Q =>
                           Q(12), QN => n53);
   Q_reg_11_inst : DFFR_X1 port map( D => D(11), CK => net3346, RN => n32, Q =>
                           Q(11), QN => n54);
   Q_reg_10_inst : DFFR_X1 port map( D => D(10), CK => net3346, RN => n32, Q =>
                           Q(10), QN => n55);
   Q_reg_9_inst : DFFR_X1 port map( D => D(9), CK => net3346, RN => n32, Q => 
                           Q(9), QN => n56);
   Q_reg_8_inst : DFFR_X1 port map( D => D(8), CK => net3346, RN => n32, Q => 
                           Q(8), QN => n57);
   Q_reg_7_inst : DFFR_X1 port map( D => D(7), CK => net3346, RN => n32, Q => 
                           Q(7), QN => n58);
   Q_reg_6_inst : DFFR_X1 port map( D => D(6), CK => net3346, RN => n32, Q => 
                           Q(6), QN => n59);
   Q_reg_5_inst : DFFR_X1 port map( D => D(5), CK => net3346, RN => n32, Q => 
                           Q(5), QN => n60);
   Q_reg_4_inst : DFFR_X1 port map( D => D(4), CK => net3346, RN => n32, Q => 
                           Q(4), QN => n61);
   Q_reg_3_inst : DFFR_X1 port map( D => D(3), CK => net3346, RN => n32, Q => 
                           Q(3), QN => n62);
   Q_reg_2_inst : DFFR_X1 port map( D => D(2), CK => net3346, RN => n32, Q => 
                           Q(2), QN => n63);
   Q_reg_1_inst : DFFR_X1 port map( D => D(1), CK => net3346, RN => n32, Q => 
                           Q(1), QN => n64);
   Q_reg_0_inst : DFFR_X1 port map( D => D(0), CK => net3346, RN => n32, Q => 
                           Q(0), QN => n65);
   clk_gate_Q_reg : SNPS_CLOCK_GATE_HIGH_ff32_en_SIZE32_5 port map( CLK => clk,
                           EN => en, ENCLK => net3346);
   U2 : INV_X2 port map( A => rst, ZN => n32);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity ff32_en_SIZE32_4 is

   port( D : in std_logic_vector (31 downto 0);  en, clk, rst : in std_logic;  
         Q : out std_logic_vector (31 downto 0));

end ff32_en_SIZE32_4;

architecture SYN_behavioral of ff32_en_SIZE32_4 is

   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_ff32_en_SIZE32_4
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal net3346, n32, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, 
      n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59
      , n60, n61, n62, n63, n64, n65 : std_logic;

begin
   
   Q_reg_31_inst : DFFR_X1 port map( D => D(31), CK => net3346, RN => n32, Q =>
                           Q(31), QN => n34);
   Q_reg_30_inst : DFFR_X1 port map( D => D(30), CK => net3346, RN => n32, Q =>
                           Q(30), QN => n35);
   Q_reg_29_inst : DFFR_X1 port map( D => D(29), CK => net3346, RN => n32, Q =>
                           Q(29), QN => n36);
   Q_reg_28_inst : DFFR_X1 port map( D => D(28), CK => net3346, RN => n32, Q =>
                           Q(28), QN => n37);
   Q_reg_27_inst : DFFR_X1 port map( D => D(27), CK => net3346, RN => n32, Q =>
                           Q(27), QN => n38);
   Q_reg_26_inst : DFFR_X1 port map( D => D(26), CK => net3346, RN => n32, Q =>
                           Q(26), QN => n39);
   Q_reg_25_inst : DFFR_X1 port map( D => D(25), CK => net3346, RN => n32, Q =>
                           Q(25), QN => n40);
   Q_reg_24_inst : DFFR_X1 port map( D => D(24), CK => net3346, RN => n32, Q =>
                           Q(24), QN => n41);
   Q_reg_23_inst : DFFR_X1 port map( D => D(23), CK => net3346, RN => n32, Q =>
                           Q(23), QN => n42);
   Q_reg_22_inst : DFFR_X1 port map( D => D(22), CK => net3346, RN => n32, Q =>
                           Q(22), QN => n43);
   Q_reg_21_inst : DFFR_X1 port map( D => D(21), CK => net3346, RN => n32, Q =>
                           Q(21), QN => n44);
   Q_reg_20_inst : DFFR_X1 port map( D => D(20), CK => net3346, RN => n32, Q =>
                           Q(20), QN => n45);
   Q_reg_19_inst : DFFR_X1 port map( D => D(19), CK => net3346, RN => n32, Q =>
                           Q(19), QN => n46);
   Q_reg_18_inst : DFFR_X1 port map( D => D(18), CK => net3346, RN => n32, Q =>
                           Q(18), QN => n47);
   Q_reg_17_inst : DFFR_X1 port map( D => D(17), CK => net3346, RN => n32, Q =>
                           Q(17), QN => n48);
   Q_reg_16_inst : DFFR_X1 port map( D => D(16), CK => net3346, RN => n32, Q =>
                           Q(16), QN => n49);
   Q_reg_15_inst : DFFR_X1 port map( D => D(15), CK => net3346, RN => n32, Q =>
                           Q(15), QN => n50);
   Q_reg_14_inst : DFFR_X1 port map( D => D(14), CK => net3346, RN => n32, Q =>
                           Q(14), QN => n51);
   Q_reg_13_inst : DFFR_X1 port map( D => D(13), CK => net3346, RN => n32, Q =>
                           Q(13), QN => n52);
   Q_reg_12_inst : DFFR_X1 port map( D => D(12), CK => net3346, RN => n32, Q =>
                           Q(12), QN => n53);
   Q_reg_11_inst : DFFR_X1 port map( D => D(11), CK => net3346, RN => n32, Q =>
                           Q(11), QN => n54);
   Q_reg_10_inst : DFFR_X1 port map( D => D(10), CK => net3346, RN => n32, Q =>
                           Q(10), QN => n55);
   Q_reg_9_inst : DFFR_X1 port map( D => D(9), CK => net3346, RN => n32, Q => 
                           Q(9), QN => n56);
   Q_reg_8_inst : DFFR_X1 port map( D => D(8), CK => net3346, RN => n32, Q => 
                           Q(8), QN => n57);
   Q_reg_7_inst : DFFR_X1 port map( D => D(7), CK => net3346, RN => n32, Q => 
                           Q(7), QN => n58);
   Q_reg_6_inst : DFFR_X1 port map( D => D(6), CK => net3346, RN => n32, Q => 
                           Q(6), QN => n59);
   Q_reg_5_inst : DFFR_X1 port map( D => D(5), CK => net3346, RN => n32, Q => 
                           Q(5), QN => n60);
   Q_reg_4_inst : DFFR_X1 port map( D => D(4), CK => net3346, RN => n32, Q => 
                           Q(4), QN => n61);
   Q_reg_3_inst : DFFR_X1 port map( D => D(3), CK => net3346, RN => n32, Q => 
                           Q(3), QN => n62);
   Q_reg_2_inst : DFFR_X1 port map( D => D(2), CK => net3346, RN => n32, Q => 
                           Q(2), QN => n63);
   Q_reg_1_inst : DFFR_X1 port map( D => D(1), CK => net3346, RN => n32, Q => 
                           Q(1), QN => n64);
   Q_reg_0_inst : DFFR_X1 port map( D => D(0), CK => net3346, RN => n32, Q => 
                           Q(0), QN => n65);
   clk_gate_Q_reg : SNPS_CLOCK_GATE_HIGH_ff32_en_SIZE32_4 port map( CLK => clk,
                           EN => en, ENCLK => net3346);
   U2 : INV_X2 port map( A => rst, ZN => n32);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity ff32_en_SIZE32_3 is

   port( D : in std_logic_vector (31 downto 0);  en, clk, rst : in std_logic;  
         Q : out std_logic_vector (31 downto 0));

end ff32_en_SIZE32_3;

architecture SYN_behavioral of ff32_en_SIZE32_3 is

   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n32, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, 
      n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60
      , n61, n62, n63, n64 : std_logic;

begin
   
   Q_reg_31_inst : DFFR_X1 port map( D => D(31), CK => clk, RN => n32, Q => 
                           Q(31), QN => n34);
   Q_reg_30_inst : DFFR_X1 port map( D => D(30), CK => clk, RN => n32, Q => 
                           Q(30), QN => n35);
   Q_reg_29_inst : DFFR_X1 port map( D => D(29), CK => clk, RN => n32, Q => 
                           Q(29), QN => n36);
   Q_reg_28_inst : DFFR_X1 port map( D => D(28), CK => clk, RN => n32, Q => 
                           Q(28), QN => n37);
   Q_reg_27_inst : DFFR_X1 port map( D => D(27), CK => clk, RN => n32, Q => 
                           Q(27), QN => n38);
   Q_reg_26_inst : DFFR_X1 port map( D => D(26), CK => clk, RN => n32, Q => 
                           Q(26), QN => n39);
   Q_reg_25_inst : DFFR_X1 port map( D => D(25), CK => clk, RN => n32, Q => 
                           Q(25), QN => n40);
   Q_reg_24_inst : DFFR_X1 port map( D => D(24), CK => clk, RN => n32, Q => 
                           Q(24), QN => n41);
   Q_reg_23_inst : DFFR_X1 port map( D => D(23), CK => clk, RN => n32, Q => 
                           Q(23), QN => n42);
   Q_reg_22_inst : DFFR_X1 port map( D => D(22), CK => clk, RN => n32, Q => 
                           Q(22), QN => n43);
   Q_reg_21_inst : DFFR_X1 port map( D => D(21), CK => clk, RN => n32, Q => 
                           Q(21), QN => n44);
   Q_reg_20_inst : DFFR_X1 port map( D => D(20), CK => clk, RN => n32, Q => 
                           Q(20), QN => n45);
   Q_reg_19_inst : DFFR_X1 port map( D => D(19), CK => clk, RN => n32, Q => 
                           Q(19), QN => n46);
   Q_reg_18_inst : DFFR_X1 port map( D => D(18), CK => clk, RN => n32, Q => 
                           Q(18), QN => n47);
   Q_reg_17_inst : DFFR_X1 port map( D => D(17), CK => clk, RN => n32, Q => 
                           Q(17), QN => n48);
   Q_reg_16_inst : DFFR_X1 port map( D => D(16), CK => clk, RN => n32, Q => 
                           Q(16), QN => n49);
   Q_reg_15_inst : DFFR_X1 port map( D => D(15), CK => clk, RN => n32, Q => 
                           Q(15), QN => n50);
   Q_reg_14_inst : DFFR_X1 port map( D => D(14), CK => clk, RN => n32, Q => 
                           Q(14), QN => n51);
   Q_reg_13_inst : DFFR_X1 port map( D => D(13), CK => clk, RN => n32, Q => 
                           Q(13), QN => n52);
   Q_reg_12_inst : DFFR_X1 port map( D => D(12), CK => clk, RN => n32, Q => 
                           Q(12), QN => n53);
   Q_reg_11_inst : DFFR_X1 port map( D => D(11), CK => clk, RN => n32, Q => 
                           Q(11), QN => n54);
   Q_reg_10_inst : DFFR_X1 port map( D => D(10), CK => clk, RN => n32, Q => 
                           Q(10), QN => n55);
   Q_reg_9_inst : DFFR_X1 port map( D => D(9), CK => clk, RN => n32, Q => Q(9),
                           QN => n56);
   Q_reg_8_inst : DFFR_X1 port map( D => D(8), CK => clk, RN => n32, Q => Q(8),
                           QN => n57);
   Q_reg_7_inst : DFFR_X1 port map( D => D(7), CK => clk, RN => n32, Q => Q(7),
                           QN => n58);
   Q_reg_6_inst : DFFR_X1 port map( D => D(6), CK => clk, RN => n32, Q => Q(6),
                           QN => n59);
   Q_reg_5_inst : DFFR_X1 port map( D => D(5), CK => clk, RN => n32, Q => Q(5),
                           QN => n60);
   Q_reg_4_inst : DFFR_X1 port map( D => D(4), CK => clk, RN => n32, Q => Q(4),
                           QN => n61);
   Q_reg_3_inst : DFFR_X1 port map( D => D(3), CK => clk, RN => n32, Q => Q(3),
                           QN => n62);
   Q_reg_2_inst : DFFR_X1 port map( D => D(2), CK => clk, RN => n32, Q => Q(2),
                           QN => n63);
   Q_reg_1_inst : DFFR_X1 port map( D => D(1), CK => clk, RN => n32, Q => Q(1),
                           QN => n64);
   Q_reg_0_inst : DFFR_X1 port map( D => D(0), CK => clk, RN => n32, Q => Q(0),
                           QN => n1);
   U2 : INV_X2 port map( A => rst, ZN => n32);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity ff32_en_SIZE32_2 is

   port( D : in std_logic_vector (31 downto 0);  en, clk, rst : in std_logic;  
         Q : out std_logic_vector (31 downto 0));

end ff32_en_SIZE32_2;

architecture SYN_behavioral of ff32_en_SIZE32_2 is

   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
      n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62
      , n63, n64, n65, n66 : std_logic;

begin
   
   Q_reg_31_inst : DFFR_X1 port map( D => D(31), CK => clk, RN => n34, Q => 
                           Q(31), QN => n35);
   Q_reg_30_inst : DFFR_X1 port map( D => D(30), CK => clk, RN => n34, Q => 
                           Q(30), QN => n36);
   Q_reg_29_inst : DFFR_X1 port map( D => D(29), CK => clk, RN => n34, Q => 
                           Q(29), QN => n37);
   Q_reg_28_inst : DFFR_X1 port map( D => D(28), CK => clk, RN => n34, Q => 
                           Q(28), QN => n38);
   Q_reg_27_inst : DFFR_X1 port map( D => D(27), CK => clk, RN => n34, Q => 
                           Q(27), QN => n39);
   Q_reg_26_inst : DFFR_X1 port map( D => D(26), CK => clk, RN => n34, Q => 
                           Q(26), QN => n40);
   Q_reg_25_inst : DFFR_X1 port map( D => D(25), CK => clk, RN => n34, Q => 
                           Q(25), QN => n41);
   Q_reg_24_inst : DFFR_X1 port map( D => D(24), CK => clk, RN => n34, Q => 
                           Q(24), QN => n42);
   Q_reg_23_inst : DFFR_X1 port map( D => D(23), CK => clk, RN => n34, Q => 
                           Q(23), QN => n43);
   Q_reg_22_inst : DFFR_X1 port map( D => D(22), CK => clk, RN => n34, Q => 
                           Q(22), QN => n44);
   Q_reg_21_inst : DFFR_X1 port map( D => D(21), CK => clk, RN => n34, Q => 
                           Q(21), QN => n45);
   Q_reg_20_inst : DFFR_X1 port map( D => D(20), CK => clk, RN => n34, Q => 
                           Q(20), QN => n46);
   Q_reg_19_inst : DFFR_X1 port map( D => D(19), CK => clk, RN => n34, Q => 
                           Q(19), QN => n47);
   Q_reg_18_inst : DFFR_X1 port map( D => D(18), CK => clk, RN => n34, Q => 
                           Q(18), QN => n48);
   Q_reg_17_inst : DFFR_X1 port map( D => D(17), CK => clk, RN => n34, Q => 
                           Q(17), QN => n49);
   Q_reg_16_inst : DFFR_X1 port map( D => D(16), CK => clk, RN => n34, Q => 
                           Q(16), QN => n50);
   Q_reg_15_inst : DFFR_X1 port map( D => D(15), CK => clk, RN => n34, Q => 
                           Q(15), QN => n51);
   Q_reg_14_inst : DFFR_X1 port map( D => D(14), CK => clk, RN => n34, Q => 
                           Q(14), QN => n52);
   Q_reg_13_inst : DFFR_X1 port map( D => D(13), CK => clk, RN => n34, Q => 
                           Q(13), QN => n53);
   Q_reg_12_inst : DFFR_X1 port map( D => D(12), CK => clk, RN => n34, Q => 
                           Q(12), QN => n54);
   Q_reg_11_inst : DFFR_X1 port map( D => D(11), CK => clk, RN => n34, Q => 
                           Q(11), QN => n55);
   Q_reg_10_inst : DFFR_X1 port map( D => D(10), CK => clk, RN => n34, Q => 
                           Q(10), QN => n56);
   Q_reg_9_inst : DFFR_X1 port map( D => D(9), CK => clk, RN => n34, Q => Q(9),
                           QN => n57);
   Q_reg_8_inst : DFFR_X1 port map( D => D(8), CK => clk, RN => n34, Q => Q(8),
                           QN => n58);
   Q_reg_7_inst : DFFR_X1 port map( D => D(7), CK => clk, RN => n34, Q => Q(7),
                           QN => n59);
   Q_reg_6_inst : DFFR_X1 port map( D => D(6), CK => clk, RN => n34, Q => Q(6),
                           QN => n60);
   Q_reg_5_inst : DFFR_X1 port map( D => D(5), CK => clk, RN => n34, Q => Q(5),
                           QN => n61);
   Q_reg_4_inst : DFFR_X1 port map( D => D(4), CK => clk, RN => n34, Q => Q(4),
                           QN => n62);
   Q_reg_3_inst : DFFR_X1 port map( D => D(3), CK => clk, RN => n34, Q => Q(3),
                           QN => n63);
   Q_reg_2_inst : DFFR_X1 port map( D => D(2), CK => clk, RN => n34, Q => Q(2),
                           QN => n64);
   Q_reg_1_inst : DFFR_X1 port map( D => D(1), CK => clk, RN => n34, Q => Q(1),
                           QN => n65);
   Q_reg_0_inst : DFFR_X1 port map( D => D(0), CK => clk, RN => n34, Q => Q(0),
                           QN => n66);
   U2 : INV_X2 port map( A => rst, ZN => n34);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity ff32_en_SIZE32_1 is

   port( D : in std_logic_vector (31 downto 0);  en, clk, rst : in std_logic;  
         Q : out std_logic_vector (31 downto 0));

end ff32_en_SIZE32_1;

architecture SYN_behavioral of ff32_en_SIZE32_1 is

   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_ff32_en_SIZE32_1
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal net3346, n32, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, 
      n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59
      , n60, n61, n62, n63, n64, n65 : std_logic;

begin
   
   Q_reg_31_inst : DFFR_X1 port map( D => D(31), CK => net3346, RN => n32, Q =>
                           Q(31), QN => n34);
   Q_reg_30_inst : DFFR_X1 port map( D => D(30), CK => net3346, RN => n32, Q =>
                           Q(30), QN => n35);
   Q_reg_29_inst : DFFR_X1 port map( D => D(29), CK => net3346, RN => n32, Q =>
                           Q(29), QN => n36);
   Q_reg_28_inst : DFFR_X1 port map( D => D(28), CK => net3346, RN => n32, Q =>
                           Q(28), QN => n37);
   Q_reg_27_inst : DFFR_X1 port map( D => D(27), CK => net3346, RN => n32, Q =>
                           Q(27), QN => n38);
   Q_reg_26_inst : DFFR_X1 port map( D => D(26), CK => net3346, RN => n32, Q =>
                           Q(26), QN => n39);
   Q_reg_25_inst : DFFR_X1 port map( D => D(25), CK => net3346, RN => n32, Q =>
                           Q(25), QN => n40);
   Q_reg_24_inst : DFFR_X1 port map( D => D(24), CK => net3346, RN => n32, Q =>
                           Q(24), QN => n41);
   Q_reg_23_inst : DFFR_X1 port map( D => D(23), CK => net3346, RN => n32, Q =>
                           Q(23), QN => n42);
   Q_reg_22_inst : DFFR_X1 port map( D => D(22), CK => net3346, RN => n32, Q =>
                           Q(22), QN => n43);
   Q_reg_21_inst : DFFR_X1 port map( D => D(21), CK => net3346, RN => n32, Q =>
                           Q(21), QN => n44);
   Q_reg_20_inst : DFFR_X1 port map( D => D(20), CK => net3346, RN => n32, Q =>
                           Q(20), QN => n45);
   Q_reg_19_inst : DFFR_X1 port map( D => D(19), CK => net3346, RN => n32, Q =>
                           Q(19), QN => n46);
   Q_reg_18_inst : DFFR_X1 port map( D => D(18), CK => net3346, RN => n32, Q =>
                           Q(18), QN => n47);
   Q_reg_17_inst : DFFR_X1 port map( D => D(17), CK => net3346, RN => n32, Q =>
                           Q(17), QN => n48);
   Q_reg_16_inst : DFFR_X1 port map( D => D(16), CK => net3346, RN => n32, Q =>
                           Q(16), QN => n49);
   Q_reg_15_inst : DFFR_X1 port map( D => D(15), CK => net3346, RN => n32, Q =>
                           Q(15), QN => n50);
   Q_reg_14_inst : DFFR_X1 port map( D => D(14), CK => net3346, RN => n32, Q =>
                           Q(14), QN => n51);
   Q_reg_13_inst : DFFR_X1 port map( D => D(13), CK => net3346, RN => n32, Q =>
                           Q(13), QN => n52);
   Q_reg_12_inst : DFFR_X1 port map( D => D(12), CK => net3346, RN => n32, Q =>
                           Q(12), QN => n53);
   Q_reg_11_inst : DFFR_X1 port map( D => D(11), CK => net3346, RN => n32, Q =>
                           Q(11), QN => n54);
   Q_reg_10_inst : DFFR_X1 port map( D => D(10), CK => net3346, RN => n32, Q =>
                           Q(10), QN => n55);
   Q_reg_9_inst : DFFR_X1 port map( D => D(9), CK => net3346, RN => n32, Q => 
                           Q(9), QN => n56);
   Q_reg_8_inst : DFFR_X1 port map( D => D(8), CK => net3346, RN => n32, Q => 
                           Q(8), QN => n57);
   Q_reg_7_inst : DFFR_X1 port map( D => D(7), CK => net3346, RN => n32, Q => 
                           Q(7), QN => n58);
   Q_reg_6_inst : DFFR_X1 port map( D => D(6), CK => net3346, RN => n32, Q => 
                           Q(6), QN => n59);
   Q_reg_5_inst : DFFR_X1 port map( D => D(5), CK => net3346, RN => n32, Q => 
                           Q(5), QN => n60);
   Q_reg_4_inst : DFFR_X1 port map( D => D(4), CK => net3346, RN => n32, Q => 
                           Q(4), QN => n61);
   Q_reg_3_inst : DFFR_X1 port map( D => D(3), CK => net3346, RN => n32, Q => 
                           Q(3), QN => n62);
   Q_reg_2_inst : DFFR_X1 port map( D => D(2), CK => net3346, RN => n32, Q => 
                           Q(2), QN => n63);
   Q_reg_1_inst : DFFR_X1 port map( D => D(1), CK => net3346, RN => n32, Q => 
                           Q(1), QN => n64);
   Q_reg_0_inst : DFFR_X1 port map( D => D(0), CK => net3346, RN => n32, Q => 
                           Q(0), QN => n65);
   clk_gate_Q_reg : SNPS_CLOCK_GATE_HIGH_ff32_en_SIZE32_1 port map( CLK => clk,
                           EN => en, ENCLK => net3346);
   U2 : INV_X2 port map( A => rst, ZN => n32);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity mux41_MUX_SIZE32_2 is

   port( IN0, IN1, IN2, IN3 : in std_logic_vector (31 downto 0);  CTRL : in 
         std_logic_vector (1 downto 0);  OUT1 : out std_logic_vector (31 downto
         0));

end mux41_MUX_SIZE32_2;

architecture SYN_bhe of mux41_MUX_SIZE32_2 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X4
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, 
      n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98
      , n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, 
      n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, 
      n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, 
      n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146 : 
      std_logic;

begin
   
   U87 : AOI22_X1 port map( A1 => n142, A2 => IN1(12), B1 => n73, B2 => IN0(12)
                           , ZN => n86);
   U63 : AOI22_X1 port map( A1 => n142, A2 => IN1(1), B1 => n73, B2 => IN0(1), 
                           ZN => n102);
   U98 : AOI22_X1 port map( A1 => n142, A2 => IN1(0), B1 => n73, B2 => IN0(0), 
                           ZN => n80);
   U21 : AOI22_X1 port map( A1 => n75, A2 => IN1(3), B1 => n72, B2 => IN0(3), 
                           ZN => n130);
   U30 : AOI22_X1 port map( A1 => n74, A2 => IN1(2), B1 => n72, B2 => IN0(2), 
                           ZN => n124);
   U12 : AOI22_X1 port map( A1 => n75, A2 => IN1(6), B1 => n72, B2 => IN0(6), 
                           ZN => n136);
   U11 : AOI22_X1 port map( A1 => n2, A2 => IN3(6), B1 => n1, B2 => IN2(6), ZN 
                           => n135);
   U9 : AOI22_X1 port map( A1 => n75, A2 => IN1(7), B1 => n72, B2 => IN0(7), ZN
                           => n138);
   U8 : AOI22_X1 port map( A1 => n2, A2 => IN3(7), B1 => n1, B2 => IN2(7), ZN 
                           => n137);
   U15 : AOI22_X1 port map( A1 => n75, A2 => IN1(5), B1 => n72, B2 => IN0(5), 
                           ZN => n134);
   U14 : AOI22_X1 port map( A1 => n2, A2 => IN3(5), B1 => n1, B2 => IN2(5), ZN 
                           => n133);
   U18 : AOI22_X1 port map( A1 => n75, A2 => IN1(4), B1 => n72, B2 => IN0(4), 
                           ZN => n132);
   U17 : AOI22_X1 port map( A1 => n2, A2 => IN3(4), B1 => n1, B2 => IN2(4), ZN 
                           => n131);
   U90 : AOI22_X1 port map( A1 => n75, A2 => IN1(11), B1 => n73, B2 => IN0(11),
                           ZN => n84);
   U93 : AOI22_X1 port map( A1 => n142, A2 => IN1(10), B1 => n73, B2 => IN0(10)
                           , ZN => n82);
   U3 : AOI22_X1 port map( A1 => n75, A2 => IN1(9), B1 => n72, B2 => IN0(9), ZN
                           => n146);
   U2 : AOI22_X1 port map( A1 => n2, A2 => IN3(9), B1 => n1, B2 => IN2(9), ZN 
                           => n145);
   U6 : AOI22_X1 port map( A1 => n75, A2 => IN1(8), B1 => n72, B2 => IN0(8), ZN
                           => n140);
   U5 : AOI22_X1 port map( A1 => n2, A2 => IN3(8), B1 => n1, B2 => IN2(8), ZN 
                           => n139);
   U81 : AOI22_X1 port map( A1 => n142, A2 => IN1(14), B1 => n73, B2 => IN0(14)
                           , ZN => n90);
   U84 : AOI22_X1 port map( A1 => n142, A2 => IN1(13), B1 => n73, B2 => IN0(13)
                           , ZN => n88);
   U78 : AOI22_X1 port map( A1 => n75, A2 => IN1(15), B1 => n73, B2 => IN0(15),
                           ZN => n92);
   U75 : AOI22_X1 port map( A1 => n142, A2 => IN1(16), B1 => n73, B2 => IN0(16)
                           , ZN => n94);
   U73 : NAND2_X1 port map( A1 => n94, A2 => n93, ZN => OUT1(16));
   U51 : AOI22_X1 port map( A1 => n74, A2 => IN1(23), B1 => n72, B2 => IN0(23),
                           ZN => n110);
   U49 : NAND2_X1 port map( A1 => n110, A2 => n109, ZN => OUT1(23));
   U60 : AOI22_X1 port map( A1 => n74, A2 => IN1(20), B1 => n72, B2 => IN0(20),
                           ZN => n104);
   U59 : AOI22_X1 port map( A1 => n2, A2 => IN3(20), B1 => n1, B2 => IN2(20), 
                           ZN => n103);
   U58 : NAND2_X1 port map( A1 => n104, A2 => n103, ZN => OUT1(20));
   U57 : AOI22_X1 port map( A1 => n74, A2 => IN1(21), B1 => n72, B2 => IN0(21),
                           ZN => n106);
   U55 : NAND2_X1 port map( A1 => n106, A2 => n105, ZN => OUT1(21));
   U54 : AOI22_X1 port map( A1 => n74, A2 => IN1(22), B1 => n72, B2 => IN0(22),
                           ZN => n108);
   U52 : NAND2_X1 port map( A1 => n108, A2 => n107, ZN => OUT1(22));
   U69 : AOI22_X1 port map( A1 => n142, A2 => IN1(18), B1 => n73, B2 => IN0(18)
                           , ZN => n98);
   U67 : NAND2_X1 port map( A1 => n98, A2 => n97, ZN => OUT1(18));
   U66 : AOI22_X1 port map( A1 => n142, A2 => IN1(19), B1 => n73, B2 => IN0(19)
                           , ZN => n100);
   U64 : NAND2_X1 port map( A1 => n100, A2 => n99, ZN => OUT1(19));
   U72 : AOI22_X1 port map( A1 => n75, A2 => IN1(17), B1 => n73, B2 => IN0(17),
                           ZN => n96);
   U70 : NAND2_X1 port map( A1 => n96, A2 => n95, ZN => OUT1(17));
   U24 : AOI22_X1 port map( A1 => n75, A2 => IN1(31), B1 => n72, B2 => IN0(31),
                           ZN => n128);
   U23 : AOI22_X1 port map( A1 => n2, A2 => IN3(31), B1 => n1, B2 => IN2(31), 
                           ZN => n127);
   U22 : NAND2_X1 port map( A1 => n128, A2 => n127, ZN => OUT1(31));
   U36 : AOI22_X1 port map( A1 => n74, A2 => IN1(28), B1 => n72, B2 => IN0(28),
                           ZN => n120);
   U35 : AOI22_X1 port map( A1 => n2, A2 => IN3(28), B1 => n1, B2 => IN2(28), 
                           ZN => n119);
   U34 : NAND2_X1 port map( A1 => n120, A2 => n119, ZN => OUT1(28));
   U33 : AOI22_X1 port map( A1 => n74, A2 => IN1(29), B1 => n72, B2 => IN0(29),
                           ZN => n122);
   U32 : AOI22_X1 port map( A1 => n2, A2 => IN3(29), B1 => n1, B2 => IN2(29), 
                           ZN => n121);
   U31 : NAND2_X1 port map( A1 => n122, A2 => n121, ZN => OUT1(29));
   U27 : AOI22_X1 port map( A1 => n74, A2 => IN1(30), B1 => n72, B2 => IN0(30),
                           ZN => n126);
   U26 : AOI22_X1 port map( A1 => n2, A2 => IN3(30), B1 => n1, B2 => IN2(30), 
                           ZN => n125);
   U25 : NAND2_X1 port map( A1 => n126, A2 => n125, ZN => OUT1(30));
   U39 : AOI22_X1 port map( A1 => n74, A2 => IN1(27), B1 => n72, B2 => IN0(27),
                           ZN => n118);
   U37 : NAND2_X1 port map( A1 => n118, A2 => n117, ZN => OUT1(27));
   U42 : AOI22_X1 port map( A1 => n74, A2 => IN1(26), B1 => n72, B2 => IN0(26),
                           ZN => n116);
   U41 : AOI22_X1 port map( A1 => n2, A2 => IN3(26), B1 => n1, B2 => IN2(26), 
                           ZN => n115);
   U40 : NAND2_X1 port map( A1 => n116, A2 => n115, ZN => OUT1(26));
   U45 : AOI22_X1 port map( A1 => n74, A2 => IN1(25), B1 => n72, B2 => IN0(25),
                           ZN => n114);
   U43 : NAND2_X1 port map( A1 => n114, A2 => n113, ZN => OUT1(25));
   U48 : AOI22_X1 port map( A1 => n74, A2 => IN1(24), B1 => n72, B2 => IN0(24),
                           ZN => n112);
   U47 : AOI22_X1 port map( A1 => n2, A2 => IN3(24), B1 => n1, B2 => IN2(24), 
                           ZN => n111);
   U46 : NAND2_X1 port map( A1 => n112, A2 => n111, ZN => OUT1(24));
   U28 : NAND2_X1 port map( A1 => n124, A2 => n123, ZN => OUT1(2));
   U10 : NAND2_X1 port map( A1 => n136, A2 => n135, ZN => OUT1(6));
   U13 : NAND2_X1 port map( A1 => n134, A2 => n133, ZN => OUT1(5));
   U16 : NAND2_X1 port map( A1 => n132, A2 => n131, ZN => OUT1(4));
   U88 : NAND2_X1 port map( A1 => n84, A2 => n83, ZN => OUT1(11));
   U91 : NAND2_X1 port map( A1 => n82, A2 => n81, ZN => OUT1(10));
   U1 : NAND2_X1 port map( A1 => n146, A2 => n145, ZN => OUT1(9));
   U79 : NAND2_X1 port map( A1 => n90, A2 => n89, ZN => OUT1(14));
   U82 : NAND2_X1 port map( A1 => n88, A2 => n87, ZN => OUT1(13));
   U85 : NAND2_X1 port map( A1 => n86, A2 => n85, ZN => OUT1(12));
   U61 : NAND2_X1 port map( A1 => n102, A2 => n101, ZN => OUT1(1));
   U19 : NAND2_X1 port map( A1 => n130, A2 => n129, ZN => OUT1(3));
   U7 : NAND2_X1 port map( A1 => n138, A2 => n137, ZN => OUT1(7));
   U4 : NAND2_X1 port map( A1 => n140, A2 => n139, ZN => OUT1(8));
   U76 : NAND2_X1 port map( A1 => n92, A2 => n91, ZN => OUT1(15));
   U20 : BUF_X4 port map( A => n143, Z => n1);
   U29 : AND2_X2 port map( A1 => n78, A2 => CTRL(0), ZN => n142);
   U38 : BUF_X2 port map( A => n142, Z => n75);
   U44 : BUF_X1 port map( A => n142, Z => n74);
   U50 : BUF_X2 port map( A => n144, Z => n2);
   U53 : BUF_X1 port map( A => n144, Z => n77);
   U56 : BUF_X1 port map( A => n141, Z => n73);
   U62 : BUF_X2 port map( A => n141, Z => n72);
   U65 : BUF_X2 port map( A => n143, Z => n76);
   U68 : INV_X1 port map( A => CTRL(1), ZN => n78);
   U71 : AND2_X1 port map( A1 => CTRL(0), A2 => CTRL(1), ZN => n144);
   U74 : AOI22_X1 port map( A1 => n2, A2 => IN3(23), B1 => n1, B2 => IN2(23), 
                           ZN => n109);
   U77 : AOI22_X1 port map( A1 => n2, A2 => IN3(21), B1 => n1, B2 => IN2(21), 
                           ZN => n105);
   U80 : AOI22_X1 port map( A1 => n2, A2 => IN3(22), B1 => n1, B2 => IN2(22), 
                           ZN => n107);
   U83 : AOI22_X1 port map( A1 => n2, A2 => IN3(2), B1 => n1, B2 => IN2(2), ZN 
                           => n123);
   U86 : AOI22_X1 port map( A1 => n2, A2 => IN3(27), B1 => n1, B2 => IN2(27), 
                           ZN => n117);
   U89 : AOI22_X1 port map( A1 => n2, A2 => IN3(25), B1 => n1, B2 => IN2(25), 
                           ZN => n113);
   U92 : AOI22_X1 port map( A1 => n2, A2 => IN3(3), B1 => n1, B2 => IN2(3), ZN 
                           => n129);
   U94 : NAND2_X1 port map( A1 => n80, A2 => n79, ZN => OUT1(0));
   U95 : AOI22_X1 port map( A1 => n77, A2 => IN3(16), B1 => n76, B2 => IN2(16),
                           ZN => n93);
   U96 : AOI22_X1 port map( A1 => n77, A2 => IN3(12), B1 => n76, B2 => IN2(12),
                           ZN => n85);
   U97 : AOI22_X1 port map( A1 => n77, A2 => IN3(18), B1 => n76, B2 => IN2(18),
                           ZN => n97);
   U99 : AOI22_X1 port map( A1 => n77, A2 => IN3(10), B1 => n76, B2 => IN2(10),
                           ZN => n81);
   U100 : AOI22_X1 port map( A1 => n77, A2 => IN3(14), B1 => n76, B2 => IN2(14)
                           , ZN => n89);
   U101 : AOI22_X1 port map( A1 => n77, A2 => IN3(13), B1 => n76, B2 => IN2(13)
                           , ZN => n87);
   U102 : AOI22_X1 port map( A1 => n77, A2 => IN3(19), B1 => n76, B2 => IN2(19)
                           , ZN => n99);
   U103 : AOI22_X1 port map( A1 => n77, A2 => IN3(17), B1 => n76, B2 => IN2(17)
                           , ZN => n95);
   U104 : AOI22_X1 port map( A1 => n77, A2 => IN3(1), B1 => n76, B2 => IN2(1), 
                           ZN => n101);
   U105 : AOI22_X1 port map( A1 => n77, A2 => IN3(15), B1 => n76, B2 => IN2(15)
                           , ZN => n91);
   U106 : AOI22_X1 port map( A1 => n77, A2 => IN3(11), B1 => n76, B2 => IN2(11)
                           , ZN => n83);
   U107 : AOI22_X1 port map( A1 => n77, A2 => IN3(0), B1 => n76, B2 => IN2(0), 
                           ZN => n79);
   U108 : NOR2_X1 port map( A1 => CTRL(1), A2 => CTRL(0), ZN => n141);
   U109 : NOR2_X1 port map( A1 => CTRL(0), A2 => n78, ZN => n143);

end SYN_bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity mux41_MUX_SIZE32_1 is

   port( IN0, IN1, IN2, IN3 : in std_logic_vector (31 downto 0);  CTRL : in 
         std_logic_vector (1 downto 0);  OUT1 : out std_logic_vector (31 downto
         0));

end mux41_MUX_SIZE32_1;

architecture SYN_bhe of mux41_MUX_SIZE32_1 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X3
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n47, n48, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, 
      n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93
      , n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
      n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, 
      n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, 
      n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, 
      n143, n144, n145, n146, n147 : std_logic;

begin
   
   U25 : NAND2_X1 port map( A1 => n128, A2 => n127, ZN => OUT1(30));
   U22 : NAND2_X1 port map( A1 => n130, A2 => n129, ZN => OUT1(31));
   U46 : NAND2_X1 port map( A1 => n114, A2 => n113, ZN => OUT1(24));
   U1 : BUF_X1 port map( A => n69, Z => n2);
   U2 : CLKBUF_X3 port map( A => n69, Z => n1);
   U3 : BUF_X1 port map( A => n69, Z => n47);
   U4 : NOR2_X1 port map( A1 => n48, A2 => CTRL(0), ZN => n69);
   U5 : BUF_X2 port map( A => n144, Z => n79);
   U6 : AND2_X2 port map( A1 => n48, A2 => CTRL(0), ZN => n144);
   U7 : BUF_X1 port map( A => n144, Z => n74);
   U8 : BUF_X1 port map( A => n145, Z => n82);
   U9 : BUF_X1 port map( A => n145, Z => n84);
   U10 : BUF_X2 port map( A => n144, Z => n80);
   U11 : BUF_X2 port map( A => n144, Z => n81);
   U12 : BUF_X2 port map( A => n144, Z => n75);
   U13 : BUF_X2 port map( A => n143, Z => n78);
   U14 : BUF_X2 port map( A => n143, Z => n77);
   U15 : BUF_X2 port map( A => n143, Z => n76);
   U16 : BUF_X2 port map( A => n145, Z => n83);
   U17 : AND2_X1 port map( A1 => CTRL(1), A2 => CTRL(0), ZN => n145);
   U18 : INV_X1 port map( A => CTRL(1), ZN => n48);
   U19 : NAND2_X1 port map( A1 => n1, A2 => IN2(1), ZN => n70);
   U20 : NAND2_X1 port map( A1 => n1, A2 => IN2(0), ZN => n72);
   U21 : AOI22_X1 port map( A1 => n84, A2 => IN3(6), B1 => n47, B2 => IN2(6), 
                           ZN => n137);
   U23 : AOI22_X1 port map( A1 => n82, A2 => IN3(18), B1 => n1, B2 => IN2(18), 
                           ZN => n101);
   U24 : AOI22_X1 port map( A1 => n82, A2 => IN3(13), B1 => n2, B2 => IN2(13), 
                           ZN => n91);
   U26 : AOI22_X1 port map( A1 => n82, A2 => IN3(15), B1 => n1, B2 => IN2(15), 
                           ZN => n95);
   U27 : AOI22_X1 port map( A1 => n83, A2 => IN3(23), B1 => n2, B2 => IN2(23), 
                           ZN => n111);
   U28 : NAND2_X1 port map( A1 => n72, A2 => n73, ZN => OUT1(0));
   U29 : NOR2_X1 port map( A1 => CTRL(0), A2 => CTRL(1), ZN => n143);
   U30 : AOI22_X1 port map( A1 => n79, A2 => IN1(1), B1 => n78, B2 => IN0(1), 
                           ZN => n71);
   U31 : NAND2_X1 port map( A1 => n71, A2 => n70, ZN => OUT1(1));
   U32 : AOI22_X1 port map( A1 => n79, A2 => IN1(0), B1 => n78, B2 => IN0(0), 
                           ZN => n73);
   U33 : NAND2_X1 port map( A1 => n2, A2 => IN2(19), ZN => n103);
   U34 : NAND2_X1 port map( A1 => n131, A2 => n132, ZN => OUT1(3));
   U35 : NAND2_X1 port map( A1 => n106, A2 => n105, ZN => OUT1(20));
   U36 : NAND2_X1 port map( A1 => n124, A2 => n123, ZN => OUT1(29));
   U37 : NAND2_X1 port map( A1 => n120, A2 => n119, ZN => OUT1(27));
   U38 : NAND2_X1 port map( A1 => n90, A2 => n89, ZN => OUT1(12));
   U39 : NAND2_X1 port map( A1 => n98, A2 => n97, ZN => OUT1(16));
   U40 : NAND2_X1 port map( A1 => n118, A2 => n117, ZN => OUT1(26));
   U41 : NAND2_X1 port map( A1 => n142, A2 => n141, ZN => OUT1(8));
   U42 : NAND2_X1 port map( A1 => n138, A2 => n137, ZN => OUT1(6));
   U43 : NAND2_X1 port map( A1 => n134, A2 => n133, ZN => OUT1(4));
   U44 : NAND2_X1 port map( A1 => n122, A2 => n121, ZN => OUT1(28));
   U45 : NAND2_X1 port map( A1 => n86, A2 => n85, ZN => OUT1(10));
   U47 : NAND2_X1 port map( A1 => n109, A2 => n110, ZN => OUT1(22));
   U48 : NAND2_X1 port map( A1 => n104, A2 => n103, ZN => OUT1(19));
   U49 : NAND2_X1 port map( A1 => n107, A2 => n108, ZN => OUT1(21));
   U50 : NAND2_X1 port map( A1 => n96, A2 => n95, ZN => OUT1(15));
   U51 : NAND2_X1 port map( A1 => n147, A2 => n146, ZN => OUT1(9));
   U52 : NAND2_X1 port map( A1 => n100, A2 => n99, ZN => OUT1(17));
   U53 : NAND2_X1 port map( A1 => n102, A2 => n101, ZN => OUT1(18));
   U54 : AOI22_X1 port map( A1 => n74, A2 => IN1(30), B1 => n77, B2 => IN0(30),
                           ZN => n128);
   U55 : AOI22_X1 port map( A1 => n75, A2 => IN1(29), B1 => n77, B2 => IN0(29),
                           ZN => n124);
   U56 : AOI22_X1 port map( A1 => n75, A2 => IN1(25), B1 => n77, B2 => IN0(25),
                           ZN => n116);
   U57 : AOI22_X1 port map( A1 => n81, A2 => IN1(24), B1 => n76, B2 => IN0(24),
                           ZN => n114);
   U58 : AOI22_X1 port map( A1 => n74, A2 => IN1(27), B1 => n76, B2 => IN0(27),
                           ZN => n120);
   U59 : AOI22_X1 port map( A1 => n80, A2 => IN1(26), B1 => n77, B2 => IN0(26),
                           ZN => n118);
   U60 : AOI22_X1 port map( A1 => n81, A2 => IN1(20), B1 => n76, B2 => IN0(20),
                           ZN => n106);
   U61 : AOI22_X1 port map( A1 => n81, A2 => IN1(2), B1 => n76, B2 => IN0(2), 
                           ZN => n126);
   U62 : AOI22_X1 port map( A1 => n75, A2 => IN1(22), B1 => n76, B2 => IN0(22),
                           ZN => n110);
   U63 : AOI22_X1 port map( A1 => n74, A2 => IN1(23), B1 => n76, B2 => IN0(23),
                           ZN => n112);
   U64 : AOI22_X1 port map( A1 => n74, A2 => IN1(28), B1 => n77, B2 => IN0(28),
                           ZN => n122);
   U65 : AOI22_X1 port map( A1 => n74, A2 => IN1(21), B1 => n77, B2 => IN0(21),
                           ZN => n108);
   U66 : NAND2_X1 port map( A1 => n112, A2 => n111, ZN => OUT1(23));
   U67 : AOI22_X1 port map( A1 => n80, A2 => IN1(31), B1 => n76, B2 => IN0(31),
                           ZN => n130);
   U68 : AOI22_X1 port map( A1 => n79, A2 => IN1(3), B1 => n78, B2 => IN0(3), 
                           ZN => n132);
   U69 : AOI22_X1 port map( A1 => n75, A2 => IN1(6), B1 => n77, B2 => IN0(6), 
                           ZN => n138);
   U70 : AOI22_X1 port map( A1 => n81, A2 => IN1(8), B1 => n77, B2 => IN0(8), 
                           ZN => n142);
   U71 : AOI22_X1 port map( A1 => n80, A2 => IN1(4), B1 => n77, B2 => IN0(4), 
                           ZN => n134);
   U72 : AOI22_X1 port map( A1 => n79, A2 => IN1(7), B1 => n76, B2 => IN0(7), 
                           ZN => n140);
   U73 : AOI22_X1 port map( A1 => n81, A2 => IN1(5), B1 => n76, B2 => IN0(5), 
                           ZN => n136);
   U74 : AOI22_X1 port map( A1 => n74, A2 => IN1(9), B1 => n76, B2 => IN0(9), 
                           ZN => n147);
   U75 : NAND2_X1 port map( A1 => n92, A2 => n91, ZN => OUT1(13));
   U76 : AOI22_X1 port map( A1 => n84, A2 => IN3(31), B1 => n47, B2 => IN2(31),
                           ZN => n129);
   U77 : AOI22_X1 port map( A1 => n84, A2 => IN3(3), B1 => n2, B2 => IN2(3), ZN
                           => n131);
   U78 : AOI22_X1 port map( A1 => n84, A2 => IN3(4), B1 => n47, B2 => IN2(4), 
                           ZN => n133);
   U79 : AOI22_X1 port map( A1 => n84, A2 => IN3(7), B1 => n2, B2 => IN2(7), ZN
                           => n139);
   U80 : AOI22_X1 port map( A1 => n84, A2 => IN3(5), B1 => n47, B2 => IN2(5), 
                           ZN => n135);
   U81 : AOI22_X1 port map( A1 => n84, A2 => IN3(8), B1 => n47, B2 => IN2(8), 
                           ZN => n141);
   U82 : AOI22_X1 port map( A1 => n84, A2 => IN3(9), B1 => n47, B2 => IN2(9), 
                           ZN => n146);
   U83 : NAND2_X1 port map( A1 => n125, A2 => n126, ZN => OUT1(2));
   U84 : NAND2_X1 port map( A1 => n116, A2 => n115, ZN => OUT1(25));
   U85 : NAND2_X1 port map( A1 => n88, A2 => n87, ZN => OUT1(11));
   U86 : NAND2_X1 port map( A1 => n94, A2 => n93, ZN => OUT1(14));
   U87 : NAND2_X1 port map( A1 => n140, A2 => n139, ZN => OUT1(7));
   U88 : AOI22_X1 port map( A1 => n83, A2 => IN3(30), B1 => n2, B2 => IN2(30), 
                           ZN => n127);
   U89 : AOI22_X1 port map( A1 => n83, A2 => IN3(29), B1 => n47, B2 => IN2(29),
                           ZN => n123);
   U90 : AOI22_X1 port map( A1 => n83, A2 => IN3(24), B1 => n2, B2 => IN2(24), 
                           ZN => n113);
   U91 : AOI22_X1 port map( A1 => n83, A2 => IN3(27), B1 => n1, B2 => IN2(27), 
                           ZN => n119);
   U92 : AOI22_X1 port map( A1 => n83, A2 => IN3(26), B1 => n2, B2 => IN2(26), 
                           ZN => n117);
   U93 : AOI22_X1 port map( A1 => n83, A2 => IN3(28), B1 => n1, B2 => IN2(28), 
                           ZN => n121);
   U94 : AOI22_X1 port map( A1 => n83, A2 => IN3(20), B1 => n2, B2 => IN2(20), 
                           ZN => n105);
   U95 : AOI22_X1 port map( A1 => n83, A2 => IN3(25), B1 => n47, B2 => IN2(25),
                           ZN => n115);
   U96 : AOI22_X1 port map( A1 => n83, A2 => IN3(22), B1 => n1, B2 => IN2(22), 
                           ZN => n109);
   U97 : AOI22_X1 port map( A1 => n83, A2 => IN3(2), B1 => IN2(2), B2 => n2, ZN
                           => n125);
   U98 : AOI22_X1 port map( A1 => n83, A2 => IN3(21), B1 => n1, B2 => IN2(21), 
                           ZN => n107);
   U99 : AOI22_X1 port map( A1 => n81, A2 => IN1(16), B1 => n76, B2 => IN0(16),
                           ZN => n98);
   U100 : AOI22_X1 port map( A1 => n81, A2 => IN1(19), B1 => n78, B2 => IN0(19)
                           , ZN => n104);
   U101 : AOI22_X1 port map( A1 => n75, A2 => IN1(12), B1 => n77, B2 => IN0(12)
                           , ZN => n90);
   U102 : AOI22_X1 port map( A1 => n80, A2 => IN1(18), B1 => n78, B2 => IN0(18)
                           , ZN => n102);
   U103 : AOI22_X1 port map( A1 => n80, A2 => IN1(11), B1 => n76, B2 => IN0(11)
                           , ZN => n88);
   U104 : AOI22_X1 port map( A1 => n79, A2 => IN1(10), B1 => n77, B2 => IN0(10)
                           , ZN => n86);
   U105 : AOI22_X1 port map( A1 => n80, A2 => IN1(14), B1 => n77, B2 => IN0(14)
                           , ZN => n94);
   U106 : AOI22_X1 port map( A1 => n74, A2 => IN1(15), B1 => n77, B2 => IN0(15)
                           , ZN => n96);
   U107 : AOI22_X1 port map( A1 => n75, A2 => IN1(17), B1 => n78, B2 => IN0(17)
                           , ZN => n100);
   U108 : AOI22_X1 port map( A1 => n75, A2 => IN1(13), B1 => n76, B2 => IN0(13)
                           , ZN => n92);
   U109 : NAND2_X1 port map( A1 => n136, A2 => n135, ZN => OUT1(5));
   U110 : AOI22_X1 port map( A1 => n82, A2 => IN3(16), B1 => n2, B2 => IN2(16),
                           ZN => n97);
   U111 : AOI22_X1 port map( A1 => n82, A2 => IN3(12), B1 => n1, B2 => IN2(12),
                           ZN => n89);
   U112 : AOI22_X1 port map( A1 => n82, A2 => IN3(11), B1 => n47, B2 => IN2(11)
                           , ZN => n87);
   U113 : AOI22_X1 port map( A1 => n82, A2 => IN3(10), B1 => n1, B2 => IN2(10),
                           ZN => n85);
   U114 : AOI22_X1 port map( A1 => n82, A2 => IN3(17), B1 => n1, B2 => IN2(17),
                           ZN => n99);
   U115 : AOI22_X1 port map( A1 => n82, A2 => IN3(14), B1 => n47, B2 => IN2(14)
                           , ZN => n93);

end SYN_bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity mux21_4 is

   port( IN0, IN1 : in std_logic_vector (31 downto 0);  CTRL : in std_logic;  
         OUT1 : out std_logic_vector (31 downto 0));

end mux21_4;

architecture SYN_Bhe of mux21_4 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => IN0(9), B => IN1(9), S => CTRL, Z => OUT1(9));
   U2 : MUX2_X1 port map( A => IN0(8), B => IN1(8), S => CTRL, Z => OUT1(8));
   U3 : MUX2_X1 port map( A => IN0(7), B => IN1(7), S => CTRL, Z => OUT1(7));
   U4 : MUX2_X1 port map( A => IN0(6), B => IN1(6), S => CTRL, Z => OUT1(6));
   U5 : MUX2_X1 port map( A => IN0(5), B => IN1(5), S => CTRL, Z => OUT1(5));
   U6 : MUX2_X1 port map( A => IN0(4), B => IN1(4), S => CTRL, Z => OUT1(4));
   U7 : MUX2_X1 port map( A => IN0(3), B => IN1(3), S => CTRL, Z => OUT1(3));
   U8 : MUX2_X1 port map( A => IN0(31), B => IN1(31), S => CTRL, Z => OUT1(31))
                           ;
   U9 : MUX2_X1 port map( A => IN0(30), B => IN1(30), S => CTRL, Z => OUT1(30))
                           ;
   U10 : MUX2_X1 port map( A => IN0(2), B => IN1(2), S => CTRL, Z => OUT1(2));
   U11 : MUX2_X1 port map( A => IN0(29), B => IN1(29), S => CTRL, Z => OUT1(29)
                           );
   U12 : MUX2_X1 port map( A => IN0(28), B => IN1(28), S => CTRL, Z => OUT1(28)
                           );
   U16 : MUX2_X1 port map( A => IN0(24), B => IN1(24), S => CTRL, Z => OUT1(24)
                           );
   U17 : MUX2_X1 port map( A => IN0(23), B => IN1(23), S => CTRL, Z => OUT1(23)
                           );
   U18 : MUX2_X1 port map( A => IN0(22), B => IN1(22), S => CTRL, Z => OUT1(22)
                           );
   U19 : MUX2_X1 port map( A => IN0(21), B => IN1(21), S => CTRL, Z => OUT1(21)
                           );
   U20 : MUX2_X1 port map( A => IN0(20), B => IN1(20), S => CTRL, Z => OUT1(20)
                           );
   U21 : MUX2_X1 port map( A => IN0(1), B => IN1(1), S => CTRL, Z => OUT1(1));
   U22 : MUX2_X1 port map( A => IN0(19), B => IN1(19), S => CTRL, Z => OUT1(19)
                           );
   U23 : MUX2_X1 port map( A => IN0(18), B => IN1(18), S => CTRL, Z => OUT1(18)
                           );
   U24 : MUX2_X1 port map( A => IN0(17), B => IN1(17), S => CTRL, Z => OUT1(17)
                           );
   U25 : MUX2_X1 port map( A => IN0(16), B => IN1(16), S => CTRL, Z => OUT1(16)
                           );
   U26 : MUX2_X1 port map( A => IN0(15), B => IN1(15), S => CTRL, Z => OUT1(15)
                           );
   U27 : MUX2_X1 port map( A => IN0(14), B => IN1(14), S => CTRL, Z => OUT1(14)
                           );
   U28 : MUX2_X1 port map( A => IN0(13), B => IN1(13), S => CTRL, Z => OUT1(13)
                           );
   U29 : MUX2_X1 port map( A => IN0(12), B => IN1(12), S => CTRL, Z => OUT1(12)
                           );
   U30 : MUX2_X1 port map( A => IN0(11), B => IN1(11), S => CTRL, Z => OUT1(11)
                           );
   U31 : MUX2_X1 port map( A => IN0(10), B => IN1(10), S => CTRL, Z => OUT1(10)
                           );
   U32 : MUX2_X1 port map( A => IN0(0), B => IN1(0), S => CTRL, Z => OUT1(0));
   U13 : MUX2_X1 port map( A => IN0(27), B => IN1(27), S => CTRL, Z => OUT1(27)
                           );
   U14 : MUX2_X1 port map( A => IN0(26), B => IN1(26), S => CTRL, Z => OUT1(26)
                           );
   U15 : MUX2_X1 port map( A => IN0(25), B => IN1(25), S => CTRL, Z => OUT1(25)
                           );

end SYN_Bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity mux21_3 is

   port( IN0, IN1 : in std_logic_vector (31 downto 0);  CTRL : in std_logic;  
         OUT1 : out std_logic_vector (31 downto 0));

end mux21_3;

architecture SYN_Bhe of mux21_3 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X2
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n3, n4, n5, n6, n7 : std_logic;

begin
   
   U2 : MUX2_X1 port map( A => IN0(8), B => IN1(8), S => CTRL, Z => OUT1(8));
   U8 : MUX2_X1 port map( A => IN0(31), B => IN1(31), S => CTRL, Z => OUT1(31))
                           ;
   U9 : MUX2_X1 port map( A => IN0(30), B => IN1(30), S => CTRL, Z => OUT1(30))
                           ;
   U11 : MUX2_X1 port map( A => IN0(29), B => IN1(29), S => CTRL, Z => OUT1(29)
                           );
   U13 : MUX2_X1 port map( A => IN0(27), B => IN1(27), S => CTRL, Z => OUT1(27)
                           );
   U14 : MUX2_X1 port map( A => IN0(26), B => IN1(26), S => CTRL, Z => OUT1(26)
                           );
   U16 : MUX2_X1 port map( A => IN0(24), B => IN1(24), S => CTRL, Z => OUT1(24)
                           );
   U20 : MUX2_X1 port map( A => IN0(20), B => IN1(20), S => CTRL, Z => OUT1(20)
                           );
   U1 : MUX2_X1 port map( A => IN0(18), B => IN1(18), S => CTRL, Z => OUT1(18))
                           ;
   U3 : AOI22_X1 port map( A1 => CTRL, A2 => IN1(6), B1 => n3, B2 => IN0(6), ZN
                           => n1);
   U4 : INV_X1 port map( A => n1, ZN => OUT1(6));
   U5 : MUX2_X1 port map( A => IN0(2), B => IN1(2), S => CTRL, Z => OUT1(2));
   U6 : MUX2_X2 port map( A => IN0(4), B => IN1(4), S => CTRL, Z => OUT1(4));
   U7 : NAND2_X1 port map( A1 => IN0(13), A2 => n3, ZN => n4);
   U10 : NAND2_X1 port map( A1 => IN1(13), A2 => CTRL, ZN => n5);
   U12 : NAND2_X2 port map( A1 => n4, A2 => n5, ZN => OUT1(13));
   U15 : INV_X1 port map( A => CTRL, ZN => n3);
   U17 : MUX2_X1 port map( A => IN0(25), B => IN1(25), S => CTRL, Z => OUT1(25)
                           );
   U18 : MUX2_X1 port map( A => IN0(28), B => IN1(28), S => CTRL, Z => OUT1(28)
                           );
   U19 : MUX2_X1 port map( A => IN0(23), B => IN1(23), S => CTRL, Z => OUT1(23)
                           );
   U21 : MUX2_X1 port map( A => IN0(22), B => IN1(22), S => CTRL, Z => OUT1(22)
                           );
   U22 : MUX2_X1 port map( A => IN0(16), B => IN1(16), S => CTRL, Z => OUT1(16)
                           );
   U23 : MUX2_X1 port map( A => IN0(9), B => IN1(9), S => CTRL, Z => OUT1(9));
   U24 : MUX2_X1 port map( A => IN0(10), B => IN1(10), S => CTRL, Z => OUT1(10)
                           );
   U25 : MUX2_X1 port map( A => IN0(3), B => IN1(3), S => CTRL, Z => OUT1(3));
   U26 : MUX2_X1 port map( A => IN0(12), B => IN1(12), S => CTRL, Z => OUT1(12)
                           );
   U27 : NAND2_X1 port map( A1 => n6, A2 => n7, ZN => OUT1(0));
   U28 : MUX2_X1 port map( A => IN0(1), B => IN1(1), S => CTRL, Z => OUT1(1));
   U29 : NAND2_X1 port map( A1 => IN1(0), A2 => CTRL, ZN => n7);
   U30 : NAND2_X1 port map( A1 => IN0(0), A2 => n3, ZN => n6);
   U31 : MUX2_X1 port map( A => IN0(19), B => IN1(19), S => CTRL, Z => OUT1(19)
                           );
   U32 : MUX2_X1 port map( A => IN0(7), B => IN1(7), S => CTRL, Z => OUT1(7));
   U33 : MUX2_X1 port map( A => IN0(17), B => IN1(17), S => CTRL, Z => OUT1(17)
                           );
   U34 : MUX2_X1 port map( A => IN0(21), B => IN1(21), S => CTRL, Z => OUT1(21)
                           );
   U35 : MUX2_X1 port map( A => IN0(14), B => IN1(14), S => CTRL, Z => OUT1(14)
                           );
   U36 : MUX2_X1 port map( A => IN0(11), B => IN1(11), S => CTRL, Z => OUT1(11)
                           );
   U37 : MUX2_X1 port map( A => IN0(15), B => IN1(15), S => CTRL, Z => OUT1(15)
                           );
   U38 : MUX2_X1 port map( A => IN0(5), B => IN1(5), S => CTRL, Z => OUT1(5));

end SYN_Bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity mux21_2 is

   port( IN0, IN1 : in std_logic_vector (31 downto 0);  OUT1 : out 
         std_logic_vector (31 downto 0);  CTRL_BAR : in std_logic);

end mux21_2;

architecture SYN_Bhe of mux21_2 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : MUX2_X1 port map( A => IN0(9), B => IN1(9), S => n3, Z => OUT1(9));
   U2 : MUX2_X1 port map( A => IN0(8), B => IN1(8), S => n3, Z => OUT1(8));
   U3 : MUX2_X1 port map( A => IN0(7), B => IN1(7), S => n3, Z => OUT1(7));
   U4 : MUX2_X1 port map( A => IN0(6), B => IN1(6), S => n3, Z => OUT1(6));
   U5 : MUX2_X1 port map( A => IN0(5), B => IN1(5), S => n3, Z => OUT1(5));
   U6 : MUX2_X1 port map( A => IN0(4), B => IN1(4), S => n3, Z => OUT1(4));
   U7 : MUX2_X1 port map( A => IN0(3), B => IN1(3), S => n3, Z => OUT1(3));
   U8 : MUX2_X1 port map( A => IN0(31), B => IN1(31), S => n3, Z => OUT1(31));
   U9 : MUX2_X1 port map( A => IN0(30), B => IN1(30), S => n3, Z => OUT1(30));
   U10 : MUX2_X1 port map( A => IN0(2), B => IN1(2), S => n3, Z => OUT1(2));
   U11 : MUX2_X1 port map( A => IN0(29), B => IN1(29), S => n3, Z => OUT1(29));
   U12 : MUX2_X1 port map( A => IN0(28), B => IN1(28), S => n3, Z => OUT1(28));
   U13 : MUX2_X1 port map( A => IN0(27), B => IN1(27), S => n2, Z => OUT1(27));
   U14 : MUX2_X1 port map( A => IN0(26), B => IN1(26), S => n2, Z => OUT1(26));
   U15 : MUX2_X1 port map( A => IN0(25), B => IN1(25), S => n2, Z => OUT1(25));
   U16 : MUX2_X1 port map( A => IN0(24), B => IN1(24), S => n2, Z => OUT1(24));
   U17 : MUX2_X1 port map( A => IN0(23), B => IN1(23), S => n2, Z => OUT1(23));
   U18 : MUX2_X1 port map( A => IN0(22), B => IN1(22), S => n2, Z => OUT1(22));
   U19 : MUX2_X1 port map( A => IN0(21), B => IN1(21), S => n2, Z => OUT1(21));
   U20 : MUX2_X1 port map( A => IN0(20), B => IN1(20), S => n2, Z => OUT1(20));
   U21 : MUX2_X1 port map( A => IN0(1), B => IN1(1), S => n2, Z => OUT1(1));
   U22 : MUX2_X1 port map( A => IN0(19), B => IN1(19), S => n2, Z => OUT1(19));
   U23 : MUX2_X1 port map( A => IN0(18), B => IN1(18), S => n2, Z => OUT1(18));
   U24 : MUX2_X1 port map( A => IN0(17), B => IN1(17), S => n2, Z => OUT1(17));
   U25 : MUX2_X1 port map( A => IN0(16), B => IN1(16), S => n1, Z => OUT1(16));
   U26 : MUX2_X1 port map( A => IN0(15), B => IN1(15), S => n1, Z => OUT1(15));
   U27 : MUX2_X1 port map( A => IN0(14), B => IN1(14), S => n1, Z => OUT1(14));
   U28 : MUX2_X1 port map( A => IN0(13), B => IN1(13), S => n1, Z => OUT1(13));
   U29 : MUX2_X1 port map( A => IN0(12), B => IN1(12), S => n1, Z => OUT1(12));
   U30 : MUX2_X1 port map( A => IN0(11), B => IN1(11), S => n1, Z => OUT1(11));
   U31 : MUX2_X1 port map( A => IN0(10), B => IN1(10), S => n1, Z => OUT1(10));
   U32 : MUX2_X1 port map( A => IN0(0), B => IN1(0), S => n1, Z => OUT1(0));
   U33 : INV_X1 port map( A => CTRL_BAR, ZN => n1);
   U34 : INV_X1 port map( A => CTRL_BAR, ZN => n2);
   U35 : INV_X1 port map( A => CTRL_BAR, ZN => n3);

end SYN_Bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity mux21_1 is

   port( IN0, IN1 : in std_logic_vector (31 downto 0);  CTRL : in std_logic;  
         OUT1 : out std_logic_vector (31 downto 0));

end mux21_1;

architecture SYN_Bhe of mux21_1 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : MUX2_X1 port map( A => IN0(9), B => IN1(9), S => CTRL, Z => OUT1(9));
   U2 : MUX2_X1 port map( A => IN0(8), B => IN1(8), S => CTRL, Z => OUT1(8));
   U3 : MUX2_X1 port map( A => IN0(7), B => IN1(7), S => CTRL, Z => OUT1(7));
   U4 : MUX2_X1 port map( A => IN0(6), B => IN1(6), S => CTRL, Z => OUT1(6));
   U6 : MUX2_X1 port map( A => IN0(4), B => IN1(4), S => CTRL, Z => OUT1(4));
   U7 : MUX2_X1 port map( A => IN0(3), B => IN1(3), S => CTRL, Z => OUT1(3));
   U8 : MUX2_X1 port map( A => IN0(31), B => IN1(31), S => CTRL, Z => OUT1(31))
                           ;
   U9 : MUX2_X1 port map( A => IN0(30), B => IN1(30), S => CTRL, Z => OUT1(30))
                           ;
   U10 : MUX2_X1 port map( A => IN0(2), B => IN1(2), S => CTRL, Z => OUT1(2));
   U11 : MUX2_X1 port map( A => IN0(29), B => IN1(29), S => CTRL, Z => OUT1(29)
                           );
   U12 : MUX2_X1 port map( A => IN0(28), B => IN1(28), S => CTRL, Z => OUT1(28)
                           );
   U13 : MUX2_X1 port map( A => IN0(27), B => IN1(27), S => CTRL, Z => OUT1(27)
                           );
   U14 : MUX2_X1 port map( A => IN0(26), B => IN1(26), S => CTRL, Z => OUT1(26)
                           );
   U15 : MUX2_X1 port map( A => IN0(25), B => IN1(25), S => CTRL, Z => OUT1(25)
                           );
   U16 : MUX2_X1 port map( A => IN0(24), B => IN1(24), S => CTRL, Z => OUT1(24)
                           );
   U17 : MUX2_X1 port map( A => IN0(23), B => IN1(23), S => CTRL, Z => OUT1(23)
                           );
   U18 : MUX2_X1 port map( A => IN0(22), B => IN1(22), S => CTRL, Z => OUT1(22)
                           );
   U19 : MUX2_X1 port map( A => IN0(21), B => IN1(21), S => CTRL, Z => OUT1(21)
                           );
   U20 : MUX2_X1 port map( A => IN0(20), B => IN1(20), S => CTRL, Z => OUT1(20)
                           );
   U21 : MUX2_X1 port map( A => IN0(1), B => IN1(1), S => CTRL, Z => OUT1(1));
   U22 : MUX2_X1 port map( A => IN0(19), B => IN1(19), S => CTRL, Z => OUT1(19)
                           );
   U23 : MUX2_X1 port map( A => IN0(18), B => IN1(18), S => CTRL, Z => OUT1(18)
                           );
   U24 : MUX2_X1 port map( A => IN0(17), B => IN1(17), S => CTRL, Z => OUT1(17)
                           );
   U25 : MUX2_X1 port map( A => IN0(16), B => IN1(16), S => CTRL, Z => OUT1(16)
                           );
   U26 : MUX2_X1 port map( A => IN0(15), B => IN1(15), S => CTRL, Z => OUT1(15)
                           );
   U27 : MUX2_X1 port map( A => IN0(14), B => IN1(14), S => CTRL, Z => OUT1(14)
                           );
   U28 : MUX2_X1 port map( A => IN0(13), B => IN1(13), S => CTRL, Z => OUT1(13)
                           );
   U29 : MUX2_X1 port map( A => IN0(12), B => IN1(12), S => CTRL, Z => OUT1(12)
                           );
   U30 : MUX2_X1 port map( A => IN0(11), B => IN1(11), S => CTRL, Z => OUT1(11)
                           );
   U31 : MUX2_X1 port map( A => IN0(10), B => IN1(10), S => CTRL, Z => OUT1(10)
                           );
   U5 : MUX2_X1 port map( A => IN0(5), B => IN1(5), S => CTRL, Z => OUT1(5));
   U32 : INV_X1 port map( A => IN0(0), ZN => n1);
   U33 : NOR2_X1 port map( A1 => CTRL, A2 => n1, ZN => OUT1(0));

end SYN_Bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity p4add_N32_logN5_1 is

   port( A, B : in std_logic_vector (31 downto 0);  Cin, sign : in std_logic;  
         S : out std_logic_vector (31 downto 0);  Cout_BAR : out std_logic);

end p4add_N32_logN5_1;

architecture SYN_STRUCTURAL of p4add_N32_logN5_1 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component sum_gen_N32_1
      port( A, B : in std_logic_vector (31 downto 0);  Cin : in 
            std_logic_vector (8 downto 0);  S : out std_logic_vector (31 downto
            0));
   end component;
   
   component carry_tree_N32_logN5_1
      port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  
            Cout_7_BAR, Cout_6_port, Cout_5_port, Cout_4_port, Cout_3_port, 
            Cout_2_port, Cout_1_port, Cout_0_port : out std_logic);
   end component;
   
   component xor_gen_N32_1
      port( A : in std_logic_vector (31 downto 0);  B : in std_logic;  S : out 
            std_logic_vector (31 downto 0));
   end component;
   
   signal new_B_31_port, new_B_30_port, new_B_29_port, new_B_28_port, 
      new_B_27_port, new_B_26_port, new_B_25_port, new_B_24_port, new_B_23_port
      , new_B_22_port, new_B_21_port, new_B_20_port, new_B_19_port, 
      new_B_18_port, new_B_17_port, new_B_16_port, new_B_15_port, new_B_14_port
      , new_B_13_port, new_B_12_port, new_B_11_port, new_B_10_port, 
      new_B_9_port, new_B_8_port, new_B_7_port, new_B_6_port, new_B_5_port, 
      new_B_4_port, new_B_3_port, new_B_2_port, new_B_0_port, carry_pro_7_port,
      carry_pro_6_port, carry_pro_5_port, carry_pro_4_port, carry_pro_3_port, 
      carry_pro_2_port, carry_pro_1_port, n1, n3, n4, n5, n6, n7, n8, n9, n10, 
      n11, n12, n13, n14 : std_logic;

begin
   
   xor32 : xor_gen_N32_1 port map( A(31) => B(31), A(30) => B(30), A(29) => 
                           B(29), A(28) => B(28), A(27) => B(27), A(26) => 
                           B(26), A(25) => B(25), A(24) => B(24), A(23) => 
                           B(23), A(22) => B(22), A(21) => B(21), A(20) => 
                           B(20), A(19) => B(19), A(18) => B(18), A(17) => 
                           B(17), A(16) => B(16), A(15) => B(15), A(14) => 
                           B(14), A(13) => B(13), A(12) => B(12), A(11) => 
                           B(11), A(10) => B(10), A(9) => B(9), A(8) => B(8), 
                           A(7) => B(7), A(6) => B(6), A(5) => B(5), A(4) => 
                           B(4), A(3) => B(3), A(2) => B(2), A(1) => B(1), A(0)
                           => B(0), B => sign, S(31) => new_B_31_port, S(30) =>
                           new_B_30_port, S(29) => new_B_29_port, S(28) => 
                           new_B_28_port, S(27) => new_B_27_port, S(26) => 
                           new_B_26_port, S(25) => new_B_25_port, S(24) => 
                           new_B_24_port, S(23) => new_B_23_port, S(22) => 
                           new_B_22_port, S(21) => new_B_21_port, S(20) => 
                           new_B_20_port, S(19) => new_B_19_port, S(18) => 
                           new_B_18_port, S(17) => new_B_17_port, S(16) => 
                           new_B_16_port, S(15) => new_B_15_port, S(14) => 
                           new_B_14_port, S(13) => new_B_13_port, S(12) => 
                           new_B_12_port, S(11) => new_B_11_port, S(10) => 
                           new_B_10_port, S(9) => new_B_9_port, S(8) => 
                           new_B_8_port, S(7) => new_B_7_port, S(6) => 
                           new_B_6_port, S(5) => new_B_5_port, S(4) => 
                           new_B_4_port, S(3) => new_B_3_port, S(2) => 
                           new_B_2_port, S(1) => n1, S(0) => new_B_0_port);
   ct : carry_tree_N32_logN5_1 port map( A(31) => A(31), A(30) => A(30), A(29) 
                           => A(29), A(28) => A(28), A(27) => A(27), A(26) => 
                           A(26), A(25) => A(25), A(24) => A(24), A(23) => 
                           A(23), A(22) => A(22), A(21) => A(21), A(20) => 
                           A(20), A(19) => A(19), A(18) => A(18), A(17) => 
                           A(17), A(16) => A(16), A(15) => A(15), A(14) => 
                           A(14), A(13) => A(13), A(12) => A(12), A(11) => 
                           A(11), A(10) => A(10), A(9) => A(9), A(8) => A(8), 
                           A(7) => A(7), A(6) => A(6), A(5) => A(5), A(4) => 
                           A(4), A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(31) => new_B_31_port, B(30) => 
                           new_B_30_port, B(29) => new_B_29_port, B(28) => 
                           new_B_28_port, B(27) => new_B_27_port, B(26) => 
                           new_B_26_port, B(25) => new_B_25_port, B(24) => 
                           new_B_24_port, B(23) => new_B_23_port, B(22) => 
                           new_B_22_port, B(21) => new_B_21_port, B(20) => 
                           new_B_20_port, B(19) => new_B_19_port, B(18) => 
                           new_B_18_port, B(17) => new_B_17_port, B(16) => 
                           new_B_16_port, B(15) => new_B_15_port, B(14) => 
                           new_B_14_port, B(13) => new_B_13_port, B(12) => 
                           new_B_12_port, B(11) => new_B_11_port, B(10) => 
                           new_B_10_port, B(9) => new_B_9_port, B(8) => 
                           new_B_8_port, B(7) => new_B_7_port, B(6) => 
                           new_B_6_port, B(5) => new_B_5_port, B(4) => 
                           new_B_4_port, B(3) => new_B_3_port, B(2) => 
                           new_B_2_port, B(1) => n1, B(0) => new_B_0_port, Cin 
                           => sign, Cout_7_BAR => Cout_BAR, Cout_6_port => 
                           carry_pro_7_port, Cout_5_port => carry_pro_6_port, 
                           Cout_4_port => carry_pro_5_port, Cout_3_port => 
                           carry_pro_4_port, Cout_2_port => carry_pro_3_port, 
                           Cout_1_port => carry_pro_2_port, Cout_0_port => 
                           carry_pro_1_port);
   add : sum_gen_N32_1 port map( A(31) => A(31), A(30) => A(30), A(29) => A(29)
                           , A(28) => A(28), A(27) => A(27), A(26) => A(26), 
                           A(25) => A(25), A(24) => A(24), A(23) => A(23), 
                           A(22) => A(22), A(21) => A(21), A(20) => A(20), 
                           A(19) => A(19), A(18) => A(18), A(17) => A(17), 
                           A(16) => A(16), A(15) => A(15), A(14) => A(14), 
                           A(13) => A(13), A(12) => A(12), A(11) => A(11), 
                           A(10) => A(10), A(9) => A(9), A(8) => A(8), A(7) => 
                           A(7), A(6) => A(6), A(5) => A(5), A(4) => A(4), A(3)
                           => A(3), A(2) => A(2), A(1) => A(1), A(0) => A(0), 
                           B(31) => new_B_31_port, B(30) => new_B_30_port, 
                           B(29) => new_B_29_port, B(28) => new_B_28_port, 
                           B(27) => new_B_27_port, B(26) => new_B_26_port, 
                           B(25) => new_B_25_port, B(24) => new_B_24_port, 
                           B(23) => n6, B(22) => new_B_22_port, B(21) => n3, 
                           B(20) => new_B_20_port, B(19) => new_B_19_port, 
                           B(18) => new_B_18_port, B(17) => n9, B(16) => 
                           new_B_16_port, B(15) => n5, B(14) => new_B_14_port, 
                           B(13) => n13, B(12) => n7, B(11) => new_B_11_port, 
                           B(10) => n8, B(9) => n11, B(8) => new_B_8_port, B(7)
                           => new_B_7_port, B(6) => n4, B(5) => n12, B(4) => 
                           new_B_4_port, B(3) => new_B_3_port, B(2) => 
                           new_B_2_port, B(1) => n1, B(0) => n10, Cin(8) => n14
                           , Cin(7) => carry_pro_7_port, Cin(6) => 
                           carry_pro_6_port, Cin(5) => carry_pro_5_port, Cin(4)
                           => carry_pro_4_port, Cin(3) => carry_pro_3_port, 
                           Cin(2) => carry_pro_2_port, Cin(1) => 
                           carry_pro_1_port, Cin(0) => sign, S(31) => S(31), 
                           S(30) => S(30), S(29) => S(29), S(28) => S(28), 
                           S(27) => S(27), S(26) => S(26), S(25) => S(25), 
                           S(24) => S(24), S(23) => S(23), S(22) => S(22), 
                           S(21) => S(21), S(20) => S(20), S(19) => S(19), 
                           S(18) => S(18), S(17) => S(17), S(16) => S(16), 
                           S(15) => S(15), S(14) => S(14), S(13) => S(13), 
                           S(12) => S(12), S(11) => S(11), S(10) => S(10), S(9)
                           => S(9), S(8) => S(8), S(7) => S(7), S(6) => S(6), 
                           S(5) => S(5), S(4) => S(4), S(3) => S(3), S(2) => 
                           S(2), S(1) => S(1), S(0) => S(0));
   U1 : BUF_X1 port map( A => new_B_12_port, Z => n7);
   U2 : BUF_X1 port map( A => new_B_9_port, Z => n11);
   U3 : BUF_X1 port map( A => new_B_17_port, Z => n9);
   U4 : BUF_X1 port map( A => new_B_15_port, Z => n5);
   U5 : BUF_X1 port map( A => new_B_5_port, Z => n12);
   U6 : BUF_X1 port map( A => new_B_21_port, Z => n3);
   U7 : BUF_X1 port map( A => new_B_6_port, Z => n4);
   U8 : CLKBUF_X1 port map( A => new_B_23_port, Z => n6);
   U9 : CLKBUF_X1 port map( A => new_B_13_port, Z => n13);
   U10 : CLKBUF_X1 port map( A => new_B_0_port, Z => n10);
   U11 : CLKBUF_X1 port map( A => new_B_10_port, Z => n8);
   n14 <= '0';

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity predictor_2_15 is

   port( clock, reset, enable, taken_i : in std_logic;  prediction_o : out 
         std_logic);

end predictor_2_15;

architecture SYN_bhe of predictor_2_15 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal prediction_o_port, next_STATE_1_port, next_STATE_0_port, N11, N12, n1
      , n2, n5, n7, n8, n9, n10, net48732 : std_logic;

begin
   prediction_o <= prediction_o_port;
   
   next_STATE_reg_0_inst : DLH_X1 port map( G => enable, D => N11, Q => 
                           next_STATE_0_port);
   STATE_reg_0_inst : DFFR_X1 port map( D => n7, CK => clock, RN => n2, Q => n1
                           , QN => n5);
   next_STATE_reg_1_inst : DLH_X1 port map( G => enable, D => N12, Q => 
                           next_STATE_1_port);
   STATE_reg_1_inst : DFFR_X1 port map( D => n8, CK => clock, RN => n2, Q => 
                           prediction_o_port, QN => net48732);
   U2 : MUX2_X1 port map( A => prediction_o_port, B => next_STATE_1_port, S => 
                           enable, Z => n8);
   U4 : MUX2_X1 port map( A => n1, B => next_STATE_0_port, S => enable, Z => n7
                           );
   U9 : NOR2_X1 port map( A1 => prediction_o_port, A2 => taken_i, ZN => n10);
   U7 : NAND2_X1 port map( A1 => prediction_o_port, A2 => taken_i, ZN => n9);
   U6 : OAI21_X1 port map( B1 => n10, B2 => n1, A => n9, ZN => N11);
   U5 : OAI21_X1 port map( B1 => n5, B2 => n10, A => n9, ZN => N12);
   U3 : INV_X1 port map( A => reset, ZN => n2);

end SYN_bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity predictor_2_14 is

   port( clock, reset, enable, taken_i : in std_logic;  prediction_o : out 
         std_logic);

end predictor_2_14;

architecture SYN_bhe of predictor_2_14 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal prediction_o_port, next_STATE_1_port, next_STATE_0_port, N11, N12, n1
      , n2, n5, n7, n8, n9, n10, net48731 : std_logic;

begin
   prediction_o <= prediction_o_port;
   
   next_STATE_reg_0_inst : DLH_X1 port map( G => enable, D => N11, Q => 
                           next_STATE_0_port);
   STATE_reg_0_inst : DFFR_X1 port map( D => n7, CK => clock, RN => n2, Q => n1
                           , QN => n5);
   next_STATE_reg_1_inst : DLH_X1 port map( G => enable, D => N12, Q => 
                           next_STATE_1_port);
   STATE_reg_1_inst : DFFR_X1 port map( D => n8, CK => clock, RN => n2, Q => 
                           prediction_o_port, QN => net48731);
   U2 : MUX2_X1 port map( A => prediction_o_port, B => next_STATE_1_port, S => 
                           enable, Z => n8);
   U4 : MUX2_X1 port map( A => n1, B => next_STATE_0_port, S => enable, Z => n7
                           );
   U9 : NOR2_X1 port map( A1 => prediction_o_port, A2 => taken_i, ZN => n10);
   U7 : NAND2_X1 port map( A1 => prediction_o_port, A2 => taken_i, ZN => n9);
   U6 : OAI21_X1 port map( B1 => n10, B2 => n1, A => n9, ZN => N11);
   U5 : OAI21_X1 port map( B1 => n5, B2 => n10, A => n9, ZN => N12);
   U3 : INV_X1 port map( A => reset, ZN => n2);

end SYN_bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity predictor_2_13 is

   port( clock, reset, enable, taken_i : in std_logic;  prediction_o : out 
         std_logic);

end predictor_2_13;

architecture SYN_bhe of predictor_2_13 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal prediction_o_port, next_STATE_1_port, next_STATE_0_port, N11, N12, n1
      , n2, n5, n7, n8, n9, n10, net48730 : std_logic;

begin
   prediction_o <= prediction_o_port;
   
   next_STATE_reg_0_inst : DLH_X1 port map( G => enable, D => N11, Q => 
                           next_STATE_0_port);
   STATE_reg_0_inst : DFFR_X1 port map( D => n7, CK => clock, RN => n2, Q => n1
                           , QN => n5);
   next_STATE_reg_1_inst : DLH_X1 port map( G => enable, D => N12, Q => 
                           next_STATE_1_port);
   STATE_reg_1_inst : DFFR_X1 port map( D => n8, CK => clock, RN => n2, Q => 
                           prediction_o_port, QN => net48730);
   U2 : MUX2_X1 port map( A => prediction_o_port, B => next_STATE_1_port, S => 
                           enable, Z => n8);
   U4 : MUX2_X1 port map( A => n1, B => next_STATE_0_port, S => enable, Z => n7
                           );
   U9 : NOR2_X1 port map( A1 => prediction_o_port, A2 => taken_i, ZN => n10);
   U7 : NAND2_X1 port map( A1 => prediction_o_port, A2 => taken_i, ZN => n9);
   U5 : OAI21_X1 port map( B1 => n5, B2 => n10, A => n9, ZN => N12);
   U6 : OAI21_X1 port map( B1 => n10, B2 => n1, A => n9, ZN => N11);
   U3 : INV_X1 port map( A => reset, ZN => n2);

end SYN_bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity predictor_2_12 is

   port( clock, reset, enable, taken_i : in std_logic;  prediction_o : out 
         std_logic);

end predictor_2_12;

architecture SYN_bhe of predictor_2_12 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal prediction_o_port, next_STATE_1_port, next_STATE_0_port, N11, N12, n1
      , n2, n5, n7, n8, n9, n10, net48729 : std_logic;

begin
   prediction_o <= prediction_o_port;
   
   next_STATE_reg_0_inst : DLH_X1 port map( G => enable, D => N11, Q => 
                           next_STATE_0_port);
   STATE_reg_0_inst : DFFR_X1 port map( D => n7, CK => clock, RN => n2, Q => n1
                           , QN => n5);
   next_STATE_reg_1_inst : DLH_X1 port map( G => enable, D => N12, Q => 
                           next_STATE_1_port);
   STATE_reg_1_inst : DFFR_X1 port map( D => n8, CK => clock, RN => n2, Q => 
                           prediction_o_port, QN => net48729);
   U2 : MUX2_X1 port map( A => prediction_o_port, B => next_STATE_1_port, S => 
                           enable, Z => n8);
   U4 : MUX2_X1 port map( A => n1, B => next_STATE_0_port, S => enable, Z => n7
                           );
   U9 : NOR2_X1 port map( A1 => prediction_o_port, A2 => taken_i, ZN => n10);
   U7 : NAND2_X1 port map( A1 => prediction_o_port, A2 => taken_i, ZN => n9);
   U5 : OAI21_X1 port map( B1 => n5, B2 => n10, A => n9, ZN => N12);
   U6 : OAI21_X1 port map( B1 => n10, B2 => n1, A => n9, ZN => N11);
   U3 : INV_X1 port map( A => reset, ZN => n2);

end SYN_bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity predictor_2_11 is

   port( clock, reset, enable, taken_i : in std_logic;  prediction_o : out 
         std_logic);

end predictor_2_11;

architecture SYN_bhe of predictor_2_11 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal prediction_o_port, next_STATE_1_port, next_STATE_0_port, N11, N12, n1
      , n2, n5, n7, n8, n9, n10, net48728 : std_logic;

begin
   prediction_o <= prediction_o_port;
   
   next_STATE_reg_0_inst : DLH_X1 port map( G => enable, D => N11, Q => 
                           next_STATE_0_port);
   STATE_reg_0_inst : DFFR_X1 port map( D => n7, CK => clock, RN => n2, Q => n1
                           , QN => n5);
   next_STATE_reg_1_inst : DLH_X1 port map( G => enable, D => N12, Q => 
                           next_STATE_1_port);
   STATE_reg_1_inst : DFFR_X1 port map( D => n8, CK => clock, RN => n2, Q => 
                           prediction_o_port, QN => net48728);
   U2 : MUX2_X1 port map( A => prediction_o_port, B => next_STATE_1_port, S => 
                           enable, Z => n8);
   U4 : MUX2_X1 port map( A => n1, B => next_STATE_0_port, S => enable, Z => n7
                           );
   U9 : NOR2_X1 port map( A1 => prediction_o_port, A2 => taken_i, ZN => n10);
   U7 : NAND2_X1 port map( A1 => prediction_o_port, A2 => taken_i, ZN => n9);
   U5 : OAI21_X1 port map( B1 => n5, B2 => n10, A => n9, ZN => N12);
   U6 : OAI21_X1 port map( B1 => n10, B2 => n1, A => n9, ZN => N11);
   U3 : INV_X1 port map( A => reset, ZN => n2);

end SYN_bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity predictor_2_10 is

   port( clock, reset, enable, taken_i : in std_logic;  prediction_o : out 
         std_logic);

end predictor_2_10;

architecture SYN_bhe of predictor_2_10 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal prediction_o_port, next_STATE_1_port, next_STATE_0_port, N11, N12, n1
      , n2, n5, n7, n8, n9, n10, net48727 : std_logic;

begin
   prediction_o <= prediction_o_port;
   
   next_STATE_reg_0_inst : DLH_X1 port map( G => enable, D => N11, Q => 
                           next_STATE_0_port);
   STATE_reg_0_inst : DFFR_X1 port map( D => n7, CK => clock, RN => n2, Q => n1
                           , QN => n5);
   next_STATE_reg_1_inst : DLH_X1 port map( G => enable, D => N12, Q => 
                           next_STATE_1_port);
   STATE_reg_1_inst : DFFR_X1 port map( D => n8, CK => clock, RN => n2, Q => 
                           prediction_o_port, QN => net48727);
   U2 : MUX2_X1 port map( A => prediction_o_port, B => next_STATE_1_port, S => 
                           enable, Z => n8);
   U4 : MUX2_X1 port map( A => n1, B => next_STATE_0_port, S => enable, Z => n7
                           );
   U9 : NOR2_X1 port map( A1 => prediction_o_port, A2 => taken_i, ZN => n10);
   U7 : NAND2_X1 port map( A1 => prediction_o_port, A2 => taken_i, ZN => n9);
   U6 : OAI21_X1 port map( B1 => n10, B2 => n1, A => n9, ZN => N11);
   U5 : OAI21_X1 port map( B1 => n5, B2 => n10, A => n9, ZN => N12);
   U3 : INV_X1 port map( A => reset, ZN => n2);

end SYN_bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity predictor_2_9 is

   port( clock, reset, enable, taken_i : in std_logic;  prediction_o : out 
         std_logic);

end predictor_2_9;

architecture SYN_bhe of predictor_2_9 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal prediction_o_port, next_STATE_1_port, next_STATE_0_port, N11, N12, n1
      , n2, n5, n7, n8, n9, n10, net48726 : std_logic;

begin
   prediction_o <= prediction_o_port;
   
   next_STATE_reg_0_inst : DLH_X1 port map( G => enable, D => N11, Q => 
                           next_STATE_0_port);
   STATE_reg_0_inst : DFFR_X1 port map( D => n7, CK => clock, RN => n2, Q => n1
                           , QN => n5);
   next_STATE_reg_1_inst : DLH_X1 port map( G => enable, D => N12, Q => 
                           next_STATE_1_port);
   STATE_reg_1_inst : DFFR_X1 port map( D => n8, CK => clock, RN => n2, Q => 
                           prediction_o_port, QN => net48726);
   U2 : MUX2_X1 port map( A => prediction_o_port, B => next_STATE_1_port, S => 
                           enable, Z => n8);
   U4 : MUX2_X1 port map( A => n1, B => next_STATE_0_port, S => enable, Z => n7
                           );
   U9 : NOR2_X1 port map( A1 => prediction_o_port, A2 => taken_i, ZN => n10);
   U7 : NAND2_X1 port map( A1 => prediction_o_port, A2 => taken_i, ZN => n9);
   U6 : OAI21_X1 port map( B1 => n10, B2 => n1, A => n9, ZN => N11);
   U5 : OAI21_X1 port map( B1 => n5, B2 => n10, A => n9, ZN => N12);
   U3 : INV_X1 port map( A => reset, ZN => n2);

end SYN_bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity predictor_2_8 is

   port( clock, reset, enable, taken_i : in std_logic;  prediction_o : out 
         std_logic);

end predictor_2_8;

architecture SYN_bhe of predictor_2_8 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal prediction_o_port, next_STATE_1_port, next_STATE_0_port, N11, N12, n1
      , n2, n5, n7, n8, n9, n10, net48725 : std_logic;

begin
   prediction_o <= prediction_o_port;
   
   next_STATE_reg_0_inst : DLH_X1 port map( G => enable, D => N11, Q => 
                           next_STATE_0_port);
   STATE_reg_0_inst : DFFR_X1 port map( D => n7, CK => clock, RN => n2, Q => n1
                           , QN => n5);
   next_STATE_reg_1_inst : DLH_X1 port map( G => enable, D => N12, Q => 
                           next_STATE_1_port);
   STATE_reg_1_inst : DFFR_X1 port map( D => n8, CK => clock, RN => n2, Q => 
                           prediction_o_port, QN => net48725);
   U2 : MUX2_X1 port map( A => prediction_o_port, B => next_STATE_1_port, S => 
                           enable, Z => n8);
   U4 : MUX2_X1 port map( A => n1, B => next_STATE_0_port, S => enable, Z => n7
                           );
   U9 : NOR2_X1 port map( A1 => prediction_o_port, A2 => taken_i, ZN => n10);
   U7 : NAND2_X1 port map( A1 => prediction_o_port, A2 => taken_i, ZN => n9);
   U5 : OAI21_X1 port map( B1 => n5, B2 => n10, A => n9, ZN => N12);
   U6 : OAI21_X1 port map( B1 => n10, B2 => n1, A => n9, ZN => N11);
   U3 : INV_X1 port map( A => reset, ZN => n2);

end SYN_bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity predictor_2_7 is

   port( clock, reset, enable, taken_i : in std_logic;  prediction_o : out 
         std_logic);

end predictor_2_7;

architecture SYN_bhe of predictor_2_7 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal prediction_o_port, next_STATE_1_port, next_STATE_0_port, N11, N12, n1
      , n2, n5, n7, n8, n9, n10, net48724 : std_logic;

begin
   prediction_o <= prediction_o_port;
   
   next_STATE_reg_0_inst : DLH_X1 port map( G => enable, D => N11, Q => 
                           next_STATE_0_port);
   STATE_reg_0_inst : DFFR_X1 port map( D => n7, CK => clock, RN => n2, Q => n1
                           , QN => n5);
   next_STATE_reg_1_inst : DLH_X1 port map( G => enable, D => N12, Q => 
                           next_STATE_1_port);
   STATE_reg_1_inst : DFFR_X1 port map( D => n8, CK => clock, RN => n2, Q => 
                           prediction_o_port, QN => net48724);
   U2 : MUX2_X1 port map( A => prediction_o_port, B => next_STATE_1_port, S => 
                           enable, Z => n8);
   U4 : MUX2_X1 port map( A => n1, B => next_STATE_0_port, S => enable, Z => n7
                           );
   U9 : NOR2_X1 port map( A1 => prediction_o_port, A2 => taken_i, ZN => n10);
   U7 : NAND2_X1 port map( A1 => prediction_o_port, A2 => taken_i, ZN => n9);
   U6 : OAI21_X1 port map( B1 => n10, B2 => n1, A => n9, ZN => N11);
   U5 : OAI21_X1 port map( B1 => n5, B2 => n10, A => n9, ZN => N12);
   U3 : INV_X1 port map( A => reset, ZN => n2);

end SYN_bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity predictor_2_6 is

   port( clock, reset, enable, taken_i : in std_logic;  prediction_o : out 
         std_logic);

end predictor_2_6;

architecture SYN_bhe of predictor_2_6 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal prediction_o_port, next_STATE_1_port, next_STATE_0_port, N11, N12, n1
      , n2, n5, n7, n8, n9, n10, net48723 : std_logic;

begin
   prediction_o <= prediction_o_port;
   
   next_STATE_reg_0_inst : DLH_X1 port map( G => enable, D => N11, Q => 
                           next_STATE_0_port);
   STATE_reg_0_inst : DFFR_X1 port map( D => n7, CK => clock, RN => n2, Q => n1
                           , QN => n5);
   next_STATE_reg_1_inst : DLH_X1 port map( G => enable, D => N12, Q => 
                           next_STATE_1_port);
   STATE_reg_1_inst : DFFR_X1 port map( D => n8, CK => clock, RN => n2, Q => 
                           prediction_o_port, QN => net48723);
   U2 : MUX2_X1 port map( A => prediction_o_port, B => next_STATE_1_port, S => 
                           enable, Z => n8);
   U4 : MUX2_X1 port map( A => n1, B => next_STATE_0_port, S => enable, Z => n7
                           );
   U9 : NOR2_X1 port map( A1 => prediction_o_port, A2 => taken_i, ZN => n10);
   U7 : NAND2_X1 port map( A1 => prediction_o_port, A2 => taken_i, ZN => n9);
   U5 : OAI21_X1 port map( B1 => n5, B2 => n10, A => n9, ZN => N12);
   U6 : OAI21_X1 port map( B1 => n10, B2 => n1, A => n9, ZN => N11);
   U3 : INV_X1 port map( A => reset, ZN => n2);

end SYN_bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity predictor_2_5 is

   port( clock, reset, enable, taken_i : in std_logic;  prediction_o : out 
         std_logic);

end predictor_2_5;

architecture SYN_bhe of predictor_2_5 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal prediction_o_port, next_STATE_1_port, next_STATE_0_port, N11, N12, n1
      , n2, n5, n7, n8, n9, n10, net48722 : std_logic;

begin
   prediction_o <= prediction_o_port;
   
   next_STATE_reg_0_inst : DLH_X1 port map( G => enable, D => N11, Q => 
                           next_STATE_0_port);
   STATE_reg_0_inst : DFFR_X1 port map( D => n7, CK => clock, RN => n2, Q => n1
                           , QN => n5);
   next_STATE_reg_1_inst : DLH_X1 port map( G => enable, D => N12, Q => 
                           next_STATE_1_port);
   STATE_reg_1_inst : DFFR_X1 port map( D => n8, CK => clock, RN => n2, Q => 
                           prediction_o_port, QN => net48722);
   U2 : MUX2_X1 port map( A => prediction_o_port, B => next_STATE_1_port, S => 
                           enable, Z => n8);
   U4 : MUX2_X1 port map( A => n1, B => next_STATE_0_port, S => enable, Z => n7
                           );
   U9 : NOR2_X1 port map( A1 => prediction_o_port, A2 => taken_i, ZN => n10);
   U7 : NAND2_X1 port map( A1 => prediction_o_port, A2 => taken_i, ZN => n9);
   U5 : OAI21_X1 port map( B1 => n5, B2 => n10, A => n9, ZN => N12);
   U6 : OAI21_X1 port map( B1 => n10, B2 => n1, A => n9, ZN => N11);
   U3 : INV_X1 port map( A => reset, ZN => n2);

end SYN_bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity predictor_2_4 is

   port( clock, reset, enable, taken_i : in std_logic;  prediction_o : out 
         std_logic);

end predictor_2_4;

architecture SYN_bhe of predictor_2_4 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal prediction_o_port, next_STATE_1_port, next_STATE_0_port, N11, N12, n1
      , n2, n5, n7, n8, n9, n10, net48721 : std_logic;

begin
   prediction_o <= prediction_o_port;
   
   next_STATE_reg_0_inst : DLH_X1 port map( G => enable, D => N11, Q => 
                           next_STATE_0_port);
   STATE_reg_0_inst : DFFR_X1 port map( D => n7, CK => clock, RN => n2, Q => n1
                           , QN => n5);
   next_STATE_reg_1_inst : DLH_X1 port map( G => enable, D => N12, Q => 
                           next_STATE_1_port);
   STATE_reg_1_inst : DFFR_X1 port map( D => n8, CK => clock, RN => n2, Q => 
                           prediction_o_port, QN => net48721);
   U2 : MUX2_X1 port map( A => prediction_o_port, B => next_STATE_1_port, S => 
                           enable, Z => n8);
   U4 : MUX2_X1 port map( A => n1, B => next_STATE_0_port, S => enable, Z => n7
                           );
   U9 : NOR2_X1 port map( A1 => prediction_o_port, A2 => taken_i, ZN => n10);
   U7 : NAND2_X1 port map( A1 => prediction_o_port, A2 => taken_i, ZN => n9);
   U5 : OAI21_X1 port map( B1 => n5, B2 => n10, A => n9, ZN => N12);
   U6 : OAI21_X1 port map( B1 => n10, B2 => n1, A => n9, ZN => N11);
   U3 : INV_X1 port map( A => reset, ZN => n2);

end SYN_bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity predictor_2_3 is

   port( clock, reset, enable, taken_i : in std_logic;  prediction_o : out 
         std_logic);

end predictor_2_3;

architecture SYN_bhe of predictor_2_3 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal prediction_o_port, next_STATE_1_port, next_STATE_0_port, N11, N12, n1
      , n2, n5, n7, n8, n9, n10, net48720 : std_logic;

begin
   prediction_o <= prediction_o_port;
   
   next_STATE_reg_0_inst : DLH_X1 port map( G => enable, D => N11, Q => 
                           next_STATE_0_port);
   STATE_reg_0_inst : DFFR_X1 port map( D => n7, CK => clock, RN => n2, Q => n1
                           , QN => n5);
   next_STATE_reg_1_inst : DLH_X1 port map( G => enable, D => N12, Q => 
                           next_STATE_1_port);
   STATE_reg_1_inst : DFFR_X1 port map( D => n8, CK => clock, RN => n2, Q => 
                           prediction_o_port, QN => net48720);
   U2 : MUX2_X1 port map( A => prediction_o_port, B => next_STATE_1_port, S => 
                           enable, Z => n8);
   U4 : MUX2_X1 port map( A => n1, B => next_STATE_0_port, S => enable, Z => n7
                           );
   U9 : NOR2_X1 port map( A1 => prediction_o_port, A2 => taken_i, ZN => n10);
   U7 : NAND2_X1 port map( A1 => prediction_o_port, A2 => taken_i, ZN => n9);
   U6 : OAI21_X1 port map( B1 => n10, B2 => n1, A => n9, ZN => N11);
   U5 : OAI21_X1 port map( B1 => n5, B2 => n10, A => n9, ZN => N12);
   U3 : INV_X1 port map( A => reset, ZN => n2);

end SYN_bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity predictor_2_2 is

   port( clock, reset, enable, taken_i : in std_logic;  prediction_o : out 
         std_logic);

end predictor_2_2;

architecture SYN_bhe of predictor_2_2 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal prediction_o_port, next_STATE_1_port, next_STATE_0_port, N11, N12, n1
      , n2, n5, n7, n8, n9, n10, net48719 : std_logic;

begin
   prediction_o <= prediction_o_port;
   
   next_STATE_reg_0_inst : DLH_X1 port map( G => enable, D => N11, Q => 
                           next_STATE_0_port);
   STATE_reg_0_inst : DFFR_X1 port map( D => n7, CK => clock, RN => n2, Q => n1
                           , QN => n5);
   next_STATE_reg_1_inst : DLH_X1 port map( G => enable, D => N12, Q => 
                           next_STATE_1_port);
   STATE_reg_1_inst : DFFR_X1 port map( D => n8, CK => clock, RN => n2, Q => 
                           prediction_o_port, QN => net48719);
   U2 : MUX2_X1 port map( A => prediction_o_port, B => next_STATE_1_port, S => 
                           enable, Z => n8);
   U4 : MUX2_X1 port map( A => n1, B => next_STATE_0_port, S => enable, Z => n7
                           );
   U9 : NOR2_X1 port map( A1 => prediction_o_port, A2 => taken_i, ZN => n10);
   U7 : NAND2_X1 port map( A1 => prediction_o_port, A2 => taken_i, ZN => n9);
   U6 : OAI21_X1 port map( B1 => n10, B2 => n1, A => n9, ZN => N11);
   U5 : OAI21_X1 port map( B1 => n5, B2 => n10, A => n9, ZN => N12);
   U3 : INV_X1 port map( A => reset, ZN => n2);

end SYN_bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity predictor_2_1 is

   port( clock, reset, enable, taken_i : in std_logic;  prediction_o : out 
         std_logic);

end predictor_2_1;

architecture SYN_bhe of predictor_2_1 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal prediction_o_port, next_STATE_1_port, next_STATE_0_port, N11, N12, n1
      , n2, n5, n7, n8, n9, n10, net48718 : std_logic;

begin
   prediction_o <= prediction_o_port;
   
   next_STATE_reg_0_inst : DLH_X1 port map( G => enable, D => N11, Q => 
                           next_STATE_0_port);
   STATE_reg_0_inst : DFFR_X1 port map( D => n7, CK => clock, RN => n2, Q => n1
                           , QN => n5);
   next_STATE_reg_1_inst : DLH_X1 port map( G => enable, D => N12, Q => 
                           next_STATE_1_port);
   STATE_reg_1_inst : DFFR_X1 port map( D => n8, CK => clock, RN => n2, Q => 
                           prediction_o_port, QN => net48718);
   U2 : MUX2_X1 port map( A => prediction_o_port, B => next_STATE_1_port, S => 
                           enable, Z => n8);
   U4 : MUX2_X1 port map( A => n1, B => next_STATE_0_port, S => enable, Z => n7
                           );
   U9 : NOR2_X1 port map( A1 => prediction_o_port, A2 => taken_i, ZN => n10);
   U7 : NAND2_X1 port map( A1 => prediction_o_port, A2 => taken_i, ZN => n9);
   U6 : OAI21_X1 port map( B1 => n10, B2 => n1, A => n9, ZN => N11);
   U5 : OAI21_X1 port map( B1 => n5, B2 => n10, A => n9, ZN => N12);
   U3 : INV_X1 port map( A => reset, ZN => n2);

end SYN_bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity mux41_1 is

   port( IN0, IN1, IN2, IN3 : in std_logic_vector (31 downto 0);  CTRL : in 
         std_logic_vector (1 downto 0);  OUT1 : out std_logic_vector (31 downto
         0));

end mux41_1;

architecture SYN_bhe of mux41_1 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X3
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n6, n7, n8, n21, n22, n23, n24, n27, n28, n29, n30, n39, n40, n71
      , n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, 
      n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, 
      n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, 
      n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, 
      n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, 
      n136, n137, n138 : std_logic;

begin
   
   U1 : AOI22_X1 port map( A1 => IN1(28), A2 => n71, B1 => IN0(28), B2 => n73, 
                           ZN => n1);
   U2 : NAND2_X1 port map( A1 => n8, A2 => n1, ZN => OUT1(28));
   U3 : BUF_X2 port map( A => n83, Z => n73);
   U4 : BUF_X2 port map( A => n83, Z => n74);
   U5 : BUF_X2 port map( A => n82, Z => n71);
   U6 : CLKBUF_X3 port map( A => n83, Z => n75);
   U7 : CLKBUF_X3 port map( A => n82, Z => n72);
   U8 : BUF_X2 port map( A => n82, Z => n40);
   U9 : BUF_X2 port map( A => n84, Z => n78);
   U10 : BUF_X2 port map( A => n6, Z => n79);
   U11 : BUF_X2 port map( A => n6, Z => n80);
   U12 : BUF_X2 port map( A => n6, Z => n7);
   U13 : BUF_X2 port map( A => n84, Z => n76);
   U14 : BUF_X2 port map( A => n84, Z => n77);
   U15 : AND2_X1 port map( A1 => CTRL(1), A2 => n81, ZN => n6);
   U16 : AND2_X1 port map( A1 => CTRL(1), A2 => CTRL(0), ZN => n84);
   U17 : INV_X1 port map( A => CTRL(0), ZN => n81);
   U18 : AOI22_X1 port map( A1 => n77, A2 => IN3(23), B1 => n79, B2 => IN2(23),
                           ZN => n23);
   U19 : AOI22_X1 port map( A1 => n80, A2 => IN2(30), B1 => n78, B2 => IN3(30),
                           ZN => n28);
   U20 : AOI22_X1 port map( A1 => n76, A2 => IN3(10), B1 => n80, B2 => IN2(10),
                           ZN => n87);
   U21 : AOI22_X1 port map( A1 => n76, A2 => IN3(17), B1 => n79, B2 => IN2(17),
                           ZN => n101);
   U22 : AOI22_X1 port map( A1 => n77, A2 => IN3(4), B1 => n7, B2 => IN2(4), ZN
                           => n127);
   U23 : AOI22_X1 port map( A1 => n77, A2 => IN3(24), B1 => n80, B2 => IN2(24),
                           ZN => n115);
   U24 : AOI22_X1 port map( A1 => n77, A2 => IN3(21), B1 => n79, B2 => IN2(21),
                           ZN => n111);
   U25 : AOI22_X1 port map( A1 => n77, A2 => IN3(3), B1 => n79, B2 => IN2(3), 
                           ZN => n125);
   U26 : AOI22_X1 port map( A1 => n78, A2 => IN3(9), B1 => n79, B2 => IN2(9), 
                           ZN => n137);
   U27 : AOI22_X1 port map( A1 => n76, A2 => IN3(13), B1 => n80, B2 => IN2(13),
                           ZN => n93);
   U28 : AOI22_X1 port map( A1 => n76, A2 => IN3(14), B1 => n7, B2 => IN2(14), 
                           ZN => n95);
   U29 : NAND3_X1 port map( A1 => n23, A2 => n22, A3 => n21, ZN => OUT1(23));
   U30 : AOI22_X1 port map( A1 => n80, A2 => IN2(28), B1 => n78, B2 => IN3(28),
                           ZN => n8);
   U31 : NAND2_X1 port map( A1 => n74, A2 => IN0(23), ZN => n22);
   U32 : NAND2_X1 port map( A1 => n40, A2 => IN1(23), ZN => n21);
   U33 : NAND2_X1 port map( A1 => n27, A2 => n24, ZN => OUT1(29));
   U34 : NAND2_X1 port map( A1 => n29, A2 => n28, ZN => OUT1(30));
   U35 : NAND2_X1 port map( A1 => n39, A2 => n30, ZN => OUT1(31));
   U36 : NOR2_X1 port map( A1 => CTRL(1), A2 => CTRL(0), ZN => n83);
   U37 : AOI22_X1 port map( A1 => n72, A2 => IN1(29), B1 => n73, B2 => IN0(29),
                           ZN => n27);
   U38 : AOI22_X1 port map( A1 => n7, A2 => IN2(29), B1 => n78, B2 => IN3(29), 
                           ZN => n24);
   U39 : AOI22_X1 port map( A1 => n72, A2 => IN1(30), B1 => n74, B2 => IN0(30),
                           ZN => n29);
   U40 : AOI22_X1 port map( A1 => n71, A2 => IN1(31), B1 => n75, B2 => IN0(31),
                           ZN => n39);
   U41 : AOI22_X1 port map( A1 => n7, A2 => IN2(31), B1 => n78, B2 => IN3(31), 
                           ZN => n30);
   U42 : NAND2_X1 port map( A1 => n93, A2 => n94, ZN => OUT1(13));
   U43 : NAND2_X1 port map( A1 => n96, A2 => n95, ZN => OUT1(14));
   U44 : NAND2_X1 port map( A1 => n98, A2 => n97, ZN => OUT1(15));
   U45 : NAND2_X1 port map( A1 => n86, A2 => n85, ZN => OUT1(0));
   U46 : NAND2_X1 port map( A1 => n100, A2 => n99, ZN => OUT1(16));
   U47 : NAND2_X1 port map( A1 => n122, A2 => n121, ZN => OUT1(27));
   U48 : NAND2_X1 port map( A1 => n92, A2 => n91, ZN => OUT1(12));
   U49 : NAND2_X1 port map( A1 => n90, A2 => n89, ZN => OUT1(11));
   U50 : NAND2_X1 port map( A1 => n87, A2 => n88, ZN => OUT1(10));
   U51 : NAND2_X1 port map( A1 => n118, A2 => n117, ZN => OUT1(25));
   U52 : NAND2_X1 port map( A1 => n112, A2 => n111, ZN => OUT1(21));
   U53 : NAND2_X1 port map( A1 => n108, A2 => n107, ZN => OUT1(1));
   U54 : NAND2_X1 port map( A1 => n120, A2 => n119, ZN => OUT1(26));
   U55 : NAND2_X1 port map( A1 => n116, A2 => n115, ZN => OUT1(24));
   U56 : NAND2_X1 port map( A1 => n114, A2 => n113, ZN => OUT1(22));
   U57 : NAND2_X1 port map( A1 => n110, A2 => n109, ZN => OUT1(20));
   U58 : NAND2_X1 port map( A1 => n102, A2 => n101, ZN => OUT1(17));
   U59 : NAND2_X1 port map( A1 => n106, A2 => n105, ZN => OUT1(19));
   U60 : NAND2_X1 port map( A1 => n138, A2 => n137, ZN => OUT1(9));
   U61 : NAND2_X1 port map( A1 => n134, A2 => n133, ZN => OUT1(7));
   U62 : NAND2_X1 port map( A1 => n130, A2 => n129, ZN => OUT1(5));
   U63 : NAND2_X1 port map( A1 => n126, A2 => n125, ZN => OUT1(3));
   U64 : NAND2_X1 port map( A1 => n136, A2 => n135, ZN => OUT1(8));
   U65 : NAND2_X1 port map( A1 => n132, A2 => n131, ZN => OUT1(6));
   U66 : NAND2_X1 port map( A1 => n128, A2 => n127, ZN => OUT1(4));
   U67 : AOI22_X1 port map( A1 => n71, A2 => IN1(11), B1 => n73, B2 => IN0(11),
                           ZN => n90);
   U68 : AOI22_X1 port map( A1 => n40, A2 => IN1(10), B1 => n74, B2 => IN0(10),
                           ZN => n88);
   U69 : AOI22_X1 port map( A1 => n71, A2 => IN1(15), B1 => n75, B2 => IN0(15),
                           ZN => n98);
   U70 : AOI22_X1 port map( A1 => n40, A2 => IN1(13), B1 => n73, B2 => IN0(13),
                           ZN => n94);
   U71 : AOI22_X1 port map( A1 => n71, A2 => IN1(0), B1 => n74, B2 => IN0(0), 
                           ZN => n86);
   U72 : AOI22_X1 port map( A1 => n40, A2 => IN1(12), B1 => n73, B2 => IN0(12),
                           ZN => n92);
   U73 : AOI22_X1 port map( A1 => n71, A2 => IN1(14), B1 => n74, B2 => IN0(14),
                           ZN => n96);
   U74 : AOI22_X1 port map( A1 => n40, A2 => IN1(16), B1 => n73, B2 => IN0(16),
                           ZN => n100);
   U75 : AOI22_X1 port map( A1 => n76, A2 => IN3(0), B1 => n80, B2 => IN2(0), 
                           ZN => n85);
   U76 : AOI22_X1 port map( A1 => n76, A2 => IN3(12), B1 => n79, B2 => IN2(12),
                           ZN => n91);
   U77 : AOI22_X1 port map( A1 => n76, A2 => IN3(15), B1 => n80, B2 => IN2(15),
                           ZN => n97);
   U78 : AOI22_X1 port map( A1 => n76, A2 => IN3(11), B1 => n79, B2 => IN2(11),
                           ZN => n89);
   U79 : AOI22_X1 port map( A1 => n76, A2 => IN3(16), B1 => n7, B2 => IN2(16), 
                           ZN => n99);
   U80 : AOI22_X1 port map( A1 => n40, A2 => IN1(2), B1 => n75, B2 => IN0(2), 
                           ZN => n124);
   U81 : AOI22_X1 port map( A1 => n72, A2 => IN1(9), B1 => n75, B2 => IN0(9), 
                           ZN => n138);
   U82 : AOI22_X1 port map( A1 => n40, A2 => IN1(6), B1 => n75, B2 => IN0(6), 
                           ZN => n132);
   U83 : AOI22_X1 port map( A1 => n72, A2 => IN1(7), B1 => n73, B2 => IN0(7), 
                           ZN => n134);
   U84 : AOI22_X1 port map( A1 => n71, A2 => IN1(8), B1 => n75, B2 => IN0(8), 
                           ZN => n136);
   U85 : AOI22_X1 port map( A1 => n71, A2 => IN1(5), B1 => n75, B2 => IN0(5), 
                           ZN => n130);
   U86 : AOI22_X1 port map( A1 => n72, A2 => IN1(3), B1 => n74, B2 => IN0(3), 
                           ZN => n126);
   U87 : AOI22_X1 port map( A1 => n71, A2 => IN1(4), B1 => n73, B2 => IN0(4), 
                           ZN => n128);
   U88 : AOI22_X1 port map( A1 => n40, A2 => IN1(18), B1 => n75, B2 => IN0(18),
                           ZN => n104);
   U89 : AOI22_X1 port map( A1 => n71, A2 => IN1(1), B1 => n73, B2 => IN0(1), 
                           ZN => n108);
   U90 : AOI22_X1 port map( A1 => n40, A2 => IN1(27), B1 => n75, B2 => IN0(27),
                           ZN => n122);
   U91 : AOI22_X1 port map( A1 => n72, A2 => IN1(25), B1 => n73, B2 => IN0(25),
                           ZN => n118);
   U92 : AOI22_X1 port map( A1 => n72, A2 => IN1(17), B1 => n74, B2 => IN0(17),
                           ZN => n102);
   U93 : AOI22_X1 port map( A1 => n40, A2 => IN1(21), B1 => n74, B2 => IN0(21),
                           ZN => n112);
   U94 : AOI22_X1 port map( A1 => n72, A2 => IN1(19), B1 => n75, B2 => IN0(19),
                           ZN => n106);
   U95 : AOI22_X1 port map( A1 => n72, A2 => IN1(24), B1 => n75, B2 => IN0(24),
                           ZN => n116);
   U96 : AOI22_X1 port map( A1 => n72, A2 => IN1(26), B1 => n73, B2 => IN0(26),
                           ZN => n120);
   U97 : AOI22_X1 port map( A1 => n72, A2 => IN1(20), B1 => n74, B2 => IN0(20),
                           ZN => n110);
   U98 : AOI22_X1 port map( A1 => n40, A2 => IN1(22), B1 => n74, B2 => IN0(22),
                           ZN => n114);
   U99 : NOR2_X1 port map( A1 => n81, A2 => CTRL(1), ZN => n82);
   U100 : NAND2_X1 port map( A1 => n104, A2 => n103, ZN => OUT1(18));
   U101 : NAND2_X1 port map( A1 => n124, A2 => n123, ZN => OUT1(2));
   U102 : AOI22_X1 port map( A1 => n76, A2 => IN3(1), B1 => n80, B2 => IN2(1), 
                           ZN => n107);
   U103 : AOI22_X1 port map( A1 => n76, A2 => IN3(19), B1 => n7, B2 => IN2(19),
                           ZN => n105);
   U104 : AOI22_X1 port map( A1 => n77, A2 => IN3(27), B1 => n80, B2 => IN2(27)
                           , ZN => n121);
   U105 : AOI22_X1 port map( A1 => n77, A2 => IN3(25), B1 => n80, B2 => IN2(25)
                           , ZN => n117);
   U106 : AOI22_X1 port map( A1 => n76, A2 => IN3(18), B1 => n7, B2 => IN2(18),
                           ZN => n103);
   U107 : AOI22_X1 port map( A1 => n77, A2 => IN3(20), B1 => n7, B2 => IN2(20),
                           ZN => n109);
   U108 : AOI22_X1 port map( A1 => n77, A2 => IN3(22), B1 => n79, B2 => IN2(22)
                           , ZN => n113);
   U109 : AOI22_X1 port map( A1 => n77, A2 => IN3(26), B1 => n7, B2 => IN2(26),
                           ZN => n119);
   U110 : AOI22_X1 port map( A1 => n78, A2 => IN3(7), B1 => n80, B2 => IN2(7), 
                           ZN => n133);
   U111 : AOI22_X1 port map( A1 => n77, A2 => IN3(5), B1 => n7, B2 => IN2(5), 
                           ZN => n129);
   U112 : AOI22_X1 port map( A1 => n77, A2 => IN3(2), B1 => n7, B2 => IN2(2), 
                           ZN => n123);
   U113 : AOI22_X1 port map( A1 => n78, A2 => IN3(8), B1 => n80, B2 => IN2(8), 
                           ZN => n135);
   U114 : AOI22_X1 port map( A1 => n78, A2 => IN3(6), B1 => n7, B2 => IN2(6), 
                           ZN => n131);

end SYN_bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity ff32_en_1 is

   port( D : in std_logic_vector (31 downto 0);  en, clk, rst : in std_logic;  
         Q : out std_logic_vector (31 downto 0));

end ff32_en_1;

architecture SYN_behavioral of ff32_en_1 is

   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_ff32_en_1
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal net3606, n32, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, 
      n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59
      , n60, n61, n62, n63, n64, n65 : std_logic;

begin
   
   Q_reg_31_inst : DFFR_X1 port map( D => D(31), CK => net3606, RN => n32, Q =>
                           Q(31), QN => n34);
   Q_reg_30_inst : DFFR_X1 port map( D => D(30), CK => net3606, RN => n32, Q =>
                           Q(30), QN => n35);
   Q_reg_29_inst : DFFR_X1 port map( D => D(29), CK => net3606, RN => n32, Q =>
                           Q(29), QN => n36);
   Q_reg_28_inst : DFFR_X1 port map( D => D(28), CK => net3606, RN => n32, Q =>
                           Q(28), QN => n37);
   Q_reg_27_inst : DFFR_X1 port map( D => D(27), CK => net3606, RN => n32, Q =>
                           Q(27), QN => n38);
   Q_reg_26_inst : DFFR_X1 port map( D => D(26), CK => net3606, RN => n32, Q =>
                           Q(26), QN => n39);
   Q_reg_25_inst : DFFR_X1 port map( D => D(25), CK => net3606, RN => n32, Q =>
                           Q(25), QN => n40);
   Q_reg_24_inst : DFFR_X1 port map( D => D(24), CK => net3606, RN => n32, Q =>
                           Q(24), QN => n41);
   Q_reg_23_inst : DFFR_X1 port map( D => D(23), CK => net3606, RN => n32, Q =>
                           Q(23), QN => n42);
   Q_reg_22_inst : DFFR_X1 port map( D => D(22), CK => net3606, RN => n32, Q =>
                           Q(22), QN => n43);
   Q_reg_21_inst : DFFR_X1 port map( D => D(21), CK => net3606, RN => n32, Q =>
                           Q(21), QN => n44);
   Q_reg_20_inst : DFFR_X1 port map( D => D(20), CK => net3606, RN => n32, Q =>
                           Q(20), QN => n45);
   Q_reg_19_inst : DFFR_X1 port map( D => D(19), CK => net3606, RN => n32, Q =>
                           Q(19), QN => n46);
   Q_reg_18_inst : DFFR_X1 port map( D => D(18), CK => net3606, RN => n32, Q =>
                           Q(18), QN => n47);
   Q_reg_17_inst : DFFR_X1 port map( D => D(17), CK => net3606, RN => n32, Q =>
                           Q(17), QN => n48);
   Q_reg_16_inst : DFFR_X1 port map( D => D(16), CK => net3606, RN => n32, Q =>
                           Q(16), QN => n49);
   Q_reg_15_inst : DFFR_X1 port map( D => D(15), CK => net3606, RN => n32, Q =>
                           Q(15), QN => n50);
   Q_reg_14_inst : DFFR_X1 port map( D => D(14), CK => net3606, RN => n32, Q =>
                           Q(14), QN => n51);
   Q_reg_13_inst : DFFR_X1 port map( D => D(13), CK => net3606, RN => n32, Q =>
                           Q(13), QN => n52);
   Q_reg_12_inst : DFFR_X1 port map( D => D(12), CK => net3606, RN => n32, Q =>
                           Q(12), QN => n53);
   Q_reg_11_inst : DFFR_X1 port map( D => D(11), CK => net3606, RN => n32, Q =>
                           Q(11), QN => n54);
   Q_reg_10_inst : DFFR_X1 port map( D => D(10), CK => net3606, RN => n32, Q =>
                           Q(10), QN => n55);
   Q_reg_9_inst : DFFR_X1 port map( D => D(9), CK => net3606, RN => n32, Q => 
                           Q(9), QN => n56);
   Q_reg_8_inst : DFFR_X1 port map( D => D(8), CK => net3606, RN => n32, Q => 
                           Q(8), QN => n57);
   Q_reg_7_inst : DFFR_X1 port map( D => D(7), CK => net3606, RN => n32, Q => 
                           Q(7), QN => n58);
   Q_reg_6_inst : DFFR_X1 port map( D => D(6), CK => net3606, RN => n32, Q => 
                           Q(6), QN => n59);
   Q_reg_5_inst : DFFR_X1 port map( D => D(5), CK => net3606, RN => n32, Q => 
                           Q(5), QN => n60);
   Q_reg_4_inst : DFFR_X1 port map( D => D(4), CK => net3606, RN => n32, Q => 
                           Q(4), QN => n61);
   Q_reg_3_inst : DFFR_X1 port map( D => D(3), CK => net3606, RN => n32, Q => 
                           Q(3), QN => n62);
   Q_reg_2_inst : DFFR_X1 port map( D => D(2), CK => net3606, RN => n32, Q => 
                           Q(2), QN => n63);
   Q_reg_1_inst : DFFR_X1 port map( D => D(1), CK => net3606, RN => n32, Q => 
                           Q(1), QN => n64);
   Q_reg_0_inst : DFFR_X1 port map( D => D(0), CK => net3606, RN => n32, Q => 
                           Q(0), QN => n65);
   clk_gate_Q_reg : SNPS_CLOCK_GATE_HIGH_ff32_en_1 port map( CLK => clk, EN => 
                           en, ENCLK => net3606);
   U2 : INV_X2 port map( A => rst, ZN => n32);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_0 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_0;

architecture SYN_BEHAVIORAL of FA_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => S);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity mux21_SIZE4_0 is

   port( IN0, IN1 : in std_logic_vector (3 downto 0);  CTRL : in std_logic;  
         OUT1 : out std_logic_vector (3 downto 0));

end mux21_SIZE4_0;

architecture SYN_Bhe of mux21_SIZE4_0 is

begin
   OUT1 <= ( IN0(3), IN0(2), IN0(1), IN0(0) );

end SYN_Bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity RCA_N4_0 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_0;

architecture SYN_STRUCTURAL of RCA_N4_0 is

   component FA_125
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_126
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_127
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_0
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal n1, CTMP_3_port, CTMP_2_port, CTMP_1_port, net48717 : std_logic;

begin
   
   FAI_1 : FA_0 port map( A => A(0), B => B(0), Ci => n1, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_127 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_126 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_125 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => net48717);
   n1 <= '0';

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity shift_thirdLevel is

   port( sel : in std_logic_vector (2 downto 0);  A : in std_logic_vector (38 
         downto 0);  Y : out std_logic_vector (31 downto 0));

end shift_thirdLevel;

architecture SYN_behav of shift_thirdLevel is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, 
      n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32
      , n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, 
      n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61
      , n62, n63, n64, n65, n66, n67, n68, n69, n70, n1, n3, n71, n72, n73, n74
      , n75, n76 : std_logic;

begin
   
   U7 : MUX2_X1 port map( A => n7, B => n6, S => n71, Z => Y(30));
   U10 : MUX2_X1 port map( A => n6, B => n9, S => n71, Z => Y(29));
   U13 : MUX2_X1 port map( A => n9, B => n11, S => sel(0), Z => Y(28));
   U16 : MUX2_X1 port map( A => n11, B => n13, S => n71, Z => Y(27));
   U19 : MUX2_X1 port map( A => n13, B => n15, S => n71, Z => Y(26));
   U22 : MUX2_X1 port map( A => n15, B => n17, S => n3, Z => Y(25));
   U25 : MUX2_X1 port map( A => n17, B => n19, S => n3, Z => Y(24));
   U28 : MUX2_X1 port map( A => n19, B => n21, S => n3, Z => Y(23));
   U31 : MUX2_X1 port map( A => n21, B => n23, S => sel(0), Z => Y(22));
   U34 : MUX2_X1 port map( A => n23, B => n25, S => sel(0), Z => Y(21));
   U37 : MUX2_X1 port map( A => n25, B => n27, S => sel(0), Z => Y(20));
   U40 : MUX2_X1 port map( A => n27, B => n29, S => n71, Z => Y(19));
   U43 : MUX2_X1 port map( A => n29, B => n31, S => n3, Z => Y(18));
   U46 : MUX2_X1 port map( A => n31, B => n33, S => n3, Z => Y(17));
   U49 : MUX2_X1 port map( A => n33, B => n35, S => n3, Z => Y(16));
   U52 : MUX2_X1 port map( A => n35, B => n37, S => n3, Z => Y(15));
   U55 : MUX2_X1 port map( A => n37, B => n39, S => n3, Z => Y(14));
   U58 : MUX2_X1 port map( A => n39, B => n41, S => n3, Z => Y(13));
   U61 : MUX2_X1 port map( A => n41, B => n43, S => n3, Z => Y(12));
   U64 : MUX2_X1 port map( A => n43, B => n45, S => n3, Z => Y(11));
   U67 : MUX2_X1 port map( A => n45, B => n47, S => n3, Z => Y(10));
   U70 : MUX2_X1 port map( A => n47, B => n49, S => n3, Z => Y(9));
   U73 : MUX2_X1 port map( A => n49, B => n51, S => n3, Z => Y(8));
   U76 : MUX2_X1 port map( A => n51, B => n53, S => n3, Z => Y(7));
   U79 : MUX2_X1 port map( A => n53, B => n55, S => n71, Z => Y(6));
   U82 : MUX2_X1 port map( A => n55, B => n57, S => n71, Z => Y(5));
   U85 : MUX2_X1 port map( A => n57, B => n59, S => n71, Z => Y(4));
   U88 : MUX2_X1 port map( A => n59, B => n61, S => n71, Z => Y(3));
   U92 : MUX2_X1 port map( A => n63, B => n64, S => n71, Z => Y(1));
   U97 : MUX2_X1 port map( A => n64, B => n67, S => n71, Z => Y(0));
   U102 : MUX2_X1 port map( A => n70, B => n7, S => n71, Z => Y(31));
   U93 : AOI22_X1 port map( A1 => n75, A2 => A(1), B1 => A(5), B2 => n74, ZN =>
                           n65);
   U86 : AOI22_X1 port map( A1 => n75, A2 => A(3), B1 => A(7), B2 => n74, ZN =>
                           n60);
   U94 : AOI22_X1 port map( A1 => n73, A2 => n65, B1 => n60, B2 => n1, ZN => 
                           n64);
   U95 : AOI22_X1 port map( A1 => n75, A2 => A(0), B1 => A(4), B2 => n74, ZN =>
                           n66);
   U89 : AOI22_X1 port map( A1 => n75, A2 => A(2), B1 => A(6), B2 => n74, ZN =>
                           n62);
   U96 : AOI22_X1 port map( A1 => n73, A2 => n66, B1 => n62, B2 => n1, ZN => 
                           n67);
   U71 : AOI22_X1 port map( A1 => n75, A2 => A(8), B1 => A(12), B2 => n74, ZN 
                           => n50);
   U65 : AOI22_X1 port map( A1 => n75, A2 => A(10), B1 => A(14), B2 => n74, ZN 
                           => n46);
   U72 : AOI22_X1 port map( A1 => n73, A2 => n50, B1 => n46, B2 => n1, ZN => 
                           n51);
   U74 : AOI22_X1 port map( A1 => n76, A2 => A(7), B1 => A(11), B2 => n74, ZN 
                           => n52);
   U68 : AOI22_X1 port map( A1 => n75, A2 => A(9), B1 => A(13), B2 => n74, ZN 
                           => n48);
   U75 : AOI22_X1 port map( A1 => n73, A2 => n52, B1 => n48, B2 => n1, ZN => 
                           n53);
   U5 : AOI22_X1 port map( A1 => n75, A2 => A(30), B1 => A(34), B2 => n74, ZN 
                           => n5);
   U2 : AOI22_X1 port map( A1 => sel(2), A2 => A(32), B1 => A(36), B2 => n74, 
                           ZN => n2);
   U6 : AOI22_X1 port map( A1 => n73, A2 => n5, B1 => n2, B2 => n72, ZN => n6);
   U8 : AOI22_X1 port map( A1 => sel(2), A2 => A(29), B1 => A(33), B2 => n74, 
                           ZN => n8);
   U4 : AOI22_X1 port map( A1 => sel(2), A2 => A(31), B1 => A(35), B2 => n74, 
                           ZN => n4);
   U9 : AOI22_X1 port map( A1 => n73, A2 => n8, B1 => n4, B2 => n72, ZN => n9);
   U23 : AOI22_X1 port map( A1 => n76, A2 => A(24), B1 => A(28), B2 => n74, ZN 
                           => n18);
   U17 : AOI22_X1 port map( A1 => n76, A2 => A(26), B1 => A(30), B2 => n74, ZN 
                           => n14);
   U24 : AOI22_X1 port map( A1 => n73, A2 => n18, B1 => n14, B2 => n72, ZN => 
                           n19);
   U26 : AOI22_X1 port map( A1 => n75, A2 => A(23), B1 => A(27), B2 => n74, ZN 
                           => n20);
   U20 : AOI22_X1 port map( A1 => n76, A2 => A(25), B1 => A(29), B2 => n74, ZN 
                           => n16);
   U27 : AOI22_X1 port map( A1 => n73, A2 => n20, B1 => n16, B2 => n72, ZN => 
                           n21);
   U47 : AOI22_X1 port map( A1 => n76, A2 => A(16), B1 => A(20), B2 => n74, ZN 
                           => n34);
   U41 : AOI22_X1 port map( A1 => n76, A2 => A(18), B1 => A(22), B2 => n74, ZN 
                           => n30);
   U48 : AOI22_X1 port map( A1 => n73, A2 => n34, B1 => n30, B2 => n1, ZN => 
                           n35);
   U50 : AOI22_X1 port map( A1 => n76, A2 => A(15), B1 => A(19), B2 => n74, ZN 
                           => n36);
   U44 : AOI22_X1 port map( A1 => n76, A2 => A(17), B1 => A(21), B2 => n74, ZN 
                           => n32);
   U51 : AOI22_X1 port map( A1 => n73, A2 => n36, B1 => n32, B2 => n1, ZN => 
                           n37);
   U35 : AOI22_X1 port map( A1 => n76, A2 => A(20), B1 => A(24), B2 => n74, ZN 
                           => n26);
   U29 : AOI22_X1 port map( A1 => n76, A2 => A(22), B1 => A(26), B2 => n74, ZN 
                           => n22);
   U36 : AOI22_X1 port map( A1 => n73, A2 => n26, B1 => n22, B2 => n72, ZN => 
                           n27);
   U38 : AOI22_X1 port map( A1 => n76, A2 => A(19), B1 => A(23), B2 => n74, ZN 
                           => n28);
   U32 : AOI22_X1 port map( A1 => n76, A2 => A(21), B1 => A(25), B2 => n74, ZN 
                           => n24);
   U39 : AOI22_X1 port map( A1 => n73, A2 => n28, B1 => n24, B2 => n72, ZN => 
                           n29);
   U42 : AOI22_X1 port map( A1 => n73, A2 => n30, B1 => n26, B2 => n1, ZN => 
                           n31);
   U45 : AOI22_X1 port map( A1 => n73, A2 => n32, B1 => n28, B2 => n1, ZN => 
                           n33);
   U11 : AOI22_X1 port map( A1 => sel(2), A2 => A(28), B1 => A(32), B2 => n74, 
                           ZN => n10);
   U18 : AOI22_X1 port map( A1 => n73, A2 => n14, B1 => n10, B2 => n72, ZN => 
                           n15);
   U14 : AOI22_X1 port map( A1 => n76, A2 => A(27), B1 => A(31), B2 => n74, ZN 
                           => n12);
   U21 : AOI22_X1 port map( A1 => n73, A2 => n16, B1 => n12, B2 => n72, ZN => 
                           n17);
   U12 : AOI22_X1 port map( A1 => n73, A2 => n10, B1 => n5, B2 => n72, ZN => 
                           n11);
   U15 : AOI22_X1 port map( A1 => n73, A2 => n12, B1 => n8, B2 => n72, ZN => 
                           n13);
   U98 : AOI22_X1 port map( A1 => n75, A2 => A(33), B1 => A(37), B2 => n74, ZN 
                           => n68);
   U99 : AOI22_X1 port map( A1 => n73, A2 => n4, B1 => n68, B2 => n1, ZN => n7)
                           ;
   U30 : AOI22_X1 port map( A1 => n73, A2 => n22, B1 => n18, B2 => n72, ZN => 
                           n23);
   U33 : AOI22_X1 port map( A1 => n73, A2 => n24, B1 => n20, B2 => n72, ZN => 
                           n25);
   U100 : AOI22_X1 port map( A1 => n75, A2 => A(34), B1 => A(38), B2 => n74, ZN
                           => n69);
   U101 : AOI22_X1 port map( A1 => sel(1), A2 => n2, B1 => n69, B2 => n1, ZN =>
                           n70);
   U53 : AOI22_X1 port map( A1 => n76, A2 => A(14), B1 => A(18), B2 => n74, ZN 
                           => n38);
   U54 : AOI22_X1 port map( A1 => n73, A2 => n38, B1 => n34, B2 => n1, ZN => 
                           n39);
   U83 : AOI22_X1 port map( A1 => n76, A2 => A(4), B1 => A(8), B2 => n74, ZN =>
                           n58);
   U77 : AOI22_X1 port map( A1 => n76, A2 => A(6), B1 => A(10), B2 => n74, ZN 
                           => n54);
   U84 : AOI22_X1 port map( A1 => n73, A2 => n58, B1 => n54, B2 => n1, ZN => 
                           n59);
   U80 : AOI22_X1 port map( A1 => n75, A2 => A(5), B1 => A(9), B2 => n74, ZN =>
                           n56);
   U87 : AOI22_X1 port map( A1 => n73, A2 => n60, B1 => n56, B2 => n1, ZN => 
                           n61);
   U56 : AOI22_X1 port map( A1 => n76, A2 => A(13), B1 => A(17), B2 => n74, ZN 
                           => n40);
   U57 : AOI22_X1 port map( A1 => n73, A2 => n40, B1 => n36, B2 => n1, ZN => 
                           n41);
   U59 : AOI22_X1 port map( A1 => n75, A2 => A(12), B1 => A(16), B2 => n74, ZN 
                           => n42);
   U60 : AOI22_X1 port map( A1 => sel(1), A2 => n42, B1 => n38, B2 => n1, ZN =>
                           n43);
   U62 : AOI22_X1 port map( A1 => n75, A2 => A(11), B1 => A(15), B2 => n74, ZN 
                           => n44);
   U63 : AOI22_X1 port map( A1 => sel(1), A2 => n44, B1 => n40, B2 => n1, ZN =>
                           n45);
   U66 : AOI22_X1 port map( A1 => sel(1), A2 => n46, B1 => n42, B2 => n1, ZN =>
                           n47);
   U69 : AOI22_X1 port map( A1 => n73, A2 => n48, B1 => n44, B2 => n1, ZN => 
                           n49);
   U90 : AOI22_X1 port map( A1 => n73, A2 => n62, B1 => n58, B2 => n1, ZN => 
                           n63);
   U78 : AOI22_X1 port map( A1 => sel(1), A2 => n54, B1 => n50, B2 => n1, ZN =>
                           n55);
   U81 : AOI22_X1 port map( A1 => sel(1), A2 => n56, B1 => n52, B2 => n1, ZN =>
                           n57);
   U1 : MUX2_X1 port map( A => n61, B => n63, S => n71, Z => Y(2));
   U3 : INV_X2 port map( A => sel(2), ZN => n74);
   U91 : INV_X2 port map( A => n73, ZN => n1);
   U103 : BUF_X1 port map( A => sel(0), Z => n71);
   U104 : BUF_X1 port map( A => sel(0), Z => n3);
   U105 : BUF_X1 port map( A => sel(2), Z => n75);
   U106 : BUF_X1 port map( A => sel(2), Z => n76);
   U107 : BUF_X2 port map( A => sel(1), Z => n73);
   U108 : INV_X1 port map( A => n73, ZN => n72);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity shift_secondLevel is

   port( sel : in std_logic_vector (1 downto 0);  mask00, mask08, mask16 : in 
         std_logic_vector (38 downto 0);  Y : out std_logic_vector (38 downto 
         0));

end shift_secondLevel;

architecture SYN_behav of shift_secondLevel is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X4
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n42, n43, n44, n45, n46, n48, n49, n50, n51, n52, n53, n54, n55, n56,
      n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71
      , n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n1, n3
      , n4, n12 : std_logic;

begin
   
   U57 : AOI222_X1 port map( A1 => n4, A2 => mask00(1), B1 => n44, B2 => 
                           mask16(1), C1 => n3, C2 => mask08(1), ZN => n72);
   U11 : AOI222_X1 port map( A1 => n4, A2 => mask00(5), B1 => n44, B2 => 
                           mask16(5), C1 => n3, C2 => mask08(5), ZN => n49);
   U15 : AOI222_X1 port map( A1 => n4, A2 => mask00(3), B1 => n44, B2 => 
                           mask16(3), C1 => n3, C2 => mask08(3), ZN => n51);
   U79 : AOI222_X1 port map( A1 => n4, A2 => mask00(0), B1 => n44, B2 => 
                           mask16(0), C1 => n3, C2 => mask08(0), ZN => n83);
   U13 : AOI222_X1 port map( A1 => n4, A2 => mask00(4), B1 => n44, B2 => 
                           mask16(4), C1 => n3, C2 => mask08(4), ZN => n50);
   U35 : AOI222_X1 port map( A1 => n12, A2 => mask00(2), B1 => n44, B2 => 
                           mask16(2), C1 => n45, C2 => mask08(2), ZN => n61);
   U9 : AOI222_X1 port map( A1 => n4, A2 => mask00(6), B1 => n44, B2 => 
                           mask16(6), C1 => n3, C2 => mask08(6), ZN => n48);
   U5 : AOI222_X1 port map( A1 => n4, A2 => mask00(8), B1 => n44, B2 => 
                           mask16(8), C1 => n3, C2 => mask08(8), ZN => n46);
   U73 : AOI222_X1 port map( A1 => n4, A2 => mask00(12), B1 => n44, B2 => 
                           mask16(12), C1 => n3, C2 => mask08(12), ZN => n80);
   U77 : AOI222_X1 port map( A1 => n4, A2 => mask00(10), B1 => n44, B2 => 
                           mask16(10), C1 => n3, C2 => mask08(10), ZN => n82);
   U69 : AOI222_X1 port map( A1 => n4, A2 => mask00(14), B1 => n44, B2 => 
                           mask16(14), C1 => n3, C2 => mask08(14), ZN => n78);
   U75 : AOI222_X1 port map( A1 => n4, A2 => mask00(11), B1 => n44, B2 => 
                           mask16(11), C1 => n3, C2 => mask08(11), ZN => n81);
   U3 : AOI222_X1 port map( A1 => n12, A2 => mask00(9), B1 => n44, B2 => 
                           mask16(9), C1 => n45, C2 => mask08(9), ZN => n42);
   U71 : AOI222_X1 port map( A1 => n4, A2 => mask00(13), B1 => n44, B2 => 
                           mask16(13), C1 => n3, C2 => mask08(13), ZN => n79);
   U33 : AOI222_X1 port map( A1 => n12, A2 => mask00(30), B1 => n44, B2 => 
                           mask16(30), C1 => n45, C2 => mask08(30), ZN => n60);
   U25 : AOI222_X1 port map( A1 => n4, A2 => mask00(34), B1 => n44, B2 => 
                           mask16(34), C1 => n3, C2 => mask08(34), ZN => n56);
   U29 : AOI222_X1 port map( A1 => n4, A2 => mask00(32), B1 => n44, B2 => 
                           mask16(32), C1 => n3, C2 => mask08(32), ZN => n58);
   U21 : AOI222_X1 port map( A1 => n4, A2 => mask00(36), B1 => n44, B2 => 
                           mask16(36), C1 => n3, C2 => mask08(36), ZN => n54);
   U37 : AOI222_X1 port map( A1 => n12, A2 => mask00(29), B1 => n44, B2 => 
                           mask16(29), C1 => n45, C2 => mask08(29), ZN => n62);
   U27 : AOI222_X1 port map( A1 => n4, A2 => mask00(33), B1 => n44, B2 => 
                           mask16(33), C1 => n3, C2 => mask08(33), ZN => n57);
   U31 : AOI222_X1 port map( A1 => n4, A2 => mask00(31), B1 => n44, B2 => 
                           mask16(31), C1 => n3, C2 => mask08(31), ZN => n59);
   U23 : AOI222_X1 port map( A1 => n4, A2 => mask00(35), B1 => n44, B2 => 
                           mask16(35), C1 => n3, C2 => mask08(35), ZN => n55);
   U47 : AOI222_X1 port map( A1 => n12, A2 => mask00(24), B1 => n44, B2 => 
                           mask16(24), C1 => n45, C2 => mask08(24), ZN => n67);
   U39 : AOI222_X1 port map( A1 => n12, A2 => mask00(28), B1 => n44, B2 => 
                           mask16(28), C1 => n45, C2 => mask08(28), ZN => n63);
   U43 : AOI222_X1 port map( A1 => n12, A2 => mask00(26), B1 => n44, B2 => 
                           mask16(26), C1 => n45, C2 => mask08(26), ZN => n65);
   U49 : AOI222_X1 port map( A1 => n12, A2 => mask00(23), B1 => n44, B2 => 
                           mask16(23), C1 => n45, C2 => mask08(23), ZN => n68);
   U41 : AOI222_X1 port map( A1 => n12, A2 => mask00(27), B1 => n44, B2 => 
                           mask16(27), C1 => n45, C2 => mask08(27), ZN => n64);
   U45 : AOI222_X1 port map( A1 => n12, A2 => mask00(25), B1 => n44, B2 => 
                           mask16(25), C1 => n45, C2 => mask08(25), ZN => n66);
   U65 : AOI222_X1 port map( A1 => n4, A2 => mask00(16), B1 => n44, B2 => 
                           mask16(16), C1 => n3, C2 => mask08(16), ZN => n76);
   U55 : AOI222_X1 port map( A1 => n12, A2 => mask00(20), B1 => n44, B2 => 
                           mask16(20), C1 => n45, C2 => mask08(20), ZN => n71);
   U61 : AOI222_X1 port map( A1 => n4, A2 => mask00(18), B1 => n44, B2 => 
                           mask16(18), C1 => n3, C2 => mask08(18), ZN => n74);
   U51 : AOI222_X1 port map( A1 => n12, A2 => mask00(22), B1 => n44, B2 => 
                           mask16(22), C1 => n45, C2 => mask08(22), ZN => n69);
   U67 : AOI222_X1 port map( A1 => n4, A2 => mask00(15), B1 => n44, B2 => 
                           mask16(15), C1 => n3, C2 => mask08(15), ZN => n77);
   U59 : AOI222_X1 port map( A1 => n4, A2 => mask00(19), B1 => n44, B2 => 
                           mask16(19), C1 => n3, C2 => mask08(19), ZN => n73);
   U63 : AOI222_X1 port map( A1 => n4, A2 => mask00(17), B1 => n44, B2 => 
                           mask16(17), C1 => n3, C2 => mask08(17), ZN => n75);
   U53 : AOI222_X1 port map( A1 => n12, A2 => mask00(21), B1 => n44, B2 => 
                           mask16(21), C1 => n45, C2 => mask08(21), ZN => n70);
   U19 : AOI222_X1 port map( A1 => n4, A2 => mask00(37), B1 => n44, B2 => 
                           mask16(37), C1 => n3, C2 => mask08(37), ZN => n53);
   U17 : AOI222_X1 port map( A1 => n4, A2 => mask00(38), B1 => n44, B2 => 
                           mask16(38), C1 => n3, C2 => mask08(38), ZN => n52);
   U82 : INV_X1 port map( A => sel(0), ZN => n84);
   U56 : INV_X1 port map( A => n72, ZN => Y(1));
   U10 : INV_X1 port map( A => n49, ZN => Y(5));
   U14 : INV_X1 port map( A => n51, ZN => Y(3));
   U78 : INV_X1 port map( A => n83, ZN => Y(0));
   U12 : INV_X1 port map( A => n50, ZN => Y(4));
   U34 : INV_X1 port map( A => n61, ZN => Y(2));
   U8 : INV_X1 port map( A => n48, ZN => Y(6));
   U4 : INV_X1 port map( A => n46, ZN => Y(8));
   U72 : INV_X1 port map( A => n80, ZN => Y(12));
   U76 : INV_X1 port map( A => n82, ZN => Y(10));
   U68 : INV_X1 port map( A => n78, ZN => Y(14));
   U74 : INV_X1 port map( A => n81, ZN => Y(11));
   U2 : INV_X1 port map( A => n42, ZN => Y(9));
   U70 : INV_X1 port map( A => n79, ZN => Y(13));
   U32 : INV_X1 port map( A => n60, ZN => Y(30));
   U24 : INV_X1 port map( A => n56, ZN => Y(34));
   U28 : INV_X1 port map( A => n58, ZN => Y(32));
   U20 : INV_X1 port map( A => n54, ZN => Y(36));
   U36 : INV_X1 port map( A => n62, ZN => Y(29));
   U26 : INV_X1 port map( A => n57, ZN => Y(33));
   U30 : INV_X1 port map( A => n59, ZN => Y(31));
   U22 : INV_X1 port map( A => n55, ZN => Y(35));
   U46 : INV_X1 port map( A => n67, ZN => Y(24));
   U38 : INV_X1 port map( A => n63, ZN => Y(28));
   U42 : INV_X1 port map( A => n65, ZN => Y(26));
   U48 : INV_X1 port map( A => n68, ZN => Y(23));
   U40 : INV_X1 port map( A => n64, ZN => Y(27));
   U44 : INV_X1 port map( A => n66, ZN => Y(25));
   U64 : INV_X1 port map( A => n76, ZN => Y(16));
   U54 : INV_X1 port map( A => n71, ZN => Y(20));
   U60 : INV_X1 port map( A => n74, ZN => Y(18));
   U50 : INV_X1 port map( A => n69, ZN => Y(22));
   U66 : INV_X1 port map( A => n77, ZN => Y(15));
   U58 : INV_X1 port map( A => n73, ZN => Y(19));
   U62 : INV_X1 port map( A => n75, ZN => Y(17));
   U52 : INV_X1 port map( A => n70, ZN => Y(21));
   U18 : INV_X1 port map( A => n53, ZN => Y(37));
   U16 : INV_X1 port map( A => n52, ZN => Y(38));
   U6 : AOI222_X1 port map( A1 => mask00(7), A2 => n4, B1 => mask08(7), B2 => 
                           n3, C1 => mask16(7), C2 => n44, ZN => n1);
   U7 : INV_X1 port map( A => n1, ZN => Y(7));
   U80 : NOR2_X2 port map( A1 => sel(1), A2 => n84, ZN => n45);
   U81 : AND2_X4 port map( A1 => n84, A2 => sel(1), ZN => n44);
   U83 : BUF_X1 port map( A => n45, Z => n3);
   U84 : BUF_X1 port map( A => n43, Z => n12);
   U85 : BUF_X2 port map( A => n43, Z => n4);
   U86 : NOR2_X1 port map( A1 => sel(1), A2 => sel(0), ZN => n43);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity shift_firstLevel is

   port( A : in std_logic_vector (31 downto 0);  sel : in std_logic_vector (1 
         downto 0);  mask00, mask08, mask16 : out std_logic_vector (38 downto 
         0));

end shift_firstLevel;

architecture SYN_behav of shift_firstLevel is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal mask08_38_port, mask08_37_port, mask08_36_port, mask08_35_port, 
      mask08_34_port, mask08_33_port, mask08_32_port, mask08_31_port, 
      mask08_23_port, mask08_22_port, mask08_21_port, mask08_20_port, 
      mask08_19_port, mask08_18_port, mask08_17_port, mask08_16_port, 
      mask08_15_port, mask08_7_port, mask08_6_port, mask08_5_port, 
      mask08_4_port, mask08_3_port, mask08_2_port, mask08_1_port, mask08_0_port
      , mask16_38_port, mask16_37_port, mask16_36_port, mask16_35_port, 
      mask16_34_port, mask16_33_port, mask16_32_port, mask16_31_port, 
      mask16_30_port, mask16_29_port, mask16_28_port, mask16_27_port, 
      mask16_26_port, mask16_25_port, mask16_24_port, mask16_23_port, 
      mask16_15_port, mask16_14_port, mask16_13_port, mask16_12_port, 
      mask16_11_port, mask16_10_port, mask16_9_port, mask16_8_port, 
      mask16_7_port, mask16_6_port, mask16_5_port, mask16_4_port, mask16_3_port
      , mask16_2_port, mask16_1_port, mask16_0_port, n37, n38, n39, n40, 
      mask16_17_port, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, 
      n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67
      , n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, 
      n82, n83, n84, n85, n86, n89, n90, n91, n92, n93, n94, n95, n96, n1, n2, 
      n3 : std_logic;

begin
   mask08 <= ( mask08_38_port, mask08_37_port, mask08_36_port, mask08_35_port, 
      mask08_34_port, mask08_33_port, mask08_32_port, mask08_31_port, 
      mask16_38_port, mask16_37_port, mask16_36_port, mask16_35_port, 
      mask16_34_port, mask16_33_port, mask16_32_port, mask08_23_port, 
      mask08_22_port, mask08_21_port, mask08_20_port, mask08_19_port, 
      mask08_18_port, mask08_17_port, mask08_16_port, mask08_15_port, 
      mask16_6_port, mask16_5_port, mask16_4_port, mask16_3_port, mask16_2_port
      , mask16_1_port, mask16_0_port, mask08_7_port, mask08_6_port, 
      mask08_5_port, mask08_4_port, mask08_3_port, mask08_2_port, mask08_1_port
      , mask08_0_port );
   mask16 <= ( mask16_38_port, mask16_37_port, mask16_36_port, mask16_35_port, 
      mask16_34_port, mask16_33_port, mask16_32_port, mask16_31_port, 
      mask16_30_port, mask16_29_port, mask16_28_port, mask16_27_port, 
      mask16_26_port, mask16_25_port, mask16_24_port, mask16_23_port, 
      mask16_17_port, mask16_17_port, mask16_17_port, mask16_17_port, 
      mask16_17_port, mask16_17_port, mask16_17_port, mask16_15_port, 
      mask16_14_port, mask16_13_port, mask16_12_port, mask16_11_port, 
      mask16_10_port, mask16_9_port, mask16_8_port, mask16_7_port, 
      mask16_6_port, mask16_5_port, mask16_4_port, mask16_3_port, mask16_2_port
      , mask16_1_port, mask16_0_port );
   
   U134 : NAND2_X1 port map( A1 => sel(0), A2 => A(17), ZN => n55);
   U59 : NAND2_X1 port map( A1 => sel(0), A2 => A(9), ZN => n79);
   U122 : NAND2_X1 port map( A1 => sel(0), A2 => A(21), ZN => n81);
   U146 : NAND2_X1 port map( A1 => sel(0), A2 => A(13), ZN => n59);
   U129 : NAND2_X1 port map( A1 => sel(0), A2 => A(19), ZN => n83);
   U152 : NAND2_X1 port map( A1 => sel(0), A2 => A(11), ZN => n61);
   U157 : NOR2_X1 port map( A1 => sel(0), A2 => sel(1), ZN => n86);
   U116 : NAND2_X1 port map( A1 => sel(0), A2 => A(23), ZN => n39);
   U140 : NAND2_X1 port map( A1 => sel(0), A2 => A(15), ZN => n57);
   U137 : NAND2_X1 port map( A1 => sel(0), A2 => A(16), ZN => n56);
   U62 : NAND2_X1 port map( A1 => sel(0), A2 => A(8), ZN => n85);
   U125 : NAND2_X1 port map( A1 => sel(0), A2 => A(20), ZN => n82);
   U149 : NAND2_X1 port map( A1 => sel(0), A2 => A(12), ZN => n60);
   U131 : NAND2_X1 port map( A1 => sel(0), A2 => A(18), ZN => n84);
   U155 : NAND2_X1 port map( A1 => sel(0), A2 => A(10), ZN => n71);
   U119 : NAND2_X1 port map( A1 => sel(0), A2 => A(22), ZN => n80);
   U143 : NAND2_X1 port map( A1 => sel(0), A2 => A(14), ZN => n58);
   U63 : NAND2_X1 port map( A1 => n2, A2 => A(1), ZN => n48);
   U61 : NAND2_X1 port map( A1 => n48, A2 => n85, ZN => mask00(8));
   U113 : NAND2_X1 port map( A1 => sel(0), A2 => A(24), ZN => n38);
   U150 : NAND2_X1 port map( A1 => n2, A2 => A(5), ZN => n44);
   U148 : NAND2_X1 port map( A1 => n44, A2 => n60, ZN => mask00(12));
   U101 : NAND2_X1 port map( A1 => sel(0), A2 => A(28), ZN => n52);
   U156 : NAND2_X1 port map( A1 => n86, A2 => A(3), ZN => n46);
   U154 : NAND2_X1 port map( A1 => n46, A2 => n71, ZN => mask00(10));
   U107 : NAND2_X1 port map( A1 => sel(0), A2 => A(26), ZN => n54);
   U144 : NAND2_X1 port map( A1 => n2, A2 => A(7), ZN => n42);
   U142 : NAND2_X1 port map( A1 => n42, A2 => n58, ZN => mask00(14));
   U94 : NAND2_X1 port map( A1 => sel(0), A2 => A(30), ZN => n50);
   U153 : NAND2_X1 port map( A1 => n2, A2 => A(4), ZN => n45);
   U151 : NAND2_X1 port map( A1 => n45, A2 => n61, ZN => mask00(11));
   U104 : NAND2_X1 port map( A1 => sel(0), A2 => A(27), ZN => n53);
   U60 : NAND2_X1 port map( A1 => n2, A2 => A(2), ZN => n47);
   U58 : NAND2_X1 port map( A1 => n47, A2 => n79, ZN => mask00(9));
   U110 : NAND2_X1 port map( A1 => sel(0), A2 => A(25), ZN => n37);
   U147 : NAND2_X1 port map( A1 => n2, A2 => A(6), ZN => n43);
   U145 : NAND2_X1 port map( A1 => n43, A2 => n59, ZN => mask00(13));
   U98 : NAND2_X1 port map( A1 => sel(0), A2 => A(29), ZN => n51);
   U93 : NAND2_X1 port map( A1 => n2, A2 => A(23), ZN => n62);
   U92 : NAND2_X1 port map( A1 => n50, A2 => n62, ZN => mask00(30));
   U91 : NAND2_X1 port map( A1 => sel(0), A2 => A(31), ZN => n78);
   U6 : NAND2_X1 port map( A1 => n42, A2 => n3, ZN => mask16_30_port);
   U118 : NAND2_X1 port map( A1 => n86, A2 => A(15), ZN => n70);
   U34 : NAND2_X1 port map( A1 => n70, A2 => n3, ZN => mask16_38_port);
   U81 : AOI21_X1 port map( B1 => A(27), B2 => n2, A => mask16_17_port, ZN => 
                           n93);
   U132 : NAND2_X1 port map( A1 => n86, A2 => A(11), ZN => n75);
   U39 : NAND2_X1 port map( A1 => n75, A2 => n3, ZN => mask16_34_port);
   U106 : NAND2_X1 port map( A1 => n2, A2 => A(19), ZN => n66);
   U30 : NAND2_X1 port map( A1 => n66, A2 => n3, ZN => mask08_34_port);
   U85 : AOI21_X1 port map( B1 => A(25), B2 => n2, A => mask16_17_port, ZN => 
                           n95);
   U138 : NAND2_X1 port map( A1 => n2, A2 => A(9), ZN => n77);
   U41 : NAND2_X1 port map( A1 => n77, A2 => n3, ZN => mask16_32_port);
   U112 : NAND2_X1 port map( A1 => n2, A2 => A(17), ZN => n68);
   U32 : NAND2_X1 port map( A1 => n68, A2 => n3, ZN => mask08_32_port);
   U77 : AOI21_X1 port map( B1 => A(29), B2 => n2, A => mask16_17_port, ZN => 
                           n91);
   U124 : NAND2_X1 port map( A1 => n86, A2 => A(13), ZN => n73);
   U37 : NAND2_X1 port map( A1 => n73, A2 => n3, ZN => mask16_36_port);
   U100 : NAND2_X1 port map( A1 => n2, A2 => A(21), ZN => n64);
   U28 : NAND2_X1 port map( A1 => n64, A2 => n3, ZN => mask08_36_port);
   U97 : NAND2_X1 port map( A1 => n2, A2 => A(22), ZN => n63);
   U96 : NAND2_X1 port map( A1 => n51, A2 => n63, ZN => mask00(29));
   U7 : NAND2_X1 port map( A1 => n43, A2 => n3, ZN => mask16_29_port);
   U121 : NAND2_X1 port map( A1 => n86, A2 => A(14), ZN => n72);
   U36 : NAND2_X1 port map( A1 => n72, A2 => n3, ZN => mask16_37_port);
   U83 : AOI21_X1 port map( B1 => A(26), B2 => n2, A => mask16_17_port, ZN => 
                           n94);
   U135 : NAND2_X1 port map( A1 => n2, A2 => A(10), ZN => n76);
   U40 : NAND2_X1 port map( A1 => n76, A2 => n3, ZN => mask16_33_port);
   U109 : NAND2_X1 port map( A1 => n2, A2 => A(18), ZN => n67);
   U31 : NAND2_X1 port map( A1 => n67, A2 => n3, ZN => mask08_33_port);
   U89 : AOI21_X1 port map( B1 => A(24), B2 => n2, A => mask16_15_port, ZN => 
                           n96);
   U141 : NAND2_X1 port map( A1 => n2, A2 => A(8), ZN => n40);
   U5 : NAND2_X1 port map( A1 => n40, A2 => n3, ZN => mask16_31_port);
   U115 : NAND2_X1 port map( A1 => n2, A2 => A(16), ZN => n69);
   U33 : NAND2_X1 port map( A1 => n69, A2 => n3, ZN => mask08_31_port);
   U79 : AOI21_X1 port map( B1 => A(28), B2 => n2, A => mask16_17_port, ZN => 
                           n92);
   U128 : NAND2_X1 port map( A1 => n86, A2 => A(12), ZN => n74);
   U38 : NAND2_X1 port map( A1 => n74, A2 => n3, ZN => mask16_35_port);
   U103 : NAND2_X1 port map( A1 => n2, A2 => A(20), ZN => n65);
   U29 : NAND2_X1 port map( A1 => n65, A2 => n3, ZN => mask08_35_port);
   U111 : NAND2_X1 port map( A1 => n38, A2 => n68, ZN => mask00(24));
   U12 : NAND2_X1 port map( A1 => n3, A2 => n48, ZN => mask16_24_port);
   U99 : NAND2_X1 port map( A1 => n52, A2 => n64, ZN => mask00(28));
   U8 : NAND2_X1 port map( A1 => n44, A2 => n3, ZN => mask16_28_port);
   U105 : NAND2_X1 port map( A1 => n54, A2 => n66, ZN => mask00(26));
   U10 : NAND2_X1 port map( A1 => n46, A2 => n3, ZN => mask16_26_port);
   U114 : NAND2_X1 port map( A1 => n39, A2 => n69, ZN => mask00(23));
   U13 : NAND2_X1 port map( A1 => n3, A2 => n49, ZN => mask16_23_port);
   U42 : NAND2_X1 port map( A1 => n40, A2 => n78, ZN => mask08_23_port);
   U102 : NAND2_X1 port map( A1 => n53, A2 => n65, ZN => mask00(27));
   U9 : NAND2_X1 port map( A1 => n45, A2 => n3, ZN => mask16_27_port);
   U108 : NAND2_X1 port map( A1 => n37, A2 => n67, ZN => mask00(25));
   U11 : NAND2_X1 port map( A1 => n3, A2 => n47, ZN => mask16_25_port);
   U136 : NAND2_X1 port map( A1 => n77, A2 => n56, ZN => mask00(16));
   U50 : NAND2_X1 port map( A1 => n38, A2 => n48, ZN => mask08_16_port);
   U123 : NAND2_X1 port map( A1 => n82, A2 => n73, ZN => mask00(20));
   U45 : NAND2_X1 port map( A1 => n44, A2 => n52, ZN => mask08_20_port);
   U130 : NAND2_X1 port map( A1 => n75, A2 => n84, ZN => mask00(18));
   U48 : NAND2_X1 port map( A1 => n46, A2 => n54, ZN => mask08_18_port);
   U117 : NAND2_X1 port map( A1 => n80, A2 => n70, ZN => mask00(22));
   U43 : NAND2_X1 port map( A1 => n42, A2 => n50, ZN => mask08_22_port);
   U139 : NAND2_X1 port map( A1 => n40, A2 => n57, ZN => mask00(15));
   U51 : NAND2_X1 port map( A1 => n39, A2 => n49, ZN => mask08_15_port);
   U127 : NAND2_X1 port map( A1 => n83, A2 => n74, ZN => mask00(19));
   U47 : NAND2_X1 port map( A1 => n45, A2 => n53, ZN => mask08_19_port);
   U133 : NAND2_X1 port map( A1 => n76, A2 => n55, ZN => mask00(17));
   U49 : NAND2_X1 port map( A1 => n37, A2 => n47, ZN => mask08_17_port);
   U120 : NAND2_X1 port map( A1 => n81, A2 => n72, ZN => mask00(21));
   U44 : NAND2_X1 port map( A1 => n43, A2 => n51, ZN => mask08_21_port);
   U75 : AOI21_X1 port map( B1 => A(30), B2 => n2, A => mask16_17_port, ZN => 
                           n90);
   U27 : NAND2_X1 port map( A1 => n63, A2 => n3, ZN => mask08_37_port);
   U73 : AOI21_X1 port map( B1 => A(31), B2 => n2, A => mask16_17_port, ZN => 
                           n89);
   U26 : NAND2_X1 port map( A1 => n62, A2 => n3, ZN => mask08_38_port);
   U126 : AND2_X1 port map( A1 => sel(0), A2 => A(1), ZN => mask00(1));
   U19 : INV_X1 port map( A => n55, ZN => mask16_1_port);
   U46 : INV_X1 port map( A => n79, ZN => mask08_1_port);
   U69 : AND2_X1 port map( A1 => sel(0), A2 => A(5), ZN => mask00(5));
   U53 : INV_X1 port map( A => n81, ZN => mask16_5_port);
   U23 : INV_X1 port map( A => n59, ZN => mask08_5_port);
   U71 : AND2_X1 port map( A1 => sel(0), A2 => A(3), ZN => mask00(3));
   U55 : INV_X1 port map( A => n83, ZN => mask16_3_port);
   U25 : INV_X1 port map( A => n61, ZN => mask08_3_port);
   U20 : INV_X1 port map( A => n56, ZN => mask16_0_port);
   U57 : INV_X1 port map( A => n85, ZN => mask08_0_port);
   U70 : AND2_X1 port map( A1 => sel(0), A2 => A(4), ZN => mask00(4));
   U54 : INV_X1 port map( A => n82, ZN => mask16_4_port);
   U24 : INV_X1 port map( A => n60, ZN => mask08_4_port);
   U95 : AND2_X1 port map( A1 => sel(0), A2 => A(2), ZN => mask00(2));
   U56 : INV_X1 port map( A => n84, ZN => mask16_2_port);
   U35 : INV_X1 port map( A => n71, ZN => mask08_2_port);
   U68 : AND2_X1 port map( A1 => sel(0), A2 => A(6), ZN => mask00(6));
   U52 : INV_X1 port map( A => n80, ZN => mask16_6_port);
   U22 : INV_X1 port map( A => n58, ZN => mask08_6_port);
   U3 : INV_X1 port map( A => n38, ZN => mask16_8_port);
   U16 : INV_X1 port map( A => n52, ZN => mask16_12_port);
   U18 : INV_X1 port map( A => n54, ZN => mask16_10_port);
   U14 : INV_X1 port map( A => n50, ZN => mask16_14_port);
   U17 : INV_X1 port map( A => n53, ZN => mask16_11_port);
   U2 : INV_X1 port map( A => n37, ZN => mask16_9_port);
   U15 : INV_X1 port map( A => n51, ZN => mask16_13_port);
   U90 : INV_X1 port map( A => n78, ZN => mask16_15_port);
   U80 : INV_X1 port map( A => n93, ZN => mask00(34));
   U84 : INV_X1 port map( A => n95, ZN => mask00(32));
   U76 : INV_X1 port map( A => n91, ZN => mask00(36));
   U82 : INV_X1 port map( A => n94, ZN => mask00(33));
   U88 : INV_X1 port map( A => n96, ZN => mask00(31));
   U78 : INV_X1 port map( A => n92, ZN => mask00(35));
   U74 : INV_X1 port map( A => n90, ZN => mask00(37));
   U72 : INV_X1 port map( A => n89, ZN => mask00(38));
   U4 : INV_X1 port map( A => n57, ZN => mask08_7_port);
   U21 : INV_X1 port map( A => n39, ZN => mask16_7_port);
   U64 : NAND2_X1 port map( A1 => sel(0), A2 => A(7), ZN => n1);
   U65 : NAND2_X1 port map( A1 => n49, A2 => n1, ZN => mask00(7));
   U66 : AND2_X2 port map( A1 => sel(1), A2 => mask16_15_port, ZN => 
                           mask16_17_port);
   U67 : INV_X2 port map( A => mask16_17_port, ZN => n3);
   U86 : BUF_X1 port map( A => n86, Z => n2);
   U87 : AND2_X1 port map( A1 => sel(0), A2 => A(0), ZN => mask00(0));
   U158 : NAND2_X1 port map( A1 => n2, A2 => A(0), ZN => n49);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_simple_booth_add_ext_N16 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_simple_booth_add_ext_N16;

architecture SYN_USE_DEFA_ARCH_NAME of 
   SNPS_CLOCK_GATE_HIGH_simple_booth_add_ext_N16 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net3325 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net3325);
   main_gate : AND2_X1 port map( A1 => net3325, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity piso_r_2_N32 is

   port( Clock, ALOAD : in std_logic;  D : in std_logic_vector (31 downto 0);  
         SO : out std_logic_vector (31 downto 0));

end piso_r_2_N32;

architecture SYN_archi of piso_r_2_N32 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component SDFF_X1
      port( D, SI, SE, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal SO_31_port, SO_30_port, SO_29_port, SO_28_port, SO_27_port, 
      SO_26_port, SO_25_port, SO_24_port, SO_23_port, SO_22_port, SO_21_port, 
      SO_20_port, SO_19_port, SO_18_port, SO_17_port, SO_16_port, SO_15_port, 
      SO_14_port, SO_13_port, SO_12_port, SO_11_port, SO_10_port, SO_9_port, 
      SO_8_port, SO_7_port, SO_6_port, SO_5_port, SO_4_port, SO_3_port, 
      SO_2_port, SO_1_port, SO_0_port, N3, N4, n2, n3_port, n4_port, n5, n6, n7
      , n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22
      , n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33 : std_logic;

begin
   SO <= ( SO_31_port, SO_30_port, SO_29_port, SO_28_port, SO_27_port, 
      SO_26_port, SO_25_port, SO_24_port, SO_23_port, SO_22_port, SO_21_port, 
      SO_20_port, SO_19_port, SO_18_port, SO_17_port, SO_16_port, SO_15_port, 
      SO_14_port, SO_13_port, SO_12_port, SO_11_port, SO_10_port, SO_9_port, 
      SO_8_port, SO_7_port, SO_6_port, SO_5_port, SO_4_port, SO_3_port, 
      SO_2_port, SO_1_port, SO_0_port );
   
   tmp_reg_1_inst : DFF_X1 port map( D => N4, CK => Clock, Q => SO_1_port, QN 
                           => n33);
   tmp_reg_3_inst : SDFF_X1 port map( D => SO_1_port, SI => D(3), SE => ALOAD, 
                           CK => Clock, Q => SO_3_port, QN => n32);
   tmp_reg_5_inst : SDFF_X1 port map( D => SO_3_port, SI => D(5), SE => ALOAD, 
                           CK => Clock, Q => SO_5_port, QN => n31);
   tmp_reg_7_inst : SDFF_X1 port map( D => SO_5_port, SI => D(7), SE => ALOAD, 
                           CK => Clock, Q => SO_7_port, QN => n30);
   tmp_reg_9_inst : SDFF_X1 port map( D => SO_7_port, SI => D(9), SE => ALOAD, 
                           CK => Clock, Q => SO_9_port, QN => n29);
   tmp_reg_11_inst : SDFF_X1 port map( D => SO_9_port, SI => D(11), SE => ALOAD
                           , CK => Clock, Q => SO_11_port, QN => n28);
   tmp_reg_13_inst : SDFF_X1 port map( D => SO_11_port, SI => D(13), SE => 
                           ALOAD, CK => Clock, Q => SO_13_port, QN => n27);
   tmp_reg_15_inst : SDFF_X1 port map( D => SO_13_port, SI => D(15), SE => 
                           ALOAD, CK => Clock, Q => SO_15_port, QN => n26);
   tmp_reg_17_inst : SDFF_X1 port map( D => SO_15_port, SI => D(17), SE => 
                           ALOAD, CK => Clock, Q => SO_17_port, QN => n25);
   tmp_reg_19_inst : SDFF_X1 port map( D => SO_17_port, SI => D(19), SE => 
                           ALOAD, CK => Clock, Q => SO_19_port, QN => n24);
   tmp_reg_21_inst : SDFF_X1 port map( D => SO_19_port, SI => D(21), SE => 
                           ALOAD, CK => Clock, Q => SO_21_port, QN => n23);
   tmp_reg_23_inst : SDFF_X1 port map( D => SO_21_port, SI => D(23), SE => 
                           ALOAD, CK => Clock, Q => SO_23_port, QN => n22);
   tmp_reg_25_inst : SDFF_X1 port map( D => SO_23_port, SI => D(25), SE => 
                           ALOAD, CK => Clock, Q => SO_25_port, QN => n21);
   tmp_reg_27_inst : SDFF_X1 port map( D => SO_25_port, SI => D(27), SE => 
                           ALOAD, CK => Clock, Q => SO_27_port, QN => n20);
   tmp_reg_29_inst : SDFF_X1 port map( D => SO_27_port, SI => D(29), SE => 
                           ALOAD, CK => Clock, Q => SO_29_port, QN => n19);
   tmp_reg_31_inst : SDFF_X1 port map( D => SO_29_port, SI => D(31), SE => 
                           ALOAD, CK => Clock, Q => SO_31_port, QN => n18);
   tmp_reg_0_inst : DFF_X1 port map( D => N3, CK => Clock, Q => SO_0_port, QN 
                           => n17);
   tmp_reg_2_inst : SDFF_X1 port map( D => SO_0_port, SI => D(2), SE => ALOAD, 
                           CK => Clock, Q => SO_2_port, QN => n16);
   tmp_reg_4_inst : SDFF_X1 port map( D => SO_2_port, SI => D(4), SE => ALOAD, 
                           CK => Clock, Q => SO_4_port, QN => n15);
   tmp_reg_6_inst : SDFF_X1 port map( D => SO_4_port, SI => D(6), SE => ALOAD, 
                           CK => Clock, Q => SO_6_port, QN => n14);
   tmp_reg_8_inst : SDFF_X1 port map( D => SO_6_port, SI => D(8), SE => ALOAD, 
                           CK => Clock, Q => SO_8_port, QN => n13);
   tmp_reg_10_inst : SDFF_X1 port map( D => SO_8_port, SI => D(10), SE => ALOAD
                           , CK => Clock, Q => SO_10_port, QN => n12);
   tmp_reg_12_inst : SDFF_X1 port map( D => SO_10_port, SI => D(12), SE => 
                           ALOAD, CK => Clock, Q => SO_12_port, QN => n11);
   tmp_reg_14_inst : SDFF_X1 port map( D => SO_12_port, SI => D(14), SE => 
                           ALOAD, CK => Clock, Q => SO_14_port, QN => n10);
   tmp_reg_16_inst : SDFF_X1 port map( D => SO_14_port, SI => D(16), SE => 
                           ALOAD, CK => Clock, Q => SO_16_port, QN => n9);
   tmp_reg_18_inst : SDFF_X1 port map( D => SO_16_port, SI => D(18), SE => 
                           ALOAD, CK => Clock, Q => SO_18_port, QN => n8);
   tmp_reg_20_inst : SDFF_X1 port map( D => SO_18_port, SI => D(20), SE => 
                           ALOAD, CK => Clock, Q => SO_20_port, QN => n7);
   tmp_reg_22_inst : SDFF_X1 port map( D => SO_20_port, SI => D(22), SE => 
                           ALOAD, CK => Clock, Q => SO_22_port, QN => n6);
   tmp_reg_24_inst : SDFF_X1 port map( D => SO_22_port, SI => D(24), SE => 
                           ALOAD, CK => Clock, Q => SO_24_port, QN => n5);
   tmp_reg_26_inst : SDFF_X1 port map( D => SO_24_port, SI => D(26), SE => 
                           ALOAD, CK => Clock, Q => SO_26_port, QN => n4_port);
   tmp_reg_28_inst : SDFF_X1 port map( D => SO_26_port, SI => D(28), SE => 
                           ALOAD, CK => Clock, Q => SO_28_port, QN => n3_port);
   tmp_reg_30_inst : SDFF_X1 port map( D => SO_28_port, SI => D(30), SE => 
                           ALOAD, CK => Clock, Q => SO_30_port, QN => n2);
   U3 : AND2_X1 port map( A1 => ALOAD, A2 => D(1), ZN => N4);
   U4 : AND2_X1 port map( A1 => ALOAD, A2 => D(0), ZN => N3);

end SYN_archi;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity shift_N9_0 is

   port( Clock, ALOAD : in std_logic;  D : in std_logic_vector (8 downto 0);  
         SO : out std_logic);

end shift_N9_0;

architecture SYN_archi of shift_N9_0 is

   component SDFF_X2
      port( D, SI, SE, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component SDFF_X1
      port( D, SI, SE, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal tmp_8_port, tmp_7_port, tmp_6_port, tmp_5_port, tmp_4_port, 
      tmp_3_port, tmp_2_port, tmp_1_port, N11, n3, n4, n5, n6, n7, n8, n9, n10,
      n1 : std_logic;

begin
   
   tmp_reg_8_inst : DFF_X1 port map( D => N11, CK => Clock, Q => tmp_8_port, QN
                           => n10);
   tmp_reg_7_inst : SDFF_X1 port map( D => tmp_8_port, SI => D(7), SE => ALOAD,
                           CK => Clock, Q => tmp_7_port, QN => n9);
   tmp_reg_6_inst : SDFF_X1 port map( D => tmp_7_port, SI => D(6), SE => ALOAD,
                           CK => Clock, Q => tmp_6_port, QN => n8);
   tmp_reg_5_inst : SDFF_X1 port map( D => tmp_6_port, SI => D(5), SE => ALOAD,
                           CK => Clock, Q => tmp_5_port, QN => n7);
   tmp_reg_4_inst : SDFF_X1 port map( D => tmp_5_port, SI => D(4), SE => ALOAD,
                           CK => Clock, Q => tmp_4_port, QN => n6);
   tmp_reg_3_inst : SDFF_X1 port map( D => tmp_4_port, SI => D(3), SE => ALOAD,
                           CK => Clock, Q => tmp_3_port, QN => n5);
   tmp_reg_2_inst : SDFF_X1 port map( D => tmp_3_port, SI => D(2), SE => ALOAD,
                           CK => Clock, Q => tmp_2_port, QN => n4);
   tmp_reg_1_inst : SDFF_X1 port map( D => tmp_2_port, SI => D(1), SE => ALOAD,
                           CK => Clock, Q => tmp_1_port, QN => n3);
   U3 : AND2_X1 port map( A1 => ALOAD, A2 => D(8), ZN => N11);
   tmp_reg_0_inst : SDFF_X2 port map( D => tmp_1_port, SI => D(0), SE => ALOAD,
                           CK => Clock, Q => SO, QN => n1);

end SYN_archi;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity booth_encoder_0 is

   port( B_in : in std_logic_vector (2 downto 0);  A_out : out std_logic_vector
         (2 downto 0));

end booth_encoder_0;

architecture SYN_bhe of booth_encoder_0 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal A_out_2_port, A_out_0_port, n3, n4 : std_logic;

begin
   A_out <= ( A_out_2_port, B_in(2), A_out_0_port );
   
   U3 : INV_X1 port map( A => B_in(1), ZN => n3);
   U4 : INV_X1 port map( A => B_in(2), ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n3, ZN => A_out_2_port);
   U6 : NOR2_X1 port map( A1 => B_in(1), A2 => n4, ZN => A_out_0_port);

end SYN_bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity carry_sel_gen_N4_0 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end carry_sel_gen_N4_0;

architecture SYN_STRUCTURAL of carry_sel_gen_N4_0 is

   component mux21_SIZE4_0
      port( IN0, IN1 : in std_logic_vector (3 downto 0);  CTRL : in std_logic; 
            OUT1 : out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_N4_0
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic0_port, n5, nocarry_sum_to_mux_3_port, 
      nocarry_sum_to_mux_2_port, nocarry_sum_to_mux_1_port, 
      nocarry_sum_to_mux_0_port, n1, n2, n3, n4, net48716 : std_logic;

begin
   
   X_Logic0_port <= '0';
   rca_nocarry : RCA_N4_0 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           nocarry_sum_to_mux_3_port, S(2) => 
                           nocarry_sum_to_mux_2_port, S(1) => 
                           nocarry_sum_to_mux_1_port, S(0) => 
                           nocarry_sum_to_mux_0_port, Co => net48716);
   outmux : mux21_SIZE4_0 port map( IN0(3) => nocarry_sum_to_mux_3_port, IN0(2)
                           => nocarry_sum_to_mux_2_port, IN0(1) => 
                           nocarry_sum_to_mux_1_port, IN0(0) => 
                           nocarry_sum_to_mux_0_port, IN1(3) => n1, IN1(2) => 
                           n2, IN1(1) => n3, IN1(0) => n4, CTRL => n5, OUT1(3) 
                           => S(3), OUT1(2) => S(2), OUT1(1) => S(1), OUT1(0) 
                           => S(0));
   n1 <= '0';
   n2 <= '0';
   n3 <= '0';
   n4 <= '0';
   n5 <= '0';

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_0 is

   port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic);

end pg_0;

architecture SYN_beh of pg_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U3 : AOI21_X1 port map( B1 => g_prec, B2 => p, A => g, ZN => n2);
   U1 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);
   U2 : INV_X1 port map( A => n2, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity g_0 is

   port( g, p, g_prec : in std_logic;  g_out : out std_logic);

end g_0;

architecture SYN_beh of g_0 is

begin
   g_out <= g;

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_0 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_0;

architecture SYN_beh of pg_net_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity logic_unit_SIZE32 is

   port( IN1, IN2 : in std_logic_vector (31 downto 0);  CTRL : in 
         std_logic_vector (1 downto 0);  OUT1 : out std_logic_vector (31 downto
         0));

end logic_unit_SIZE32;

architecture SYN_Bhe of logic_unit_SIZE32 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X4
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, 
      n18, n19, n20, n21, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34
      , n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, 
      n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63
      , n64, n65, n1, n2, n22, n23 : std_logic;

begin
   
   U8 : AOI21_X1 port map( B1 => n3, B2 => n8, A => n9, ZN => OUT1(7));
   U32 : AOI21_X1 port map( B1 => n3, B2 => n24, A => n25, ZN => OUT1(29));
   U50 : AOI21_X1 port map( B1 => n3, B2 => n36, A => n37, ZN => OUT1(23));
   U77 : AOI21_X1 port map( B1 => n3, B2 => n54, A => n55, ZN => OUT1(15));
   U67 : AOI21_X1 port map( B1 => IN2(19), B2 => IN1(19), A => CTRL(0), ZN => 
                           n46);
   U66 : OAI22_X1 port map( A1 => IN1(19), A2 => IN2(19), B1 => n3, B2 => n46, 
                           ZN => n47);
   U65 : AOI21_X1 port map( B1 => n3, B2 => n46, A => n47, ZN => OUT1(19));
   U70 : AOI21_X1 port map( B1 => IN2(18), B2 => IN1(18), A => CTRL(0), ZN => 
                           n48);
   U69 : OAI22_X1 port map( A1 => IN1(18), A2 => IN2(18), B1 => n3, B2 => n48, 
                           ZN => n49);
   U68 : AOI21_X1 port map( B1 => n3, B2 => n48, A => n49, ZN => OUT1(18));
   U73 : AOI21_X1 port map( B1 => IN2(17), B2 => IN1(17), A => CTRL(0), ZN => 
                           n50);
   U72 : OAI22_X1 port map( A1 => IN1(17), A2 => IN2(17), B1 => n3, B2 => n50, 
                           ZN => n51);
   U71 : AOI21_X1 port map( B1 => n3, B2 => n50, A => n51, ZN => OUT1(17));
   U46 : AOI21_X1 port map( B1 => IN2(25), B2 => IN1(25), A => CTRL(0), ZN => 
                           n32);
   U45 : OAI22_X1 port map( A1 => IN1(25), A2 => IN2(25), B1 => n3, B2 => n32, 
                           ZN => n33);
   U44 : AOI21_X1 port map( B1 => n3, B2 => n32, A => n33, ZN => OUT1(25));
   U40 : AOI21_X1 port map( B1 => IN2(27), B2 => IN1(27), A => CTRL(0), ZN => 
                           n28);
   U39 : OAI22_X1 port map( A1 => IN1(27), A2 => IN2(27), B1 => n3, B2 => n28, 
                           ZN => n29);
   U38 : AOI21_X1 port map( B1 => n3, B2 => n28, A => n29, ZN => OUT1(27));
   U43 : AOI21_X1 port map( B1 => IN2(26), B2 => IN1(26), A => CTRL(0), ZN => 
                           n30);
   U42 : OAI22_X1 port map( A1 => IN1(26), A2 => IN2(26), B1 => n3, B2 => n30, 
                           ZN => n31);
   U41 : AOI21_X1 port map( B1 => n3, B2 => n30, A => n31, ZN => OUT1(26));
   U28 : AOI21_X1 port map( B1 => IN2(30), B2 => IN1(30), A => CTRL(0), ZN => 
                           n20);
   U27 : OAI22_X1 port map( A1 => IN1(30), A2 => IN2(30), B1 => n3, B2 => n20, 
                           ZN => n21);
   U26 : AOI21_X1 port map( B1 => n3, B2 => n20, A => n21, ZN => OUT1(30));
   U49 : AOI21_X1 port map( B1 => IN2(24), B2 => IN1(24), A => CTRL(0), ZN => 
                           n34);
   U48 : OAI22_X1 port map( A1 => IN1(24), A2 => IN2(24), B1 => n3, B2 => n34, 
                           ZN => n35);
   U47 : AOI21_X1 port map( B1 => n3, B2 => n34, A => n35, ZN => OUT1(24));
   U55 : AOI21_X1 port map( B1 => IN2(22), B2 => IN1(22), A => CTRL(0), ZN => 
                           n38);
   U54 : OAI22_X1 port map( A1 => IN1(22), A2 => IN2(22), B1 => n3, B2 => n38, 
                           ZN => n39);
   U53 : AOI21_X1 port map( B1 => n3, B2 => n38, A => n39, ZN => OUT1(22));
   U58 : AOI21_X1 port map( B1 => IN2(21), B2 => IN1(21), A => CTRL(0), ZN => 
                           n40);
   U57 : OAI22_X1 port map( A1 => IN1(21), A2 => IN2(21), B1 => n3, B2 => n40, 
                           ZN => n41);
   U56 : AOI21_X1 port map( B1 => n3, B2 => n40, A => n41, ZN => OUT1(21));
   U25 : AOI21_X1 port map( B1 => IN2(31), B2 => IN1(31), A => CTRL(0), ZN => 
                           n18);
   U24 : OAI22_X1 port map( A1 => IN1(31), A2 => IN2(31), B1 => n3, B2 => n18, 
                           ZN => n19);
   U23 : AOI21_X1 port map( B1 => n3, B2 => n18, A => n19, ZN => OUT1(31));
   U61 : AOI21_X1 port map( B1 => IN2(20), B2 => IN1(20), A => CTRL(0), ZN => 
                           n42);
   U60 : OAI22_X1 port map( A1 => IN1(20), A2 => IN2(20), B1 => n3, B2 => n42, 
                           ZN => n43);
   U59 : AOI21_X1 port map( B1 => n3, B2 => n42, A => n43, ZN => OUT1(20));
   U37 : AOI21_X1 port map( B1 => IN2(28), B2 => IN1(28), A => CTRL(0), ZN => 
                           n26);
   U36 : OAI22_X1 port map( A1 => IN1(28), A2 => IN2(28), B1 => n3, B2 => n26, 
                           ZN => n27);
   U35 : AOI21_X1 port map( B1 => n3, B2 => n26, A => n27, ZN => OUT1(28));
   U82 : AOI21_X1 port map( B1 => IN2(14), B2 => IN1(14), A => CTRL(0), ZN => 
                           n56);
   U81 : OAI22_X1 port map( A1 => IN1(14), A2 => IN2(14), B1 => n3, B2 => n56, 
                           ZN => n57);
   U80 : AOI21_X1 port map( B1 => n3, B2 => n56, A => n57, ZN => OUT1(14));
   U22 : AOI21_X1 port map( B1 => IN2(3), B2 => IN1(3), A => CTRL(0), ZN => n16
                           );
   U21 : OAI22_X1 port map( A1 => IN1(3), A2 => IN2(3), B1 => n3, B2 => n16, ZN
                           => n17);
   U20 : AOI21_X1 port map( B1 => n3, B2 => n16, A => n17, ZN => OUT1(3));
   U86 : AOI21_X1 port map( B1 => n3, B2 => n60, A => n61, ZN => OUT1(12));
   U89 : AOI21_X1 port map( B1 => n3, B2 => n62, A => n63, ZN => OUT1(11));
   U76 : AOI21_X1 port map( B1 => IN2(16), B2 => IN1(16), A => CTRL(0), ZN => 
                           n52);
   U75 : OAI22_X1 port map( A1 => IN1(16), A2 => IN2(16), B1 => n3, B2 => n52, 
                           ZN => n53);
   U74 : AOI21_X1 port map( B1 => n3, B2 => n52, A => n53, ZN => OUT1(16));
   U83 : AOI21_X1 port map( B1 => n3, B2 => n58, A => n59, ZN => OUT1(13));
   U2 : AOI21_X1 port map( B1 => n3, B2 => n4, A => n5, ZN => OUT1(9));
   U11 : AOI21_X1 port map( B1 => n3, B2 => n10, A => n11, ZN => OUT1(6));
   U7 : AOI21_X1 port map( B1 => IN2(8), B2 => IN1(8), A => CTRL(0), ZN => n6);
   U6 : OAI22_X1 port map( A1 => IN1(8), A2 => IN2(8), B1 => n3, B2 => n6, ZN 
                           => n7);
   U5 : AOI21_X1 port map( B1 => n3, B2 => n6, A => n7, ZN => OUT1(8));
   U92 : AOI21_X1 port map( B1 => n3, B2 => n64, A => n65, ZN => OUT1(10));
   U14 : AOI21_X1 port map( B1 => n3, B2 => n12, A => n13, ZN => OUT1(5));
   U19 : AOI21_X1 port map( B1 => IN2(4), B2 => IN1(4), A => CTRL(0), ZN => n14
                           );
   U18 : OAI22_X1 port map( A1 => IN1(4), A2 => IN2(4), B1 => n3, B2 => n14, ZN
                           => n15);
   U17 : AOI21_X1 port map( B1 => n3, B2 => n14, A => n15, ZN => OUT1(4));
   U62 : AOI21_X1 port map( B1 => n3, B2 => n44, A => n45, ZN => OUT1(1));
   U3 : AOI21_X1 port map( B1 => IN1(0), B2 => IN2(0), A => CTRL(0), ZN => n1);
   U4 : OAI22_X1 port map( A1 => IN2(0), A2 => IN1(0), B1 => n3, B2 => n1, ZN 
                           => n2);
   U9 : AOI21_X1 port map( B1 => n3, B2 => n1, A => n2, ZN => OUT1(0));
   U10 : AOI21_X1 port map( B1 => IN1(2), B2 => IN2(2), A => CTRL(0), ZN => n22
                           );
   U12 : OAI22_X1 port map( A1 => IN2(2), A2 => IN1(2), B1 => n3, B2 => n22, ZN
                           => n23);
   U13 : AOI21_X1 port map( B1 => n3, B2 => n22, A => n23, ZN => OUT1(2));
   U15 : INV_X4 port map( A => CTRL(1), ZN => n3);
   U16 : OAI22_X1 port map( A1 => IN1(10), A2 => IN2(10), B1 => n3, B2 => n64, 
                           ZN => n65);
   U29 : AOI21_X1 port map( B1 => IN2(10), B2 => IN1(10), A => CTRL(0), ZN => 
                           n64);
   U30 : OAI22_X1 port map( A1 => IN1(29), A2 => IN2(29), B1 => n3, B2 => n24, 
                           ZN => n25);
   U31 : AOI21_X1 port map( B1 => IN2(29), B2 => IN1(29), A => CTRL(0), ZN => 
                           n24);
   U33 : OAI22_X1 port map( A1 => IN1(12), A2 => IN2(12), B1 => n3, B2 => n60, 
                           ZN => n61);
   U34 : AOI21_X1 port map( B1 => IN2(12), B2 => IN1(12), A => CTRL(0), ZN => 
                           n60);
   U51 : OAI22_X1 port map( A1 => IN1(23), A2 => IN2(23), B1 => n3, B2 => n36, 
                           ZN => n37);
   U52 : AOI21_X1 port map( B1 => IN2(23), B2 => IN1(23), A => CTRL(0), ZN => 
                           n36);
   U63 : OAI22_X1 port map( A1 => IN1(11), A2 => IN2(11), B1 => n3, B2 => n62, 
                           ZN => n63);
   U64 : AOI21_X1 port map( B1 => IN2(11), B2 => IN1(11), A => CTRL(0), ZN => 
                           n62);
   U78 : OAI22_X1 port map( A1 => IN1(15), A2 => IN2(15), B1 => n3, B2 => n54, 
                           ZN => n55);
   U79 : AOI21_X1 port map( B1 => IN2(15), B2 => IN1(15), A => CTRL(0), ZN => 
                           n54);
   U84 : OAI22_X1 port map( A1 => IN1(7), A2 => IN2(7), B1 => n3, B2 => n8, ZN 
                           => n9);
   U85 : AOI21_X1 port map( B1 => IN2(7), B2 => IN1(7), A => CTRL(0), ZN => n8)
                           ;
   U87 : OAI22_X1 port map( A1 => IN1(6), A2 => IN2(6), B1 => n3, B2 => n10, ZN
                           => n11);
   U88 : AOI21_X1 port map( B1 => IN2(6), B2 => IN1(6), A => CTRL(0), ZN => n10
                           );
   U90 : OAI22_X1 port map( A1 => IN1(9), A2 => IN2(9), B1 => n3, B2 => n4, ZN 
                           => n5);
   U91 : AOI21_X1 port map( B1 => IN2(9), B2 => IN1(9), A => CTRL(0), ZN => n4)
                           ;
   U93 : OAI22_X1 port map( A1 => IN1(13), A2 => IN2(13), B1 => n3, B2 => n58, 
                           ZN => n59);
   U94 : AOI21_X1 port map( B1 => IN2(13), B2 => IN1(13), A => CTRL(0), ZN => 
                           n58);
   U95 : OAI22_X1 port map( A1 => IN1(5), A2 => IN2(5), B1 => n3, B2 => n12, ZN
                           => n13);
   U96 : AOI21_X1 port map( B1 => IN2(5), B2 => IN1(5), A => CTRL(0), ZN => n12
                           );
   U97 : OAI22_X1 port map( A1 => IN1(1), A2 => IN2(1), B1 => n3, B2 => n44, ZN
                           => n45);
   U98 : AOI21_X1 port map( B1 => IN2(1), B2 => IN1(1), A => CTRL(0), ZN => n44
                           );

end SYN_Bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity shifter is

   port( A : in std_logic_vector (31 downto 0);  B : in std_logic_vector (4 
         downto 0);  LOGIC_ARITH, LEFT_RIGHT : in std_logic;  OUTPUT : out 
         std_logic_vector (31 downto 0));

end shifter;

architecture SYN_struct of shifter is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component shift_thirdLevel
      port( sel : in std_logic_vector (2 downto 0);  A : in std_logic_vector 
            (38 downto 0);  Y : out std_logic_vector (31 downto 0));
   end component;
   
   component shift_secondLevel
      port( sel : in std_logic_vector (1 downto 0);  mask00, mask08, mask16 : 
            in std_logic_vector (38 downto 0);  Y : out std_logic_vector (38 
            downto 0));
   end component;
   
   component shift_firstLevel
      port( A : in std_logic_vector (31 downto 0);  sel : in std_logic_vector 
            (1 downto 0);  mask00, mask08, mask16 : out std_logic_vector (38 
            downto 0));
   end component;
   
   signal s3_2_port, s3_1_port, s3_0_port, m0_38_port, m0_37_port, m0_36_port, 
      m0_35_port, m0_34_port, m0_33_port, m0_32_port, m0_31_port, m0_30_port, 
      m0_29_port, m0_28_port, m0_27_port, m0_26_port, m0_25_port, m0_24_port, 
      m0_23_port, m0_22_port, m0_21_port, m0_20_port, m0_19_port, m0_18_port, 
      m0_17_port, m0_16_port, m0_15_port, m0_14_port, m0_13_port, m0_12_port, 
      m0_11_port, m0_10_port, m0_9_port, m0_8_port, m0_7_port, m0_6_port, 
      m0_5_port, m0_4_port, m0_3_port, m0_2_port, m0_1_port, m0_0_port, 
      m8_38_port, m8_37_port, m8_36_port, m8_35_port, m8_34_port, m8_33_port, 
      m8_32_port, m8_31_port, m8_30_port, m8_29_port, m8_28_port, m8_27_port, 
      m8_26_port, m8_25_port, m8_24_port, m8_23_port, m8_22_port, m8_21_port, 
      m8_20_port, m8_19_port, m8_18_port, m8_17_port, m8_16_port, m8_15_port, 
      m8_14_port, m8_13_port, m8_12_port, m8_11_port, m8_10_port, m8_9_port, 
      m8_8_port, m8_7_port, m8_6_port, m8_5_port, m8_4_port, m8_3_port, 
      m8_2_port, m8_1_port, m8_0_port, m16_38_port, m16_37_port, m16_36_port, 
      m16_35_port, m16_34_port, m16_33_port, m16_32_port, m16_31_port, 
      m16_30_port, m16_29_port, m16_28_port, m16_27_port, m16_26_port, 
      m16_25_port, m16_24_port, m16_23_port, m16_15_port, m16_14_port, 
      m16_13_port, m16_12_port, m16_11_port, m16_10_port, m16_9_port, 
      m16_8_port, m16_7_port, m16_6_port, m16_5_port, m16_4_port, m16_3_port, 
      m16_2_port, m16_1_port, m16_0_port, y_38_port, y_37_port, y_36_port, 
      y_35_port, y_34_port, y_33_port, y_32_port, y_31_port, y_30_port, 
      y_29_port, y_28_port, y_27_port, y_26_port, y_25_port, y_24_port, 
      y_23_port, y_22_port, y_21_port, y_20_port, y_19_port, y_18_port, 
      y_17_port, y_16_port, y_15_port, y_14_port, y_13_port, y_12_port, 
      y_11_port, y_10_port, y_9_port, y_8_port, y_7_port, y_6_port, y_5_port, 
      y_4_port, y_3_port, y_2_port, y_1_port, y_0_port, n6, n8, n9, n10, n2, n3
      , n4, n5, n7, n11, n12, n13 : std_logic;

begin
   
   IL : shift_firstLevel port map( A(31) => A(31), A(30) => A(30), A(29) => 
                           A(29), A(28) => A(28), A(27) => A(27), A(26) => 
                           A(26), A(25) => A(25), A(24) => A(24), A(23) => 
                           A(23), A(22) => A(22), A(21) => A(21), A(20) => 
                           A(20), A(19) => A(19), A(18) => A(18), A(17) => 
                           A(17), A(16) => A(16), A(15) => A(15), A(14) => 
                           A(14), A(13) => A(13), A(12) => A(12), A(11) => 
                           A(11), A(10) => A(10), A(9) => A(9), A(8) => A(8), 
                           A(7) => A(7), A(6) => A(6), A(5) => A(5), A(4) => 
                           A(4), A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), sel(1) => LOGIC_ARITH, sel(0) => LEFT_RIGHT
                           , mask00(38) => m0_38_port, mask00(37) => m0_37_port
                           , mask00(36) => m0_36_port, mask00(35) => m0_35_port
                           , mask00(34) => m0_34_port, mask00(33) => m0_33_port
                           , mask00(32) => m0_32_port, mask00(31) => m0_31_port
                           , mask00(30) => m0_30_port, mask00(29) => m0_29_port
                           , mask00(28) => m0_28_port, mask00(27) => m0_27_port
                           , mask00(26) => m0_26_port, mask00(25) => m0_25_port
                           , mask00(24) => m0_24_port, mask00(23) => m0_23_port
                           , mask00(22) => m0_22_port, mask00(21) => m0_21_port
                           , mask00(20) => m0_20_port, mask00(19) => m0_19_port
                           , mask00(18) => m0_18_port, mask00(17) => m0_17_port
                           , mask00(16) => m0_16_port, mask00(15) => m0_15_port
                           , mask00(14) => m0_14_port, mask00(13) => m0_13_port
                           , mask00(12) => m0_12_port, mask00(11) => m0_11_port
                           , mask00(10) => m0_10_port, mask00(9) => m0_9_port, 
                           mask00(8) => m0_8_port, mask00(7) => m0_7_port, 
                           mask00(6) => m0_6_port, mask00(5) => m0_5_port, 
                           mask00(4) => m0_4_port, mask00(3) => m0_3_port, 
                           mask00(2) => m0_2_port, mask00(1) => m0_1_port, 
                           mask00(0) => m0_0_port, mask08(38) => m8_38_port, 
                           mask08(37) => m8_37_port, mask08(36) => m8_36_port, 
                           mask08(35) => m8_35_port, mask08(34) => m8_34_port, 
                           mask08(33) => m8_33_port, mask08(32) => m8_32_port, 
                           mask08(31) => m8_31_port, mask08(30) => m8_30_port, 
                           mask08(29) => m8_29_port, mask08(28) => m8_28_port, 
                           mask08(27) => m8_27_port, mask08(26) => m8_26_port, 
                           mask08(25) => m8_25_port, mask08(24) => m8_24_port, 
                           mask08(23) => m8_23_port, mask08(22) => m8_22_port, 
                           mask08(21) => m8_21_port, mask08(20) => m8_20_port, 
                           mask08(19) => m8_19_port, mask08(18) => m8_18_port, 
                           mask08(17) => m8_17_port, mask08(16) => m8_16_port, 
                           mask08(15) => m8_15_port, mask08(14) => m8_14_port, 
                           mask08(13) => m8_13_port, mask08(12) => m8_12_port, 
                           mask08(11) => m8_11_port, mask08(10) => m8_10_port, 
                           mask08(9) => m8_9_port, mask08(8) => m8_8_port, 
                           mask08(7) => m8_7_port, mask08(6) => m8_6_port, 
                           mask08(5) => m8_5_port, mask08(4) => m8_4_port, 
                           mask08(3) => m8_3_port, mask08(2) => m8_2_port, 
                           mask08(1) => m8_1_port, mask08(0) => m8_0_port, 
                           mask16(38) => m16_38_port, mask16(37) => m16_37_port
                           , mask16(36) => m16_36_port, mask16(35) => 
                           m16_35_port, mask16(34) => m16_34_port, mask16(33) 
                           => m16_33_port, mask16(32) => m16_32_port, 
                           mask16(31) => m16_31_port, mask16(30) => m16_30_port
                           , mask16(29) => m16_29_port, mask16(28) => 
                           m16_28_port, mask16(27) => m16_27_port, mask16(26) 
                           => m16_26_port, mask16(25) => m16_25_port, 
                           mask16(24) => m16_24_port, mask16(23) => m16_23_port
                           , mask16(22) => n4, mask16(21) => n3, mask16(20) => 
                           n5, mask16(19) => n7, mask16(18) => n11, mask16(17) 
                           => n12, mask16(16) => n2, mask16(15) => m16_15_port,
                           mask16(14) => m16_14_port, mask16(13) => m16_13_port
                           , mask16(12) => m16_12_port, mask16(11) => 
                           m16_11_port, mask16(10) => m16_10_port, mask16(9) =>
                           m16_9_port, mask16(8) => m16_8_port, mask16(7) => 
                           m16_7_port, mask16(6) => m16_6_port, mask16(5) => 
                           m16_5_port, mask16(4) => m16_4_port, mask16(3) => 
                           m16_3_port, mask16(2) => m16_2_port, mask16(1) => 
                           m16_1_port, mask16(0) => m16_0_port);
   IIL : shift_secondLevel port map( sel(1) => B(4), sel(0) => B(3), mask00(38)
                           => m0_38_port, mask00(37) => m0_37_port, mask00(36) 
                           => m0_36_port, mask00(35) => m0_35_port, mask00(34) 
                           => m0_34_port, mask00(33) => m0_33_port, mask00(32) 
                           => m0_32_port, mask00(31) => m0_31_port, mask00(30) 
                           => m0_30_port, mask00(29) => m0_29_port, mask00(28) 
                           => m0_28_port, mask00(27) => m0_27_port, mask00(26) 
                           => m0_26_port, mask00(25) => m0_25_port, mask00(24) 
                           => m0_24_port, mask00(23) => m0_23_port, mask00(22) 
                           => m0_22_port, mask00(21) => m0_21_port, mask00(20) 
                           => m0_20_port, mask00(19) => m0_19_port, mask00(18) 
                           => m0_18_port, mask00(17) => m0_17_port, mask00(16) 
                           => m0_16_port, mask00(15) => m0_15_port, mask00(14) 
                           => m0_14_port, mask00(13) => m0_13_port, mask00(12) 
                           => m0_12_port, mask00(11) => m0_11_port, mask00(10) 
                           => m0_10_port, mask00(9) => m0_9_port, mask00(8) => 
                           m0_8_port, mask00(7) => m0_7_port, mask00(6) => 
                           m0_6_port, mask00(5) => m0_5_port, mask00(4) => 
                           m0_4_port, mask00(3) => m0_3_port, mask00(2) => 
                           m0_2_port, mask00(1) => m0_1_port, mask00(0) => 
                           m0_0_port, mask08(38) => m8_38_port, mask08(37) => 
                           m8_37_port, mask08(36) => m8_36_port, mask08(35) => 
                           m8_35_port, mask08(34) => m8_34_port, mask08(33) => 
                           m8_33_port, mask08(32) => m8_32_port, mask08(31) => 
                           m8_31_port, mask08(30) => m8_30_port, mask08(29) => 
                           m8_29_port, mask08(28) => m8_28_port, mask08(27) => 
                           m8_27_port, mask08(26) => m8_26_port, mask08(25) => 
                           m8_25_port, mask08(24) => m8_24_port, mask08(23) => 
                           m8_23_port, mask08(22) => m8_22_port, mask08(21) => 
                           m8_21_port, mask08(20) => m8_20_port, mask08(19) => 
                           m8_19_port, mask08(18) => m8_18_port, mask08(17) => 
                           m8_17_port, mask08(16) => m8_16_port, mask08(15) => 
                           m8_15_port, mask08(14) => m8_14_port, mask08(13) => 
                           m8_13_port, mask08(12) => m8_12_port, mask08(11) => 
                           m8_11_port, mask08(10) => m8_10_port, mask08(9) => 
                           m8_9_port, mask08(8) => m8_8_port, mask08(7) => 
                           m8_7_port, mask08(6) => m8_6_port, mask08(5) => 
                           m8_5_port, mask08(4) => m8_4_port, mask08(3) => 
                           m8_3_port, mask08(2) => m8_2_port, mask08(1) => 
                           m8_1_port, mask08(0) => m8_0_port, mask16(38) => 
                           m16_38_port, mask16(37) => m16_37_port, mask16(36) 
                           => m16_36_port, mask16(35) => m16_35_port, 
                           mask16(34) => m16_34_port, mask16(33) => m16_33_port
                           , mask16(32) => m16_32_port, mask16(31) => 
                           m16_31_port, mask16(30) => m16_30_port, mask16(29) 
                           => m16_29_port, mask16(28) => m16_28_port, 
                           mask16(27) => m16_27_port, mask16(26) => m16_26_port
                           , mask16(25) => m16_25_port, mask16(24) => 
                           m16_24_port, mask16(23) => m16_23_port, mask16(22) 
                           => n4, mask16(21) => n3, mask16(20) => n5, 
                           mask16(19) => n7, mask16(18) => n11, mask16(17) => 
                           n12, mask16(16) => n2, mask16(15) => m16_15_port, 
                           mask16(14) => m16_14_port, mask16(13) => m16_13_port
                           , mask16(12) => m16_12_port, mask16(11) => 
                           m16_11_port, mask16(10) => m16_10_port, mask16(9) =>
                           m16_9_port, mask16(8) => m16_8_port, mask16(7) => 
                           m16_7_port, mask16(6) => m16_6_port, mask16(5) => 
                           m16_5_port, mask16(4) => m16_4_port, mask16(3) => 
                           m16_3_port, mask16(2) => m16_2_port, mask16(1) => 
                           m16_1_port, mask16(0) => m16_0_port, Y(38) => 
                           y_38_port, Y(37) => y_37_port, Y(36) => y_36_port, 
                           Y(35) => y_35_port, Y(34) => y_34_port, Y(33) => 
                           y_33_port, Y(32) => y_32_port, Y(31) => y_31_port, 
                           Y(30) => y_30_port, Y(29) => y_29_port, Y(28) => 
                           y_28_port, Y(27) => y_27_port, Y(26) => y_26_port, 
                           Y(25) => y_25_port, Y(24) => y_24_port, Y(23) => 
                           y_23_port, Y(22) => y_22_port, Y(21) => y_21_port, 
                           Y(20) => y_20_port, Y(19) => y_19_port, Y(18) => 
                           y_18_port, Y(17) => y_17_port, Y(16) => y_16_port, 
                           Y(15) => y_15_port, Y(14) => y_14_port, Y(13) => 
                           y_13_port, Y(12) => y_12_port, Y(11) => y_11_port, 
                           Y(10) => y_10_port, Y(9) => y_9_port, Y(8) => 
                           y_8_port, Y(7) => y_7_port, Y(6) => y_6_port, Y(5) 
                           => y_5_port, Y(4) => y_4_port, Y(3) => y_3_port, 
                           Y(2) => y_2_port, Y(1) => y_1_port, Y(0) => y_0_port
                           );
   IIIL : shift_thirdLevel port map( sel(2) => s3_2_port, sel(1) => s3_1_port, 
                           sel(0) => s3_0_port, A(38) => y_38_port, A(37) => 
                           y_37_port, A(36) => y_36_port, A(35) => y_35_port, 
                           A(34) => y_34_port, A(33) => y_33_port, A(32) => 
                           y_32_port, A(31) => y_31_port, A(30) => y_30_port, 
                           A(29) => y_29_port, A(28) => y_28_port, A(27) => 
                           y_27_port, A(26) => y_26_port, A(25) => y_25_port, 
                           A(24) => y_24_port, A(23) => y_23_port, A(22) => 
                           y_22_port, A(21) => y_21_port, A(20) => y_20_port, 
                           A(19) => y_19_port, A(18) => y_18_port, A(17) => 
                           y_17_port, A(16) => y_16_port, A(15) => y_15_port, 
                           A(14) => y_14_port, A(13) => y_13_port, A(12) => 
                           y_12_port, A(11) => y_11_port, A(10) => y_10_port, 
                           A(9) => y_9_port, A(8) => y_8_port, A(7) => y_7_port
                           , A(6) => y_6_port, A(5) => y_5_port, A(4) => 
                           y_4_port, A(3) => y_3_port, A(2) => y_2_port, A(1) 
                           => y_1_port, A(0) => y_0_port, Y(31) => OUTPUT(31), 
                           Y(30) => OUTPUT(30), Y(29) => OUTPUT(29), Y(28) => 
                           OUTPUT(28), Y(27) => OUTPUT(27), Y(26) => OUTPUT(26)
                           , Y(25) => OUTPUT(25), Y(24) => OUTPUT(24), Y(23) =>
                           OUTPUT(23), Y(22) => OUTPUT(22), Y(21) => OUTPUT(21)
                           , Y(20) => OUTPUT(20), Y(19) => OUTPUT(19), Y(18) =>
                           OUTPUT(18), Y(17) => OUTPUT(17), Y(16) => OUTPUT(16)
                           , Y(15) => OUTPUT(15), Y(14) => OUTPUT(14), Y(13) =>
                           OUTPUT(13), Y(12) => OUTPUT(12), Y(11) => OUTPUT(11)
                           , Y(10) => OUTPUT(10), Y(9) => OUTPUT(9), Y(8) => 
                           OUTPUT(8), Y(7) => OUTPUT(7), Y(6) => OUTPUT(6), 
                           Y(5) => OUTPUT(5), Y(4) => OUTPUT(4), Y(3) => 
                           OUTPUT(3), Y(2) => OUTPUT(2), Y(1) => OUTPUT(1), 
                           Y(0) => OUTPUT(0));
   U8 : OR2_X1 port map( A1 => LOGIC_ARITH, A2 => LEFT_RIGHT, ZN => n6);
   U1 : INV_X1 port map( A => B(0), ZN => n10);
   U2 : INV_X1 port map( A => B(2), ZN => n8);
   U3 : INV_X1 port map( A => B(1), ZN => n9);
   U4 : INV_X1 port map( A => LEFT_RIGHT, ZN => n13);
   U5 : AOI22_X1 port map( A1 => B(1), A2 => n6, B1 => n13, B2 => n9, ZN => 
                           s3_1_port);
   U6 : AOI22_X1 port map( A1 => B(2), A2 => n6, B1 => n13, B2 => n8, ZN => 
                           s3_2_port);
   U7 : AOI22_X1 port map( A1 => B(0), A2 => n6, B1 => n13, B2 => n10, ZN => 
                           s3_0_port);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity comparator_M32 is

   port( V : in std_logic;  SUM : in std_logic_vector (31 downto 0);  sel : in 
         std_logic_vector (2 downto 0);  sign : in std_logic;  S : out 
         std_logic;  C_BAR : in std_logic);

end comparator_M32;

architecture SYN_BEHAVIORAL of comparator_M32 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n8, n6, n1, n2, n3, n4, n5, n7, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40 : std_logic;

begin
   
   U1 : NOR4_X1 port map( A1 => SUM(6), A2 => SUM(5), A3 => SUM(3), A4 => 
                           SUM(4), ZN => n25);
   U2 : AND2_X1 port map( A1 => n16, A2 => n17, ZN => n1);
   U3 : CLKBUF_X1 port map( A => SUM(31), Z => n2);
   U4 : INV_X1 port map( A => n40, ZN => n14);
   U5 : INV_X1 port map( A => sel(2), ZN => n13);
   U6 : INV_X1 port map( A => n12, ZN => n11);
   U7 : INV_X1 port map( A => sign, ZN => n18);
   U8 : OR2_X1 port map( A1 => n6, A2 => sel(0), ZN => n15);
   U9 : AND4_X1 port map( A1 => n23, A2 => n25, A3 => n24, A4 => n26, ZN => n39
                           );
   U10 : INV_X1 port map( A => SUM(9), ZN => n26);
   U11 : INV_X1 port map( A => SUM(31), ZN => n23);
   U12 : INV_X1 port map( A => SUM(0), ZN => n38);
   U13 : INV_X1 port map( A => SUM(10), ZN => n37);
   U14 : NOR2_X1 port map( A1 => n40, A2 => n10, ZN => n9);
   U15 : NOR2_X1 port map( A1 => sel(0), A2 => sel(2), ZN => n10);
   U16 : OAI21_X1 port map( B1 => sel(1), B2 => sel(0), A => sel(2), ZN => n12)
                           ;
   U17 : NAND2_X1 port map( A1 => C_BAR, A2 => n18, ZN => n17);
   U18 : NOR2_X1 port map( A1 => sel(1), A2 => sel(2), ZN => n40);
   U19 : NOR4_X1 port map( A1 => SUM(25), A2 => SUM(24), A3 => SUM(26), A4 => 
                           SUM(27), ZN => n22);
   U20 : NOR4_X1 port map( A1 => SUM(29), A2 => SUM(30), A3 => SUM(28), A4 => 
                           SUM(2), ZN => n21);
   U21 : NAND4_X1 port map( A1 => n20, A2 => n39, A3 => n21, A4 => n22, ZN => 
                           n6);
   U22 : XNOR2_X1 port map( A => n6, B => n11, ZN => n7);
   U23 : NAND3_X1 port map( A1 => n8, A2 => n13, A3 => n14, ZN => n4);
   U24 : NAND2_X1 port map( A1 => n7, A2 => n9, ZN => n5);
   U25 : NAND3_X1 port map( A1 => n15, A2 => n40, A3 => n1, ZN => n3);
   U26 : NAND3_X1 port map( A1 => n5, A2 => n3, A3 => n4, ZN => S);
   U27 : NAND2_X1 port map( A1 => V, A2 => n2, ZN => n19);
   U28 : OAI211_X1 port map( C1 => V, C2 => n2, A => n19, B => sign, ZN => n16)
                           ;
   U29 : NAND2_X1 port map( A1 => n16, A2 => n17, ZN => n8);
   U30 : NAND3_X1 port map( A1 => n33, A2 => n34, A3 => n35, ZN => n27);
   U31 : NAND2_X1 port map( A1 => n37, A2 => n38, ZN => n36);
   U32 : NOR2_X1 port map( A1 => SUM(22), A2 => SUM(23), ZN => n29);
   U33 : NAND4_X1 port map( A1 => n30, A2 => n29, A3 => n31, A4 => n32, ZN => 
                           n28);
   U34 : NOR3_X1 port map( A1 => SUM(12), A2 => SUM(11), A3 => n36, ZN => n33);
   U35 : NOR2_X1 port map( A1 => SUM(21), A2 => SUM(20), ZN => n30);
   U36 : NOR2_X1 port map( A1 => SUM(18), A2 => SUM(17), ZN => n31);
   U37 : NOR2_X1 port map( A1 => SUM(19), A2 => SUM(1), ZN => n32);
   U38 : NOR2_X1 port map( A1 => SUM(14), A2 => SUM(13), ZN => n34);
   U39 : NOR2_X1 port map( A1 => SUM(15), A2 => SUM(16), ZN => n35);
   U40 : NOR2_X1 port map( A1 => n28, A2 => n27, ZN => n20);
   U41 : NOR2_X1 port map( A1 => SUM(7), A2 => SUM(8), ZN => n24);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity simple_booth_add_ext_N16 is

   port( Clock, Reset, sign, enable : in std_logic;  valid : out std_logic;  A,
         B : in std_logic_vector (15 downto 0);  A_to_add, B_to_add : out 
         std_logic_vector (31 downto 0);  sign_to_add : out std_logic;  
         final_out : out std_logic_vector (31 downto 0);  ACC_from_add : in 
         std_logic_vector (31 downto 0));

end simple_booth_add_ext_N16;

architecture SYN_struct of simple_booth_add_ext_N16 is

   component NAND3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X4
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_simple_booth_add_ext_N16
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component ff32_en_SIZE32_1
      port( D : in std_logic_vector (31 downto 0);  en, clk, rst : in std_logic
            ;  Q : out std_logic_vector (31 downto 0));
   end component;
   
   component mux21_1
      port( IN0, IN1 : in std_logic_vector (31 downto 0);  CTRL : in std_logic;
            OUT1 : out std_logic_vector (31 downto 0));
   end component;
   
   component piso_r_2_N32
      port( Clock, ALOAD : in std_logic;  D : in std_logic_vector (31 downto 0)
            ;  SO : out std_logic_vector (31 downto 0));
   end component;
   
   component shift_N9_1
      port( Clock, ALOAD : in std_logic;  D : in std_logic_vector (8 downto 0);
            SO : out std_logic);
   end component;
   
   component shift_N9_2
      port( Clock, ALOAD : in std_logic;  D : in std_logic_vector (8 downto 0);
            SO : out std_logic);
   end component;
   
   component shift_N9_0
      port( Clock, ALOAD : in std_logic;  D : in std_logic_vector (8 downto 0);
            SO : out std_logic);
   end component;
   
   component booth_encoder_1
      port( B_in : in std_logic_vector (2 downto 0);  A_out : out 
            std_logic_vector (2 downto 0));
   end component;
   
   component booth_encoder_2
      port( B_in : in std_logic_vector (2 downto 0);  A_out : out 
            std_logic_vector (2 downto 0));
   end component;
   
   component booth_encoder_3
      port( B_in : in std_logic_vector (2 downto 0);  A_out : out 
            std_logic_vector (2 downto 0));
   end component;
   
   component booth_encoder_4
      port( B_in : in std_logic_vector (2 downto 0);  A_out : out 
            std_logic_vector (2 downto 0));
   end component;
   
   component booth_encoder_5
      port( B_in : in std_logic_vector (2 downto 0);  A_out : out 
            std_logic_vector (2 downto 0));
   end component;
   
   component booth_encoder_6
      port( B_in : in std_logic_vector (2 downto 0);  A_out : out 
            std_logic_vector (2 downto 0));
   end component;
   
   component booth_encoder_7
      port( B_in : in std_logic_vector (2 downto 0);  A_out : out 
            std_logic_vector (2 downto 0));
   end component;
   
   component booth_encoder_8
      port( B_in : in std_logic_vector (2 downto 0);  A_out : out 
            std_logic_vector (2 downto 0));
   end component;
   
   component booth_encoder_0
      port( B_in : in std_logic_vector (2 downto 0);  A_out : out 
            std_logic_vector (2 downto 0));
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFS_X1
      port( D, CK, SN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal X_Logic0_port, valid_port, A_to_add_31_port, A_to_add_30_port, 
      A_to_add_29_port, A_to_add_28_port, A_to_add_27_port, A_to_add_26_port, 
      A_to_add_25_port, A_to_add_24_port, A_to_add_23_port, A_to_add_22_port, 
      A_to_add_21_port, A_to_add_20_port, A_to_add_19_port, A_to_add_18_port, 
      A_to_add_17_port, A_to_add_16_port, A_to_add_15_port, A_to_add_14_port, 
      A_to_add_13_port, A_to_add_12_port, A_to_add_11_port, A_to_add_10_port, 
      A_to_add_9_port, A_to_add_8_port, A_to_add_7_port, A_to_add_6_port, 
      A_to_add_5_port, A_to_add_4_port, A_to_add_3_port, A_to_add_2_port, 
      A_to_add_1_port, A_to_add_0_port, enc_N2_in_2_port, piso_0_in_8_port, 
      piso_0_in_7_port, piso_0_in_6_port, piso_0_in_5_port, piso_0_in_4_port, 
      piso_0_in_3_port, piso_0_in_2_port, piso_0_in_1_port, piso_0_in_0_port, 
      piso_1_in_8_port, piso_1_in_7_port, piso_1_in_6_port, piso_1_in_5_port, 
      piso_1_in_4_port, piso_1_in_3_port, piso_1_in_2_port, piso_1_in_1_port, 
      piso_1_in_0_port, piso_2_in_8_port, piso_2_in_7_port, piso_2_in_6_port, 
      piso_2_in_5_port, piso_2_in_4_port, piso_2_in_3_port, piso_2_in_2_port, 
      piso_2_in_1_port, piso_2_in_0_port, extend_vector_15_port, 
      A_to_mux_31_port, A_to_mux_30_port, A_to_mux_29_port, A_to_mux_28_port, 
      A_to_mux_27_port, A_to_mux_26_port, A_to_mux_25_port, A_to_mux_24_port, 
      A_to_mux_23_port, A_to_mux_22_port, A_to_mux_21_port, A_to_mux_20_port, 
      A_to_mux_19_port, A_to_mux_18_port, A_to_mux_17_port, A_to_mux_16_port, 
      A_to_mux_15_port, A_to_mux_14_port, A_to_mux_13_port, A_to_mux_12_port, 
      A_to_mux_11_port, A_to_mux_10_port, A_to_mux_9_port, A_to_mux_8_port, 
      A_to_mux_7_port, A_to_mux_6_port, A_to_mux_5_port, A_to_mux_4_port, 
      A_to_mux_3_port, A_to_mux_2_port, A_to_mux_1_port, A_to_mux_0_port, 
      input_mux_sel_2_port, input_mux_sel_0, next_accumulate_31_port, 
      next_accumulate_30_port, next_accumulate_29_port, next_accumulate_28_port
      , next_accumulate_27_port, next_accumulate_26_port, 
      next_accumulate_25_port, next_accumulate_24_port, next_accumulate_23_port
      , next_accumulate_22_port, next_accumulate_21_port, 
      next_accumulate_20_port, next_accumulate_19_port, next_accumulate_18_port
      , next_accumulate_17_port, next_accumulate_16_port, 
      next_accumulate_15_port, next_accumulate_14_port, next_accumulate_13_port
      , next_accumulate_12_port, next_accumulate_11_port, 
      next_accumulate_10_port, next_accumulate_9_port, next_accumulate_8_port, 
      next_accumulate_7_port, next_accumulate_6_port, next_accumulate_5_port, 
      next_accumulate_4_port, next_accumulate_3_port, next_accumulate_2_port, 
      next_accumulate_1_port, next_accumulate_0_port, reg_enable, count_4_port,
      count_3_port, count_2_port, count_1_port, count_0_port, N23, N37, N39, 
      N41, N43, N44, N45, net3331, n2, n3, n5, n8, n9, n10, n11, n1, n4, n6, n7
      , n12, n13, n14, n16, n17, n18, n19 : std_logic;

begin
   valid <= valid_port;
   A_to_add <= ( A_to_add_31_port, A_to_add_30_port, A_to_add_29_port, 
      A_to_add_28_port, A_to_add_27_port, A_to_add_26_port, A_to_add_25_port, 
      A_to_add_24_port, A_to_add_23_port, A_to_add_22_port, A_to_add_21_port, 
      A_to_add_20_port, A_to_add_19_port, A_to_add_18_port, A_to_add_17_port, 
      A_to_add_16_port, A_to_add_15_port, A_to_add_14_port, A_to_add_13_port, 
      A_to_add_12_port, A_to_add_11_port, A_to_add_10_port, A_to_add_9_port, 
      A_to_add_8_port, A_to_add_7_port, A_to_add_6_port, A_to_add_5_port, 
      A_to_add_4_port, A_to_add_3_port, A_to_add_2_port, A_to_add_1_port, 
      A_to_add_0_port );
   
   X_Logic0_port <= '0';
   count_reg_0_inst : DFFS_X1 port map( D => N37, CK => net3331, SN => n19, Q 
                           => count_0_port, QN => n13);
   count_reg_1_inst : DFFR_X1 port map( D => N39, CK => net3331, RN => n19, Q 
                           => count_1_port, QN => n5);
   count_reg_2_inst : DFFR_X1 port map( D => N41, CK => net3331, RN => n19, Q 
                           => count_2_port, QN => n14);
   count_reg_3_inst : DFFS_X1 port map( D => N43, CK => net3331, SN => n19, Q 
                           => count_3_port, QN => n3);
   count_reg_4_inst : DFFR_X1 port map( D => N45, CK => net3331, RN => n19, Q 
                           => count_4_port, QN => n2);
   U51 : MUX2_X1 port map( A => A_to_add_9_port, B => ACC_from_add(9), S => 
                           input_mux_sel_2_port, Z => final_out(9));
   U52 : MUX2_X1 port map( A => A_to_add_8_port, B => ACC_from_add(8), S => 
                           input_mux_sel_2_port, Z => final_out(8));
   U53 : MUX2_X1 port map( A => A_to_add_7_port, B => ACC_from_add(7), S => 
                           input_mux_sel_2_port, Z => final_out(7));
   U54 : MUX2_X1 port map( A => A_to_add_6_port, B => ACC_from_add(6), S => 
                           input_mux_sel_2_port, Z => final_out(6));
   U55 : MUX2_X1 port map( A => A_to_add_5_port, B => ACC_from_add(5), S => 
                           input_mux_sel_2_port, Z => final_out(5));
   U56 : MUX2_X1 port map( A => A_to_add_4_port, B => ACC_from_add(4), S => 
                           input_mux_sel_2_port, Z => final_out(4));
   U57 : MUX2_X1 port map( A => A_to_add_3_port, B => ACC_from_add(3), S => 
                           input_mux_sel_2_port, Z => final_out(3));
   U58 : MUX2_X1 port map( A => A_to_add_31_port, B => ACC_from_add(31), S => 
                           input_mux_sel_2_port, Z => final_out(31));
   U59 : MUX2_X1 port map( A => A_to_add_30_port, B => ACC_from_add(30), S => 
                           input_mux_sel_2_port, Z => final_out(30));
   U61 : MUX2_X1 port map( A => A_to_add_29_port, B => ACC_from_add(29), S => 
                           input_mux_sel_2_port, Z => final_out(29));
   U62 : MUX2_X1 port map( A => A_to_add_28_port, B => ACC_from_add(28), S => 
                           input_mux_sel_2_port, Z => final_out(28));
   U63 : MUX2_X1 port map( A => A_to_add_27_port, B => ACC_from_add(27), S => 
                           input_mux_sel_2_port, Z => final_out(27));
   U64 : MUX2_X1 port map( A => A_to_add_26_port, B => ACC_from_add(26), S => 
                           input_mux_sel_2_port, Z => final_out(26));
   U65 : MUX2_X1 port map( A => A_to_add_25_port, B => ACC_from_add(25), S => 
                           input_mux_sel_2_port, Z => final_out(25));
   U66 : MUX2_X1 port map( A => A_to_add_24_port, B => ACC_from_add(24), S => 
                           input_mux_sel_2_port, Z => final_out(24));
   U67 : MUX2_X1 port map( A => A_to_add_23_port, B => ACC_from_add(23), S => 
                           input_mux_sel_2_port, Z => final_out(23));
   U68 : MUX2_X1 port map( A => A_to_add_22_port, B => ACC_from_add(22), S => 
                           input_mux_sel_2_port, Z => final_out(22));
   U69 : MUX2_X1 port map( A => A_to_add_21_port, B => ACC_from_add(21), S => 
                           input_mux_sel_2_port, Z => final_out(21));
   U70 : MUX2_X1 port map( A => A_to_add_20_port, B => ACC_from_add(20), S => 
                           input_mux_sel_2_port, Z => final_out(20));
   U71 : MUX2_X1 port map( A => A_to_add_1_port, B => ACC_from_add(1), S => 
                           input_mux_sel_2_port, Z => final_out(1));
   U72 : MUX2_X1 port map( A => A_to_add_19_port, B => ACC_from_add(19), S => 
                           input_mux_sel_2_port, Z => final_out(19));
   U73 : MUX2_X1 port map( A => A_to_add_18_port, B => ACC_from_add(18), S => 
                           input_mux_sel_2_port, Z => final_out(18));
   U74 : MUX2_X1 port map( A => A_to_add_17_port, B => ACC_from_add(17), S => 
                           input_mux_sel_2_port, Z => final_out(17));
   U75 : MUX2_X1 port map( A => A_to_add_16_port, B => ACC_from_add(16), S => 
                           input_mux_sel_2_port, Z => final_out(16));
   U76 : MUX2_X1 port map( A => A_to_add_15_port, B => ACC_from_add(15), S => 
                           input_mux_sel_2_port, Z => final_out(15));
   U77 : MUX2_X1 port map( A => A_to_add_14_port, B => ACC_from_add(14), S => 
                           input_mux_sel_2_port, Z => final_out(14));
   U78 : MUX2_X1 port map( A => A_to_add_13_port, B => ACC_from_add(13), S => 
                           input_mux_sel_2_port, Z => final_out(13));
   U79 : MUX2_X1 port map( A => A_to_add_12_port, B => ACC_from_add(12), S => 
                           input_mux_sel_2_port, Z => final_out(12));
   U80 : MUX2_X1 port map( A => A_to_add_11_port, B => ACC_from_add(11), S => 
                           input_mux_sel_2_port, Z => final_out(11));
   U81 : MUX2_X1 port map( A => A_to_add_10_port, B => ACC_from_add(10), S => 
                           input_mux_sel_2_port, Z => final_out(10));
   encod_0_0 : booth_encoder_0 port map( B_in(2) => B(1), B_in(1) => B(0), 
                           B_in(0) => X_Logic0_port, A_out(2) => 
                           piso_2_in_0_port, A_out(1) => piso_1_in_0_port, 
                           A_out(0) => piso_0_in_0_port);
   encod_i_1 : booth_encoder_8 port map( B_in(2) => B(3), B_in(1) => B(2), 
                           B_in(0) => B(1), A_out(2) => piso_2_in_1_port, 
                           A_out(1) => piso_1_in_1_port, A_out(0) => 
                           piso_0_in_1_port);
   encod_i_2 : booth_encoder_7 port map( B_in(2) => B(5), B_in(1) => B(4), 
                           B_in(0) => B(3), A_out(2) => piso_2_in_2_port, 
                           A_out(1) => piso_1_in_2_port, A_out(0) => 
                           piso_0_in_2_port);
   encod_i_3 : booth_encoder_6 port map( B_in(2) => B(7), B_in(1) => B(6), 
                           B_in(0) => B(5), A_out(2) => piso_2_in_3_port, 
                           A_out(1) => piso_1_in_3_port, A_out(0) => 
                           piso_0_in_3_port);
   encod_i_4 : booth_encoder_5 port map( B_in(2) => B(9), B_in(1) => B(8), 
                           B_in(0) => B(7), A_out(2) => piso_2_in_4_port, 
                           A_out(1) => piso_1_in_4_port, A_out(0) => 
                           piso_0_in_4_port);
   encod_i_5 : booth_encoder_4 port map( B_in(2) => B(11), B_in(1) => B(10), 
                           B_in(0) => B(9), A_out(2) => piso_2_in_5_port, 
                           A_out(1) => piso_1_in_5_port, A_out(0) => 
                           piso_0_in_5_port);
   encod_i_6 : booth_encoder_3 port map( B_in(2) => B(13), B_in(1) => B(12), 
                           B_in(0) => B(11), A_out(2) => piso_2_in_6_port, 
                           A_out(1) => piso_1_in_6_port, A_out(0) => 
                           piso_0_in_6_port);
   encod_i_7 : booth_encoder_2 port map( B_in(2) => B(15), B_in(1) => B(14), 
                           B_in(0) => B(13), A_out(2) => piso_2_in_7_port, 
                           A_out(1) => piso_1_in_7_port, A_out(0) => 
                           piso_0_in_7_port);
   encod_i_8 : booth_encoder_1 port map( B_in(2) => enc_N2_in_2_port, B_in(1) 
                           => enc_N2_in_2_port, B_in(0) => B(15), A_out(2) => 
                           piso_2_in_8_port, A_out(1) => piso_1_in_8_port, 
                           A_out(0) => piso_0_in_8_port);
   piso_0 : shift_N9_0 port map( Clock => Clock, ALOAD => n18, D(8) => 
                           piso_0_in_8_port, D(7) => piso_0_in_7_port, D(6) => 
                           piso_0_in_6_port, D(5) => piso_0_in_5_port, D(4) => 
                           piso_0_in_4_port, D(3) => piso_0_in_3_port, D(2) => 
                           piso_0_in_2_port, D(1) => piso_0_in_1_port, D(0) => 
                           piso_0_in_0_port, SO => input_mux_sel_0);
   piso_1 : shift_N9_2 port map( Clock => Clock, ALOAD => n18, D(8) => 
                           piso_1_in_8_port, D(7) => piso_1_in_7_port, D(6) => 
                           piso_1_in_6_port, D(5) => piso_1_in_5_port, D(4) => 
                           piso_1_in_4_port, D(3) => piso_1_in_3_port, D(2) => 
                           piso_1_in_2_port, D(1) => piso_1_in_1_port, D(0) => 
                           piso_1_in_0_port, SO => sign_to_add);
   piso_2 : shift_N9_1 port map( Clock => Clock, ALOAD => n18, D(8) => 
                           piso_2_in_8_port, D(7) => piso_2_in_7_port, D(6) => 
                           piso_2_in_6_port, D(5) => piso_2_in_5_port, D(4) => 
                           piso_2_in_4_port, D(3) => piso_2_in_3_port, D(2) => 
                           piso_2_in_2_port, D(1) => piso_2_in_1_port, D(0) => 
                           piso_2_in_0_port, SO => input_mux_sel_2_port);
   A_reg : piso_r_2_N32 port map( Clock => Clock, ALOAD => n18, D(31) => 
                           extend_vector_15_port, D(30) => 
                           extend_vector_15_port, D(29) => 
                           extend_vector_15_port, D(28) => 
                           extend_vector_15_port, D(27) => 
                           extend_vector_15_port, D(26) => 
                           extend_vector_15_port, D(25) => 
                           extend_vector_15_port, D(24) => 
                           extend_vector_15_port, D(23) => 
                           extend_vector_15_port, D(22) => 
                           extend_vector_15_port, D(21) => 
                           extend_vector_15_port, D(20) => 
                           extend_vector_15_port, D(19) => 
                           extend_vector_15_port, D(18) => 
                           extend_vector_15_port, D(17) => 
                           extend_vector_15_port, D(16) => 
                           extend_vector_15_port, D(15) => A(15), D(14) => 
                           A(14), D(13) => A(13), D(12) => A(12), D(11) => 
                           A(11), D(10) => A(10), D(9) => A(9), D(8) => A(8), 
                           D(7) => A(7), D(6) => A(6), D(5) => A(5), D(4) => 
                           A(4), D(3) => A(3), D(2) => A(2), D(1) => A(1), D(0)
                           => A(0), SO(31) => A_to_mux_31_port, SO(30) => 
                           A_to_mux_30_port, SO(29) => A_to_mux_29_port, SO(28)
                           => A_to_mux_28_port, SO(27) => A_to_mux_27_port, 
                           SO(26) => A_to_mux_26_port, SO(25) => 
                           A_to_mux_25_port, SO(24) => A_to_mux_24_port, SO(23)
                           => A_to_mux_23_port, SO(22) => A_to_mux_22_port, 
                           SO(21) => A_to_mux_21_port, SO(20) => 
                           A_to_mux_20_port, SO(19) => A_to_mux_19_port, SO(18)
                           => A_to_mux_18_port, SO(17) => A_to_mux_17_port, 
                           SO(16) => A_to_mux_16_port, SO(15) => 
                           A_to_mux_15_port, SO(14) => A_to_mux_14_port, SO(13)
                           => A_to_mux_13_port, SO(12) => A_to_mux_12_port, 
                           SO(11) => A_to_mux_11_port, SO(10) => 
                           A_to_mux_10_port, SO(9) => A_to_mux_9_port, SO(8) =>
                           A_to_mux_8_port, SO(7) => A_to_mux_7_port, SO(6) => 
                           A_to_mux_6_port, SO(5) => A_to_mux_5_port, SO(4) => 
                           A_to_mux_4_port, SO(3) => A_to_mux_3_port, SO(2) => 
                           A_to_mux_2_port, SO(1) => A_to_mux_1_port, SO(0) => 
                           A_to_mux_0_port);
   INPUTMUX : mux21_1 port map( IN0(31) => A_to_mux_31_port, IN0(30) => 
                           A_to_mux_30_port, IN0(29) => A_to_mux_29_port, 
                           IN0(28) => A_to_mux_28_port, IN0(27) => 
                           A_to_mux_27_port, IN0(26) => A_to_mux_26_port, 
                           IN0(25) => A_to_mux_25_port, IN0(24) => 
                           A_to_mux_24_port, IN0(23) => A_to_mux_23_port, 
                           IN0(22) => A_to_mux_22_port, IN0(21) => 
                           A_to_mux_21_port, IN0(20) => A_to_mux_20_port, 
                           IN0(19) => A_to_mux_19_port, IN0(18) => 
                           A_to_mux_18_port, IN0(17) => A_to_mux_17_port, 
                           IN0(16) => A_to_mux_16_port, IN0(15) => 
                           A_to_mux_15_port, IN0(14) => A_to_mux_14_port, 
                           IN0(13) => A_to_mux_13_port, IN0(12) => 
                           A_to_mux_12_port, IN0(11) => A_to_mux_11_port, 
                           IN0(10) => A_to_mux_10_port, IN0(9) => 
                           A_to_mux_9_port, IN0(8) => A_to_mux_8_port, IN0(7) 
                           => A_to_mux_7_port, IN0(6) => A_to_mux_6_port, 
                           IN0(5) => A_to_mux_5_port, IN0(4) => A_to_mux_4_port
                           , IN0(3) => A_to_mux_3_port, IN0(2) => 
                           A_to_mux_2_port, IN0(1) => A_to_mux_1_port, IN0(0) 
                           => A_to_mux_0_port, IN1(31) => A_to_mux_30_port, 
                           IN1(30) => A_to_mux_29_port, IN1(29) => 
                           A_to_mux_28_port, IN1(28) => A_to_mux_27_port, 
                           IN1(27) => A_to_mux_26_port, IN1(26) => 
                           A_to_mux_25_port, IN1(25) => A_to_mux_24_port, 
                           IN1(24) => A_to_mux_23_port, IN1(23) => 
                           A_to_mux_22_port, IN1(22) => A_to_mux_21_port, 
                           IN1(21) => A_to_mux_20_port, IN1(20) => 
                           A_to_mux_19_port, IN1(19) => A_to_mux_18_port, 
                           IN1(18) => A_to_mux_17_port, IN1(17) => 
                           A_to_mux_16_port, IN1(16) => A_to_mux_15_port, 
                           IN1(15) => A_to_mux_14_port, IN1(14) => 
                           A_to_mux_13_port, IN1(13) => A_to_mux_12_port, 
                           IN1(12) => A_to_mux_11_port, IN1(11) => 
                           A_to_mux_10_port, IN1(10) => A_to_mux_9_port, IN1(9)
                           => A_to_mux_8_port, IN1(8) => A_to_mux_7_port, 
                           IN1(7) => A_to_mux_6_port, IN1(6) => A_to_mux_5_port
                           , IN1(5) => A_to_mux_4_port, IN1(4) => 
                           A_to_mux_3_port, IN1(3) => A_to_mux_2_port, IN1(2) 
                           => A_to_mux_1_port, IN1(1) => A_to_mux_0_port, 
                           IN1(0) => X_Logic0_port, CTRL => input_mux_sel_0, 
                           OUT1(31) => B_to_add(31), OUT1(30) => B_to_add(30), 
                           OUT1(29) => B_to_add(29), OUT1(28) => B_to_add(28), 
                           OUT1(27) => B_to_add(27), OUT1(26) => B_to_add(26), 
                           OUT1(25) => B_to_add(25), OUT1(24) => B_to_add(24), 
                           OUT1(23) => B_to_add(23), OUT1(22) => B_to_add(22), 
                           OUT1(21) => B_to_add(21), OUT1(20) => B_to_add(20), 
                           OUT1(19) => B_to_add(19), OUT1(18) => B_to_add(18), 
                           OUT1(17) => B_to_add(17), OUT1(16) => B_to_add(16), 
                           OUT1(15) => B_to_add(15), OUT1(14) => B_to_add(14), 
                           OUT1(13) => B_to_add(13), OUT1(12) => B_to_add(12), 
                           OUT1(11) => B_to_add(11), OUT1(10) => B_to_add(10), 
                           OUT1(9) => B_to_add(9), OUT1(8) => B_to_add(8), 
                           OUT1(7) => B_to_add(7), OUT1(6) => B_to_add(6), 
                           OUT1(5) => B_to_add(5), OUT1(4) => B_to_add(4), 
                           OUT1(3) => B_to_add(3), OUT1(2) => B_to_add(2), 
                           OUT1(1) => B_to_add(1), OUT1(0) => B_to_add(0));
   ACCUMULATOR : ff32_en_SIZE32_1 port map( D(31) => next_accumulate_31_port, 
                           D(30) => next_accumulate_30_port, D(29) => 
                           next_accumulate_29_port, D(28) => 
                           next_accumulate_28_port, D(27) => 
                           next_accumulate_27_port, D(26) => 
                           next_accumulate_26_port, D(25) => 
                           next_accumulate_25_port, D(24) => 
                           next_accumulate_24_port, D(23) => 
                           next_accumulate_23_port, D(22) => 
                           next_accumulate_22_port, D(21) => 
                           next_accumulate_21_port, D(20) => 
                           next_accumulate_20_port, D(19) => 
                           next_accumulate_19_port, D(18) => 
                           next_accumulate_18_port, D(17) => 
                           next_accumulate_17_port, D(16) => 
                           next_accumulate_16_port, D(15) => 
                           next_accumulate_15_port, D(14) => 
                           next_accumulate_14_port, D(13) => 
                           next_accumulate_13_port, D(12) => 
                           next_accumulate_12_port, D(11) => 
                           next_accumulate_11_port, D(10) => 
                           next_accumulate_10_port, D(9) => 
                           next_accumulate_9_port, D(8) => 
                           next_accumulate_8_port, D(7) => 
                           next_accumulate_7_port, D(6) => 
                           next_accumulate_6_port, D(5) => 
                           next_accumulate_5_port, D(4) => 
                           next_accumulate_4_port, D(3) => 
                           next_accumulate_3_port, D(2) => 
                           next_accumulate_2_port, D(1) => 
                           next_accumulate_1_port, D(0) => 
                           next_accumulate_0_port, en => reg_enable, clk => 
                           Clock, rst => Reset, Q(31) => A_to_add_31_port, 
                           Q(30) => A_to_add_30_port, Q(29) => A_to_add_29_port
                           , Q(28) => A_to_add_28_port, Q(27) => 
                           A_to_add_27_port, Q(26) => A_to_add_26_port, Q(25) 
                           => A_to_add_25_port, Q(24) => A_to_add_24_port, 
                           Q(23) => A_to_add_23_port, Q(22) => A_to_add_22_port
                           , Q(21) => A_to_add_21_port, Q(20) => 
                           A_to_add_20_port, Q(19) => A_to_add_19_port, Q(18) 
                           => A_to_add_18_port, Q(17) => A_to_add_17_port, 
                           Q(16) => A_to_add_16_port, Q(15) => A_to_add_15_port
                           , Q(14) => A_to_add_14_port, Q(13) => 
                           A_to_add_13_port, Q(12) => A_to_add_12_port, Q(11) 
                           => A_to_add_11_port, Q(10) => A_to_add_10_port, Q(9)
                           => A_to_add_9_port, Q(8) => A_to_add_8_port, Q(7) =>
                           A_to_add_7_port, Q(6) => A_to_add_6_port, Q(5) => 
                           A_to_add_5_port, Q(4) => A_to_add_4_port, Q(3) => 
                           A_to_add_3_port, Q(2) => A_to_add_2_port, Q(1) => 
                           A_to_add_1_port, Q(0) => A_to_add_0_port);
   clk_gate_count_reg : SNPS_CLOCK_GATE_HIGH_simple_booth_add_ext_N16 port map(
                           CLK => Clock, EN => N44, ENCLK => net3331);
   U41 : OR2_X1 port map( A1 => valid_port, A2 => enable, ZN => N44);
   U48 : INV_X1 port map( A => n9, ZN => n11);
   U4 : OR2_X1 port map( A1 => n18, A2 => input_mux_sel_2_port, ZN => 
                           reg_enable);
   U17 : AND2_X1 port map( A1 => n8, A2 => ACC_from_add(27), ZN => 
                           next_accumulate_27_port);
   U7 : AND2_X1 port map( A1 => n8, A2 => ACC_from_add(7), ZN => 
                           next_accumulate_7_port);
   U13 : AND2_X1 port map( A1 => n8, A2 => ACC_from_add(30), ZN => 
                           next_accumulate_30_port);
   U15 : AND2_X1 port map( A1 => n8, A2 => ACC_from_add(29), ZN => 
                           next_accumulate_29_port);
   U18 : AND2_X1 port map( A1 => n8, A2 => ACC_from_add(26), ZN => 
                           next_accumulate_26_port);
   U19 : AND2_X1 port map( A1 => n8, A2 => ACC_from_add(25), ZN => 
                           next_accumulate_25_port);
   U30 : AND2_X1 port map( A1 => n8, A2 => ACC_from_add(15), ZN => 
                           next_accumulate_15_port);
   U31 : AND2_X1 port map( A1 => n8, A2 => ACC_from_add(14), ZN => 
                           next_accumulate_14_port);
   U11 : AND2_X1 port map( A1 => n8, A2 => ACC_from_add(3), ZN => 
                           next_accumulate_3_port);
   U21 : AND2_X1 port map( A1 => n8, A2 => ACC_from_add(23), ZN => 
                           next_accumulate_23_port);
   U33 : AND2_X1 port map( A1 => n8, A2 => ACC_from_add(12), ZN => 
                           next_accumulate_12_port);
   U26 : AND2_X1 port map( A1 => n8, A2 => ACC_from_add(19), ZN => 
                           next_accumulate_19_port);
   U27 : AND2_X1 port map( A1 => n8, A2 => ACC_from_add(18), ZN => 
                           next_accumulate_18_port);
   U28 : AND2_X1 port map( A1 => n8, A2 => ACC_from_add(17), ZN => 
                           next_accumulate_17_port);
   U29 : AND2_X1 port map( A1 => n8, A2 => ACC_from_add(16), ZN => 
                           next_accumulate_16_port);
   U34 : AND2_X1 port map( A1 => n8, A2 => ACC_from_add(11), ZN => 
                           next_accumulate_11_port);
   U8 : AND2_X1 port map( A1 => n8, A2 => ACC_from_add(6), ZN => 
                           next_accumulate_6_port);
   U5 : AND2_X1 port map( A1 => n8, A2 => ACC_from_add(9), ZN => 
                           next_accumulate_9_port);
   U6 : AND2_X1 port map( A1 => n8, A2 => ACC_from_add(8), ZN => 
                           next_accumulate_8_port);
   U35 : AND2_X1 port map( A1 => n8, A2 => ACC_from_add(10), ZN => 
                           next_accumulate_10_port);
   U14 : AND2_X1 port map( A1 => n8, A2 => ACC_from_add(2), ZN => 
                           next_accumulate_2_port);
   U9 : AND2_X1 port map( A1 => n8, A2 => ACC_from_add(5), ZN => 
                           next_accumulate_5_port);
   U25 : AND2_X1 port map( A1 => n8, A2 => ACC_from_add(1), ZN => 
                           next_accumulate_1_port);
   U10 : AND2_X1 port map( A1 => n8, A2 => ACC_from_add(4), ZN => 
                           next_accumulate_4_port);
   U36 : AND2_X1 port map( A1 => n8, A2 => ACC_from_add(0), ZN => 
                           next_accumulate_0_port);
   U38 : AND2_X1 port map( A1 => sign, A2 => A(15), ZN => extend_vector_15_port
                           );
   U45 : INV_X1 port map( A => valid_port, ZN => n10);
   U43 : AND2_X1 port map( A1 => N23, A2 => n10, ZN => N41);
   U46 : OR2_X1 port map( A1 => valid_port, A2 => n13, ZN => N37);
   U49 : NOR3_X1 port map( A1 => count_1_port, A2 => count_4_port, A3 => 
                           count_2_port, ZN => n9);
   U47 : NOR3_X1 port map( A1 => count_3_port, A2 => count_0_port, A3 => n11, 
                           ZN => valid_port);
   U3 : NOR2_X1 port map( A1 => count_3_port, A2 => n17, ZN => n1);
   U12 : OAI21_X1 port map( B1 => count_4_port, B2 => n1, A => n10, ZN => n4);
   U16 : AOI21_X1 port map( B1 => count_4_port, B2 => n1, A => n4, ZN => N45);
   U20 : MUX2_X1 port map( A => A_to_add_0_port, B => ACC_from_add(0), S => 
                           input_mux_sel_2_port, Z => final_out(0));
   U22 : AOI21_X1 port map( B1 => n17, B2 => count_3_port, A => valid_port, ZN 
                           => n6);
   U23 : OAI21_X1 port map( B1 => n17, B2 => count_3_port, A => n6, ZN => N43);
   U24 : MUX2_X1 port map( A => A_to_add_2_port, B => ACC_from_add(2), S => 
                           input_mux_sel_2_port, Z => final_out(2));
   U32 : INV_X1 port map( A => n10, ZN => n7);
   U37 : AOI21_X1 port map( B1 => count_1_port, B2 => count_0_port, A => n16, 
                           ZN => n12);
   U39 : NOR2_X1 port map( A1 => n12, A2 => n7, ZN => N39);
   U40 : INV_X4 port map( A => n8, ZN => n18);
   U42 : NOR2_X1 port map( A1 => count_0_port, A2 => count_1_port, ZN => n16);
   U44 : OR3_X1 port map( A1 => count_2_port, A2 => count_0_port, A3 => 
                           count_1_port, ZN => n17);
   U50 : OAI21_X1 port map( B1 => n16, B2 => n14, A => n17, ZN => N23);
   U60 : INV_X1 port map( A => Reset, ZN => n19);
   U82 : AND2_X1 port map( A1 => sign, A2 => B(15), ZN => enc_N2_in_2_port);
   U83 : AND2_X1 port map( A1 => n8, A2 => ACC_from_add(13), ZN => 
                           next_accumulate_13_port);
   U84 : AND2_X1 port map( A1 => n8, A2 => ACC_from_add(21), ZN => 
                           next_accumulate_21_port);
   U85 : AND2_X1 port map( A1 => n8, A2 => ACC_from_add(20), ZN => 
                           next_accumulate_20_port);
   U86 : AND2_X1 port map( A1 => n8, A2 => ACC_from_add(22), ZN => 
                           next_accumulate_22_port);
   U87 : AND2_X1 port map( A1 => n8, A2 => ACC_from_add(24), ZN => 
                           next_accumulate_24_port);
   U88 : AND2_X1 port map( A1 => n8, A2 => ACC_from_add(28), ZN => 
                           next_accumulate_28_port);
   U89 : AND2_X1 port map( A1 => n8, A2 => ACC_from_add(31), ZN => 
                           next_accumulate_31_port);
   U90 : NAND3_X2 port map( A1 => n9, A2 => count_3_port, A3 => count_0_port, 
                           ZN => n8);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_ff32_en_SIZE13 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_ff32_en_SIZE13;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_ff32_en_SIZE13 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net3370 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net3370);
   main_gate : AND2_X1 port map( A1 => net3370, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_ff32_en_SIZE5_0 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_ff32_en_SIZE5_0;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_ff32_en_SIZE5_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net3355 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net3355);
   main_gate : AND2_X1 port map( A1 => net3355, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_ff32_en_SIZE32_0 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_ff32_en_SIZE32_0;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_ff32_en_SIZE32_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net3340 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net3340);
   main_gate : AND2_X1 port map( A1 => net3340, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity sum_gen_N32_0 is

   port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic_vector 
         (8 downto 0);  S : out std_logic_vector (31 downto 0));

end sum_gen_N32_0;

architecture SYN_STRUCTURAL of sum_gen_N32_0 is

   component carry_sel_gen_N4_9
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component carry_sel_gen_N4_10
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component carry_sel_gen_N4_11
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component carry_sel_gen_N4_12
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component carry_sel_gen_N4_13
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component carry_sel_gen_N4_14
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component carry_sel_gen_N4_15
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component carry_sel_gen_N4_0
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal n1, net3145, net3146, net3147, net3148, net3149, net3150, net3151, 
      net3152 : std_logic;

begin
   
   csel_N_0 : carry_sel_gen_N4_0 port map( A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), Ci => n1, S(3) => S(3), S(2) 
                           => S(2), S(1) => S(1), S(0) => S(0), Co => net3152);
   csel_N_1 : carry_sel_gen_N4_15 port map( A(3) => A(7), A(2) => A(6), A(1) =>
                           A(5), A(0) => A(4), B(3) => B(7), B(2) => B(6), B(1)
                           => B(5), B(0) => B(4), Ci => Cin(1), S(3) => S(7), 
                           S(2) => S(6), S(1) => S(5), S(0) => S(4), Co => 
                           net3151);
   csel_N_2 : carry_sel_gen_N4_14 port map( A(3) => A(11), A(2) => A(10), A(1) 
                           => A(9), A(0) => A(8), B(3) => B(11), B(2) => B(10),
                           B(1) => B(9), B(0) => B(8), Ci => Cin(2), S(3) => 
                           S(11), S(2) => S(10), S(1) => S(9), S(0) => S(8), Co
                           => net3150);
   csel_N_3 : carry_sel_gen_N4_13 port map( A(3) => A(15), A(2) => A(14), A(1) 
                           => A(13), A(0) => A(12), B(3) => B(15), B(2) => 
                           B(14), B(1) => B(13), B(0) => B(12), Ci => Cin(3), 
                           S(3) => S(15), S(2) => S(14), S(1) => S(13), S(0) =>
                           S(12), Co => net3149);
   csel_N_4 : carry_sel_gen_N4_12 port map( A(3) => A(19), A(2) => A(18), A(1) 
                           => A(17), A(0) => A(16), B(3) => B(19), B(2) => 
                           B(18), B(1) => B(17), B(0) => B(16), Ci => Cin(4), 
                           S(3) => S(19), S(2) => S(18), S(1) => S(17), S(0) =>
                           S(16), Co => net3148);
   csel_N_5 : carry_sel_gen_N4_11 port map( A(3) => A(23), A(2) => A(22), A(1) 
                           => A(21), A(0) => A(20), B(3) => B(23), B(2) => 
                           B(22), B(1) => B(21), B(0) => B(20), Ci => Cin(5), 
                           S(3) => S(23), S(2) => S(22), S(1) => S(21), S(0) =>
                           S(20), Co => net3147);
   csel_N_6 : carry_sel_gen_N4_10 port map( A(3) => A(27), A(2) => A(26), A(1) 
                           => A(25), A(0) => A(24), B(3) => B(27), B(2) => 
                           B(26), B(1) => B(25), B(0) => B(24), Ci => Cin(6), 
                           S(3) => S(27), S(2) => S(26), S(1) => S(25), S(0) =>
                           S(24), Co => net3146);
   csel_N_7 : carry_sel_gen_N4_9 port map( A(3) => A(31), A(2) => A(30), A(1) 
                           => A(29), A(0) => A(28), B(3) => B(31), B(2) => 
                           B(30), B(1) => B(29), B(0) => B(28), Ci => Cin(7), 
                           S(3) => S(31), S(2) => S(30), S(1) => S(29), S(0) =>
                           S(28), Co => net3145);
   n1 <= '0';

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity carry_tree_N32_logN5_0 is

   port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  Cout :
         out std_logic_vector (7 downto 0));

end carry_tree_N32_logN5_0;

architecture SYN_arch of carry_tree_N32_logN5_0 is

   component pg_29
      port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic
            );
   end component;
   
   component pg_31
      port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic
            );
   end component;
   
   component pg_32
      port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic
            );
   end component;
   
   component g_12
      port( g, p, g_prec : in std_logic;  g_out : out std_logic);
   end component;
   
   component g_13
      port( g, p, g_prec : in std_logic;  g_out : out std_logic);
   end component;
   
   component g_14
      port( g, p, g_prec : in std_logic;  g_out : out std_logic);
   end component;
   
   component g_15
      port( g, p, g_prec : in std_logic;  g_out : out std_logic);
   end component;
   
   component g_16
      port( g, p, g_prec : in std_logic;  g_out : out std_logic);
   end component;
   
   component g_17
      port( g, p, g_prec : in std_logic;  g_out : out std_logic);
   end component;
   
   component pg_34
      port( p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic;  
            g_BAR : in std_logic);
   end component;
   
   component pg_35
      port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic
            );
   end component;
   
   component pg_36
      port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic
            );
   end component;
   
   component pg_37
      port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic
            );
   end component;
   
   component pg_38
      port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic
            );
   end component;
   
   component pg_39
      port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic
            );
   end component;
   
   component g_18
      port( g, p, g_prec : in std_logic;  g_out : out std_logic);
   end component;
   
   component pg_42
      port( g, p, g_prec, p_prec : in std_logic;  p_out, g_out_BAR : out 
            std_logic);
   end component;
   
   component pg_43
      port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic
            );
   end component;
   
   component pg_44
      port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic
            );
   end component;
   
   component pg_45
      port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic
            );
   end component;
   
   component pg_46
      port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic
            );
   end component;
   
   component pg_47
      port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic
            );
   end component;
   
   component pg_48
      port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic
            );
   end component;
   
   component pg_49
      port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic
            );
   end component;
   
   component pg_50
      port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic
            );
   end component;
   
   component pg_51
      port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic
            );
   end component;
   
   component pg_52
      port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic
            );
   end component;
   
   component pg_53
      port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic
            );
   end component;
   
   component pg_0
      port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic
            );
   end component;
   
   component g_19
      port( g, p, g_prec : in std_logic;  g_out : out std_logic);
   end component;
   
   component g_0
      port( g, p, g_prec : in std_logic;  g_out : out std_logic);
   end component;
   
   component pg_net_33
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_38
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_39
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_40
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_41
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_42
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_43
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_44
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_45
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_46
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_47
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_48
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_49
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_50
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_51
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_52
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_53
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_54
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_55
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_56
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_57
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_58
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_59
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_60
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_61
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_62
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_63
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_0
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   signal n2, Cout_6_port, Cout_5_port, Cout_4_port, Cout_3_port, Cout_2_port, 
      Cout_1_port, Cout_0_port, p_net_27_port, p_net_26_port, p_net_25_port, 
      p_net_24_port, p_net_23_port, p_net_22_port, p_net_21_port, p_net_20_port
      , p_net_19_port, p_net_18_port, p_net_17_port, p_net_16_port, 
      p_net_15_port, p_net_14_port, p_net_13_port, p_net_12_port, p_net_11_port
      , p_net_10_port, p_net_9_port, p_net_8_port, p_net_7_port, p_net_6_port, 
      p_net_5_port, p_net_4_port, p_net_3_port, p_net_2_port, p_net_1_port, 
      g_net_27_port, g_net_26_port, g_net_25_port, g_net_24_port, g_net_23_port
      , g_net_22_port, g_net_21_port, g_net_20_port, g_net_19_port, 
      g_net_18_port, g_net_17_port, g_net_16_port, g_net_15_port, g_net_14_port
      , g_net_13_port, g_net_12_port, g_net_11_port, g_net_10_port, 
      g_net_9_port, g_net_8_port, g_net_7_port, g_net_6_port, g_net_5_port, 
      g_net_4_port, g_net_3_port, g_net_2_port, g_net_1_port, g_net_0_port, 
      magic_pro_0_port, pg_1_13_1_port, pg_1_13_0_port, pg_1_12_1_port, 
      pg_1_12_0_port, pg_1_11_1_port, pg_1_11_0_port, pg_1_10_1_port, 
      pg_1_10_0_port, pg_1_9_1_port, pg_1_9_0_port, pg_1_8_1_port, 
      pg_1_8_0_port, pg_1_7_1_port, pg_1_7_0_port, pg_1_6_1_port, pg_1_6_0_port
      , pg_1_5_1_port, pg_1_5_0_port, pg_1_4_1_port, pg_1_4_0_port, 
      pg_1_3_1_port, pg_1_3_0_port, pg_1_2_1_port, pg_1_2_0_port, pg_1_1_1_port
      , pg_1_1_0_port, pg_1_0_0_port, pg_n_4_6_1_port, pg_n_4_6_0_port, 
      pg_n_3_5_1_port, pg_n_3_5_0_port, pg_n_3_3_1_port, pg_n_3_3_0_port, 
      pg_n_2_6_1_port, pg_n_2_6_0_port, pg_n_2_5_1_port, pg_n_2_5_0_port, 
      pg_n_2_4_1_port, pg_n_2_4_0_port, pg_n_2_3_1_port, pg_n_2_3_0_port, 
      pg_n_2_2_1_port, pg_n_2_2_0_port, pg_n_2_1_1_port, pg_n_2_1_0_port, n1, 
      net48715, n_1170 : std_logic;

begin
   Cout <= ( n_1170, Cout_6_port, Cout_5_port, Cout_4_port, Cout_3_port, 
      Cout_2_port, Cout_1_port, Cout_0_port );
   
   pg_net_x_1 : pg_net_0 port map( a => A(1), b => B(1), g_out => g_net_1_port,
                           p_out => p_net_1_port);
   pg_net_x_2 : pg_net_63 port map( a => A(2), b => B(2), g_out => g_net_2_port
                           , p_out => p_net_2_port);
   pg_net_x_3 : pg_net_62 port map( a => A(3), b => B(3), g_out => g_net_3_port
                           , p_out => p_net_3_port);
   pg_net_x_4 : pg_net_61 port map( a => A(4), b => B(4), g_out => g_net_4_port
                           , p_out => p_net_4_port);
   pg_net_x_5 : pg_net_60 port map( a => A(5), b => B(5), g_out => g_net_5_port
                           , p_out => p_net_5_port);
   pg_net_x_6 : pg_net_59 port map( a => A(6), b => B(6), g_out => g_net_6_port
                           , p_out => p_net_6_port);
   pg_net_x_7 : pg_net_58 port map( a => A(7), b => B(7), g_out => g_net_7_port
                           , p_out => p_net_7_port);
   pg_net_x_8 : pg_net_57 port map( a => A(8), b => B(8), g_out => g_net_8_port
                           , p_out => p_net_8_port);
   pg_net_x_9 : pg_net_56 port map( a => A(9), b => B(9), g_out => g_net_9_port
                           , p_out => p_net_9_port);
   pg_net_x_10 : pg_net_55 port map( a => A(10), b => B(10), g_out => 
                           g_net_10_port, p_out => p_net_10_port);
   pg_net_x_11 : pg_net_54 port map( a => A(11), b => B(11), g_out => 
                           g_net_11_port, p_out => p_net_11_port);
   pg_net_x_12 : pg_net_53 port map( a => A(12), b => B(12), g_out => 
                           g_net_12_port, p_out => p_net_12_port);
   pg_net_x_13 : pg_net_52 port map( a => A(13), b => B(13), g_out => 
                           g_net_13_port, p_out => p_net_13_port);
   pg_net_x_14 : pg_net_51 port map( a => A(14), b => B(14), g_out => 
                           g_net_14_port, p_out => p_net_14_port);
   pg_net_x_15 : pg_net_50 port map( a => A(15), b => B(15), g_out => 
                           g_net_15_port, p_out => p_net_15_port);
   pg_net_x_16 : pg_net_49 port map( a => A(16), b => B(16), g_out => 
                           g_net_16_port, p_out => p_net_16_port);
   pg_net_x_17 : pg_net_48 port map( a => A(17), b => B(17), g_out => 
                           g_net_17_port, p_out => p_net_17_port);
   pg_net_x_18 : pg_net_47 port map( a => A(18), b => B(18), g_out => 
                           g_net_18_port, p_out => p_net_18_port);
   pg_net_x_19 : pg_net_46 port map( a => A(19), b => B(19), g_out => 
                           g_net_19_port, p_out => p_net_19_port);
   pg_net_x_20 : pg_net_45 port map( a => A(20), b => B(20), g_out => 
                           g_net_20_port, p_out => p_net_20_port);
   pg_net_x_21 : pg_net_44 port map( a => A(21), b => B(21), g_out => 
                           g_net_21_port, p_out => p_net_21_port);
   pg_net_x_22 : pg_net_43 port map( a => A(22), b => B(22), g_out => 
                           g_net_22_port, p_out => p_net_22_port);
   pg_net_x_23 : pg_net_42 port map( a => A(23), b => B(23), g_out => 
                           g_net_23_port, p_out => p_net_23_port);
   pg_net_x_24 : pg_net_41 port map( a => A(24), b => B(24), g_out => 
                           g_net_24_port, p_out => p_net_24_port);
   pg_net_x_25 : pg_net_40 port map( a => A(25), b => B(25), g_out => 
                           g_net_25_port, p_out => p_net_25_port);
   pg_net_x_26 : pg_net_39 port map( a => A(26), b => B(26), g_out => 
                           g_net_26_port, p_out => p_net_26_port);
   pg_net_x_27 : pg_net_38 port map( a => A(27), b => B(27), g_out => 
                           g_net_27_port, p_out => p_net_27_port);
   pg_net_0_MAGIC : pg_net_33 port map( a => A(0), b => B(0), g_out => 
                           magic_pro_0_port, p_out => net48715);
   xG_0_0_MAGIC : g_0 port map( g => magic_pro_0_port, p => n1, g_prec => n2, 
                           g_out => g_net_0_port);
   xG_1_0 : g_19 port map( g => g_net_1_port, p => p_net_1_port, g_prec => 
                           g_net_0_port, g_out => pg_1_0_0_port);
   xPG_1_1 : pg_0 port map( g => g_net_3_port, p => p_net_3_port, g_prec => 
                           g_net_2_port, p_prec => p_net_2_port, g_out => 
                           pg_1_1_0_port, p_out => pg_1_1_1_port);
   xPG_1_2 : pg_53 port map( g => g_net_5_port, p => p_net_5_port, g_prec => 
                           g_net_4_port, p_prec => p_net_4_port, g_out => 
                           pg_1_2_0_port, p_out => pg_1_2_1_port);
   xPG_1_3 : pg_52 port map( g => g_net_7_port, p => p_net_7_port, g_prec => 
                           g_net_6_port, p_prec => p_net_6_port, g_out => 
                           pg_1_3_0_port, p_out => pg_1_3_1_port);
   xPG_1_4 : pg_51 port map( g => g_net_9_port, p => p_net_9_port, g_prec => 
                           g_net_8_port, p_prec => p_net_8_port, g_out => 
                           pg_1_4_0_port, p_out => pg_1_4_1_port);
   xPG_1_5 : pg_50 port map( g => g_net_11_port, p => p_net_11_port, g_prec => 
                           g_net_10_port, p_prec => p_net_10_port, g_out => 
                           pg_1_5_0_port, p_out => pg_1_5_1_port);
   xPG_1_6 : pg_49 port map( g => g_net_13_port, p => p_net_13_port, g_prec => 
                           g_net_12_port, p_prec => p_net_12_port, g_out => 
                           pg_1_6_0_port, p_out => pg_1_6_1_port);
   xPG_1_7 : pg_48 port map( g => g_net_15_port, p => p_net_15_port, g_prec => 
                           g_net_14_port, p_prec => p_net_14_port, g_out => 
                           pg_1_7_0_port, p_out => pg_1_7_1_port);
   xPG_1_8 : pg_47 port map( g => g_net_17_port, p => p_net_17_port, g_prec => 
                           g_net_16_port, p_prec => p_net_16_port, g_out => 
                           pg_1_8_0_port, p_out => pg_1_8_1_port);
   xPG_1_9 : pg_46 port map( g => g_net_19_port, p => p_net_19_port, g_prec => 
                           g_net_18_port, p_prec => p_net_18_port, g_out => 
                           pg_1_9_0_port, p_out => pg_1_9_1_port);
   xPG_1_10 : pg_45 port map( g => g_net_21_port, p => p_net_21_port, g_prec =>
                           g_net_20_port, p_prec => p_net_20_port, g_out => 
                           pg_1_10_0_port, p_out => pg_1_10_1_port);
   xPG_1_11 : pg_44 port map( g => g_net_23_port, p => p_net_23_port, g_prec =>
                           g_net_22_port, p_prec => p_net_22_port, g_out => 
                           pg_1_11_0_port, p_out => pg_1_11_1_port);
   xPG_1_12 : pg_43 port map( g => g_net_25_port, p => p_net_25_port, g_prec =>
                           g_net_24_port, p_prec => p_net_24_port, g_out => 
                           pg_1_12_0_port, p_out => pg_1_12_1_port);
   xPG_1_13 : pg_42 port map( g => g_net_27_port, p => p_net_27_port, g_prec =>
                           g_net_26_port, p_prec => p_net_26_port, p_out => 
                           pg_1_13_1_port, g_out_BAR => pg_1_13_0_port);
   xG_2_0 : g_18 port map( g => pg_1_1_0_port, p => pg_1_1_1_port, g_prec => 
                           pg_1_0_0_port, g_out => Cout_0_port);
   xPG_2_1 : pg_39 port map( g => pg_1_3_0_port, p => pg_1_3_1_port, g_prec => 
                           pg_1_2_0_port, p_prec => pg_1_2_1_port, g_out => 
                           pg_n_2_1_0_port, p_out => pg_n_2_1_1_port);
   xPG_2_2 : pg_38 port map( g => pg_1_5_0_port, p => pg_1_5_1_port, g_prec => 
                           pg_1_4_0_port, p_prec => pg_1_4_1_port, g_out => 
                           pg_n_2_2_0_port, p_out => pg_n_2_2_1_port);
   xPG_2_3 : pg_37 port map( g => pg_1_7_0_port, p => pg_1_7_1_port, g_prec => 
                           pg_1_6_0_port, p_prec => pg_1_6_1_port, g_out => 
                           pg_n_2_3_0_port, p_out => pg_n_2_3_1_port);
   xPG_2_4 : pg_36 port map( g => pg_1_9_0_port, p => pg_1_9_1_port, g_prec => 
                           pg_1_8_0_port, p_prec => pg_1_8_1_port, g_out => 
                           pg_n_2_4_0_port, p_out => pg_n_2_4_1_port);
   xPG_2_5 : pg_35 port map( g => pg_1_11_0_port, p => pg_1_11_1_port, g_prec 
                           => pg_1_10_0_port, p_prec => pg_1_10_1_port, g_out 
                           => pg_n_2_5_0_port, p_out => pg_n_2_5_1_port);
   xPG_2_6 : pg_34 port map( p => pg_1_13_1_port, g_prec => pg_1_12_0_port, 
                           p_prec => pg_1_12_1_port, g_out => pg_n_2_6_0_port, 
                           p_out => pg_n_2_6_1_port, g_BAR => pg_1_13_0_port);
   xG_3_1 : g_17 port map( g => pg_n_2_1_0_port, p => pg_n_2_1_1_port, g_prec 
                           => Cout_0_port, g_out => Cout_1_port);
   xG_4_2 : g_16 port map( g => pg_n_2_2_0_port, p => pg_n_2_2_1_port, g_prec 
                           => Cout_1_port, g_out => Cout_2_port);
   xG_4_3 : g_15 port map( g => pg_n_3_3_0_port, p => pg_n_3_3_1_port, g_prec 
                           => Cout_1_port, g_out => Cout_3_port);
   xG_5_4 : g_14 port map( g => pg_n_2_4_0_port, p => pg_n_2_4_1_port, g_prec 
                           => Cout_3_port, g_out => Cout_4_port);
   xG_5_5 : g_13 port map( g => pg_n_3_5_0_port, p => pg_n_3_5_1_port, g_prec 
                           => Cout_3_port, g_out => Cout_5_port);
   xG_5_6 : g_12 port map( g => pg_n_4_6_0_port, p => pg_n_4_6_1_port, g_prec 
                           => Cout_3_port, g_out => Cout_6_port);
   xPG_3_3 : pg_32 port map( g => pg_n_2_3_0_port, p => pg_n_2_3_1_port, g_prec
                           => pg_n_2_2_0_port, p_prec => pg_n_2_2_1_port, g_out
                           => pg_n_3_3_0_port, p_out => pg_n_3_3_1_port);
   xPG_3_5 : pg_31 port map( g => pg_n_2_5_0_port, p => pg_n_2_5_1_port, g_prec
                           => pg_n_2_4_0_port, p_prec => pg_n_2_4_1_port, g_out
                           => pg_n_3_5_0_port, p_out => pg_n_3_5_1_port);
   xPG_4_6 : pg_29 port map( g => pg_n_2_6_0_port, p => pg_n_2_6_1_port, g_prec
                           => pg_n_3_5_0_port, p_prec => pg_n_3_5_1_port, g_out
                           => pg_n_4_6_0_port, p_out => pg_n_4_6_1_port);
   n1 <= '0';
   n2 <= '0';

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity xor_gen_N32_0 is

   port( A : in std_logic_vector (31 downto 0);  B : in std_logic;  S : out 
         std_logic_vector (31 downto 0));

end xor_gen_N32_0;

architecture SYN_bhe of xor_gen_N32_0 is

begin
   S <= ( A(31), A(30), A(29), A(28), A(27), A(26), A(25), A(24), A(23), A(22),
      A(21), A(20), A(19), A(18), A(17), A(16), A(15), A(14), A(13), A(12), 
      A(11), A(10), A(9), A(8), A(7), A(6), A(5), A(4), A(3), A(2), A(1), A(0) 
      );

end SYN_bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_ff32_en_IR is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_ff32_en_IR;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_ff32_en_IR is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net3585 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net3585);
   main_gate : AND2_X1 port map( A1 => net3585, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_ff32_en_0 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_ff32_en_0;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_ff32_en_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net3600 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net3600);
   main_gate : AND2_X1 port map( A1 => net3600, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity ff32_SIZE5 is

   port( D : in std_logic_vector (4 downto 0);  clk, rst : in std_logic;  Q : 
         out std_logic_vector (4 downto 0));

end ff32_SIZE5;

architecture SYN_behavioral of ff32_SIZE5 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n6, n2, n3, n4, n9 : std_logic;

begin
   
   Q_reg_4_inst : DFFR_X1 port map( D => D(4), CK => clk, RN => n9, Q => Q(4), 
                           QN => n6);
   Q_reg_0_inst : DFFR_X1 port map( D => D(0), CK => clk, RN => n9, Q => Q(0), 
                           QN => n1);
   Q_reg_3_inst : DFFR_X1 port map( D => D(3), CK => clk, RN => n9, Q => Q(3), 
                           QN => n4);
   Q_reg_2_inst : DFFR_X1 port map( D => D(2), CK => clk, RN => n9, Q => Q(2), 
                           QN => n3);
   Q_reg_1_inst : DFFR_X1 port map( D => D(1), CK => clk, RN => n9, Q => Q(1), 
                           QN => n2);
   U3 : INV_X1 port map( A => rst, ZN => n9);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity ff32_SIZE32 is

   port( D : in std_logic_vector (31 downto 0);  clk, rst : in std_logic;  Q : 
         out std_logic_vector (31 downto 0));

end ff32_SIZE32;

architecture SYN_behavioral of ff32_SIZE32 is

   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n33, n32 : std_logic;

begin
   
   Q_reg_31_inst : DFFR_X1 port map( D => D(31), CK => clk, RN => n32, Q => 
                           Q(31), QN => n33);
   Q_reg_30_inst : DFFR_X1 port map( D => D(30), CK => clk, RN => n32, Q => 
                           Q(30), QN => n31);
   Q_reg_29_inst : DFFR_X1 port map( D => D(29), CK => clk, RN => n32, Q => 
                           Q(29), QN => n30);
   Q_reg_28_inst : DFFR_X1 port map( D => D(28), CK => clk, RN => n32, Q => 
                           Q(28), QN => n29);
   Q_reg_27_inst : DFFR_X1 port map( D => D(27), CK => clk, RN => n32, Q => 
                           Q(27), QN => n28);
   Q_reg_26_inst : DFFR_X1 port map( D => D(26), CK => clk, RN => n32, Q => 
                           Q(26), QN => n27);
   Q_reg_25_inst : DFFR_X1 port map( D => D(25), CK => clk, RN => n32, Q => 
                           Q(25), QN => n26);
   Q_reg_24_inst : DFFR_X1 port map( D => D(24), CK => clk, RN => n32, Q => 
                           Q(24), QN => n25);
   Q_reg_23_inst : DFFR_X1 port map( D => D(23), CK => clk, RN => n32, Q => 
                           Q(23), QN => n24);
   Q_reg_22_inst : DFFR_X1 port map( D => D(22), CK => clk, RN => n32, Q => 
                           Q(22), QN => n23);
   Q_reg_21_inst : DFFR_X1 port map( D => D(21), CK => clk, RN => n32, Q => 
                           Q(21), QN => n22);
   Q_reg_20_inst : DFFR_X1 port map( D => D(20), CK => clk, RN => n32, Q => 
                           Q(20), QN => n21);
   Q_reg_19_inst : DFFR_X1 port map( D => D(19), CK => clk, RN => n32, Q => 
                           Q(19), QN => n20);
   Q_reg_18_inst : DFFR_X1 port map( D => D(18), CK => clk, RN => n32, Q => 
                           Q(18), QN => n19);
   Q_reg_17_inst : DFFR_X1 port map( D => D(17), CK => clk, RN => n32, Q => 
                           Q(17), QN => n18);
   Q_reg_16_inst : DFFR_X1 port map( D => D(16), CK => clk, RN => n32, Q => 
                           Q(16), QN => n17);
   Q_reg_15_inst : DFFR_X1 port map( D => D(15), CK => clk, RN => n32, Q => 
                           Q(15), QN => n16);
   Q_reg_14_inst : DFFR_X1 port map( D => D(14), CK => clk, RN => n32, Q => 
                           Q(14), QN => n15);
   Q_reg_13_inst : DFFR_X1 port map( D => D(13), CK => clk, RN => n32, Q => 
                           Q(13), QN => n14);
   Q_reg_12_inst : DFFR_X1 port map( D => D(12), CK => clk, RN => n32, Q => 
                           Q(12), QN => n13);
   Q_reg_11_inst : DFFR_X1 port map( D => D(11), CK => clk, RN => n32, Q => 
                           Q(11), QN => n12);
   Q_reg_10_inst : DFFR_X1 port map( D => D(10), CK => clk, RN => n32, Q => 
                           Q(10), QN => n11);
   Q_reg_9_inst : DFFR_X1 port map( D => D(9), CK => clk, RN => n32, Q => Q(9),
                           QN => n10);
   Q_reg_8_inst : DFFR_X1 port map( D => D(8), CK => clk, RN => n32, Q => Q(8),
                           QN => n9);
   Q_reg_7_inst : DFFR_X1 port map( D => D(7), CK => clk, RN => n32, Q => Q(7),
                           QN => n8);
   Q_reg_6_inst : DFFR_X1 port map( D => D(6), CK => clk, RN => n32, Q => Q(6),
                           QN => n7);
   Q_reg_5_inst : DFFR_X1 port map( D => D(5), CK => clk, RN => n32, Q => Q(5),
                           QN => n6);
   Q_reg_4_inst : DFFR_X1 port map( D => D(4), CK => clk, RN => n32, Q => Q(4),
                           QN => n5);
   Q_reg_3_inst : DFFR_X1 port map( D => D(3), CK => clk, RN => n32, Q => Q(3),
                           QN => n4);
   Q_reg_2_inst : DFFR_X1 port map( D => D(2), CK => clk, RN => n32, Q => Q(2),
                           QN => n3);
   Q_reg_1_inst : DFFR_X1 port map( D => D(1), CK => clk, RN => n32, Q => Q(1),
                           QN => n2);
   Q_reg_0_inst : DFFR_X1 port map( D => D(0), CK => clk, RN => n32, Q => Q(0),
                           QN => n1);
   U3 : INV_X2 port map( A => rst, ZN => n32);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity mux41_MUX_SIZE5 is

   port( IN0, IN1, IN2, IN3 : in std_logic_vector (4 downto 0);  CTRL : in 
         std_logic_vector (1 downto 0);  OUT1 : out std_logic_vector (4 downto 
         0));

end mux41_MUX_SIZE5;

architecture SYN_bhe of mux41_MUX_SIZE5 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7, n9, n10, n11, n12, n13, n14, n15, n16, n17 : 
      std_logic;

begin
   
   U7 : NAND2_X1 port map( A1 => n11, A2 => n12, ZN => OUT1(2));
   U17 : AOI22_X1 port map( A1 => n6, A2 => IN2(0), B1 => n7, B2 => IN1(0), ZN 
                           => n15);
   U4 : NAND2_X1 port map( A1 => n9, A2 => n10, ZN => OUT1(3));
   U10 : NAND2_X1 port map( A1 => n13, A2 => n14, ZN => OUT1(1));
   U20 : INV_X1 port map( A => CTRL(1), ZN => n17);
   U18 : AND2_X1 port map( A1 => n17, A2 => CTRL(0), ZN => n7);
   U19 : NOR2_X1 port map( A1 => CTRL(0), A2 => n17, ZN => n6);
   U16 : AND2_X1 port map( A1 => CTRL(0), A2 => CTRL(1), ZN => n5);
   U13 : NAND2_X1 port map( A1 => n15, A2 => n16, ZN => OUT1(0));
   U1 : INV_X1 port map( A => n5, ZN => n16);
   U2 : AOI21_X1 port map( B1 => n6, B2 => IN2(1), A => n5, ZN => n14);
   U3 : NAND2_X1 port map( A1 => n7, A2 => IN1(1), ZN => n13);
   U5 : AOI21_X1 port map( B1 => n6, B2 => IN2(2), A => n5, ZN => n12);
   U6 : NAND2_X1 port map( A1 => n7, A2 => IN1(2), ZN => n11);
   U8 : AOI21_X1 port map( B1 => n6, B2 => IN2(3), A => n5, ZN => n10);
   U9 : NAND2_X1 port map( A1 => n7, A2 => IN1(3), ZN => n9);
   U11 : AOI21_X1 port map( B1 => n6, B2 => IN2(4), A => n5, ZN => n4);
   U12 : NAND2_X1 port map( A1 => n7, A2 => IN1(4), ZN => n3);
   U14 : NAND2_X1 port map( A1 => n3, A2 => n4, ZN => OUT1(4));

end SYN_bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity real_alu_DATA_SIZE32 is

   port( IN1, IN2 : in std_logic_vector (31 downto 0);  ALUW_i : in 
         std_logic_vector (12 downto 0);  DOUT : out std_logic_vector (31 
         downto 0);  stall_o : out std_logic;  Clock, Reset : in std_logic);

end real_alu_DATA_SIZE32;

architecture SYN_Bhe of real_alu_DATA_SIZE32 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X4
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X2
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component logic_unit_SIZE32
      port( IN1, IN2 : in std_logic_vector (31 downto 0);  CTRL : in 
            std_logic_vector (1 downto 0);  OUT1 : out std_logic_vector (31 
            downto 0));
   end component;
   
   component shifter
      port( A : in std_logic_vector (31 downto 0);  B : in std_logic_vector (4 
            downto 0);  LOGIC_ARITH, LEFT_RIGHT : in std_logic;  OUTPUT : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component comparator_M32
      port( V : in std_logic;  SUM : in std_logic_vector (31 downto 0);  sel : 
            in std_logic_vector (2 downto 0);  sign : in std_logic;  S : out 
            std_logic;  C_BAR : in std_logic);
   end component;
   
   component p4add_N32_logN5_1
      port( A, B : in std_logic_vector (31 downto 0);  Cin, sign : in std_logic
            ;  S : out std_logic_vector (31 downto 0);  Cout_BAR : out 
            std_logic);
   end component;
   
   component simple_booth_add_ext_N16
      port( Clock, Reset, sign, enable : in std_logic;  valid : out std_logic; 
            A, B : in std_logic_vector (15 downto 0);  A_to_add, B_to_add : out
            std_logic_vector (31 downto 0);  sign_to_add : out std_logic;  
            final_out : out std_logic_vector (31 downto 0);  ACC_from_add : in 
            std_logic_vector (31 downto 0));
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal X_Logic0_port, mux_A_31_port, mux_A_30_port, mux_A_29_port, 
      mux_A_28_port, mux_A_27_port, mux_A_26_port, mux_A_25_port, mux_A_24_port
      , mux_A_23_port, mux_A_22_port, mux_A_21_port, mux_A_20_port, 
      mux_A_19_port, mux_A_18_port, mux_A_17_port, mux_A_16_port, mux_A_15_port
      , mux_A_14_port, mux_A_13_port, mux_A_12_port, mux_A_11_port, 
      mux_A_10_port, mux_A_9_port, mux_A_8_port, mux_A_7_port, mux_A_6_port, 
      mux_A_5_port, mux_A_4_port, mux_A_3_port, mux_A_2_port, mux_A_1_port, 
      mux_A_0_port, A_booth_to_add_31_port, A_booth_to_add_30_port, 
      A_booth_to_add_29_port, A_booth_to_add_28_port, A_booth_to_add_27_port, 
      A_booth_to_add_26_port, A_booth_to_add_25_port, A_booth_to_add_24_port, 
      A_booth_to_add_23_port, A_booth_to_add_22_port, A_booth_to_add_21_port, 
      A_booth_to_add_20_port, A_booth_to_add_19_port, A_booth_to_add_18_port, 
      A_booth_to_add_17_port, A_booth_to_add_16_port, A_booth_to_add_15_port, 
      A_booth_to_add_14_port, A_booth_to_add_13_port, A_booth_to_add_12_port, 
      A_booth_to_add_11_port, A_booth_to_add_10_port, A_booth_to_add_9_port, 
      A_booth_to_add_8_port, A_booth_to_add_7_port, A_booth_to_add_6_port, 
      A_booth_to_add_5_port, A_booth_to_add_4_port, A_booth_to_add_3_port, 
      A_booth_to_add_2_port, A_booth_to_add_1_port, A_booth_to_add_0_port, 
      mux_B_31_port, mux_B_30_port, mux_B_29_port, mux_B_28_port, mux_B_27_port
      , mux_B_26_port, mux_B_25_port, mux_B_24_port, mux_B_23_port, 
      mux_B_22_port, mux_B_21_port, mux_B_20_port, mux_B_19_port, mux_B_18_port
      , mux_B_17_port, mux_B_16_port, mux_B_15_port, mux_B_14_port, 
      mux_B_13_port, mux_B_12_port, mux_B_11_port, mux_B_10_port, mux_B_9_port,
      mux_B_8_port, mux_B_7_port, mux_B_6_port, mux_B_5_port, mux_B_4_port, 
      mux_B_3_port, mux_B_2_port, mux_B_1_port, mux_B_0_port, 
      B_booth_to_add_31_port, B_booth_to_add_30_port, B_booth_to_add_29_port, 
      B_booth_to_add_28_port, B_booth_to_add_27_port, B_booth_to_add_26_port, 
      B_booth_to_add_25_port, B_booth_to_add_24_port, B_booth_to_add_23_port, 
      B_booth_to_add_22_port, B_booth_to_add_21_port, B_booth_to_add_20_port, 
      B_booth_to_add_19_port, B_booth_to_add_18_port, B_booth_to_add_17_port, 
      B_booth_to_add_16_port, B_booth_to_add_15_port, B_booth_to_add_14_port, 
      B_booth_to_add_13_port, B_booth_to_add_12_port, B_booth_to_add_11_port, 
      B_booth_to_add_10_port, B_booth_to_add_9_port, B_booth_to_add_8_port, 
      B_booth_to_add_7_port, B_booth_to_add_6_port, B_booth_to_add_5_port, 
      B_booth_to_add_4_port, B_booth_to_add_3_port, B_booth_to_add_2_port, 
      B_booth_to_add_1_port, B_booth_to_add_0_port, mux_sign, sign_booth_to_add
      , valid_from_booth, mult_out_31_port, mult_out_30_port, mult_out_29_port,
      mult_out_28_port, mult_out_27_port, mult_out_26_port, mult_out_25_port, 
      mult_out_24_port, mult_out_23_port, mult_out_22_port, mult_out_21_port, 
      mult_out_20_port, mult_out_19_port, mult_out_18_port, mult_out_17_port, 
      mult_out_16_port, mult_out_15_port, mult_out_14_port, mult_out_13_port, 
      mult_out_12_port, mult_out_11_port, mult_out_10_port, mult_out_9_port, 
      mult_out_8_port, mult_out_7_port, mult_out_6_port, mult_out_5_port, 
      mult_out_4_port, mult_out_3_port, mult_out_2_port, mult_out_1_port, 
      mult_out_0_port, sum_out_31_port, sum_out_30_port, sum_out_29_port, 
      sum_out_28_port, sum_out_27_port, sum_out_26_port, sum_out_25_port, 
      sum_out_24_port, sum_out_23_port, sum_out_22_port, sum_out_21_port, 
      sum_out_20_port, sum_out_19_port, sum_out_18_port, sum_out_17_port, 
      sum_out_16_port, sum_out_15_port, sum_out_14_port, sum_out_13_port, 
      sum_out_12_port, sum_out_11_port, sum_out_10_port, sum_out_9_port, 
      sum_out_8_port, sum_out_7_port, sum_out_6_port, sum_out_5_port, 
      sum_out_4_port, sum_out_3_port, sum_out_2_port, sum_out_1_port, 
      sum_out_0_port, carry_from_adder, overflow, comp_out, shift_out_31_port, 
      shift_out_30_port, shift_out_29_port, shift_out_28_port, 
      shift_out_27_port, shift_out_26_port, shift_out_25_port, 
      shift_out_24_port, shift_out_23_port, shift_out_22_port, 
      shift_out_21_port, shift_out_20_port, shift_out_19_port, 
      shift_out_18_port, shift_out_17_port, shift_out_16_port, 
      shift_out_15_port, shift_out_14_port, shift_out_13_port, 
      shift_out_12_port, shift_out_11_port, shift_out_10_port, shift_out_9_port
      , shift_out_8_port, shift_out_7_port, shift_out_6_port, shift_out_5_port,
      shift_out_4_port, shift_out_3_port, shift_out_2_port, shift_out_1_port, 
      shift_out_0_port, lu_out_31_port, lu_out_30_port, lu_out_29_port, 
      lu_out_28_port, lu_out_27_port, lu_out_26_port, lu_out_25_port, 
      lu_out_24_port, lu_out_23_port, lu_out_22_port, lu_out_21_port, 
      lu_out_20_port, lu_out_19_port, lu_out_18_port, lu_out_17_port, 
      lu_out_16_port, lu_out_15_port, lu_out_14_port, lu_out_13_port, 
      lu_out_12_port, lu_out_11_port, lu_out_10_port, lu_out_9_port, 
      lu_out_8_port, lu_out_7_port, lu_out_6_port, lu_out_5_port, lu_out_4_port
      , lu_out_3_port, lu_out_2_port, lu_out_1_port, lu_out_0_port, n9, n11, 
      n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27
      , n28, n29, n30, n31, n32, n33, n34, n35, n36, n39, n40, n41, n42, n43, 
      n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58
      , n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, 
      n73, n74, n75, n76, n77, n78, n79, n80, n84, n85, n1, n2, n3, n4, n5, n6,
      n7, n8, n10, n12, n37, n38, n81, n83, n86, n87, n88, n89, n90, n91, n92, 
      n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, 
      n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, 
      n118, n119 : std_logic;

begin
   
   X_Logic0_port <= '0';
   U120 : MUX2_X1 port map( A => B_booth_to_add_31_port, B => IN2(31), S => n9,
                           Z => mux_B_31_port);
   U121 : MUX2_X1 port map( A => B_booth_to_add_30_port, B => IN2(30), S => n9,
                           Z => mux_B_30_port);
   U123 : MUX2_X1 port map( A => B_booth_to_add_29_port, B => IN2(29), S => n9,
                           Z => mux_B_29_port);
   U124 : MUX2_X1 port map( A => B_booth_to_add_28_port, B => IN2(28), S => n9,
                           Z => mux_B_28_port);
   U125 : MUX2_X1 port map( A => B_booth_to_add_27_port, B => IN2(27), S => n9,
                           Z => mux_B_27_port);
   U126 : MUX2_X1 port map( A => B_booth_to_add_26_port, B => IN2(26), S => n9,
                           Z => mux_B_26_port);
   U128 : MUX2_X1 port map( A => B_booth_to_add_24_port, B => IN2(24), S => n9,
                           Z => mux_B_24_port);
   U132 : MUX2_X1 port map( A => B_booth_to_add_20_port, B => IN2(20), S => n9,
                           Z => mux_B_20_port);
   U134 : MUX2_X1 port map( A => B_booth_to_add_19_port, B => IN2(19), S => n9,
                           Z => mux_B_19_port);
   U138 : MUX2_X1 port map( A => B_booth_to_add_15_port, B => IN2(15), S => n9,
                           Z => mux_B_15_port);
   U139 : MUX2_X1 port map( A => B_booth_to_add_14_port, B => IN2(14), S => n9,
                           Z => mux_B_14_port);
   U141 : MUX2_X1 port map( A => B_booth_to_add_12_port, B => IN2(12), S => n9,
                           Z => mux_B_12_port);
   U143 : MUX2_X1 port map( A => B_booth_to_add_10_port, B => IN2(10), S => n9,
                           Z => mux_B_10_port);
   U145 : MUX2_X1 port map( A => A_booth_to_add_9_port, B => IN1(9), S => n9, Z
                           => mux_A_9_port);
   U146 : MUX2_X1 port map( A => A_booth_to_add_8_port, B => IN1(8), S => n9, Z
                           => mux_A_8_port);
   U147 : MUX2_X1 port map( A => A_booth_to_add_7_port, B => IN1(7), S => n9, Z
                           => mux_A_7_port);
   U148 : MUX2_X1 port map( A => A_booth_to_add_6_port, B => IN1(6), S => n9, Z
                           => mux_A_6_port);
   U150 : MUX2_X1 port map( A => A_booth_to_add_4_port, B => IN1(4), S => n9, Z
                           => mux_A_4_port);
   U152 : MUX2_X1 port map( A => A_booth_to_add_31_port, B => IN1(31), S => n9,
                           Z => mux_A_31_port);
   U153 : MUX2_X1 port map( A => A_booth_to_add_30_port, B => IN1(30), S => n9,
                           Z => mux_A_30_port);
   U154 : MUX2_X1 port map( A => A_booth_to_add_2_port, B => IN1(2), S => n9, Z
                           => mux_A_2_port);
   U155 : MUX2_X1 port map( A => A_booth_to_add_29_port, B => IN1(29), S => n9,
                           Z => mux_A_29_port);
   U156 : MUX2_X1 port map( A => A_booth_to_add_28_port, B => IN1(28), S => n9,
                           Z => mux_A_28_port);
   U157 : MUX2_X1 port map( A => A_booth_to_add_27_port, B => IN1(27), S => n9,
                           Z => mux_A_27_port);
   U158 : MUX2_X1 port map( A => A_booth_to_add_26_port, B => IN1(26), S => n9,
                           Z => mux_A_26_port);
   U159 : MUX2_X1 port map( A => A_booth_to_add_25_port, B => IN1(25), S => n9,
                           Z => mux_A_25_port);
   U160 : MUX2_X1 port map( A => A_booth_to_add_24_port, B => IN1(24), S => n9,
                           Z => mux_A_24_port);
   U161 : MUX2_X1 port map( A => A_booth_to_add_23_port, B => IN1(23), S => n9,
                           Z => mux_A_23_port);
   U162 : MUX2_X1 port map( A => A_booth_to_add_22_port, B => IN1(22), S => n9,
                           Z => mux_A_22_port);
   U163 : MUX2_X1 port map( A => A_booth_to_add_21_port, B => IN1(21), S => n9,
                           Z => mux_A_21_port);
   U164 : MUX2_X1 port map( A => A_booth_to_add_20_port, B => IN1(20), S => n9,
                           Z => mux_A_20_port);
   U166 : MUX2_X1 port map( A => A_booth_to_add_19_port, B => IN1(19), S => n9,
                           Z => mux_A_19_port);
   U167 : MUX2_X1 port map( A => A_booth_to_add_18_port, B => IN1(18), S => n9,
                           Z => mux_A_18_port);
   U168 : MUX2_X1 port map( A => A_booth_to_add_17_port, B => IN1(17), S => n9,
                           Z => mux_A_17_port);
   U169 : MUX2_X1 port map( A => A_booth_to_add_16_port, B => IN1(16), S => n9,
                           Z => mux_A_16_port);
   U170 : MUX2_X1 port map( A => A_booth_to_add_15_port, B => IN1(15), S => n9,
                           Z => mux_A_15_port);
   U171 : MUX2_X1 port map( A => A_booth_to_add_14_port, B => IN1(14), S => n9,
                           Z => mux_A_14_port);
   U172 : MUX2_X1 port map( A => A_booth_to_add_13_port, B => IN1(13), S => n9,
                           Z => mux_A_13_port);
   U173 : MUX2_X1 port map( A => A_booth_to_add_12_port, B => IN1(12), S => n9,
                           Z => mux_A_12_port);
   U174 : MUX2_X1 port map( A => A_booth_to_add_11_port, B => IN1(11), S => n9,
                           Z => mux_A_11_port);
   U175 : MUX2_X1 port map( A => A_booth_to_add_10_port, B => IN1(10), S => n9,
                           Z => mux_A_10_port);
   U178 : NAND3_X1 port map( A1 => n84, A2 => n85, A3 => ALUW_i(12), ZN => n32)
                           ;
   MULT : simple_booth_add_ext_N16 port map( Clock => Clock, Reset => Reset, 
                           sign => ALUW_i(0), enable => ALUW_i(1), valid => 
                           valid_from_booth, A(15) => IN1(15), A(14) => IN1(14)
                           , A(13) => IN1(13), A(12) => IN1(12), A(11) => 
                           IN1(11), A(10) => IN1(10), A(9) => IN1(9), A(8) => 
                           IN1(8), A(7) => IN1(7), A(6) => IN1(6), A(5) => 
                           IN1(5), A(4) => IN1(4), A(3) => IN1(3), A(2) => 
                           IN1(2), A(1) => IN1(1), A(0) => n108, B(15) => n112,
                           B(14) => n110, B(13) => IN2(13), B(12) => IN2(12), 
                           B(11) => n111, B(10) => IN2(10), B(9) => n113, B(8) 
                           => IN2(8), B(7) => n107, B(6) => IN2(6), B(5) => 
                           n114, B(4) => IN2(4), B(3) => n117, B(2) => n81, 
                           B(1) => n115, B(0) => n116, A_to_add(31) => 
                           A_booth_to_add_31_port, A_to_add(30) => 
                           A_booth_to_add_30_port, A_to_add(29) => 
                           A_booth_to_add_29_port, A_to_add(28) => 
                           A_booth_to_add_28_port, A_to_add(27) => 
                           A_booth_to_add_27_port, A_to_add(26) => 
                           A_booth_to_add_26_port, A_to_add(25) => 
                           A_booth_to_add_25_port, A_to_add(24) => 
                           A_booth_to_add_24_port, A_to_add(23) => 
                           A_booth_to_add_23_port, A_to_add(22) => 
                           A_booth_to_add_22_port, A_to_add(21) => 
                           A_booth_to_add_21_port, A_to_add(20) => 
                           A_booth_to_add_20_port, A_to_add(19) => 
                           A_booth_to_add_19_port, A_to_add(18) => 
                           A_booth_to_add_18_port, A_to_add(17) => 
                           A_booth_to_add_17_port, A_to_add(16) => 
                           A_booth_to_add_16_port, A_to_add(15) => 
                           A_booth_to_add_15_port, A_to_add(14) => 
                           A_booth_to_add_14_port, A_to_add(13) => 
                           A_booth_to_add_13_port, A_to_add(12) => 
                           A_booth_to_add_12_port, A_to_add(11) => 
                           A_booth_to_add_11_port, A_to_add(10) => 
                           A_booth_to_add_10_port, A_to_add(9) => 
                           A_booth_to_add_9_port, A_to_add(8) => 
                           A_booth_to_add_8_port, A_to_add(7) => 
                           A_booth_to_add_7_port, A_to_add(6) => 
                           A_booth_to_add_6_port, A_to_add(5) => 
                           A_booth_to_add_5_port, A_to_add(4) => 
                           A_booth_to_add_4_port, A_to_add(3) => 
                           A_booth_to_add_3_port, A_to_add(2) => 
                           A_booth_to_add_2_port, A_to_add(1) => 
                           A_booth_to_add_1_port, A_to_add(0) => 
                           A_booth_to_add_0_port, B_to_add(31) => 
                           B_booth_to_add_31_port, B_to_add(30) => 
                           B_booth_to_add_30_port, B_to_add(29) => 
                           B_booth_to_add_29_port, B_to_add(28) => 
                           B_booth_to_add_28_port, B_to_add(27) => 
                           B_booth_to_add_27_port, B_to_add(26) => 
                           B_booth_to_add_26_port, B_to_add(25) => 
                           B_booth_to_add_25_port, B_to_add(24) => 
                           B_booth_to_add_24_port, B_to_add(23) => 
                           B_booth_to_add_23_port, B_to_add(22) => 
                           B_booth_to_add_22_port, B_to_add(21) => 
                           B_booth_to_add_21_port, B_to_add(20) => 
                           B_booth_to_add_20_port, B_to_add(19) => 
                           B_booth_to_add_19_port, B_to_add(18) => 
                           B_booth_to_add_18_port, B_to_add(17) => 
                           B_booth_to_add_17_port, B_to_add(16) => 
                           B_booth_to_add_16_port, B_to_add(15) => 
                           B_booth_to_add_15_port, B_to_add(14) => 
                           B_booth_to_add_14_port, B_to_add(13) => 
                           B_booth_to_add_13_port, B_to_add(12) => 
                           B_booth_to_add_12_port, B_to_add(11) => 
                           B_booth_to_add_11_port, B_to_add(10) => 
                           B_booth_to_add_10_port, B_to_add(9) => 
                           B_booth_to_add_9_port, B_to_add(8) => 
                           B_booth_to_add_8_port, B_to_add(7) => 
                           B_booth_to_add_7_port, B_to_add(6) => 
                           B_booth_to_add_6_port, B_to_add(5) => 
                           B_booth_to_add_5_port, B_to_add(4) => 
                           B_booth_to_add_4_port, B_to_add(3) => 
                           B_booth_to_add_3_port, B_to_add(2) => 
                           B_booth_to_add_2_port, B_to_add(1) => 
                           B_booth_to_add_1_port, B_to_add(0) => 
                           B_booth_to_add_0_port, sign_to_add => 
                           sign_booth_to_add, final_out(31) => mult_out_31_port
                           , final_out(30) => mult_out_30_port, final_out(29) 
                           => mult_out_29_port, final_out(28) => 
                           mult_out_28_port, final_out(27) => mult_out_27_port,
                           final_out(26) => mult_out_26_port, final_out(25) => 
                           mult_out_25_port, final_out(24) => mult_out_24_port,
                           final_out(23) => mult_out_23_port, final_out(22) => 
                           mult_out_22_port, final_out(21) => mult_out_21_port,
                           final_out(20) => mult_out_20_port, final_out(19) => 
                           mult_out_19_port, final_out(18) => mult_out_18_port,
                           final_out(17) => mult_out_17_port, final_out(16) => 
                           mult_out_16_port, final_out(15) => mult_out_15_port,
                           final_out(14) => mult_out_14_port, final_out(13) => 
                           mult_out_13_port, final_out(12) => mult_out_12_port,
                           final_out(11) => mult_out_11_port, final_out(10) => 
                           mult_out_10_port, final_out(9) => mult_out_9_port, 
                           final_out(8) => mult_out_8_port, final_out(7) => 
                           mult_out_7_port, final_out(6) => mult_out_6_port, 
                           final_out(5) => mult_out_5_port, final_out(4) => 
                           mult_out_4_port, final_out(3) => mult_out_3_port, 
                           final_out(2) => mult_out_2_port, final_out(1) => 
                           mult_out_1_port, final_out(0) => mult_out_0_port, 
                           ACC_from_add(31) => sum_out_31_port, 
                           ACC_from_add(30) => sum_out_30_port, 
                           ACC_from_add(29) => sum_out_29_port, 
                           ACC_from_add(28) => sum_out_28_port, 
                           ACC_from_add(27) => sum_out_27_port, 
                           ACC_from_add(26) => sum_out_26_port, 
                           ACC_from_add(25) => sum_out_25_port, 
                           ACC_from_add(24) => sum_out_24_port, 
                           ACC_from_add(23) => n87, ACC_from_add(22) => n86, 
                           ACC_from_add(21) => n38, ACC_from_add(20) => n88, 
                           ACC_from_add(19) => sum_out_19_port, 
                           ACC_from_add(18) => sum_out_18_port, 
                           ACC_from_add(17) => sum_out_17_port, 
                           ACC_from_add(16) => sum_out_16_port, 
                           ACC_from_add(15) => sum_out_15_port, 
                           ACC_from_add(14) => sum_out_14_port, 
                           ACC_from_add(13) => sum_out_13_port, 
                           ACC_from_add(12) => sum_out_12_port, 
                           ACC_from_add(11) => sum_out_11_port, 
                           ACC_from_add(10) => sum_out_10_port, ACC_from_add(9)
                           => sum_out_9_port, ACC_from_add(8) => sum_out_8_port
                           , ACC_from_add(7) => sum_out_7_port, ACC_from_add(6)
                           => sum_out_6_port, ACC_from_add(5) => sum_out_5_port
                           , ACC_from_add(4) => sum_out_4_port, ACC_from_add(3)
                           => sum_out_3_port, ACC_from_add(2) => sum_out_2_port
                           , ACC_from_add(1) => sum_out_1_port, ACC_from_add(0)
                           => sum_out_0_port);
   ADDER : p4add_N32_logN5_1 port map( A(31) => mux_A_31_port, A(30) => 
                           mux_A_30_port, A(29) => mux_A_29_port, A(28) => 
                           mux_A_28_port, A(27) => mux_A_27_port, A(26) => 
                           mux_A_26_port, A(25) => mux_A_25_port, A(24) => 
                           mux_A_24_port, A(23) => mux_A_23_port, A(22) => 
                           mux_A_22_port, A(21) => mux_A_21_port, A(20) => 
                           mux_A_20_port, A(19) => mux_A_19_port, A(18) => 
                           mux_A_18_port, A(17) => mux_A_17_port, A(16) => 
                           mux_A_16_port, A(15) => mux_A_15_port, A(14) => 
                           mux_A_14_port, A(13) => mux_A_13_port, A(12) => 
                           mux_A_12_port, A(11) => mux_A_11_port, A(10) => 
                           mux_A_10_port, A(9) => mux_A_9_port, A(8) => 
                           mux_A_8_port, A(7) => mux_A_7_port, A(6) => 
                           mux_A_6_port, A(5) => mux_A_5_port, A(4) => 
                           mux_A_4_port, A(3) => mux_A_3_port, A(2) => 
                           mux_A_2_port, A(1) => mux_A_1_port, A(0) => 
                           mux_A_0_port, B(31) => mux_B_31_port, B(30) => 
                           mux_B_30_port, B(29) => mux_B_29_port, B(28) => 
                           mux_B_28_port, B(27) => mux_B_27_port, B(26) => 
                           mux_B_26_port, B(25) => mux_B_25_port, B(24) => 
                           mux_B_24_port, B(23) => mux_B_23_port, B(22) => 
                           mux_B_22_port, B(21) => mux_B_21_port, B(20) => 
                           mux_B_20_port, B(19) => mux_B_19_port, B(18) => 
                           mux_B_18_port, B(17) => mux_B_17_port, B(16) => 
                           mux_B_16_port, B(15) => mux_B_15_port, B(14) => 
                           mux_B_14_port, B(13) => mux_B_13_port, B(12) => 
                           mux_B_12_port, B(11) => mux_B_11_port, B(10) => 
                           mux_B_10_port, B(9) => mux_B_9_port, B(8) => 
                           mux_B_8_port, B(7) => mux_B_7_port, B(6) => 
                           mux_B_6_port, B(5) => mux_B_5_port, B(4) => 
                           mux_B_4_port, B(3) => mux_B_3_port, B(2) => 
                           mux_B_2_port, B(1) => mux_B_1_port, B(0) => 
                           mux_B_0_port, Cin => X_Logic0_port, sign => mux_sign
                           , S(31) => sum_out_31_port, S(30) => sum_out_30_port
                           , S(29) => sum_out_29_port, S(28) => sum_out_28_port
                           , S(27) => sum_out_27_port, S(26) => sum_out_26_port
                           , S(25) => sum_out_25_port, S(24) => sum_out_24_port
                           , S(23) => sum_out_23_port, S(22) => sum_out_22_port
                           , S(21) => sum_out_21_port, S(20) => sum_out_20_port
                           , S(19) => sum_out_19_port, S(18) => sum_out_18_port
                           , S(17) => sum_out_17_port, S(16) => sum_out_16_port
                           , S(15) => sum_out_15_port, S(14) => sum_out_14_port
                           , S(13) => sum_out_13_port, S(12) => sum_out_12_port
                           , S(11) => sum_out_11_port, S(10) => sum_out_10_port
                           , S(9) => sum_out_9_port, S(8) => sum_out_8_port, 
                           S(7) => sum_out_7_port, S(6) => sum_out_6_port, S(5)
                           => sum_out_5_port, S(4) => sum_out_4_port, S(3) => 
                           sum_out_3_port, S(2) => sum_out_2_port, S(1) => 
                           sum_out_1_port, S(0) => sum_out_0_port, Cout_BAR => 
                           carry_from_adder);
   COMP : comparator_M32 port map( V => overflow, SUM(31) => sum_out_31_port, 
                           SUM(30) => sum_out_30_port, SUM(29) => 
                           sum_out_29_port, SUM(28) => sum_out_28_port, SUM(27)
                           => sum_out_27_port, SUM(26) => sum_out_26_port, 
                           SUM(25) => sum_out_25_port, SUM(24) => 
                           sum_out_24_port, SUM(23) => sum_out_23_port, SUM(22)
                           => sum_out_22_port, SUM(21) => sum_out_21_port, 
                           SUM(20) => sum_out_20_port, SUM(19) => 
                           sum_out_19_port, SUM(18) => sum_out_18_port, SUM(17)
                           => sum_out_17_port, SUM(16) => sum_out_16_port, 
                           SUM(15) => sum_out_15_port, SUM(14) => 
                           sum_out_14_port, SUM(13) => sum_out_13_port, SUM(12)
                           => sum_out_12_port, SUM(11) => sum_out_11_port, 
                           SUM(10) => sum_out_10_port, SUM(9) => sum_out_9_port
                           , SUM(8) => sum_out_8_port, SUM(7) => sum_out_7_port
                           , SUM(6) => sum_out_6_port, SUM(5) => sum_out_5_port
                           , SUM(4) => sum_out_4_port, SUM(3) => sum_out_3_port
                           , SUM(2) => sum_out_2_port, SUM(1) => sum_out_1_port
                           , SUM(0) => sum_out_0_port, sel(2) => ALUW_i(4), 
                           sel(1) => ALUW_i(3), sel(0) => ALUW_i(2), sign => 
                           ALUW_i(0), S => comp_out, C_BAR => carry_from_adder)
                           ;
   SHIFT : shifter port map( A(31) => IN1(31), A(30) => IN1(30), A(29) => 
                           IN1(29), A(28) => IN1(28), A(27) => IN1(27), A(26) 
                           => IN1(26), A(25) => IN1(25), A(24) => IN1(24), 
                           A(23) => IN1(23), A(22) => IN1(22), A(21) => IN1(21)
                           , A(20) => IN1(20), A(19) => IN1(19), A(18) => 
                           IN1(18), A(17) => IN1(17), A(16) => IN1(16), A(15) 
                           => IN1(15), A(14) => IN1(14), A(13) => IN1(13), 
                           A(12) => IN1(12), A(11) => IN1(11), A(10) => IN1(10)
                           , A(9) => IN1(9), A(8) => IN1(8), A(7) => IN1(7), 
                           A(6) => IN1(6), A(5) => IN1(5), A(4) => IN1(4), A(3)
                           => IN1(3), A(2) => IN1(2), A(1) => IN1(1), A(0) => 
                           n108, B(4) => IN2(4), B(3) => n117, B(2) => n81, 
                           B(1) => n115, B(0) => n116, LOGIC_ARITH => ALUW_i(8)
                           , LEFT_RIGHT => ALUW_i(9), OUTPUT(31) => 
                           shift_out_31_port, OUTPUT(30) => shift_out_30_port, 
                           OUTPUT(29) => shift_out_29_port, OUTPUT(28) => 
                           shift_out_28_port, OUTPUT(27) => shift_out_27_port, 
                           OUTPUT(26) => shift_out_26_port, OUTPUT(25) => 
                           shift_out_25_port, OUTPUT(24) => shift_out_24_port, 
                           OUTPUT(23) => shift_out_23_port, OUTPUT(22) => 
                           shift_out_22_port, OUTPUT(21) => shift_out_21_port, 
                           OUTPUT(20) => shift_out_20_port, OUTPUT(19) => 
                           shift_out_19_port, OUTPUT(18) => shift_out_18_port, 
                           OUTPUT(17) => shift_out_17_port, OUTPUT(16) => 
                           shift_out_16_port, OUTPUT(15) => shift_out_15_port, 
                           OUTPUT(14) => shift_out_14_port, OUTPUT(13) => 
                           shift_out_13_port, OUTPUT(12) => shift_out_12_port, 
                           OUTPUT(11) => shift_out_11_port, OUTPUT(10) => 
                           shift_out_10_port, OUTPUT(9) => shift_out_9_port, 
                           OUTPUT(8) => shift_out_8_port, OUTPUT(7) => 
                           shift_out_7_port, OUTPUT(6) => shift_out_6_port, 
                           OUTPUT(5) => shift_out_5_port, OUTPUT(4) => 
                           shift_out_4_port, OUTPUT(3) => shift_out_3_port, 
                           OUTPUT(2) => shift_out_2_port, OUTPUT(1) => 
                           shift_out_1_port, OUTPUT(0) => shift_out_0_port);
   LU : logic_unit_SIZE32 port map( IN1(31) => IN1(31), IN1(30) => IN1(30), 
                           IN1(29) => IN1(29), IN1(28) => IN1(28), IN1(27) => 
                           IN1(27), IN1(26) => IN1(26), IN1(25) => IN1(25), 
                           IN1(24) => IN1(24), IN1(23) => IN1(23), IN1(22) => 
                           IN1(22), IN1(21) => IN1(21), IN1(20) => IN1(20), 
                           IN1(19) => IN1(19), IN1(18) => IN1(18), IN1(17) => 
                           IN1(17), IN1(16) => IN1(16), IN1(15) => IN1(15), 
                           IN1(14) => IN1(14), IN1(13) => IN1(13), IN1(12) => 
                           IN1(12), IN1(11) => IN1(11), IN1(10) => IN1(10), 
                           IN1(9) => IN1(9), IN1(8) => IN1(8), IN1(7) => IN1(7)
                           , IN1(6) => IN1(6), IN1(5) => IN1(5), IN1(4) => 
                           IN1(4), IN1(3) => IN1(3), IN1(2) => IN1(2), IN1(1) 
                           => IN1(1), IN1(0) => n108, IN2(31) => IN2(31), 
                           IN2(30) => IN2(30), IN2(29) => IN2(29), IN2(28) => 
                           IN2(28), IN2(27) => IN2(27), IN2(26) => IN2(26), 
                           IN2(25) => IN2(25), IN2(24) => IN2(24), IN2(23) => 
                           n12, IN2(22) => n109, IN2(21) => IN2(21), IN2(20) =>
                           IN2(20), IN2(19) => n106, IN2(18) => IN2(18), 
                           IN2(17) => IN2(17), IN2(16) => IN2(16), IN2(15) => 
                           n112, IN2(14) => n110, IN2(13) => IN2(13), IN2(12) 
                           => IN2(12), IN2(11) => n111, IN2(10) => IN2(10), 
                           IN2(9) => n113, IN2(8) => IN2(8), IN2(7) => n107, 
                           IN2(6) => IN2(6), IN2(5) => n114, IN2(4) => IN2(4), 
                           IN2(3) => n117, IN2(2) => n81, IN2(1) => n115, 
                           IN2(0) => n116, CTRL(1) => ALUW_i(6), CTRL(0) => 
                           ALUW_i(5), OUT1(31) => lu_out_31_port, OUT1(30) => 
                           lu_out_30_port, OUT1(29) => lu_out_29_port, OUT1(28)
                           => lu_out_28_port, OUT1(27) => lu_out_27_port, 
                           OUT1(26) => lu_out_26_port, OUT1(25) => 
                           lu_out_25_port, OUT1(24) => lu_out_24_port, OUT1(23)
                           => lu_out_23_port, OUT1(22) => lu_out_22_port, 
                           OUT1(21) => lu_out_21_port, OUT1(20) => 
                           lu_out_20_port, OUT1(19) => lu_out_19_port, OUT1(18)
                           => lu_out_18_port, OUT1(17) => lu_out_17_port, 
                           OUT1(16) => lu_out_16_port, OUT1(15) => 
                           lu_out_15_port, OUT1(14) => lu_out_14_port, OUT1(13)
                           => lu_out_13_port, OUT1(12) => lu_out_12_port, 
                           OUT1(11) => lu_out_11_port, OUT1(10) => 
                           lu_out_10_port, OUT1(9) => lu_out_9_port, OUT1(8) =>
                           lu_out_8_port, OUT1(7) => lu_out_7_port, OUT1(6) => 
                           lu_out_6_port, OUT1(5) => lu_out_5_port, OUT1(4) => 
                           lu_out_4_port, OUT1(3) => lu_out_3_port, OUT1(2) => 
                           lu_out_2_port, OUT1(1) => lu_out_1_port, OUT1(0) => 
                           lu_out_0_port);
   U114 : MUX2_X1 port map( A => B_booth_to_add_8_port, B => IN2(8), S => n9, Z
                           => mux_B_8_port);
   U137 : MUX2_X1 port map( A => B_booth_to_add_16_port, B => IN2(16), S => n9,
                           Z => mux_B_16_port);
   U13 : AOI22_X1 port map( A1 => n15, A2 => shift_out_7_port, B1 => n119, B2 
                           => sum_out_7_port, ZN => n23);
   U12 : NAND2_X1 port map( A1 => n22, A2 => n23, ZN => DOUT(7));
   U38 : AOI22_X1 port map( A1 => n83, A2 => shift_out_29_port, B1 => n119, B2 
                           => sum_out_29_port, ZN => n40);
   U37 : NAND2_X1 port map( A1 => n39, A2 => n40, ZN => DOUT(29));
   U56 : AOI22_X1 port map( A1 => n83, A2 => shift_out_23_port, B1 => n119, B2 
                           => n87, ZN => n52);
   U55 : NAND2_X1 port map( A1 => n51, A2 => n52, ZN => DOUT(23));
   U83 : AOI22_X1 port map( A1 => n83, A2 => shift_out_15_port, B1 => n119, B2 
                           => sum_out_15_port, ZN => n70);
   U82 : NAND2_X1 port map( A1 => n69, A2 => n70, ZN => DOUT(15));
   U72 : AOI222_X1 port map( A1 => n106, A2 => n17, B1 => n118, B2 => 
                           lu_out_19_port, C1 => n19, C2 => mult_out_19_port, 
                           ZN => n61);
   U71 : AOI22_X1 port map( A1 => n83, A2 => shift_out_19_port, B1 => n119, B2 
                           => sum_out_19_port, ZN => n62);
   U70 : NAND2_X1 port map( A1 => n61, A2 => n62, ZN => DOUT(19));
   U75 : AOI222_X1 port map( A1 => IN2(18), A2 => n17, B1 => n18, B2 => 
                           lu_out_18_port, C1 => n19, C2 => mult_out_18_port, 
                           ZN => n63);
   U74 : AOI22_X1 port map( A1 => n83, A2 => shift_out_18_port, B1 => n119, B2 
                           => sum_out_18_port, ZN => n64);
   U73 : NAND2_X1 port map( A1 => n63, A2 => n64, ZN => DOUT(18));
   U78 : AOI222_X1 port map( A1 => IN2(17), A2 => n17, B1 => n118, B2 => 
                           lu_out_17_port, C1 => n19, C2 => mult_out_17_port, 
                           ZN => n65);
   U77 : AOI22_X1 port map( A1 => n83, A2 => shift_out_17_port, B1 => n119, B2 
                           => sum_out_17_port, ZN => n66);
   U76 : NAND2_X1 port map( A1 => n65, A2 => n66, ZN => DOUT(17));
   U51 : AOI222_X1 port map( A1 => IN2(25), A2 => n17, B1 => n118, B2 => 
                           lu_out_25_port, C1 => n19, C2 => mult_out_25_port, 
                           ZN => n47);
   U50 : AOI22_X1 port map( A1 => n83, A2 => shift_out_25_port, B1 => n119, B2 
                           => sum_out_25_port, ZN => n48);
   U49 : NAND2_X1 port map( A1 => n47, A2 => n48, ZN => DOUT(25));
   U45 : AOI222_X1 port map( A1 => IN2(27), A2 => n17, B1 => n118, B2 => 
                           lu_out_27_port, C1 => n19, C2 => mult_out_27_port, 
                           ZN => n43);
   U44 : AOI22_X1 port map( A1 => n83, A2 => shift_out_27_port, B1 => n119, B2 
                           => sum_out_27_port, ZN => n44);
   U43 : NAND2_X1 port map( A1 => n43, A2 => n44, ZN => DOUT(27));
   U48 : AOI222_X1 port map( A1 => IN2(26), A2 => n17, B1 => n118, B2 => 
                           lu_out_26_port, C1 => n19, C2 => mult_out_26_port, 
                           ZN => n45);
   U47 : AOI22_X1 port map( A1 => n83, A2 => shift_out_26_port, B1 => n119, B2 
                           => sum_out_26_port, ZN => n46);
   U46 : NAND2_X1 port map( A1 => n45, A2 => n46, ZN => DOUT(26));
   U33 : AOI222_X1 port map( A1 => IN2(30), A2 => n17, B1 => n118, B2 => 
                           lu_out_30_port, C1 => n19, C2 => mult_out_30_port, 
                           ZN => n35);
   U32 : AOI22_X1 port map( A1 => n83, A2 => shift_out_30_port, B1 => n119, B2 
                           => sum_out_30_port, ZN => n36);
   U31 : NAND2_X1 port map( A1 => n35, A2 => n36, ZN => DOUT(30));
   U54 : AOI222_X1 port map( A1 => IN2(24), A2 => n17, B1 => n118, B2 => 
                           lu_out_24_port, C1 => n19, C2 => mult_out_24_port, 
                           ZN => n49);
   U52 : NAND2_X1 port map( A1 => n49, A2 => n50, ZN => DOUT(24));
   U60 : AOI222_X1 port map( A1 => n109, A2 => n17, B1 => n118, B2 => 
                           lu_out_22_port, C1 => n19, C2 => mult_out_22_port, 
                           ZN => n53);
   U58 : NAND2_X1 port map( A1 => n53, A2 => n54, ZN => DOUT(22));
   U63 : AOI222_X1 port map( A1 => IN2(21), A2 => n17, B1 => n118, B2 => 
                           lu_out_21_port, C1 => n19, C2 => mult_out_21_port, 
                           ZN => n55);
   U61 : NAND2_X1 port map( A1 => n55, A2 => n56, ZN => DOUT(21));
   U28 : AOI22_X1 port map( A1 => n118, A2 => lu_out_31_port, B1 => n19, B2 => 
                           mult_out_31_port, ZN => n34);
   U27 : OAI211_X1 port map( C1 => n32, C2 => n11, A => n33, B => n34, ZN => 
                           DOUT(31));
   U66 : AOI222_X1 port map( A1 => IN2(20), A2 => n17, B1 => n118, B2 => 
                           lu_out_20_port, C1 => n19, C2 => mult_out_20_port, 
                           ZN => n57);
   U64 : NAND2_X1 port map( A1 => n57, A2 => n58, ZN => DOUT(20));
   U42 : AOI222_X1 port map( A1 => IN2(28), A2 => n17, B1 => n118, B2 => 
                           lu_out_28_port, C1 => n19, C2 => mult_out_28_port, 
                           ZN => n41);
   U40 : NAND2_X1 port map( A1 => n41, A2 => n42, ZN => DOUT(28));
   U87 : AOI222_X1 port map( A1 => n110, A2 => n17, B1 => n118, B2 => 
                           lu_out_14_port, C1 => n19, C2 => mult_out_14_port, 
                           ZN => n71);
   U86 : AOI22_X1 port map( A1 => n83, A2 => shift_out_14_port, B1 => n119, B2 
                           => sum_out_14_port, ZN => n72);
   U85 : NAND2_X1 port map( A1 => n71, A2 => n72, ZN => DOUT(14));
   U26 : AOI222_X1 port map( A1 => n117, A2 => n17, B1 => n118, B2 => 
                           lu_out_3_port, C1 => n19, C2 => mult_out_3_port, ZN 
                           => n30);
   U25 : AOI22_X1 port map( A1 => n83, A2 => shift_out_3_port, B1 => n119, B2 
                           => sum_out_3_port, ZN => n31);
   U24 : NAND2_X1 port map( A1 => n30, A2 => n31, ZN => DOUT(3));
   U92 : AOI22_X1 port map( A1 => n83, A2 => shift_out_12_port, B1 => n119, B2 
                           => sum_out_12_port, ZN => n76);
   U91 : NAND2_X1 port map( A1 => n75, A2 => n76, ZN => DOUT(12));
   U95 : AOI22_X1 port map( A1 => n83, A2 => shift_out_11_port, B1 => n119, B2 
                           => sum_out_11_port, ZN => n78);
   U94 : NAND2_X1 port map( A1 => n77, A2 => n78, ZN => DOUT(11));
   U81 : AOI222_X1 port map( A1 => IN2(16), A2 => n17, B1 => n118, B2 => 
                           lu_out_16_port, C1 => n19, C2 => mult_out_16_port, 
                           ZN => n67);
   U80 : AOI22_X1 port map( A1 => n83, A2 => shift_out_16_port, B1 => n119, B2 
                           => sum_out_16_port, ZN => n68);
   U79 : NAND2_X1 port map( A1 => n67, A2 => n68, ZN => DOUT(16));
   U88 : NAND2_X1 port map( A1 => n73, A2 => n74, ZN => DOUT(13));
   U7 : AOI22_X1 port map( A1 => n15, A2 => shift_out_9_port, B1 => n119, B2 =>
                           sum_out_9_port, ZN => n14);
   U6 : NAND2_X1 port map( A1 => n13, A2 => n14, ZN => DOUT(9));
   U16 : AOI22_X1 port map( A1 => n83, A2 => shift_out_6_port, B1 => n16, B2 =>
                           sum_out_6_port, ZN => n25);
   U15 : NAND2_X1 port map( A1 => n24, A2 => n25, ZN => DOUT(6));
   U11 : AOI222_X1 port map( A1 => IN2(8), A2 => n17, B1 => n118, B2 => 
                           lu_out_8_port, C1 => n19, C2 => mult_out_8_port, ZN 
                           => n20);
   U10 : AOI22_X1 port map( A1 => n83, A2 => shift_out_8_port, B1 => n119, B2 
                           => sum_out_8_port, ZN => n21);
   U9 : NAND2_X1 port map( A1 => n20, A2 => n21, ZN => DOUT(8));
   U98 : AOI22_X1 port map( A1 => n83, A2 => shift_out_10_port, B1 => n119, B2 
                           => sum_out_10_port, ZN => n80);
   U97 : NAND2_X1 port map( A1 => n79, A2 => n80, ZN => DOUT(10));
   U19 : AOI22_X1 port map( A1 => n83, A2 => shift_out_5_port, B1 => n119, B2 
                           => sum_out_5_port, ZN => n27);
   U18 : NAND2_X1 port map( A1 => n26, A2 => n27, ZN => DOUT(5));
   U23 : AOI222_X1 port map( A1 => IN2(4), A2 => n17, B1 => n118, B2 => 
                           lu_out_4_port, C1 => n19, C2 => mult_out_4_port, ZN 
                           => n28);
   U22 : AOI22_X1 port map( A1 => n83, A2 => shift_out_4_port, B1 => n119, B2 
                           => sum_out_4_port, ZN => n29);
   U21 : NAND2_X1 port map( A1 => n28, A2 => n29, ZN => DOUT(4));
   U68 : AOI22_X1 port map( A1 => n83, A2 => shift_out_1_port, B1 => n119, B2 
                           => sum_out_1_port, ZN => n60);
   U67 : NAND2_X1 port map( A1 => n59, A2 => n60, ZN => DOUT(1));
   U108 : INV_X1 port map( A => ALUW_i(11), ZN => n84);
   U112 : MUX2_X2 port map( A => sign_booth_to_add, B => ALUW_i(7), S => n9, Z 
                           => mux_sign);
   U2 : NOR2_X1 port map( A1 => valid_from_booth, A2 => n9, ZN => stall_o);
   U3 : MUX2_X1 port map( A => B_booth_to_add_23_port, B => IN2(23), S => n9, Z
                           => mux_B_23_port);
   U4 : AOI22_X1 port map( A1 => ALUW_i(1), A2 => B_booth_to_add_5_port, B1 => 
                           n9, B2 => IN2(5), ZN => n1);
   U5 : INV_X1 port map( A => n1, ZN => mux_B_5_port);
   U8 : MUX2_X1 port map( A => B_booth_to_add_6_port, B => IN2(6), S => n9, Z 
                           => mux_B_6_port);
   U14 : MUX2_X1 port map( A => B_booth_to_add_3_port, B => IN2(3), S => n9, Z 
                           => mux_B_3_port);
   U17 : AOI222_X1 port map( A1 => sum_out_0_port, A2 => n119, B1 => n118, B2 
                           => lu_out_0_port, C1 => n116, C2 => n17, ZN => n2);
   U20 : INV_X1 port map( A => n2, ZN => n3);
   U29 : AOI21_X1 port map( B1 => n19, B2 => mult_out_0_port, A => n3, ZN => 
                           n104);
   U30 : AOI22_X1 port map( A1 => ALUW_i(1), A2 => B_booth_to_add_13_port, B1 
                           => n9, B2 => IN2(13), ZN => n4);
   U34 : INV_X1 port map( A => n4, ZN => mux_B_13_port);
   U35 : MUX2_X1 port map( A => A_booth_to_add_5_port, B => IN1(5), S => n9, Z 
                           => mux_A_5_port);
   U36 : MUX2_X1 port map( A => B_booth_to_add_7_port, B => IN2(7), S => n9, Z 
                           => mux_B_7_port);
   U39 : INV_X1 port map( A => ALUW_i(10), ZN => n5);
   U41 : NOR3_X1 port map( A1 => ALUW_i(12), A2 => n84, A3 => n5, ZN => n90);
   U53 : INV_X1 port map( A => n17, ZN => n6);
   U57 : INV_X1 port map( A => n81, ZN => n7);
   U59 : AOI22_X1 port map( A1 => mult_out_2_port, A2 => n19, B1 => 
                           lu_out_2_port, B2 => n118, ZN => n8);
   U62 : AOI22_X1 port map( A1 => sum_out_2_port, A2 => n119, B1 => 
                           shift_out_2_port, B2 => n83, ZN => n10);
   U65 : OAI211_X1 port map( C1 => n6, C2 => n7, A => n8, B => n10, ZN => 
                           DOUT(2));
   U69 : CLKBUF_X1 port map( A => IN2(23), Z => n12);
   U84 : CLKBUF_X1 port map( A => sum_out_31_port, Z => n37);
   U89 : CLKBUF_X1 port map( A => sum_out_21_port, Z => n38);
   U90 : CLKBUF_X1 port map( A => IN2(2), Z => n81);
   U93 : BUF_X1 port map( A => IN2(3), Z => n117);
   U96 : BUF_X1 port map( A => IN2(15), Z => n112);
   U99 : BUF_X1 port map( A => IN1(0), Z => n108);
   U100 : AND2_X1 port map( A1 => n105, A2 => n104, ZN => n89);
   U101 : BUF_X1 port map( A => IN2(5), Z => n114);
   U102 : BUF_X1 port map( A => IN2(14), Z => n110);
   U103 : BUF_X1 port map( A => IN2(1), Z => n115);
   U104 : BUF_X1 port map( A => IN2(9), Z => n113);
   U105 : BUF_X1 port map( A => n18, Z => n118);
   U106 : AND2_X2 port map( A1 => n32, A2 => ALUW_i(12), ZN => n19);
   U107 : BUF_X1 port map( A => n16, Z => n119);
   U109 : BUF_X2 port map( A => n15, Z => n83);
   U110 : INV_X2 port map( A => n32, ZN => n17);
   U111 : CLKBUF_X1 port map( A => sum_out_22_port, Z => n86);
   U113 : CLKBUF_X1 port map( A => sum_out_23_port, Z => n87);
   U115 : CLKBUF_X1 port map( A => sum_out_20_port, Z => n88);
   U116 : NAND2_X1 port map( A1 => n103, A2 => n89, ZN => DOUT(0));
   U117 : AOI222_X1 port map( A1 => IN2(13), A2 => n17, B1 => n18, B2 => 
                           lu_out_13_port, C1 => n19, C2 => mult_out_13_port, 
                           ZN => n73);
   U118 : NAND2_X1 port map( A1 => comp_out, A2 => n90, ZN => n103);
   U119 : CLKBUF_X1 port map( A => IN2(11), Z => n111);
   U122 : CLKBUF_X1 port map( A => IN2(22), Z => n109);
   U127 : CLKBUF_X1 port map( A => IN2(19), Z => n106);
   U129 : CLKBUF_X1 port map( A => IN2(7), Z => n107);
   U130 : CLKBUF_X1 port map( A => IN2(0), Z => n116);
   U131 : INV_X1 port map( A => ALUW_i(10), ZN => n85);
   U133 : INV_X1 port map( A => IN2(31), ZN => n11);
   U135 : OR2_X1 port map( A1 => n9, A2 => n97, ZN => n92);
   U136 : INV_X1 port map( A => B_booth_to_add_11_port, ZN => n97);
   U140 : OR2_X1 port map( A1 => n9, A2 => n99, ZN => n93);
   U142 : INV_X1 port map( A => B_booth_to_add_0_port, ZN => n99);
   U144 : OR2_X1 port map( A1 => n9, A2 => n95, ZN => n91);
   U149 : INV_X1 port map( A => B_booth_to_add_1_port, ZN => n95);
   U151 : INV_X4 port map( A => ALUW_i(1), ZN => n9);
   U165 : NOR3_X1 port map( A1 => ALUW_i(12), A2 => ALUW_i(10), A3 => n84, ZN 
                           => n15);
   U176 : NOR3_X1 port map( A1 => ALUW_i(11), A2 => ALUW_i(12), A3 => n85, ZN 
                           => n18);
   U177 : NOR3_X1 port map( A1 => ALUW_i(11), A2 => ALUW_i(12), A3 => 
                           ALUW_i(10), ZN => n16);
   U179 : AOI222_X1 port map( A1 => n115, A2 => n17, B1 => n118, B2 => 
                           lu_out_1_port, C1 => n19, C2 => mult_out_1_port, ZN 
                           => n59);
   U180 : AOI222_X1 port map( A1 => n113, A2 => n17, B1 => n18, B2 => 
                           lu_out_9_port, C1 => n19, C2 => mult_out_9_port, ZN 
                           => n13);
   U181 : AOI222_X1 port map( A1 => n111, A2 => n17, B1 => n18, B2 => 
                           lu_out_11_port, C1 => n19, C2 => mult_out_11_port, 
                           ZN => n77);
   U182 : AOI222_X1 port map( A1 => n112, A2 => n17, B1 => n118, B2 => 
                           lu_out_15_port, C1 => n19, C2 => mult_out_15_port, 
                           ZN => n69);
   U183 : AOI222_X1 port map( A1 => n12, A2 => n17, B1 => n18, B2 => 
                           lu_out_23_port, C1 => n19, C2 => mult_out_23_port, 
                           ZN => n51);
   U184 : AOI222_X1 port map( A1 => IN2(29), A2 => n17, B1 => n118, B2 => 
                           lu_out_29_port, C1 => n19, C2 => mult_out_29_port, 
                           ZN => n39);
   U185 : AOI222_X1 port map( A1 => n107, A2 => n17, B1 => n118, B2 => 
                           lu_out_7_port, C1 => n19, C2 => mult_out_7_port, ZN 
                           => n22);
   U186 : NAND2_X1 port map( A1 => shift_out_0_port, A2 => n83, ZN => n105);
   U187 : NOR2_X1 port map( A1 => n11, A2 => IN1(31), ZN => n102);
   U188 : NAND2_X1 port map( A1 => IN1(31), A2 => n11, ZN => n100);
   U189 : MUX2_X1 port map( A => B_booth_to_add_25_port, B => IN2(25), S => n9,
                           Z => mux_B_25_port);
   U190 : MUX2_X1 port map( A => B_booth_to_add_17_port, B => IN2(17), S => n9,
                           Z => mux_B_17_port);
   U191 : MUX2_X1 port map( A => B_booth_to_add_18_port, B => IN2(18), S => n9,
                           Z => mux_B_18_port);
   U192 : MUX2_X1 port map( A => B_booth_to_add_22_port, B => IN2(22), S => n9,
                           Z => mux_B_22_port);
   U193 : MUX2_X1 port map( A => B_booth_to_add_21_port, B => IN2(21), S => n9,
                           Z => mux_B_21_port);
   U194 : MUX2_X1 port map( A => B_booth_to_add_9_port, B => IN2(9), S => n9, Z
                           => mux_B_9_port);
   U195 : MUX2_X1 port map( A => B_booth_to_add_4_port, B => IN2(4), S => n9, Z
                           => mux_B_4_port);
   U196 : MUX2_X1 port map( A => B_booth_to_add_2_port, B => IN2(2), S => n9, Z
                           => mux_B_2_port);
   U197 : MUX2_X1 port map( A => A_booth_to_add_3_port, B => IN1(3), S => n9, Z
                           => mux_A_3_port);
   U198 : MUX2_X1 port map( A => A_booth_to_add_0_port, B => IN1(0), S => n9, Z
                           => mux_A_0_port);
   U199 : MUX2_X1 port map( A => A_booth_to_add_1_port, B => IN1(1), S => n9, Z
                           => mux_A_1_port);
   U200 : NAND2_X1 port map( A1 => n98, A2 => n93, ZN => mux_B_0_port);
   U201 : NAND2_X1 port map( A1 => IN2(1), A2 => n9, ZN => n94);
   U202 : NAND2_X1 port map( A1 => n94, A2 => n91, ZN => mux_B_1_port);
   U203 : NAND2_X1 port map( A1 => IN2(11), A2 => n9, ZN => n96);
   U204 : NAND2_X1 port map( A1 => n96, A2 => n92, ZN => mux_B_11_port);
   U205 : NAND2_X1 port map( A1 => IN2(0), A2 => n9, ZN => n98);
   U206 : NAND2_X1 port map( A1 => sum_out_31_port, A2 => n102, ZN => n101);
   U207 : OAI21_X1 port map( B1 => sum_out_31_port, B2 => n100, A => n101, ZN 
                           => overflow);
   U208 : AOI222_X1 port map( A1 => IN2(6), A2 => n17, B1 => n118, B2 => 
                           lu_out_6_port, C1 => n19, C2 => mult_out_6_port, ZN 
                           => n24);
   U209 : AOI222_X1 port map( A1 => IN2(10), A2 => n17, B1 => n118, B2 => 
                           lu_out_10_port, C1 => n19, C2 => mult_out_10_port, 
                           ZN => n79);
   U210 : AOI222_X1 port map( A1 => IN2(12), A2 => n17, B1 => n18, B2 => 
                           lu_out_12_port, C1 => n19, C2 => mult_out_12_port, 
                           ZN => n75);
   U211 : AOI22_X1 port map( A1 => n83, A2 => shift_out_13_port, B1 => n119, B2
                           => sum_out_13_port, ZN => n74);
   U212 : AOI222_X1 port map( A1 => n114, A2 => n17, B1 => n118, B2 => 
                           lu_out_5_port, C1 => n19, C2 => mult_out_5_port, ZN 
                           => n26);
   U213 : AOI22_X1 port map( A1 => n83, A2 => shift_out_22_port, B1 => n16, B2 
                           => n86, ZN => n54);
   U214 : AOI22_X1 port map( A1 => n83, A2 => shift_out_21_port, B1 => n16, B2 
                           => n38, ZN => n56);
   U215 : AOI22_X1 port map( A1 => n83, A2 => shift_out_28_port, B1 => n16, B2 
                           => sum_out_28_port, ZN => n42);
   U216 : AOI22_X1 port map( A1 => n83, A2 => shift_out_20_port, B1 => n88, B2 
                           => n16, ZN => n58);
   U217 : AOI22_X1 port map( A1 => n83, A2 => shift_out_24_port, B1 => n16, B2 
                           => sum_out_24_port, ZN => n50);
   U218 : AOI22_X1 port map( A1 => n83, A2 => shift_out_31_port, B1 => n119, B2
                           => n37, ZN => n33);

end SYN_Bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity ff32_en_SIZE13 is

   port( D : in std_logic_vector (12 downto 0);  en, clk, rst : in std_logic;  
         Q : out std_logic_vector (12 downto 0));

end ff32_en_SIZE13;

architecture SYN_behavioral of ff32_en_SIZE13 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X2
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_ff32_en_SIZE13
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal net3376, n1, n2, n3, n4, n5, n7, n8, n9, n11, n12, n14, n6, n10, n13 
      : std_logic;

begin
   
   Q_reg_12_inst : DFFR_X1 port map( D => D(12), CK => net3376, RN => n13, Q =>
                           Q(12), QN => n14);
   Q_reg_11_inst : DFFR_X1 port map( D => D(11), CK => net3376, RN => n13, Q =>
                           Q(11), QN => n12);
   Q_reg_10_inst : DFFR_X1 port map( D => D(10), CK => net3376, RN => n13, Q =>
                           Q(10), QN => n11);
   Q_reg_8_inst : DFFR_X1 port map( D => D(8), CK => net3376, RN => n13, Q => 
                           Q(8), QN => n9);
   Q_reg_7_inst : DFFR_X1 port map( D => D(7), CK => net3376, RN => n13, Q => 
                           Q(7), QN => n8);
   Q_reg_6_inst : DFFR_X1 port map( D => D(6), CK => net3376, RN => n13, Q => 
                           Q(6), QN => n7);
   Q_reg_4_inst : DFFR_X1 port map( D => D(4), CK => net3376, RN => n13, Q => 
                           Q(4), QN => n5);
   Q_reg_3_inst : DFFR_X1 port map( D => D(3), CK => net3376, RN => n13, Q => 
                           Q(3), QN => n4);
   Q_reg_2_inst : DFFR_X1 port map( D => D(2), CK => net3376, RN => n13, Q => 
                           Q(2), QN => n3);
   Q_reg_1_inst : DFFR_X1 port map( D => D(1), CK => net3376, RN => n13, Q => 
                           Q(1), QN => n2);
   Q_reg_0_inst : DFFR_X1 port map( D => D(0), CK => net3376, RN => n13, Q => 
                           Q(0), QN => n1);
   clk_gate_Q_reg : SNPS_CLOCK_GATE_HIGH_ff32_en_SIZE13 port map( CLK => clk, 
                           EN => en, ENCLK => net3376);
   Q_reg_9_inst : DFFR_X2 port map( D => D(9), CK => net3376, RN => n13, Q => 
                           Q(9), QN => n10);
   Q_reg_5_inst : DFFR_X2 port map( D => D(5), CK => net3376, RN => n13, Q => 
                           Q(5), QN => n6);
   U2 : INV_X1 port map( A => rst, ZN => n13);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity ff32_en_SIZE5_0 is

   port( D : in std_logic_vector (4 downto 0);  en, clk, rst : in std_logic;  Q
         : out std_logic_vector (4 downto 0));

end ff32_en_SIZE5_0;

architecture SYN_behavioral of ff32_en_SIZE5_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_ff32_en_SIZE5_0
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal net3361, n1, n2, n3, n4, n6, n5 : std_logic;

begin
   
   Q_reg_4_inst : DFFR_X1 port map( D => D(4), CK => net3361, RN => n5, Q => 
                           Q(4), QN => n6);
   Q_reg_3_inst : DFFR_X1 port map( D => D(3), CK => net3361, RN => n5, Q => 
                           Q(3), QN => n4);
   Q_reg_2_inst : DFFR_X1 port map( D => D(2), CK => net3361, RN => n5, Q => 
                           Q(2), QN => n3);
   Q_reg_1_inst : DFFR_X1 port map( D => D(1), CK => net3361, RN => n5, Q => 
                           Q(1), QN => n2);
   Q_reg_0_inst : DFFR_X1 port map( D => D(0), CK => net3361, RN => n5, Q => 
                           Q(0), QN => n1);
   clk_gate_Q_reg : SNPS_CLOCK_GATE_HIGH_ff32_en_SIZE5_0 port map( CLK => clk, 
                           EN => en, ENCLK => net3361);
   U2 : INV_X1 port map( A => rst, ZN => n5);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity ff32_en_SIZE32_0 is

   port( D : in std_logic_vector (31 downto 0);  en, clk, rst : in std_logic;  
         Q : out std_logic_vector (31 downto 0));

end ff32_en_SIZE32_0;

architecture SYN_behavioral of ff32_en_SIZE32_0 is

   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_ff32_en_SIZE32_0
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal net3346, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
      n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29
      , n30, n31, n33, n32 : std_logic;

begin
   
   Q_reg_31_inst : DFFR_X1 port map( D => D(31), CK => net3346, RN => n32, Q =>
                           Q(31), QN => n33);
   Q_reg_30_inst : DFFR_X1 port map( D => D(30), CK => net3346, RN => n32, Q =>
                           Q(30), QN => n31);
   Q_reg_29_inst : DFFR_X1 port map( D => D(29), CK => net3346, RN => n32, Q =>
                           Q(29), QN => n30);
   Q_reg_28_inst : DFFR_X1 port map( D => D(28), CK => net3346, RN => n32, Q =>
                           Q(28), QN => n29);
   Q_reg_27_inst : DFFR_X1 port map( D => D(27), CK => net3346, RN => n32, Q =>
                           Q(27), QN => n28);
   Q_reg_26_inst : DFFR_X1 port map( D => D(26), CK => net3346, RN => n32, Q =>
                           Q(26), QN => n27);
   Q_reg_25_inst : DFFR_X1 port map( D => D(25), CK => net3346, RN => n32, Q =>
                           Q(25), QN => n26);
   Q_reg_24_inst : DFFR_X1 port map( D => D(24), CK => net3346, RN => n32, Q =>
                           Q(24), QN => n25);
   Q_reg_23_inst : DFFR_X1 port map( D => D(23), CK => net3346, RN => n32, Q =>
                           Q(23), QN => n24);
   Q_reg_22_inst : DFFR_X1 port map( D => D(22), CK => net3346, RN => n32, Q =>
                           Q(22), QN => n23);
   Q_reg_21_inst : DFFR_X1 port map( D => D(21), CK => net3346, RN => n32, Q =>
                           Q(21), QN => n22);
   Q_reg_20_inst : DFFR_X1 port map( D => D(20), CK => net3346, RN => n32, Q =>
                           Q(20), QN => n21);
   Q_reg_19_inst : DFFR_X1 port map( D => D(19), CK => net3346, RN => n32, Q =>
                           Q(19), QN => n20);
   Q_reg_18_inst : DFFR_X1 port map( D => D(18), CK => net3346, RN => n32, Q =>
                           Q(18), QN => n19);
   Q_reg_17_inst : DFFR_X1 port map( D => D(17), CK => net3346, RN => n32, Q =>
                           Q(17), QN => n18);
   Q_reg_16_inst : DFFR_X1 port map( D => D(16), CK => net3346, RN => n32, Q =>
                           Q(16), QN => n17);
   Q_reg_15_inst : DFFR_X1 port map( D => D(15), CK => net3346, RN => n32, Q =>
                           Q(15), QN => n16);
   Q_reg_14_inst : DFFR_X1 port map( D => D(14), CK => net3346, RN => n32, Q =>
                           Q(14), QN => n15);
   Q_reg_13_inst : DFFR_X1 port map( D => D(13), CK => net3346, RN => n32, Q =>
                           Q(13), QN => n14);
   Q_reg_12_inst : DFFR_X1 port map( D => D(12), CK => net3346, RN => n32, Q =>
                           Q(12), QN => n13);
   Q_reg_11_inst : DFFR_X1 port map( D => D(11), CK => net3346, RN => n32, Q =>
                           Q(11), QN => n12);
   Q_reg_10_inst : DFFR_X1 port map( D => D(10), CK => net3346, RN => n32, Q =>
                           Q(10), QN => n11);
   Q_reg_9_inst : DFFR_X1 port map( D => D(9), CK => net3346, RN => n32, Q => 
                           Q(9), QN => n10);
   Q_reg_8_inst : DFFR_X1 port map( D => D(8), CK => net3346, RN => n32, Q => 
                           Q(8), QN => n9);
   Q_reg_7_inst : DFFR_X1 port map( D => D(7), CK => net3346, RN => n32, Q => 
                           Q(7), QN => n8);
   Q_reg_6_inst : DFFR_X1 port map( D => D(6), CK => net3346, RN => n32, Q => 
                           Q(6), QN => n7);
   Q_reg_5_inst : DFFR_X1 port map( D => D(5), CK => net3346, RN => n32, Q => 
                           Q(5), QN => n6);
   Q_reg_4_inst : DFFR_X1 port map( D => D(4), CK => net3346, RN => n32, Q => 
                           Q(4), QN => n5);
   Q_reg_3_inst : DFFR_X1 port map( D => D(3), CK => net3346, RN => n32, Q => 
                           Q(3), QN => n4);
   Q_reg_2_inst : DFFR_X1 port map( D => D(2), CK => net3346, RN => n32, Q => 
                           Q(2), QN => n3);
   Q_reg_1_inst : DFFR_X1 port map( D => D(1), CK => net3346, RN => n32, Q => 
                           Q(1), QN => n2);
   Q_reg_0_inst : DFFR_X1 port map( D => D(0), CK => net3346, RN => n32, Q => 
                           Q(0), QN => n1);
   clk_gate_Q_reg : SNPS_CLOCK_GATE_HIGH_ff32_en_SIZE32_0 port map( CLK => clk,
                           EN => en, ENCLK => net3346);
   U2 : INV_X2 port map( A => rst, ZN => n32);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_dlx_regfile_0 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_dlx_regfile_0;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_dlx_regfile_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net3385 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net3385);
   main_gate : AND2_X1 port map( A1 => net3385, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity 
   SNPS_CLOCK_GATE_HIGH_dlx_cu_MICROCODE_MEM_SIZE64_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE13_0 
   is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end 
   SNPS_CLOCK_GATE_HIGH_dlx_cu_MICROCODE_MEM_SIZE64_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE13_0;

architecture SYN_USE_DEFA_ARCH_NAME of 
   SNPS_CLOCK_GATE_HIGH_dlx_cu_MICROCODE_MEM_SIZE64_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE13_0 
   is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net3565 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net3565);
   main_gate : AND2_X1 port map( A1 => net3565, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity alu_ctrl is

   port( OP : in std_logic_vector (0 to 4);  ALU_WORD : out std_logic_vector 
         (12 downto 0));

end alu_ctrl;

architecture SYN_bhe of alu_ctrl is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal ALU_WORD_12_port, ALU_WORD_11_port, ALU_WORD_10_port, ALU_WORD_9_port
      , ALU_WORD_8_port, ALU_WORD_7_port, ALU_WORD_6_port, ALU_WORD_5_port, 
      ALU_WORD_4_port, ALU_WORD_3_port, ALU_WORD_2_port, ALU_WORD_1_port, 
      ALU_WORD_0_port, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, 
      N31, N32, N33, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, 
      n14, n15, n16, n17, n18, n19, n20_port, n21_port, n22_port, n23_port, 
      n24_port, n25_port, n26_port, n27_port, n28_port, n29_port, n30_port, 
      n31_port, n32_port, n33_port, n34, n35 : std_logic;

begin
   ALU_WORD <= ( ALU_WORD_12_port, ALU_WORD_11_port, ALU_WORD_10_port, 
      ALU_WORD_9_port, ALU_WORD_8_port, ALU_WORD_7_port, ALU_WORD_6_port, 
      ALU_WORD_5_port, ALU_WORD_4_port, ALU_WORD_3_port, ALU_WORD_2_port, 
      ALU_WORD_1_port, ALU_WORD_0_port );
   
   comp_sel_reg_2_inst : DLH_X1 port map( G => N32, D => N33, Q => 
                           ALU_WORD_4_port);
   comp_sel_reg_1_inst : DLH_X1 port map( G => N32, D => N31, Q => 
                           ALU_WORD_3_port);
   comp_sel_reg_0_inst : DLH_X1 port map( G => N32, D => N30, Q => 
                           ALU_WORD_2_port);
   sign_to_booth_reg : DLH_X1 port map( G => N20, D => N21, Q => 
                           ALU_WORD_0_port);
   left_right_reg : DLH_X1 port map( G => N23, D => N22, Q => ALU_WORD_9_port);
   logic_arith_reg : DLH_X1 port map( G => N23, D => N24, Q => ALU_WORD_8_port)
                           ;
   sign_to_adder_reg : DLH_X1 port map( G => N25, D => N26, Q => 
                           ALU_WORD_7_port);
   lu_ctrl_reg_1_inst : DLH_X1 port map( G => N28, D => N29, Q => 
                           ALU_WORD_6_port);
   lu_ctrl_reg_0_inst : DLH_X1 port map( G => N28, D => N27, Q => 
                           ALU_WORD_5_port);
   U53 : NAND3_X1 port map( A1 => n9, A2 => OP(3), A3 => n28_port, ZN => 
                           n30_port);
   U54 : NAND3_X1 port map( A1 => n15, A2 => n35, A3 => n22_port, ZN => n19);
   U48 : NOR3_X1 port map( A1 => OP(2), A2 => OP(4), A3 => n22_port, ZN => n10)
                           ;
   U47 : NAND2_X1 port map( A1 => OP(1), A2 => n23_port, ZN => n3);
   U45 : NOR3_X1 port map( A1 => OP(2), A2 => n35, A3 => n22_port, ZN => 
                           n33_port);
   U43 : NOR2_X1 port map( A1 => n3, A2 => n2, ZN => n32_port);
   U41 : NOR2_X1 port map( A1 => OP(4), A2 => n15, ZN => n28_port);
   U40 : NAND2_X1 port map( A1 => n28_port, A2 => n22_port, ZN => n1);
   U39 : NOR2_X1 port map( A1 => n19, A2 => OP(1), ZN => n34);
   U38 : NOR4_X1 port map( A1 => n15, A2 => n3, A3 => n35, A4 => n22_port, ZN 
                           => n8);
   U37 : AOI21_X1 port map( B1 => n34, B2 => OP(0), A => n8, ZN => n18);
   U36 : NAND2_X1 port map( A1 => n33_port, A2 => n26_port, ZN => n6);
   U35 : OAI211_X1 port map( C1 => n1, C2 => n16, A => n18, B => n6, ZN => N30)
                           ;
   U34 : AOI211_X1 port map( C1 => n26_port, C2 => n10, A => n32_port, B => N30
                           , ZN => n29_port);
   U33 : NAND2_X1 port map( A1 => OP(4), A2 => n22_port, ZN => n27_port);
   U32 : NOR2_X1 port map( A1 => n3, A2 => n27_port, ZN => n31_port);
   U31 : NAND2_X1 port map( A1 => OP(2), A2 => n31_port, ZN => n4);
   U29 : NOR2_X1 port map( A1 => OP(2), A2 => n27_port, ZN => n24_port);
   U28 : NAND2_X1 port map( A1 => n26_port, A2 => n24_port, ZN => n7);
   U27 : NAND4_X1 port map( A1 => n29_port, A2 => n4, A3 => n30_port, A4 => n7,
                           ZN => N32);
   U26 : AOI211_X1 port map( C1 => OP(4), C2 => OP(3), A => OP(2), B => n3, ZN 
                           => N28);
   U25 : NAND2_X1 port map( A1 => OP(3), A2 => n28_port, ZN => n17);
   U24 : OAI21_X1 port map( B1 => n27_port, B2 => n15, A => n17, ZN => n25_port
                           );
   U23 : NAND2_X1 port map( A1 => n25_port, A2 => n26_port, ZN => n20_port);
   U18 : NOR3_X1 port map( A1 => OP(2), A2 => n22_port, A3 => n13, ZN => N22);
   U16 : OAI21_X1 port map( B1 => n11, B2 => n13, A => n21_port, ZN => N23);
   U14 : OAI21_X1 port map( B1 => n19, B2 => n13, A => n20_port, ZN => 
                           ALU_WORD_12_port);
   U6 : NOR2_X1 port map( A1 => n3, A2 => n11, ZN => N27);
   U8 : NAND2_X1 port map( A1 => OP(2), A2 => OP(3), ZN => n12);
   U7 : OAI21_X1 port map( B1 => n12, B2 => n13, A => n14, ZN => N26);
   U11 : NOR2_X1 port map( A1 => n2, A2 => n13, ZN => N24);
   U12 : OAI211_X1 port map( C1 => n16, C2 => n17, A => n18, B => n4, ZN => N21
                           );
   U3 : NAND4_X1 port map( A1 => n4, A2 => n5, A3 => n6, A4 => n7, ZN => N31);
   U2 : AOI21_X1 port map( B1 => n1, B2 => n2, A => n3, ZN => N33);
   U9 : OAI21_X1 port map( B1 => n15, B2 => n13, A => n14, ZN => N25);
   U19 : NAND2_X1 port map( A1 => n23_port, A2 => n16, ZN => n13);
   U50 : NOR2_X1 port map( A1 => n23_port, A2 => n16, ZN => n26_port);
   U52 : INV_X1 port map( A => OP(0), ZN => n23_port);
   U51 : INV_X1 port map( A => OP(1), ZN => n16);
   U49 : INV_X1 port map( A => OP(3), ZN => n22_port);
   U46 : INV_X1 port map( A => OP(4), ZN => n35);
   U44 : INV_X1 port map( A => n33_port, ZN => n2);
   U42 : INV_X1 port map( A => OP(2), ZN => n15);
   U30 : INV_X1 port map( A => n3, ZN => n9);
   U22 : INV_X1 port map( A => n20_port, ZN => ALU_WORD_1_port);
   U21 : OR3_X1 port map( A1 => N32, A2 => N28, A3 => ALU_WORD_1_port, ZN => 
                           ALU_WORD_10_port);
   U20 : INV_X1 port map( A => n24_port, ZN => n11);
   U17 : INV_X1 port map( A => N22, ZN => n21_port);
   U15 : OR2_X1 port map( A1 => N32, A2 => N23, ZN => ALU_WORD_11_port);
   U5 : AND2_X1 port map( A1 => n9, A2 => n10, ZN => N29);
   U10 : INV_X1 port map( A => N32, ZN => n14);
   U4 : INV_X1 port map( A => n8, ZN => n5);
   U13 : OR2_X1 port map( A1 => N32, A2 => ALU_WORD_12_port, ZN => N20);

end SYN_bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity cw_mem_MICROCODE_MEM_SIZE64_OP_CODE_SIZE6_CW_SIZE13 is

   port( OPCODE_IN : in std_logic_vector (5 downto 0);  CW_OUT : out 
         std_logic_vector (12 downto 0));

end cw_mem_MICROCODE_MEM_SIZE64_OP_CODE_SIZE6_CW_SIZE13;

architecture SYN_bhe of cw_mem_MICROCODE_MEM_SIZE64_OP_CODE_SIZE6_CW_SIZE13 is

   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal CW_OUT_12_port, CW_OUT_11_port, CW_OUT_10_port, CW_OUT_9_port, 
      CW_OUT_8_port, CW_OUT_7_port, CW_OUT_5_port, CW_OUT_4, CW_OUT_3, CW_OUT_2
      , CW_OUT_1, CW_OUT_0, n7, n8, n9, n10, n11, n12, n13, n14, n17, n18, n19,
      n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n16, n15, n1, n2, n3, 
      n4, n5, n6 : std_logic;

begin
   CW_OUT <= ( CW_OUT_12_port, CW_OUT_11_port, CW_OUT_10_port, CW_OUT_9_port, 
      CW_OUT_8_port, CW_OUT_7_port, CW_OUT_5_port, CW_OUT_5_port, CW_OUT_4, 
      CW_OUT_3, CW_OUT_2, CW_OUT_1, CW_OUT_0 );
   
   U35 : NAND3_X1 port map( A1 => OPCODE_IN(3), A2 => n23, A3 => n24, ZN => n22
                           );
   U36 : NAND3_X1 port map( A1 => OPCODE_IN(4), A2 => n14, A3 => n25, ZN => n29
                           );
   U34 : NAND3_X1 port map( A1 => OPCODE_IN(3), A2 => n13, A3 => n14, ZN => n15
                           );
   U8 : NOR2_X1 port map( A1 => n10, A2 => n17, ZN => CW_OUT_8_port);
   U23 : OAI21_X1 port map( B1 => OPCODE_IN(3), B2 => n17, A => n29, ZN => 
                           CW_OUT_11_port);
   U4 : OAI22_X1 port map( A1 => OPCODE_IN(3), A2 => n11, B1 => n12, B2 => n10,
                           ZN => CW_OUT_4);
   U19 : NOR2_X1 port map( A1 => n7, A2 => n8, ZN => CW_OUT_3);
   U16 : NAND2_X1 port map( A1 => OPCODE_IN(3), A2 => OPCODE_IN(4), ZN => n20);
   U15 : NAND2_X1 port map( A1 => n23, A2 => n7, ZN => n27);
   U1 : NOR3_X1 port map( A1 => n2, A2 => n7, A3 => n8, ZN => CW_OUT_2);
   U3 : NOR2_X1 port map( A1 => n8, A2 => n10, ZN => CW_OUT_1);
   U21 : INV_X1 port map( A => OPCODE_IN(0), ZN => n7);
   U18 : NAND2_X1 port map( A1 => OPCODE_IN(0), A2 => n2, ZN => n10);
   U30 : INV_X1 port map( A => OPCODE_IN(5), ZN => n23);
   U10 : OR2_X1 port map( A1 => CW_OUT_7_port, A2 => n18, ZN => n9);
   U9 : OR2_X1 port map( A1 => CW_OUT_3, A2 => n9, ZN => CW_OUT_5_port);
   U2 : OR3_X1 port map( A1 => n9, A2 => CW_OUT_4, A3 => CW_OUT_1, ZN => 
                           CW_OUT_0);
   U5 : NOR3_X1 port map( A1 => OPCODE_IN(5), A2 => n19, A3 => n10, ZN => 
                           CW_OUT_7_port);
   U6 : INV_X1 port map( A => OPCODE_IN(3), ZN => n2);
   U7 : INV_X1 port map( A => OPCODE_IN(2), ZN => n14);
   U11 : CLKBUF_X1 port map( A => n28, Z => n5);
   U12 : INV_X1 port map( A => n16, ZN => CW_OUT_12_port);
   U13 : AND3_X1 port map( A1 => n23, A2 => n2, A3 => n6, ZN => n25);
   U14 : CLKBUF_X1 port map( A => OPCODE_IN(1), Z => n6);
   U17 : OR2_X1 port map( A1 => OPCODE_IN(0), A2 => n15, ZN => n4);
   U20 : NAND2_X1 port map( A1 => n28, A2 => n23, ZN => n12);
   U22 : NOR2_X1 port map( A1 => n19, A2 => OPCODE_IN(4), ZN => n28);
   U24 : NAND2_X1 port map( A1 => n14, A2 => OPCODE_IN(1), ZN => n19);
   U25 : OR2_X1 port map( A1 => OPCODE_IN(0), A2 => n12, ZN => n3);
   U26 : NOR3_X1 port map( A1 => OPCODE_IN(5), A2 => OPCODE_IN(1), A3 => 
                           OPCODE_IN(4), ZN => n13);
   U27 : NAND2_X1 port map( A1 => n12, A2 => n17, ZN => n1);
   U28 : NAND2_X1 port map( A1 => n1, A2 => n2, ZN => n16);
   U29 : NAND3_X1 port map( A1 => n16, A2 => n3, A3 => n4, ZN => CW_OUT_9_port)
                           ;
   U31 : NOR2_X1 port map( A1 => n12, A2 => OPCODE_IN(3), ZN => CW_OUT_10_port)
                           ;
   U32 : NAND2_X1 port map( A1 => n13, A2 => n14, ZN => n11);
   U33 : OAI211_X1 port map( C1 => n25, C2 => n26, A => OPCODE_IN(2), B => 
                           OPCODE_IN(4), ZN => n21);
   U37 : NAND2_X1 port map( A1 => OPCODE_IN(2), A2 => n13, ZN => n17);
   U38 : NAND2_X1 port map( A1 => OPCODE_IN(5), A2 => n5, ZN => n8);
   U39 : OAI211_X1 port map( C1 => n19, C2 => n20, A => n21, B => n22, ZN => 
                           n18);
   U40 : AOI21_X1 port map( B1 => n2, B2 => n27, A => n6, ZN => n26);
   U41 : OAI211_X1 port map( C1 => OPCODE_IN(4), C2 => OPCODE_IN(0), A => n6, B
                           => OPCODE_IN(2), ZN => n24);

end SYN_bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity stall_logic_FUNC_SIZE11_OP_CODE_SIZE6 is

   port( OPCODE_i : in std_logic_vector (5 downto 0);  FUNC_i : in 
         std_logic_vector (10 downto 0);  rA_i, rB_i, D1_i, D2_i : in 
         std_logic_vector (4 downto 0);  S_mem_LOAD_i, S_exe_LOAD_i, 
         S_exe_WRITE_i : in std_logic;  S_MUX_PC_BUS_i : in std_logic_vector (1
         downto 0);  mispredict_i : in std_logic;  bubble_dec_o, bubble_exe_o, 
         stall_exe_o, stall_dec_o, stall_btb_o, stall_fetch_o : out std_logic);

end stall_logic_FUNC_SIZE11_OP_CODE_SIZE6;

architecture SYN_stall_logic_hw of stall_logic_FUNC_SIZE11_OP_CODE_SIZE6 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI33_X1
      port( A1, A2, A3, B1, B2, B3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal stall_fetch_o_port, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
      n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40
      , n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, 
      n55, n56, n57, n58 : std_logic;

begin
   stall_dec_o <= stall_fetch_o_port;
   stall_btb_o <= stall_fetch_o_port;
   stall_fetch_o <= stall_fetch_o_port;
   
   U46 : OAI33_X1 port map( A1 => OPCODE_i(2), A2 => n52, A3 => n53, B1 => n50,
                           B2 => OPCODE_i(4), B3 => OPCODE_i(1), ZN => n51);
   U36 : NAND4_X1 port map( A1 => S_mem_LOAD_i, A2 => n54, A3 => n55, A4 => n56
                           , ZN => n17);
   U35 : NOR2_X1 port map( A1 => OPCODE_i(5), A2 => OPCODE_i(3), ZN => n27);
   U31 : NAND2_X1 port map( A1 => n27, A2 => n51, ZN => n18);
   U30 : OAI21_X1 port map( B1 => OPCODE_i(0), B2 => n50, A => OPCODE_i(4), ZN 
                           => n48);
   U26 : AOI21_X1 port map( B1 => n27, B2 => n46, A => n47, ZN => n34);
   U23 : XNOR2_X1 port map( A => n31, B => rA_i(4), ZN => n37);
   U22 : AOI22_X1 port map( A1 => n43, A2 => D1_i(3), B1 => D1_i(2), B2 => n44,
                           ZN => n45);
   U21 : OAI221_X1 port map( B1 => n43, B2 => D1_i(3), C1 => n44, C2 => D1_i(2)
                           , A => n45, ZN => n38);
   U20 : AOI22_X1 port map( A1 => n40, A2 => D1_i(1), B1 => D1_i(0), B2 => n41,
                           ZN => n42);
   U19 : OAI221_X1 port map( B1 => n40, B2 => D1_i(1), C1 => n41, C2 => D1_i(0)
                           , A => n42, ZN => n39);
   U18 : NOR3_X1 port map( A1 => n37, A2 => n38, A3 => n39, ZN => n36);
   U17 : OAI221_X1 port map( B1 => n34, B2 => n35, C1 => n34, C2 => 
                           S_exe_WRITE_i, A => n36, ZN => n19);
   U15 : OAI22_X1 port map( A1 => n31, A2 => rB_i(4), B1 => n32, B2 => rB_i(2),
                           ZN => n33);
   U14 : AOI221_X1 port map( B1 => n31, B2 => rB_i(4), C1 => rB_i(2), C2 => n32
                           , A => n33, ZN => n21);
   U11 : OAI22_X1 port map( A1 => n28, A2 => rB_i(0), B1 => n29, B2 => rB_i(3),
                           ZN => n30);
   U10 : AOI221_X1 port map( B1 => n28, B2 => rB_i(0), C1 => rB_i(3), C2 => n29
                           , A => n30, ZN => n22);
   U7 : OAI211_X1 port map( C1 => n25, C2 => rB_i(1), A => S_exe_LOAD_i, B => 
                           n27, ZN => n26);
   U6 : AOI21_X1 port map( B1 => n25, B2 => rB_i(1), A => n26, ZN => n24);
   U5 : NAND4_X1 port map( A1 => n21, A2 => n22, A3 => n23, A4 => n24, ZN => 
                           n20);
   U2 : NOR2_X1 port map( A1 => stall_fetch_o_port, A2 => n16, ZN => 
                           bubble_dec_o);
   U45 : INV_X1 port map( A => rA_i(3), ZN => n43);
   U44 : INV_X1 port map( A => rA_i(1), ZN => n40);
   U41 : INV_X1 port map( A => rA_i(0), ZN => n41);
   U40 : INV_X1 port map( A => rA_i(2), ZN => n44);
   U34 : INV_X1 port map( A => OPCODE_i(4), ZN => n52);
   U27 : INV_X1 port map( A => S_exe_LOAD_i, ZN => n47);
   U25 : INV_X1 port map( A => n18, ZN => n35);
   U24 : INV_X1 port map( A => D1_i(4), ZN => n31);
   U16 : INV_X1 port map( A => D1_i(2), ZN => n32);
   U13 : INV_X1 port map( A => D1_i(0), ZN => n28);
   U12 : INV_X1 port map( A => D1_i(3), ZN => n29);
   U8 : INV_X1 port map( A => D1_i(1), ZN => n25);
   U4 : OAI211_X1 port map( C1 => n17, C2 => n18, A => n19, B => n20, ZN => 
                           stall_fetch_o_port);
   U3 : AOI221_X1 port map( B1 => n41, B2 => D2_i(0), C1 => D2_i(2), C2 => n44,
                           A => n57, ZN => n55);
   U9 : INV_X1 port map( A => mispredict_i, ZN => n16);
   U28 : INV_X1 port map( A => OPCODE_i(2), ZN => n50);
   U29 : AOI221_X1 port map( B1 => n43, B2 => D2_i(3), C1 => D2_i(1), C2 => n40
                           , A => n58, ZN => n54);
   U32 : XNOR2_X1 port map( A => rA_i(4), B => D2_i(4), ZN => n56);
   U33 : OAI22_X1 port map( A1 => n41, A2 => D2_i(0), B1 => n44, B2 => D2_i(2),
                           ZN => n57);
   U37 : OAI22_X1 port map( A1 => n43, A2 => D2_i(3), B1 => n40, B2 => D2_i(1),
                           ZN => n58);
   U38 : NOR4_X1 port map( A1 => OPCODE_i(2), A2 => OPCODE_i(4), A3 => 
                           OPCODE_i(1), A4 => OPCODE_i(0), ZN => n23);
   U39 : OAI22_X1 port map( A1 => OPCODE_i(1), A2 => n48, B1 => OPCODE_i(4), B2
                           => n49, ZN => n46);
   U42 : NAND2_X1 port map( A1 => OPCODE_i(1), A2 => n50, ZN => n49);
   U43 : INV_X1 port map( A => OPCODE_i(1), ZN => n53);

end SYN_stall_logic_hw;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity mux41_MUX_SIZE32_0 is

   port( IN0, IN1, IN2, IN3 : in std_logic_vector (31 downto 0);  CTRL : in 
         std_logic_vector (1 downto 0);  OUT1 : out std_logic_vector (31 downto
         0));

end mux41_MUX_SIZE32_0;

architecture SYN_bhe of mux41_MUX_SIZE32_0 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n6, n7, n8, n15, n16, n23, n24, n31, n32, n33, n34, n39, n40,
      n41, n42, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n63
      , n64, n65, n66, n67, n68, n71, n1, n2, n5, n9, n10, n11, n12, n13, n14, 
      n17, n18, n19, n20, n21, n22, n25, n26, n27, n28, n29, n30, n35, n36, n37
      , n38, n43, n44, n45, n46, n59, n60, n61, n62, n69, n70, n72, n73, n74, 
      n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89
      , n90, n91, n92, n93, n94 : std_logic;

begin
   
   U61 : NAND2_X1 port map( A1 => n47, A2 => n48, ZN => OUT1(1));
   U64 : NAND2_X1 port map( A1 => n49, A2 => n50, ZN => OUT1(19));
   U51 : AOI22_X1 port map( A1 => n89, A2 => IN1(23), B1 => n88, B2 => IN0(23),
                           ZN => n39);
   U49 : NAND2_X1 port map( A1 => n39, A2 => n40, ZN => OUT1(23));
   U54 : AOI22_X1 port map( A1 => n91, A2 => IN1(22), B1 => n86, B2 => IN0(22),
                           ZN => n41);
   U85 : NAND2_X1 port map( A1 => n63, A2 => n64, ZN => OUT1(12));
   U88 : NAND2_X1 port map( A1 => n65, A2 => n66, ZN => OUT1(11));
   U73 : NAND2_X1 port map( A1 => n55, A2 => n56, ZN => OUT1(16));
   U76 : NAND2_X1 port map( A1 => n57, A2 => n58, ZN => OUT1(15));
   U39 : AOI22_X1 port map( A1 => n91, A2 => IN1(27), B1 => n88, B2 => IN0(27),
                           ZN => n31);
   U42 : AOI22_X1 port map( A1 => n91, A2 => IN1(26), B1 => n86, B2 => IN0(26),
                           ZN => n33);
   U3 : AOI22_X1 port map( A1 => n89, A2 => IN1(9), B1 => n87, B2 => IN0(9), ZN
                           => n3);
   U1 : NAND2_X1 port map( A1 => n3, A2 => n4, ZN => OUT1(9));
   U15 : AOI22_X1 port map( A1 => n90, A2 => IN1(5), B1 => n88, B2 => IN0(5), 
                           ZN => n15);
   U13 : NAND2_X1 port map( A1 => n15, A2 => n16, ZN => OUT1(5));
   U27 : AOI22_X1 port map( A1 => n91, A2 => IN1(30), B1 => n87, B2 => IN0(30),
                           ZN => n23);
   U2 : BUF_X2 port map( A => n8, Z => n87);
   U4 : BUF_X1 port map( A => n6, Z => n94);
   U5 : AND2_X1 port map( A1 => n71, A2 => CTRL(0), ZN => n7);
   U6 : BUF_X1 port map( A => CTRL(1), Z => n85);
   U7 : BUF_X2 port map( A => n7, Z => n91);
   U8 : BUF_X2 port map( A => n6, Z => n92);
   U9 : BUF_X2 port map( A => n6, Z => n93);
   U10 : BUF_X2 port map( A => n7, Z => n90);
   U11 : BUF_X2 port map( A => n7, Z => n89);
   U12 : BUF_X2 port map( A => n8, Z => n86);
   U14 : BUF_X2 port map( A => n8, Z => n88);
   U16 : NOR2_X1 port map( A1 => n71, A2 => CTRL(0), ZN => n6);
   U17 : NOR2_X1 port map( A1 => CTRL(0), A2 => n85, ZN => n8);
   U18 : INV_X1 port map( A => CTRL(1), ZN => n71);
   U19 : NAND2_X1 port map( A1 => n94, A2 => IN2(30), ZN => n24);
   U20 : NAND2_X1 port map( A1 => n93, A2 => IN2(5), ZN => n16);
   U21 : NAND2_X1 port map( A1 => n93, A2 => IN2(9), ZN => n4);
   U22 : NAND2_X1 port map( A1 => n94, A2 => IN2(26), ZN => n34);
   U23 : NAND2_X1 port map( A1 => n94, A2 => IN2(27), ZN => n32);
   U24 : NAND2_X1 port map( A1 => n93, A2 => IN2(15), ZN => n58);
   U25 : NAND2_X1 port map( A1 => n93, A2 => IN2(16), ZN => n56);
   U26 : NAND2_X1 port map( A1 => n92, A2 => IN2(11), ZN => n66);
   U28 : NAND2_X1 port map( A1 => n92, A2 => IN2(12), ZN => n64);
   U29 : NAND2_X1 port map( A1 => n92, A2 => IN2(22), ZN => n42);
   U30 : NAND2_X1 port map( A1 => n92, A2 => IN2(23), ZN => n40);
   U31 : NAND2_X1 port map( A1 => n92, A2 => IN2(19), ZN => n50);
   U32 : NAND2_X1 port map( A1 => n92, A2 => IN2(1), ZN => n48);
   U33 : NAND3_X1 port map( A1 => n2, A2 => n1, A3 => n5, ZN => OUT1(0));
   U34 : NAND2_X1 port map( A1 => n90, A2 => IN1(0), ZN => n2);
   U35 : NAND2_X1 port map( A1 => n88, A2 => IN0(0), ZN => n5);
   U36 : NAND2_X1 port map( A1 => n93, A2 => IN2(0), ZN => n1);
   U37 : NAND3_X1 port map( A1 => n11, A2 => n9, A3 => n10, ZN => OUT1(2));
   U38 : NAND2_X1 port map( A1 => n88, A2 => IN0(2), ZN => n9);
   U40 : NAND2_X1 port map( A1 => n91, A2 => IN1(2), ZN => n11);
   U41 : NAND2_X1 port map( A1 => n94, A2 => IN2(2), ZN => n10);
   U43 : NAND3_X1 port map( A1 => n13, A2 => n12, A3 => n14, ZN => OUT1(8));
   U44 : NAND2_X1 port map( A1 => n90, A2 => IN1(8), ZN => n13);
   U45 : NAND2_X1 port map( A1 => n88, A2 => IN0(8), ZN => n14);
   U46 : NAND2_X1 port map( A1 => n93, A2 => IN2(8), ZN => n12);
   U47 : NAND3_X1 port map( A1 => n18, A2 => n17, A3 => n19, ZN => OUT1(14));
   U48 : NAND2_X1 port map( A1 => n91, A2 => IN1(14), ZN => n18);
   U50 : NAND2_X1 port map( A1 => n88, A2 => IN0(14), ZN => n19);
   U52 : NAND2_X1 port map( A1 => n93, A2 => IN2(14), ZN => n17);
   U53 : NAND3_X1 port map( A1 => n21, A2 => n20, A3 => n22, ZN => OUT1(13));
   U55 : NAND2_X1 port map( A1 => n89, A2 => IN1(13), ZN => n21);
   U56 : NAND2_X1 port map( A1 => n87, A2 => IN0(13), ZN => n22);
   U57 : NAND2_X1 port map( A1 => n93, A2 => IN2(13), ZN => n20);
   U58 : NAND3_X1 port map( A1 => n26, A2 => n25, A3 => n27, ZN => OUT1(25));
   U59 : NAND2_X1 port map( A1 => n94, A2 => IN2(25), ZN => n26);
   U60 : NAND2_X1 port map( A1 => n87, A2 => IN0(25), ZN => n25);
   U62 : NAND2_X1 port map( A1 => n90, A2 => IN1(25), ZN => n27);
   U63 : NAND3_X1 port map( A1 => n29, A2 => n28, A3 => n30, ZN => OUT1(4));
   U65 : NAND2_X1 port map( A1 => n93, A2 => IN2(4), ZN => n29);
   U66 : NAND2_X1 port map( A1 => n89, A2 => IN1(4), ZN => n30);
   U67 : NAND2_X1 port map( A1 => n87, A2 => IN0(4), ZN => n28);
   U68 : NAND3_X1 port map( A1 => n36, A2 => n35, A3 => n37, ZN => OUT1(29));
   U69 : NAND2_X1 port map( A1 => n94, A2 => IN2(29), ZN => n36);
   U70 : NAND2_X1 port map( A1 => n87, A2 => IN0(29), ZN => n35);
   U71 : NAND2_X1 port map( A1 => n90, A2 => IN1(29), ZN => n37);
   U72 : NAND3_X1 port map( A1 => n43, A2 => n38, A3 => n44, ZN => OUT1(24));
   U74 : NAND2_X1 port map( A1 => n94, A2 => IN2(24), ZN => n43);
   U75 : NAND2_X1 port map( A1 => n87, A2 => IN0(24), ZN => n38);
   U77 : NAND2_X1 port map( A1 => n89, A2 => IN1(24), ZN => n44);
   U78 : NAND3_X1 port map( A1 => n46, A2 => n45, A3 => n59, ZN => OUT1(3));
   U79 : NAND2_X1 port map( A1 => n93, A2 => IN2(3), ZN => n46);
   U80 : NAND2_X1 port map( A1 => n90, A2 => IN1(3), ZN => n59);
   U81 : NAND2_X1 port map( A1 => n88, A2 => IN0(3), ZN => n45);
   U82 : NAND3_X1 port map( A1 => n61, A2 => n60, A3 => n62, ZN => OUT1(20));
   U83 : NAND2_X1 port map( A1 => n92, A2 => IN2(20), ZN => n61);
   U84 : NAND2_X1 port map( A1 => n87, A2 => IN0(20), ZN => n60);
   U86 : NAND2_X1 port map( A1 => n89, A2 => IN1(20), ZN => n62);
   U87 : NAND3_X1 port map( A1 => n70, A2 => n69, A3 => n72, ZN => OUT1(28));
   U89 : NAND2_X1 port map( A1 => n94, A2 => IN2(28), ZN => n70);
   U90 : NAND2_X1 port map( A1 => n88, A2 => IN0(28), ZN => n69);
   U91 : NAND2_X1 port map( A1 => n90, A2 => IN1(28), ZN => n72);
   U92 : NAND3_X1 port map( A1 => n74, A2 => n73, A3 => n75, ZN => OUT1(6));
   U93 : NAND2_X1 port map( A1 => n93, A2 => IN2(6), ZN => n74);
   U94 : NAND2_X1 port map( A1 => n91, A2 => IN1(6), ZN => n75);
   U95 : NAND2_X1 port map( A1 => n88, A2 => IN0(6), ZN => n73);
   U96 : NAND3_X1 port map( A1 => n77, A2 => n76, A3 => n78, ZN => OUT1(21));
   U97 : NAND2_X1 port map( A1 => n92, A2 => IN2(21), ZN => n77);
   U98 : NAND2_X1 port map( A1 => n88, A2 => IN0(21), ZN => n76);
   U99 : NAND2_X1 port map( A1 => n89, A2 => IN1(21), ZN => n78);
   U100 : NAND3_X1 port map( A1 => n80, A2 => n79, A3 => n81, ZN => OUT1(31));
   U101 : NAND2_X1 port map( A1 => n92, A2 => IN2(31), ZN => n80);
   U102 : NAND2_X1 port map( A1 => n89, A2 => IN1(31), ZN => n81);
   U103 : NAND2_X1 port map( A1 => n88, A2 => IN0(31), ZN => n79);
   U104 : NAND3_X1 port map( A1 => n83, A2 => n82, A3 => n84, ZN => OUT1(7));
   U105 : NAND2_X1 port map( A1 => n93, A2 => IN2(7), ZN => n83);
   U106 : NAND2_X1 port map( A1 => n91, A2 => IN1(7), ZN => n84);
   U107 : NAND2_X1 port map( A1 => n87, A2 => IN0(7), ZN => n82);
   U108 : AOI22_X1 port map( A1 => n90, A2 => IN1(1), B1 => n87, B2 => IN0(1), 
                           ZN => n47);
   U109 : AOI22_X1 port map( A1 => n89, A2 => IN1(16), B1 => n87, B2 => IN0(16)
                           , ZN => n55);
   U110 : AOI22_X1 port map( A1 => n90, A2 => IN1(12), B1 => n87, B2 => IN0(12)
                           , ZN => n63);
   U111 : AOI22_X1 port map( A1 => n90, A2 => IN1(19), B1 => n86, B2 => IN0(19)
                           , ZN => n49);
   U112 : AOI22_X1 port map( A1 => n91, A2 => IN1(15), B1 => n86, B2 => IN0(15)
                           , ZN => n57);
   U113 : AOI22_X1 port map( A1 => n91, A2 => IN1(18), B1 => n86, B2 => IN0(18)
                           , ZN => n51);
   U114 : AOI22_X1 port map( A1 => n89, A2 => IN1(11), B1 => n86, B2 => IN0(11)
                           , ZN => n65);
   U115 : AOI22_X1 port map( A1 => n90, A2 => IN1(17), B1 => n86, B2 => IN0(17)
                           , ZN => n53);
   U116 : AOI22_X1 port map( A1 => n89, A2 => IN1(10), B1 => n86, B2 => IN0(10)
                           , ZN => n67);
   U117 : NAND2_X1 port map( A1 => n53, A2 => n54, ZN => OUT1(17));
   U118 : NAND2_X1 port map( A1 => n51, A2 => n52, ZN => OUT1(18));
   U119 : NAND2_X1 port map( A1 => n23, A2 => n24, ZN => OUT1(30));
   U120 : NAND2_X1 port map( A1 => n31, A2 => n32, ZN => OUT1(27));
   U121 : NAND2_X1 port map( A1 => n67, A2 => n68, ZN => OUT1(10));
   U122 : NAND2_X1 port map( A1 => n33, A2 => n34, ZN => OUT1(26));
   U123 : NAND2_X1 port map( A1 => n92, A2 => IN2(17), ZN => n54);
   U124 : NAND2_X1 port map( A1 => n92, A2 => IN2(10), ZN => n68);
   U125 : NAND2_X1 port map( A1 => n92, A2 => IN2(18), ZN => n52);
   U126 : NAND2_X1 port map( A1 => n41, A2 => n42, ZN => OUT1(22));

end SYN_bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity zerocheck is

   port( IN0 : in std_logic_vector (31 downto 0);  CTRL : in std_logic;  OUT1 :
         out std_logic);

end zerocheck;

architecture SYN_Bhe of zerocheck is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n9, n8, n7, n6, n5, n4, n3, n2, n12, n11, n10 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n2, B => CTRL, ZN => OUT1);
   U2 : NOR2_X1 port map( A1 => n3, A2 => n4, ZN => n2);
   U3 : NOR4_X1 port map( A1 => IN0(30), A2 => IN0(2), A3 => IN0(29), A4 => 
                           IN0(28), ZN => n8);
   U4 : NOR4_X1 port map( A1 => IN0(5), A2 => IN0(4), A3 => IN0(3), A4 => 
                           IN0(31), ZN => n5);
   U5 : NOR4_X1 port map( A1 => IN0(9), A2 => IN0(8), A3 => IN0(7), A4 => 
                           IN0(6), ZN => n6);
   U6 : NOR4_X1 port map( A1 => IN0(27), A2 => IN0(26), A3 => IN0(25), A4 => 
                           IN0(24), ZN => n7);
   U7 : NOR4_X1 port map( A1 => IN0(16), A2 => IN0(15), A3 => IN0(14), A4 => 
                           IN0(13), ZN => n12);
   U8 : NOR4_X1 port map( A1 => IN0(12), A2 => IN0(11), A3 => IN0(10), A4 => 
                           IN0(0), ZN => n11);
   U9 : NOR4_X1 port map( A1 => IN0(23), A2 => IN0(22), A3 => IN0(21), A4 => 
                           IN0(20), ZN => n10);
   U10 : NOR4_X1 port map( A1 => IN0(1), A2 => IN0(19), A3 => IN0(18), A4 => 
                           IN0(17), ZN => n9);
   U11 : NAND4_X1 port map( A1 => n7, A2 => n6, A3 => n5, A4 => n8, ZN => n4);
   U12 : NAND4_X1 port map( A1 => n9, A2 => n10, A3 => n11, A4 => n12, ZN => n3
                           );

end SYN_Bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity mux21_0 is

   port( IN0, IN1 : in std_logic_vector (31 downto 0);  CTRL : in std_logic;  
         OUT1 : out std_logic_vector (31 downto 0));

end mux21_0;

architecture SYN_Bhe of mux21_0 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : MUX2_X1 port map( A => IN0(9), B => IN1(9), S => n3, Z => OUT1(9));
   U2 : MUX2_X1 port map( A => IN0(8), B => IN1(8), S => n3, Z => OUT1(8));
   U3 : MUX2_X1 port map( A => IN0(7), B => IN1(7), S => n2, Z => OUT1(7));
   U4 : MUX2_X1 port map( A => IN0(6), B => IN1(6), S => n1, Z => OUT1(6));
   U7 : MUX2_X1 port map( A => IN0(3), B => IN1(3), S => n1, Z => OUT1(3));
   U18 : MUX2_X1 port map( A => IN0(22), B => IN1(22), S => n2, Z => OUT1(22));
   U19 : MUX2_X1 port map( A => IN0(21), B => IN1(21), S => n3, Z => OUT1(21));
   U20 : MUX2_X1 port map( A => IN0(20), B => IN1(20), S => n1, Z => OUT1(20));
   U23 : MUX2_X1 port map( A => IN0(18), B => IN1(18), S => n2, Z => OUT1(18));
   U24 : MUX2_X1 port map( A => IN0(17), B => IN1(17), S => n2, Z => OUT1(17));
   U25 : MUX2_X1 port map( A => IN0(16), B => IN1(16), S => n2, Z => OUT1(16));
   U26 : MUX2_X1 port map( A => IN0(15), B => IN1(15), S => n1, Z => OUT1(15));
   U29 : MUX2_X1 port map( A => IN0(12), B => IN1(12), S => n1, Z => OUT1(12));
   U32 : MUX2_X1 port map( A => IN0(0), B => IN1(0), S => n1, Z => OUT1(0));
   U22 : MUX2_X1 port map( A => IN0(19), B => IN1(19), S => n3, Z => OUT1(19));
   U6 : MUX2_X1 port map( A => IN0(4), B => IN1(4), S => n1, Z => OUT1(4));
   U27 : MUX2_X1 port map( A => IN0(14), B => IN1(14), S => n1, Z => OUT1(14));
   U31 : MUX2_X1 port map( A => IN0(10), B => IN1(10), S => n3, Z => OUT1(10));
   U30 : MUX2_X1 port map( A => IN0(11), B => IN1(11), S => n2, Z => OUT1(11));
   U13 : MUX2_X1 port map( A => IN0(27), B => IN1(27), S => n2, Z => OUT1(27));
   U28 : MUX2_X1 port map( A => IN0(13), B => IN1(13), S => n1, Z => OUT1(13));
   U21 : MUX2_X1 port map( A => IN0(1), B => IN1(1), S => n3, Z => OUT1(1));
   U10 : MUX2_X1 port map( A => IN0(2), B => IN1(2), S => n1, Z => OUT1(2));
   U5 : MUX2_X1 port map( A => IN0(5), B => IN1(5), S => n2, Z => OUT1(5));
   U11 : MUX2_X1 port map( A => IN0(29), B => IN1(29), S => n2, Z => OUT1(29));
   U17 : MUX2_X1 port map( A => IN0(23), B => IN1(23), S => n2, Z => OUT1(23));
   U8 : MUX2_X1 port map( A => IN0(31), B => IN1(31), S => n3, Z => OUT1(31));
   U9 : BUF_X2 port map( A => CTRL, Z => n2);
   U12 : MUX2_X1 port map( A => IN0(25), B => IN1(25), S => n3, Z => OUT1(25));
   U14 : MUX2_X1 port map( A => IN0(24), B => IN1(24), S => n3, Z => OUT1(24));
   U15 : MUX2_X1 port map( A => IN0(26), B => IN1(26), S => n2, Z => OUT1(26));
   U16 : CLKBUF_X2 port map( A => CTRL, Z => n3);
   U33 : BUF_X2 port map( A => CTRL, Z => n1);
   U34 : MUX2_X1 port map( A => IN0(28), B => IN1(28), S => n3, Z => OUT1(28));
   U35 : MUX2_X1 port map( A => IN0(30), B => IN1(30), S => n3, Z => OUT1(30));

end SYN_Bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity p4add_N32_logN5_0 is

   port( A, B : in std_logic_vector (31 downto 0);  Cin, sign : in std_logic;  
         S : out std_logic_vector (31 downto 0);  Cout : out std_logic);

end p4add_N32_logN5_0;

architecture SYN_STRUCTURAL of p4add_N32_logN5_0 is

   component sum_gen_N32_0
      port( A, B : in std_logic_vector (31 downto 0);  Cin : in 
            std_logic_vector (8 downto 0);  S : out std_logic_vector (31 downto
            0));
   end component;
   
   component carry_tree_N32_logN5_0
      port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  
            Cout : out std_logic_vector (7 downto 0));
   end component;
   
   component xor_gen_N32_0
      port( A : in std_logic_vector (31 downto 0);  B : in std_logic;  S : out 
            std_logic_vector (31 downto 0));
   end component;
   
   signal n11, new_B_31_port, new_B_30_port, new_B_29_port, new_B_28_port, 
      new_B_27_port, new_B_26_port, new_B_25_port, new_B_24_port, new_B_23_port
      , new_B_22_port, new_B_21_port, new_B_20_port, new_B_19_port, 
      new_B_18_port, new_B_17_port, new_B_16_port, new_B_15_port, new_B_14_port
      , new_B_13_port, new_B_12_port, new_B_11_port, new_B_10_port, 
      new_B_9_port, new_B_8_port, new_B_7_port, new_B_6_port, new_B_5_port, 
      new_B_4_port, new_B_3_port, new_B_2_port, new_B_1_port, new_B_0_port, 
      carry_pro_7_port, carry_pro_6_port, carry_pro_5_port, carry_pro_4_port, 
      carry_pro_3_port, carry_pro_2_port, carry_pro_1_port, n1, n2, n3, n4, n5,
      n6, n7, n8, n9, n10, net48714 : std_logic;

begin
   
   xor32 : xor_gen_N32_0 port map( A(31) => B(31), A(30) => B(30), A(29) => 
                           B(29), A(28) => B(28), A(27) => B(27), A(26) => 
                           B(26), A(25) => B(25), A(24) => B(24), A(23) => 
                           B(23), A(22) => B(22), A(21) => B(21), A(20) => 
                           B(20), A(19) => B(19), A(18) => B(18), A(17) => 
                           B(17), A(16) => B(16), A(15) => B(15), A(14) => 
                           B(14), A(13) => B(13), A(12) => B(12), A(11) => 
                           B(11), A(10) => B(10), A(9) => B(9), A(8) => B(8), 
                           A(7) => B(7), A(6) => B(6), A(5) => B(5), A(4) => 
                           B(4), A(3) => B(3), A(2) => B(2), A(1) => B(1), A(0)
                           => B(0), B => n11, S(31) => new_B_31_port, S(30) => 
                           new_B_30_port, S(29) => new_B_29_port, S(28) => 
                           new_B_28_port, S(27) => new_B_27_port, S(26) => 
                           new_B_26_port, S(25) => new_B_25_port, S(24) => 
                           new_B_24_port, S(23) => new_B_23_port, S(22) => 
                           new_B_22_port, S(21) => new_B_21_port, S(20) => 
                           new_B_20_port, S(19) => new_B_19_port, S(18) => 
                           new_B_18_port, S(17) => new_B_17_port, S(16) => 
                           new_B_16_port, S(15) => new_B_15_port, S(14) => 
                           new_B_14_port, S(13) => new_B_13_port, S(12) => 
                           new_B_12_port, S(11) => new_B_11_port, S(10) => 
                           new_B_10_port, S(9) => new_B_9_port, S(8) => 
                           new_B_8_port, S(7) => new_B_7_port, S(6) => 
                           new_B_6_port, S(5) => new_B_5_port, S(4) => 
                           new_B_4_port, S(3) => new_B_3_port, S(2) => 
                           new_B_2_port, S(1) => new_B_1_port, S(0) => 
                           new_B_0_port);
   ct : carry_tree_N32_logN5_0 port map( A(31) => n2, A(30) => n3, A(29) => n4,
                           A(28) => n5, A(27) => A(27), A(26) => A(26), A(25) 
                           => A(25), A(24) => A(24), A(23) => A(23), A(22) => 
                           A(22), A(21) => A(21), A(20) => A(20), A(19) => 
                           A(19), A(18) => A(18), A(17) => A(17), A(16) => 
                           A(16), A(15) => A(15), A(14) => A(14), A(13) => 
                           A(13), A(12) => A(12), A(11) => A(11), A(10) => 
                           A(10), A(9) => A(9), A(8) => A(8), A(7) => A(7), 
                           A(6) => A(6), A(5) => A(5), A(4) => A(4), A(3) => 
                           A(3), A(2) => A(2), A(1) => A(1), A(0) => A(0), 
                           B(31) => n6, B(30) => n7, B(29) => n8, B(28) => n9, 
                           B(27) => new_B_27_port, B(26) => new_B_26_port, 
                           B(25) => new_B_25_port, B(24) => new_B_24_port, 
                           B(23) => new_B_23_port, B(22) => new_B_22_port, 
                           B(21) => new_B_21_port, B(20) => new_B_20_port, 
                           B(19) => new_B_19_port, B(18) => new_B_18_port, 
                           B(17) => new_B_17_port, B(16) => new_B_16_port, 
                           B(15) => new_B_15_port, B(14) => new_B_14_port, 
                           B(13) => new_B_13_port, B(12) => new_B_12_port, 
                           B(11) => new_B_11_port, B(10) => new_B_10_port, B(9)
                           => new_B_9_port, B(8) => new_B_8_port, B(7) => 
                           new_B_7_port, B(6) => new_B_6_port, B(5) => 
                           new_B_5_port, B(4) => new_B_4_port, B(3) => 
                           new_B_3_port, B(2) => new_B_2_port, B(1) => 
                           new_B_1_port, B(0) => new_B_0_port, Cin => n1, 
                           Cout(7) => net48714, Cout(6) => carry_pro_7_port, 
                           Cout(5) => carry_pro_6_port, Cout(4) => 
                           carry_pro_5_port, Cout(3) => carry_pro_4_port, 
                           Cout(2) => carry_pro_3_port, Cout(1) => 
                           carry_pro_2_port, Cout(0) => carry_pro_1_port);
   add : sum_gen_N32_0 port map( A(31) => A(31), A(30) => A(30), A(29) => A(29)
                           , A(28) => A(28), A(27) => A(27), A(26) => A(26), 
                           A(25) => A(25), A(24) => A(24), A(23) => A(23), 
                           A(22) => A(22), A(21) => A(21), A(20) => A(20), 
                           A(19) => A(19), A(18) => A(18), A(17) => A(17), 
                           A(16) => A(16), A(15) => A(15), A(14) => A(14), 
                           A(13) => A(13), A(12) => A(12), A(11) => A(11), 
                           A(10) => A(10), A(9) => A(9), A(8) => A(8), A(7) => 
                           A(7), A(6) => A(6), A(5) => A(5), A(4) => A(4), A(3)
                           => A(3), A(2) => A(2), A(1) => A(1), A(0) => A(0), 
                           B(31) => new_B_31_port, B(30) => new_B_30_port, 
                           B(29) => new_B_29_port, B(28) => new_B_28_port, 
                           B(27) => new_B_31_port, B(26) => new_B_26_port, 
                           B(25) => new_B_25_port, B(24) => new_B_24_port, 
                           B(23) => new_B_23_port, B(22) => new_B_22_port, 
                           B(21) => new_B_21_port, B(20) => new_B_20_port, 
                           B(19) => new_B_19_port, B(18) => new_B_18_port, 
                           B(17) => new_B_17_port, B(16) => new_B_16_port, 
                           B(15) => new_B_15_port, B(14) => new_B_14_port, 
                           B(13) => new_B_13_port, B(12) => new_B_12_port, 
                           B(11) => new_B_11_port, B(10) => new_B_10_port, B(9)
                           => new_B_9_port, B(8) => new_B_8_port, B(7) => 
                           new_B_7_port, B(6) => new_B_6_port, B(5) => 
                           new_B_5_port, B(4) => new_B_4_port, B(3) => 
                           new_B_3_port, B(2) => new_B_2_port, B(1) => 
                           new_B_1_port, B(0) => new_B_0_port, Cin(8) => n10, 
                           Cin(7) => carry_pro_7_port, Cin(6) => 
                           carry_pro_6_port, Cin(5) => carry_pro_5_port, Cin(4)
                           => carry_pro_4_port, Cin(3) => carry_pro_3_port, 
                           Cin(2) => carry_pro_2_port, Cin(1) => 
                           carry_pro_1_port, Cin(0) => n1, S(31) => S(31), 
                           S(30) => S(30), S(29) => S(29), S(28) => S(28), 
                           S(27) => S(27), S(26) => S(26), S(25) => S(25), 
                           S(24) => S(24), S(23) => S(23), S(22) => S(22), 
                           S(21) => S(21), S(20) => S(20), S(19) => S(19), 
                           S(18) => S(18), S(17) => S(17), S(16) => S(16), 
                           S(15) => S(15), S(14) => S(14), S(13) => S(13), 
                           S(12) => S(12), S(11) => S(11), S(10) => S(10), S(9)
                           => S(9), S(8) => S(8), S(7) => S(7), S(6) => S(6), 
                           S(5) => S(5), S(4) => S(4), S(3) => S(3), S(2) => 
                           S(2), S(1) => S(1), S(0) => S(0));
   n1 <= '0';
   n11 <= '0';
   n2 <= '0';
   n3 <= '0';
   n4 <= '0';
   n5 <= '0';
   n6 <= '0';
   n7 <= '0';
   n8 <= '0';
   n9 <= '0';
   n10 <= '0';

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity extender_32 is

   port( IN1 : in std_logic_vector (31 downto 0);  CTRL, SIGN : in std_logic;  
         OUT1 : out std_logic_vector (31 downto 0));

end extender_32;

architecture SYN_Bhe of extender_32 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X4
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal OUT1_31_port, OUT1_24_port, OUT1_23_port, OUT1_22_port, OUT1_21_port,
      OUT1_20_port, OUT1_19_port, OUT1_18_port, OUT1_17_port, OUT1_16_port, n4,
      n5, n6, n8, n9, n10, n13, n11, n7, n12, n1, n2, n3, n14, n15, n16, n17, 
      n18, OUT1_25_port, OUT1_28_port : std_logic;

begin
   OUT1 <= ( OUT1_28_port, OUT1_25_port, OUT1_25_port, OUT1_28_port, 
      OUT1_28_port, OUT1_28_port, OUT1_25_port, OUT1_24_port, OUT1_23_port, 
      OUT1_22_port, OUT1_21_port, OUT1_20_port, OUT1_19_port, OUT1_18_port, 
      OUT1_17_port, OUT1_16_port, IN1(15), IN1(14), IN1(13), IN1(12), IN1(11), 
      IN1(10), IN1(9), IN1(8), IN1(7), IN1(6), IN1(5), IN1(4), IN1(3), IN1(2), 
      IN1(1), IN1(0) );
   
   U2 : CLKBUF_X1 port map( A => CTRL, Z => n15);
   U3 : NAND2_X2 port map( A1 => n14, A2 => n8, ZN => OUT1_21_port);
   U4 : NAND2_X2 port map( A1 => n18, A2 => n12, ZN => OUT1_17_port);
   U5 : BUF_X4 port map( A => OUT1_31_port, Z => OUT1_28_port);
   U6 : BUF_X4 port map( A => n16, Z => OUT1_25_port);
   U7 : NAND2_X1 port map( A1 => n18, A2 => n5, ZN => OUT1_24_port);
   U8 : NAND2_X1 port map( A1 => n17, A2 => n9, ZN => OUT1_20_port);
   U9 : NAND2_X1 port map( A1 => n7, A2 => n14, ZN => OUT1_22_port);
   U10 : NAND2_X1 port map( A1 => n10, A2 => n14, ZN => OUT1_19_port);
   U11 : NAND2_X1 port map( A1 => SIGN, A2 => n1, ZN => n14);
   U12 : NAND2_X1 port map( A1 => n17, A2 => n11, ZN => OUT1_18_port);
   U13 : NAND2_X1 port map( A1 => n17, A2 => n13, ZN => OUT1_16_port);
   U14 : NAND2_X1 port map( A1 => n3, A2 => SIGN, ZN => n17);
   U15 : NAND2_X1 port map( A1 => n3, A2 => SIGN, ZN => n18);
   U16 : NOR2_X1 port map( A1 => CTRL, A2 => n2, ZN => n3);
   U17 : INV_X1 port map( A => IN1(15), ZN => n2);
   U18 : NAND2_X1 port map( A1 => CTRL, A2 => IN1(17), ZN => n12);
   U19 : NOR2_X1 port map( A1 => CTRL, A2 => n2, ZN => n1);
   U20 : NAND2_X1 port map( A1 => CTRL, A2 => IN1(22), ZN => n7);
   U21 : NAND2_X1 port map( A1 => CTRL, A2 => IN1(18), ZN => n11);
   U22 : NAND2_X1 port map( A1 => n18, A2 => n4, ZN => n16);
   U23 : NAND2_X1 port map( A1 => n15, A2 => IN1(24), ZN => n5);
   U24 : NAND2_X1 port map( A1 => n15, A2 => IN1(16), ZN => n13);
   U25 : NAND2_X1 port map( A1 => CTRL, A2 => IN1(20), ZN => n9);
   U26 : NAND2_X1 port map( A1 => CTRL, A2 => IN1(19), ZN => n10);
   U27 : NAND2_X1 port map( A1 => CTRL, A2 => IN1(23), ZN => n6);
   U28 : NAND2_X1 port map( A1 => CTRL, A2 => IN1(25), ZN => n4);
   U29 : NAND2_X1 port map( A1 => CTRL, A2 => IN1(21), ZN => n8);
   U30 : NAND2_X1 port map( A1 => n17, A2 => n6, ZN => OUT1_23_port);
   U31 : NAND2_X1 port map( A1 => n18, A2 => n4, ZN => OUT1_31_port);

end SYN_Bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity ff32_en_IR is

   port( D : in std_logic_vector (31 downto 0);  en, clk, rst : in std_logic;  
         Q : out std_logic_vector (31 downto 0));

end ff32_en_IR;

architecture SYN_behavioral of ff32_en_IR is

   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X2
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFS_X2
      port( D, CK, SN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_ff32_en_IR
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component DFFS_X1
      port( D, CK, SN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal net3591, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
      n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n33, n28
      , n29, n30, n31, n32 : std_logic;

begin
   
   Q_reg_31_inst : DFFR_X1 port map( D => D(31), CK => net3591, RN => n32, Q =>
                           Q(31), QN => n33);
   Q_reg_26_inst : DFFS_X1 port map( D => D(26), CK => net3591, SN => n32, Q =>
                           Q(26), QN => n27);
   Q_reg_25_inst : DFFR_X1 port map( D => D(25), CK => net3591, RN => n32, Q =>
                           Q(25), QN => n26);
   Q_reg_24_inst : DFFR_X1 port map( D => D(24), CK => net3591, RN => n32, Q =>
                           Q(24), QN => n25);
   Q_reg_23_inst : DFFR_X1 port map( D => D(23), CK => net3591, RN => n32, Q =>
                           Q(23), QN => n24);
   Q_reg_22_inst : DFFR_X1 port map( D => D(22), CK => net3591, RN => n32, Q =>
                           Q(22), QN => n23);
   Q_reg_21_inst : DFFR_X1 port map( D => D(21), CK => net3591, RN => n32, Q =>
                           Q(21), QN => n22);
   Q_reg_20_inst : DFFR_X1 port map( D => D(20), CK => net3591, RN => n32, Q =>
                           Q(20), QN => n21);
   Q_reg_19_inst : DFFR_X1 port map( D => D(19), CK => net3591, RN => n32, Q =>
                           Q(19), QN => n20);
   Q_reg_18_inst : DFFR_X1 port map( D => D(18), CK => net3591, RN => n32, Q =>
                           Q(18), QN => n19);
   Q_reg_17_inst : DFFR_X1 port map( D => D(17), CK => net3591, RN => n32, Q =>
                           Q(17), QN => n18);
   Q_reg_16_inst : DFFR_X1 port map( D => D(16), CK => net3591, RN => n32, Q =>
                           Q(16), QN => n17);
   Q_reg_15_inst : DFFR_X1 port map( D => D(15), CK => net3591, RN => n32, Q =>
                           Q(15), QN => n16);
   Q_reg_14_inst : DFFR_X1 port map( D => D(14), CK => net3591, RN => n32, Q =>
                           Q(14), QN => n15);
   Q_reg_13_inst : DFFR_X1 port map( D => D(13), CK => net3591, RN => n32, Q =>
                           Q(13), QN => n14);
   Q_reg_12_inst : DFFR_X1 port map( D => D(12), CK => net3591, RN => n32, Q =>
                           Q(12), QN => n13);
   Q_reg_11_inst : DFFR_X1 port map( D => D(11), CK => net3591, RN => n32, Q =>
                           Q(11), QN => n12);
   Q_reg_10_inst : DFFR_X1 port map( D => D(10), CK => net3591, RN => n32, Q =>
                           Q(10), QN => n11);
   Q_reg_9_inst : DFFR_X1 port map( D => D(9), CK => net3591, RN => n32, Q => 
                           Q(9), QN => n10);
   Q_reg_8_inst : DFFR_X1 port map( D => D(8), CK => net3591, RN => n32, Q => 
                           Q(8), QN => n9);
   Q_reg_7_inst : DFFR_X1 port map( D => D(7), CK => net3591, RN => n32, Q => 
                           Q(7), QN => n8);
   Q_reg_6_inst : DFFR_X1 port map( D => D(6), CK => net3591, RN => n32, Q => 
                           Q(6), QN => n7);
   Q_reg_5_inst : DFFR_X1 port map( D => D(5), CK => net3591, RN => n32, Q => 
                           Q(5), QN => n6);
   Q_reg_4_inst : DFFR_X1 port map( D => D(4), CK => net3591, RN => n32, Q => 
                           Q(4), QN => n5);
   Q_reg_3_inst : DFFR_X1 port map( D => D(3), CK => net3591, RN => n32, Q => 
                           Q(3), QN => n4);
   Q_reg_2_inst : DFFR_X1 port map( D => D(2), CK => net3591, RN => n32, Q => 
                           Q(2), QN => n3);
   Q_reg_1_inst : DFFR_X1 port map( D => D(1), CK => net3591, RN => n32, Q => 
                           Q(1), QN => n2);
   Q_reg_0_inst : DFFR_X1 port map( D => D(0), CK => net3591, RN => n32, Q => 
                           Q(0), QN => n1);
   clk_gate_Q_reg : SNPS_CLOCK_GATE_HIGH_ff32_en_IR port map( CLK => clk, EN =>
                           en, ENCLK => net3591);
   Q_reg_28_inst : DFFS_X2 port map( D => D(28), CK => net3591, SN => n32, Q =>
                           Q(28), QN => n31);
   Q_reg_30_inst : DFFS_X2 port map( D => D(30), CK => net3591, SN => n32, Q =>
                           Q(30), QN => n30);
   Q_reg_29_inst : DFFR_X1 port map( D => D(29), CK => net3591, RN => n32, Q =>
                           Q(29), QN => n29);
   Q_reg_27_inst : DFFR_X2 port map( D => D(27), CK => net3591, RN => n32, Q =>
                           Q(27), QN => n28);
   U2 : INV_X2 port map( A => rst, ZN => n32);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_0 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_0;

architecture SYN_USE_DEFA_ARCH_NAME of 
   SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net3615 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net3615);
   main_gate : AND2_X1 port map( A1 => net3615, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity predictor_2_0 is

   port( clock, reset, enable, taken_i : in std_logic;  prediction_o : out 
         std_logic);

end predictor_2_0;

architecture SYN_bhe of predictor_2_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal prediction_o_port, next_STATE_1_port, next_STATE_0_port, N11, N12, n3
      , n4, n6, n8, n9, n1, n2, net48713 : std_logic;

begin
   prediction_o <= prediction_o_port;
   
   next_STATE_reg_0_inst : DLH_X1 port map( G => enable, D => N11, Q => 
                           next_STATE_0_port);
   STATE_reg_0_inst : DFFR_X1 port map( D => n8, CK => clock, RN => n2, Q => n1
                           , QN => n9);
   next_STATE_reg_1_inst : DLH_X1 port map( G => enable, D => N12, Q => 
                           next_STATE_1_port);
   STATE_reg_1_inst : DFFR_X1 port map( D => n6, CK => clock, RN => n2, Q => 
                           prediction_o_port, QN => net48713);
   U2 : MUX2_X1 port map( A => prediction_o_port, B => next_STATE_1_port, S => 
                           enable, Z => n6);
   U4 : MUX2_X1 port map( A => n1, B => next_STATE_0_port, S => enable, Z => n8
                           );
   U9 : NOR2_X1 port map( A1 => prediction_o_port, A2 => taken_i, ZN => n3);
   U7 : NAND2_X1 port map( A1 => prediction_o_port, A2 => taken_i, ZN => n4);
   U5 : OAI21_X1 port map( B1 => n9, B2 => n3, A => n4, ZN => N12);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n1, A => n4, ZN => N11);
   U3 : INV_X1 port map( A => reset, ZN => n2);

end SYN_bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity mux41_0 is

   port( IN0, IN1, IN2, IN3 : in std_logic_vector (31 downto 0);  CTRL : in 
         std_logic_vector (1 downto 0);  OUT1 : out std_logic_vector (31 downto
         0));

end mux41_0;

architecture SYN_bhe of mux41_0 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n6, n7, n8, n45, n46, n51, n52, n71, n1, n2, n3, n4, n9, n10, n11
      , n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, 
      n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40
      , n41, n42, n43, n44, n47, n48, n49, n50, n53, n54, n55, n56, n57, n58, 
      n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, 
      n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, 
      n115, n116, n117, n118, n119, n120, n121 : std_logic;

begin
   
   U69 : AOI22_X1 port map( A1 => n7, A2 => IN1(18), B1 => n16, B2 => IN0(18), 
                           ZN => n51);
   U68 : AOI22_X1 port map( A1 => n5, A2 => IN3(18), B1 => n121, B2 => IN2(18),
                           ZN => n52);
   U60 : AOI22_X1 port map( A1 => n7, A2 => IN1(20), B1 => n16, B2 => IN0(20), 
                           ZN => n45);
   U101 : INV_X1 port map( A => CTRL(1), ZN => n71);
   U99 : NOR2_X1 port map( A1 => CTRL(0), A2 => CTRL(1), ZN => n8);
   U1 : NAND2_X1 port map( A1 => n86, A2 => n87, ZN => OUT1(30));
   U2 : NAND3_X2 port map( A1 => n43, A2 => n44, A3 => n47, ZN => OUT1(2));
   U3 : NAND3_X2 port map( A1 => n30, A2 => n31, A3 => n32, ZN => OUT1(4));
   U4 : NAND3_X2 port map( A1 => n35, A2 => n36, A3 => n37, ZN => OUT1(6));
   U5 : AOI222_X1 port map( A1 => n121, A2 => IN2(25), B1 => IN0(25), B2 => n16
                           , C1 => n7, C2 => IN1(25), ZN => n1);
   U6 : NAND2_X1 port map( A1 => n5, A2 => IN3(25), ZN => n2);
   U7 : NAND2_X1 port map( A1 => n1, A2 => n2, ZN => OUT1(25));
   U8 : AOI22_X1 port map( A1 => IN1(24), A2 => n7, B1 => IN3(24), B2 => n5, ZN
                           => n3);
   U9 : NAND2_X1 port map( A1 => n121, A2 => IN2(24), ZN => n4);
   U10 : NAND3_X1 port map( A1 => n4, A2 => n54, A3 => n3, ZN => OUT1(24));
   U11 : AOI22_X1 port map( A1 => IN0(31), A2 => n8, B1 => n7, B2 => IN1(31), 
                           ZN => n9);
   U12 : INV_X1 port map( A => n9, ZN => n24);
   U13 : AOI22_X1 port map( A1 => IN0(15), A2 => n16, B1 => n7, B2 => IN1(15), 
                           ZN => n10);
   U14 : INV_X1 port map( A => n10, ZN => n95);
   U15 : AOI22_X1 port map( A1 => IN0(23), A2 => n16, B1 => n7, B2 => IN1(23), 
                           ZN => n11);
   U16 : INV_X1 port map( A => n11, ZN => n50);
   U17 : AOI22_X1 port map( A1 => IN3(28), A2 => n5, B1 => IN2(28), B2 => n121,
                           ZN => n12);
   U18 : NAND3_X1 port map( A1 => n116, A2 => n117, A3 => n12, ZN => OUT1(28));
   U19 : AOI22_X1 port map( A1 => IN1(26), A2 => n7, B1 => IN3(26), B2 => n5, 
                           ZN => n13);
   U20 : NAND2_X1 port map( A1 => n121, A2 => IN2(26), ZN => n14);
   U21 : NAND3_X1 port map( A1 => n14, A2 => n53, A3 => n13, ZN => OUT1(26));
   U22 : AOI22_X1 port map( A1 => IN0(13), A2 => n16, B1 => n7, B2 => IN1(13), 
                           ZN => n15);
   U23 : INV_X1 port map( A => n15, ZN => n120);
   U24 : NAND2_X2 port map( A1 => n74, A2 => n75, ZN => OUT1(10));
   U25 : NAND3_X2 port map( A1 => n58, A2 => n59, A3 => n60, ZN => OUT1(0));
   U26 : AND2_X2 port map( A1 => CTRL(0), A2 => CTRL(1), ZN => n5);
   U27 : BUF_X1 port map( A => n6, Z => n121);
   U28 : AND2_X2 port map( A1 => n71, A2 => CTRL(0), ZN => n7);
   U29 : BUF_X2 port map( A => n8, Z => n16);
   U30 : NAND2_X2 port map( A1 => n63, A2 => n64, ZN => OUT1(17));
   U31 : NAND2_X2 port map( A1 => n81, A2 => n82, ZN => OUT1(19));
   U32 : NAND2_X2 port map( A1 => n101, A2 => n102, ZN => OUT1(14));
   U33 : NAND2_X2 port map( A1 => n91, A2 => n92, ZN => OUT1(9));
   U34 : NAND2_X2 port map( A1 => n106, A2 => n107, ZN => OUT1(12));
   U35 : NAND2_X2 port map( A1 => n76, A2 => n77, ZN => OUT1(16));
   U36 : NAND2_X2 port map( A1 => n72, A2 => n73, ZN => OUT1(7));
   U37 : NAND2_X2 port map( A1 => n33, A2 => n34, ZN => OUT1(8));
   U38 : NAND2_X2 port map( A1 => n38, A2 => n39, ZN => OUT1(21));
   U39 : NAND2_X2 port map( A1 => n111, A2 => n112, ZN => OUT1(3));
   U40 : NAND2_X2 port map( A1 => n25, A2 => n26, ZN => OUT1(22));
   U41 : NAND2_X2 port map( A1 => n48, A2 => n49, ZN => OUT1(23));
   U42 : NAND2_X2 port map( A1 => n51, A2 => n52, ZN => OUT1(18));
   U43 : NAND2_X2 port map( A1 => n45, A2 => n46, ZN => OUT1(20));
   U44 : NAND3_X2 port map( A1 => n68, A2 => n69, A3 => n70, ZN => OUT1(5));
   U45 : NAND3_X2 port map( A1 => n55, A2 => n56, A3 => n57, ZN => OUT1(1));
   U46 : NAND2_X1 port map( A1 => n118, A2 => n119, ZN => OUT1(13));
   U47 : NAND2_X1 port map( A1 => n93, A2 => n94, ZN => OUT1(15));
   U48 : NAND2_X1 port map( A1 => n17, A2 => n18, ZN => OUT1(27));
   U49 : NAND2_X1 port map( A1 => n61, A2 => n62, ZN => OUT1(11));
   U50 : NOR2_X1 port map( A1 => CTRL(0), A2 => n71, ZN => n6);
   U51 : NAND2_X1 port map( A1 => IN1(2), A2 => n7, ZN => n47);
   U52 : AOI22_X1 port map( A1 => n16, A2 => IN0(2), B1 => n121, B2 => IN2(2), 
                           ZN => n44);
   U53 : AOI21_X1 port map( B1 => IN1(3), B2 => n7, A => n113, ZN => n112);
   U54 : NAND2_X1 port map( A1 => n114, A2 => n115, ZN => n113);
   U55 : NAND2_X1 port map( A1 => n16, A2 => IN0(3), ZN => n115);
   U56 : NAND2_X1 port map( A1 => IN2(3), A2 => n6, ZN => n114);
   U57 : AOI21_X1 port map( B1 => IN2(12), B2 => n121, A => n108, ZN => n107);
   U58 : NAND2_X1 port map( A1 => n109, A2 => n110, ZN => n108);
   U59 : NAND2_X1 port map( A1 => n16, A2 => IN0(12), ZN => n110);
   U61 : NAND2_X1 port map( A1 => IN1(12), A2 => n7, ZN => n109);
   U62 : AOI21_X1 port map( B1 => IN2(13), B2 => n121, A => n120, ZN => n119);
   U63 : AOI21_X1 port map( B1 => IN2(14), B2 => n121, A => n103, ZN => n102);
   U64 : NAND2_X1 port map( A1 => n104, A2 => n105, ZN => n103);
   U65 : NAND2_X1 port map( A1 => n16, A2 => IN0(14), ZN => n105);
   U66 : NAND2_X1 port map( A1 => IN1(14), A2 => n7, ZN => n104);
   U67 : AOI21_X1 port map( B1 => IN2(15), B2 => n121, A => n95, ZN => n94);
   U70 : AOI222_X1 port map( A1 => IN1(8), A2 => n7, B1 => IN2(8), B2 => n6, C1
                           => n16, C2 => IN0(8), ZN => n34);
   U71 : AOI222_X1 port map( A1 => n7, A2 => IN1(9), B1 => IN2(9), B2 => n6, C1
                           => n16, C2 => IN0(9), ZN => n92);
   U72 : AOI21_X1 port map( B1 => IN2(22), B2 => n121, A => n27, ZN => n26);
   U73 : NAND2_X1 port map( A1 => n28, A2 => n29, ZN => n27);
   U74 : NAND2_X1 port map( A1 => n16, A2 => IN0(22), ZN => n29);
   U75 : NAND2_X1 port map( A1 => IN1(22), A2 => n7, ZN => n28);
   U76 : NAND2_X1 port map( A1 => IN1(4), A2 => n7, ZN => n32);
   U77 : AOI22_X1 port map( A1 => n6, A2 => IN2(4), B1 => n8, B2 => IN0(4), ZN 
                           => n31);
   U78 : NAND2_X1 port map( A1 => IN1(5), A2 => n7, ZN => n70);
   U79 : AOI22_X1 port map( A1 => n6, A2 => IN2(5), B1 => n8, B2 => IN0(5), ZN 
                           => n69);
   U80 : NAND2_X1 port map( A1 => IN1(6), A2 => n7, ZN => n37);
   U81 : AOI22_X1 port map( A1 => IN2(6), A2 => n6, B1 => n8, B2 => IN0(6), ZN 
                           => n36);
   U82 : AOI222_X1 port map( A1 => IN2(7), A2 => n6, B1 => n7, B2 => IN1(7), C1
                           => n16, C2 => IN0(7), ZN => n73);
   U83 : NAND2_X1 port map( A1 => IN1(0), A2 => n7, ZN => n60);
   U84 : AOI22_X1 port map( A1 => n121, A2 => IN2(0), B1 => n16, B2 => IN0(0), 
                           ZN => n59);
   U85 : NAND2_X1 port map( A1 => IN1(1), A2 => n7, ZN => n57);
   U86 : AOI22_X1 port map( A1 => n121, A2 => IN2(1), B1 => n16, B2 => IN0(1), 
                           ZN => n56);
   U87 : AOI21_X1 port map( B1 => IN2(21), B2 => n121, A => n40, ZN => n39);
   U88 : NAND2_X1 port map( A1 => n41, A2 => n42, ZN => n40);
   U89 : NAND2_X1 port map( A1 => n16, A2 => IN0(21), ZN => n42);
   U90 : NAND2_X1 port map( A1 => IN1(21), A2 => n7, ZN => n41);
   U91 : NAND2_X1 port map( A1 => n16, A2 => IN0(24), ZN => n54);
   U92 : NAND2_X1 port map( A1 => n16, A2 => IN0(26), ZN => n53);
   U93 : AOI21_X1 port map( B1 => IN2(27), B2 => n121, A => n19, ZN => n18);
   U94 : NAND2_X1 port map( A1 => n20, A2 => n21, ZN => n19);
   U95 : NAND2_X1 port map( A1 => n16, A2 => IN0(27), ZN => n21);
   U96 : NAND2_X1 port map( A1 => IN1(27), A2 => n7, ZN => n20);
   U97 : AOI21_X1 port map( B1 => IN2(30), B2 => n121, A => n88, ZN => n87);
   U98 : NAND2_X1 port map( A1 => n89, A2 => n90, ZN => n88);
   U100 : NAND2_X1 port map( A1 => n16, A2 => IN0(30), ZN => n90);
   U102 : NAND2_X1 port map( A1 => IN1(30), A2 => n7, ZN => n89);
   U103 : AOI21_X1 port map( B1 => IN2(31), B2 => n6, A => n24, ZN => n23);
   U104 : AOI222_X1 port map( A1 => IN2(10), A2 => n121, B1 => IN1(10), B2 => 
                           n7, C1 => n16, C2 => IN0(10), ZN => n75);
   U105 : AOI222_X1 port map( A1 => IN2(11), A2 => n121, B1 => IN1(11), B2 => 
                           n7, C1 => n16, C2 => IN0(11), ZN => n62);
   U106 : AOI21_X1 port map( B1 => IN2(16), B2 => n121, A => n78, ZN => n77);
   U107 : NAND2_X1 port map( A1 => n79, A2 => n80, ZN => n78);
   U108 : NAND2_X1 port map( A1 => n16, A2 => IN0(16), ZN => n80);
   U109 : NAND2_X1 port map( A1 => IN1(16), A2 => n7, ZN => n79);
   U110 : AOI21_X1 port map( B1 => IN2(17), B2 => n121, A => n65, ZN => n64);
   U111 : NAND2_X1 port map( A1 => n66, A2 => n67, ZN => n65);
   U112 : NAND2_X1 port map( A1 => n16, A2 => IN0(17), ZN => n67);
   U113 : NAND2_X1 port map( A1 => IN1(17), A2 => n7, ZN => n66);
   U114 : AOI21_X1 port map( B1 => IN2(19), B2 => n121, A => n83, ZN => n82);
   U115 : NAND2_X1 port map( A1 => n84, A2 => n85, ZN => n83);
   U116 : NAND2_X1 port map( A1 => n16, A2 => IN0(19), ZN => n85);
   U117 : NAND2_X1 port map( A1 => IN1(19), A2 => n7, ZN => n84);
   U118 : NAND2_X1 port map( A1 => n16, A2 => IN0(28), ZN => n117);
   U119 : NAND2_X1 port map( A1 => IN1(28), A2 => n7, ZN => n116);
   U120 : AOI21_X1 port map( B1 => IN2(29), B2 => n121, A => n98, ZN => n97);
   U121 : NAND2_X1 port map( A1 => n99, A2 => n100, ZN => n98);
   U122 : NAND2_X1 port map( A1 => n16, A2 => IN0(29), ZN => n100);
   U123 : NAND2_X1 port map( A1 => IN1(29), A2 => n7, ZN => n99);
   U124 : NAND2_X1 port map( A1 => n96, A2 => n97, ZN => OUT1(29));
   U125 : NAND2_X1 port map( A1 => IN3(27), A2 => n5, ZN => n17);
   U126 : NAND2_X1 port map( A1 => IN3(31), A2 => n5, ZN => n22);
   U127 : NAND2_X1 port map( A1 => n22, A2 => n23, ZN => OUT1(31));
   U128 : NAND2_X1 port map( A1 => IN3(22), A2 => n5, ZN => n25);
   U129 : NAND2_X1 port map( A1 => IN3(4), A2 => n5, ZN => n30);
   U130 : NAND2_X1 port map( A1 => IN3(8), A2 => n5, ZN => n33);
   U131 : NAND2_X1 port map( A1 => IN3(6), A2 => n5, ZN => n35);
   U132 : NAND2_X1 port map( A1 => IN3(21), A2 => n5, ZN => n38);
   U133 : NAND2_X1 port map( A1 => IN3(2), A2 => n5, ZN => n43);
   U134 : NAND2_X1 port map( A1 => IN3(23), A2 => n5, ZN => n48);
   U135 : AOI21_X1 port map( B1 => IN2(23), B2 => n121, A => n50, ZN => n49);
   U136 : NAND2_X1 port map( A1 => IN3(1), A2 => n5, ZN => n55);
   U137 : NAND2_X1 port map( A1 => IN3(0), A2 => n5, ZN => n58);
   U138 : NAND2_X1 port map( A1 => IN3(11), A2 => n5, ZN => n61);
   U139 : NAND2_X1 port map( A1 => IN3(17), A2 => n5, ZN => n63);
   U140 : NAND2_X1 port map( A1 => IN3(5), A2 => n5, ZN => n68);
   U141 : NAND2_X1 port map( A1 => IN3(7), A2 => n5, ZN => n72);
   U142 : NAND2_X1 port map( A1 => IN3(10), A2 => n5, ZN => n74);
   U143 : NAND2_X1 port map( A1 => IN3(16), A2 => n5, ZN => n76);
   U144 : NAND2_X1 port map( A1 => IN3(19), A2 => n5, ZN => n81);
   U145 : NAND2_X1 port map( A1 => IN3(30), A2 => n5, ZN => n86);
   U146 : NAND2_X1 port map( A1 => IN3(9), A2 => n5, ZN => n91);
   U147 : NAND2_X1 port map( A1 => IN3(15), A2 => n5, ZN => n93);
   U148 : NAND2_X1 port map( A1 => IN3(29), A2 => n5, ZN => n96);
   U149 : NAND2_X1 port map( A1 => IN3(14), A2 => n5, ZN => n101);
   U150 : NAND2_X1 port map( A1 => IN3(12), A2 => n5, ZN => n106);
   U151 : NAND2_X1 port map( A1 => IN3(3), A2 => n5, ZN => n111);
   U152 : NAND2_X1 port map( A1 => IN3(13), A2 => n5, ZN => n118);
   U153 : AOI22_X1 port map( A1 => n5, A2 => IN3(20), B1 => n121, B2 => IN2(20)
                           , ZN => n46);

end SYN_bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity add4 is

   port( IN1 : in std_logic_vector (31 downto 0);  OUT1 : out std_logic_vector 
         (31 downto 0));

end add4;

architecture SYN_bhe of add4 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal OUT1_31_port, OUT1_30_port, OUT1_29_port, OUT1_28_port, OUT1_27_port,
      OUT1_26_port, OUT1_25_port, OUT1_24_port, OUT1_23_port, OUT1_22_port, 
      OUT1_21_port, OUT1_20_port, OUT1_19_port, OUT1_18_port, OUT1_17_port, 
      OUT1_16_port, OUT1_15_port, OUT1_14_port, OUT1_13_port, OUT1_12_port, 
      OUT1_11_port, OUT1_10_port, OUT1_9_port, OUT1_8_port, OUT1_7_port, 
      OUT1_6_port, OUT1_5_port, OUT1_4_port, OUT1_3_port, OUT1_2_port, n1, n2, 
      n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, 
      n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33
      , n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47 : 
      std_logic;

begin
   OUT1 <= ( OUT1_31_port, OUT1_30_port, OUT1_29_port, OUT1_28_port, 
      OUT1_27_port, OUT1_26_port, OUT1_25_port, OUT1_24_port, OUT1_23_port, 
      OUT1_22_port, OUT1_21_port, OUT1_20_port, OUT1_19_port, OUT1_18_port, 
      OUT1_17_port, OUT1_16_port, OUT1_15_port, OUT1_14_port, OUT1_13_port, 
      OUT1_12_port, OUT1_11_port, OUT1_10_port, OUT1_9_port, OUT1_8_port, 
      OUT1_7_port, OUT1_6_port, OUT1_5_port, OUT1_4_port, OUT1_3_port, 
      OUT1_2_port, IN1(1), IN1(0) );
   
   U3 : NAND2_X1 port map( A1 => IN1(15), A2 => n15, ZN => n1);
   U4 : NOR4_X1 port map( A1 => n17, A2 => n16, A3 => n18, A4 => n1, ZN => n2);
   U5 : NAND3_X1 port map( A1 => n14, A2 => IN1(13), A3 => n2, ZN => n20);
   U6 : XOR2_X1 port map( A => n39, B => IN1(29), Z => OUT1_29_port);
   U7 : NAND2_X1 port map( A1 => n44, A2 => IN1(6), ZN => n3);
   U8 : XNOR2_X1 port map( A => n3, B => IN1(7), ZN => OUT1_7_port);
   U9 : NOR2_X1 port map( A1 => n8, A2 => n9, ZN => n4);
   U10 : XOR2_X1 port map( A => IN1(11), B => n4, Z => OUT1_11_port);
   U11 : NOR2_X1 port map( A1 => n18, A2 => n13, ZN => n5);
   U12 : XOR2_X1 port map( A => IN1(15), B => n5, Z => OUT1_15_port);
   U13 : XOR2_X1 port map( A => n21, B => IN1(17), Z => OUT1_17_port);
   U14 : XOR2_X1 port map( A => n24, B => IN1(19), Z => OUT1_19_port);
   U15 : XOR2_X1 port map( A => n27, B => IN1(21), Z => OUT1_21_port);
   U16 : XOR2_X1 port map( A => n30, B => IN1(23), Z => OUT1_23_port);
   U17 : XOR2_X1 port map( A => n33, B => IN1(25), Z => OUT1_25_port);
   U18 : XOR2_X1 port map( A => n36, B => IN1(27), Z => OUT1_27_port);
   U19 : INV_X1 port map( A => n40, ZN => n6);
   U20 : NAND2_X1 port map( A1 => IN1(30), A2 => n6, ZN => n7);
   U21 : XNOR2_X1 port map( A => IN1(31), B => n7, ZN => OUT1_31_port);
   U22 : NOR2_X1 port map( A1 => n45, A2 => n16, ZN => n10);
   U23 : XOR2_X1 port map( A => n8, B => n9, Z => OUT1_10_port);
   U24 : NAND4_X1 port map( A1 => IN1(8), A2 => IN1(9), A3 => IN1(10), A4 => 
                           IN1(11), ZN => n16);
   U25 : XNOR2_X1 port map( A => n10, B => n17, ZN => OUT1_12_port);
   U26 : XOR2_X1 port map( A => IN1(13), B => n12, Z => OUT1_13_port);
   U27 : XNOR2_X1 port map( A => n13, B => IN1(14), ZN => OUT1_14_port);
   U28 : XNOR2_X1 port map( A => n20, B => IN1(16), ZN => OUT1_16_port);
   U29 : XNOR2_X1 port map( A => n23, B => IN1(18), ZN => OUT1_18_port);
   U30 : XNOR2_X1 port map( A => n26, B => IN1(20), ZN => OUT1_20_port);
   U31 : XNOR2_X1 port map( A => n29, B => IN1(22), ZN => OUT1_22_port);
   U32 : XNOR2_X1 port map( A => n32, B => IN1(24), ZN => OUT1_24_port);
   U33 : XNOR2_X1 port map( A => n35, B => IN1(26), ZN => OUT1_26_port);
   U34 : XNOR2_X1 port map( A => n38, B => IN1(28), ZN => OUT1_28_port);
   U35 : XNOR2_X1 port map( A => n40, B => IN1(30), ZN => OUT1_30_port);
   U36 : XNOR2_X1 port map( A => IN1(2), B => n41, ZN => OUT1_3_port);
   U37 : XOR2_X1 port map( A => IN1(4), B => n14, Z => OUT1_4_port);
   U38 : XOR2_X1 port map( A => n42, B => n43, Z => OUT1_5_port);
   U39 : XOR2_X1 port map( A => IN1(6), B => n44, Z => OUT1_6_port);
   U40 : XOR2_X1 port map( A => n46, B => n45, Z => OUT1_8_port);
   U41 : XOR2_X1 port map( A => IN1(9), B => n47, Z => OUT1_9_port);
   U42 : NAND2_X1 port map( A1 => n14, A2 => n15, ZN => n45);
   U43 : NAND2_X1 port map( A1 => n12, A2 => IN1(13), ZN => n13);
   U44 : NOR2_X1 port map( A1 => n45, A2 => n46, ZN => n47);
   U45 : NAND2_X1 port map( A1 => n47, A2 => IN1(9), ZN => n9);
   U46 : NAND2_X1 port map( A1 => n14, A2 => IN1(4), ZN => n43);
   U47 : NOR2_X1 port map( A1 => n43, A2 => n42, ZN => n44);
   U48 : NAND2_X1 port map( A1 => n39, A2 => IN1(29), ZN => n40);
   U49 : NAND2_X1 port map( A1 => n36, A2 => IN1(27), ZN => n38);
   U50 : INV_X1 port map( A => IN1(5), ZN => n42);
   U51 : AND4_X1 port map( A1 => IN1(5), A2 => IN1(4), A3 => IN1(6), A4 => 
                           IN1(7), ZN => n15);
   U52 : INV_X1 port map( A => IN1(3), ZN => n41);
   U53 : INV_X1 port map( A => IN1(2), ZN => OUT1_2_port);
   U54 : NAND2_X1 port map( A1 => n21, A2 => IN1(17), ZN => n23);
   U55 : NAND2_X1 port map( A1 => n24, A2 => IN1(19), ZN => n26);
   U56 : NAND2_X1 port map( A1 => n27, A2 => IN1(21), ZN => n29);
   U57 : NAND2_X1 port map( A1 => n30, A2 => IN1(23), ZN => n32);
   U58 : NAND2_X1 port map( A1 => n33, A2 => IN1(25), ZN => n35);
   U59 : NOR2_X1 port map( A1 => n11, A2 => n17, ZN => n12);
   U60 : NOR2_X1 port map( A1 => n38, A2 => n37, ZN => n39);
   U61 : NOR2_X1 port map( A1 => n41, A2 => OUT1_2_port, ZN => n14);
   U62 : NOR2_X1 port map( A1 => n20, A2 => n19, ZN => n21);
   U63 : NOR2_X1 port map( A1 => n23, A2 => n22, ZN => n24);
   U64 : NOR2_X1 port map( A1 => n26, A2 => n25, ZN => n27);
   U65 : NOR2_X1 port map( A1 => n29, A2 => n28, ZN => n30);
   U66 : NOR2_X1 port map( A1 => n32, A2 => n31, ZN => n33);
   U67 : NOR2_X1 port map( A1 => n35, A2 => n34, ZN => n36);
   U68 : INV_X1 port map( A => IN1(14), ZN => n18);
   U69 : INV_X1 port map( A => IN1(12), ZN => n17);
   U70 : INV_X1 port map( A => IN1(16), ZN => n19);
   U71 : INV_X1 port map( A => IN1(18), ZN => n22);
   U72 : INV_X1 port map( A => IN1(20), ZN => n25);
   U73 : INV_X1 port map( A => IN1(22), ZN => n28);
   U74 : INV_X1 port map( A => IN1(24), ZN => n31);
   U75 : INV_X1 port map( A => IN1(26), ZN => n34);
   U76 : INV_X1 port map( A => IN1(8), ZN => n46);
   U77 : INV_X1 port map( A => IN1(28), ZN => n37);
   U78 : INV_X1 port map( A => IN1(10), ZN => n8);
   U79 : INV_X1 port map( A => n10, ZN => n11);

end SYN_bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity ff32_en_0 is

   port( D : in std_logic_vector (31 downto 0);  en, clk, rst : in std_logic;  
         Q : out std_logic_vector (31 downto 0));

end ff32_en_0;

architecture SYN_behavioral of ff32_en_0 is

   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_ff32_en_0
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal net3606, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
      n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29
      , n30, n31, n33, n32 : std_logic;

begin
   
   Q_reg_31_inst : DFFR_X1 port map( D => D(31), CK => net3606, RN => n32, Q =>
                           Q(31), QN => n33);
   Q_reg_30_inst : DFFR_X1 port map( D => D(30), CK => net3606, RN => n32, Q =>
                           Q(30), QN => n31);
   Q_reg_29_inst : DFFR_X1 port map( D => D(29), CK => net3606, RN => n32, Q =>
                           Q(29), QN => n30);
   Q_reg_28_inst : DFFR_X1 port map( D => D(28), CK => net3606, RN => n32, Q =>
                           Q(28), QN => n29);
   Q_reg_27_inst : DFFR_X1 port map( D => D(27), CK => net3606, RN => n32, Q =>
                           Q(27), QN => n28);
   Q_reg_26_inst : DFFR_X1 port map( D => D(26), CK => net3606, RN => n32, Q =>
                           Q(26), QN => n27);
   Q_reg_25_inst : DFFR_X1 port map( D => D(25), CK => net3606, RN => n32, Q =>
                           Q(25), QN => n26);
   Q_reg_24_inst : DFFR_X1 port map( D => D(24), CK => net3606, RN => n32, Q =>
                           Q(24), QN => n25);
   Q_reg_23_inst : DFFR_X1 port map( D => D(23), CK => net3606, RN => n32, Q =>
                           Q(23), QN => n24);
   Q_reg_22_inst : DFFR_X1 port map( D => D(22), CK => net3606, RN => n32, Q =>
                           Q(22), QN => n23);
   Q_reg_21_inst : DFFR_X1 port map( D => D(21), CK => net3606, RN => n32, Q =>
                           Q(21), QN => n22);
   Q_reg_20_inst : DFFR_X1 port map( D => D(20), CK => net3606, RN => n32, Q =>
                           Q(20), QN => n21);
   Q_reg_19_inst : DFFR_X1 port map( D => D(19), CK => net3606, RN => n32, Q =>
                           Q(19), QN => n20);
   Q_reg_18_inst : DFFR_X1 port map( D => D(18), CK => net3606, RN => n32, Q =>
                           Q(18), QN => n19);
   Q_reg_17_inst : DFFR_X1 port map( D => D(17), CK => net3606, RN => n32, Q =>
                           Q(17), QN => n18);
   Q_reg_16_inst : DFFR_X1 port map( D => D(16), CK => net3606, RN => n32, Q =>
                           Q(16), QN => n17);
   Q_reg_15_inst : DFFR_X1 port map( D => D(15), CK => net3606, RN => n32, Q =>
                           Q(15), QN => n16);
   Q_reg_14_inst : DFFR_X1 port map( D => D(14), CK => net3606, RN => n32, Q =>
                           Q(14), QN => n15);
   Q_reg_13_inst : DFFR_X1 port map( D => D(13), CK => net3606, RN => n32, Q =>
                           Q(13), QN => n14);
   Q_reg_12_inst : DFFR_X1 port map( D => D(12), CK => net3606, RN => n32, Q =>
                           Q(12), QN => n13);
   Q_reg_11_inst : DFFR_X1 port map( D => D(11), CK => net3606, RN => n32, Q =>
                           Q(11), QN => n12);
   Q_reg_10_inst : DFFR_X1 port map( D => D(10), CK => net3606, RN => n32, Q =>
                           Q(10), QN => n11);
   Q_reg_9_inst : DFFR_X1 port map( D => D(9), CK => net3606, RN => n32, Q => 
                           Q(9), QN => n10);
   Q_reg_8_inst : DFFR_X1 port map( D => D(8), CK => net3606, RN => n32, Q => 
                           Q(8), QN => n9);
   Q_reg_7_inst : DFFR_X1 port map( D => D(7), CK => net3606, RN => n32, Q => 
                           Q(7), QN => n8);
   Q_reg_6_inst : DFFR_X1 port map( D => D(6), CK => net3606, RN => n32, Q => 
                           Q(6), QN => n7);
   Q_reg_5_inst : DFFR_X1 port map( D => D(5), CK => net3606, RN => n32, Q => 
                           Q(5), QN => n6);
   Q_reg_4_inst : DFFR_X1 port map( D => D(4), CK => net3606, RN => n32, Q => 
                           Q(4), QN => n5);
   Q_reg_3_inst : DFFR_X1 port map( D => D(3), CK => net3606, RN => n32, Q => 
                           Q(3), QN => n4);
   Q_reg_2_inst : DFFR_X1 port map( D => D(2), CK => net3606, RN => n32, Q => 
                           Q(2), QN => n3);
   Q_reg_1_inst : DFFR_X1 port map( D => D(1), CK => net3606, RN => n32, Q => 
                           Q(1), QN => n2);
   Q_reg_0_inst : DFFR_X1 port map( D => D(0), CK => net3606, RN => n32, Q => 
                           Q(0), QN => n1);
   clk_gate_Q_reg : SNPS_CLOCK_GATE_HIGH_ff32_en_0 port map( CLK => clk, EN => 
                           en, ENCLK => net3606);
   U2 : INV_X2 port map( A => rst, ZN => n32);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity fw_logic is

   port( D1_i, rAdec_i, D2_i, D3_i, rA_i, rB_i : in std_logic_vector (4 downto 
         0);  S_mem_W, S_wb_W, S_exe_W : in std_logic;  S_FWAdec, S_FWA, S_FWB 
         : out std_logic_vector (1 downto 0);  S_mem_LOAD_BAR : in std_logic);

end fw_logic;

architecture SYN_beh of fw_logic is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal S_FWAdec_1_port, S_FWAdec_0_port, S_FWA_1_port, S_FWA_0_port, n22, 
      n23, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n51, n52, n53
      , n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n45, n44, 
      n43, n42, n41, n40, n1, n2, n3, n5, n6, n7, n8, n9, n10, n11, n12, n13, 
      n14, n15, n16, n17, n18, n19, n20, n21, n24, n25, n26, n27, n28, n46, n47
      , n48, n49, n50, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, 
      n77, n78, n79, n80, n81, n82, n83, n84, n85, n86 : std_logic;

begin
   S_FWAdec <= ( S_FWAdec_1_port, S_FWAdec_0_port );
   S_FWA <= ( S_FWA_1_port, S_FWA_0_port );
   
   U53 : XOR2_X1 port map( A => D2_i(4), B => rB_i(4), Z => n30);
   U55 : XOR2_X1 port map( A => D2_i(4), B => rA_i(4), Z => n61);
   U34 : INV_X1 port map( A => rA_i(0), ZN => n54);
   U33 : INV_X1 port map( A => rA_i(2), ZN => n55);
   U38 : INV_X1 port map( A => rA_i(3), ZN => n57);
   U37 : INV_X1 port map( A => rA_i(1), ZN => n58);
   U41 : INV_X1 port map( A => D3_i(4), ZN => n29);
   U40 : INV_X1 port map( A => rA_i(4), ZN => n60);
   U24 : INV_X1 port map( A => rAdec_i(4), ZN => n45);
   U2 : BUF_X1 port map( A => n9, Z => S_FWB(0));
   U3 : OR3_X1 port map( A1 => n42, A2 => n41, A3 => n40, ZN => n75);
   U4 : NOR3_X2 port map( A1 => n62, A2 => n63, A3 => n8, ZN => S_FWA_0_port);
   U5 : INV_X1 port map( A => D2_i(2), ZN => n1);
   U6 : OR2_X1 port map( A1 => n25, A2 => D3_i(1), ZN => n2);
   U7 : NAND2_X1 port map( A1 => n2, A2 => n26, ZN => n24);
   U8 : OR2_X1 port map( A1 => n18, A2 => D3_i(2), ZN => n3);
   U9 : NAND2_X1 port map( A1 => n3, A2 => n19, ZN => n17);
   U10 : OR3_X1 port map( A1 => n53, A2 => n52, A3 => n51, ZN => n84);
   U11 : NOR2_X1 port map( A1 => n48, A2 => n49, ZN => S_FWAdec_0_port);
   U12 : INV_X1 port map( A => n29, ZN => n5);
   U13 : INV_X1 port map( A => D2_i(1), ZN => n6);
   U14 : INV_X1 port map( A => n79, ZN => n7);
   U15 : NOR2_X1 port map( A1 => S_FWAdec_0_port, A2 => n75, ZN => 
                           S_FWAdec_1_port);
   U16 : INV_X1 port map( A => n31, ZN => n50);
   U17 : AOI21_X1 port map( B1 => n10, B2 => n11, A => n12, ZN => S_FWB(1));
   U18 : INV_X1 port map( A => D3_i(0), ZN => n20);
   U19 : INV_X1 port map( A => rB_i(2), ZN => n18);
   U20 : INV_X1 port map( A => D3_i(0), ZN => n22);
   U21 : INV_X1 port map( A => D3_i(3), ZN => n27);
   U22 : INV_X1 port map( A => rB_i(1), ZN => n25);
   U23 : INV_X1 port map( A => D3_i(3), ZN => n79);
   U25 : INV_X1 port map( A => n28, ZN => n13);
   U26 : INV_X1 port map( A => D3_i(4), ZN => n47);
   U27 : INV_X1 port map( A => n78, ZN => n11);
   U28 : OR2_X1 port map( A1 => n30, A2 => n31, ZN => n78);
   U29 : OR2_X1 port map( A1 => n38, A2 => rB_i(1), ZN => n86);
   U30 : OR2_X1 port map( A1 => n37, A2 => rB_i(3), ZN => n85);
   U31 : OR2_X1 port map( A1 => n34, A2 => rB_i(0), ZN => n82);
   U32 : OR2_X1 port map( A1 => n35, A2 => rB_i(2), ZN => n83);
   U35 : INV_X1 port map( A => D2_i(2), ZN => n35);
   U36 : NOR2_X1 port map( A1 => S_FWA_0_port, A2 => n84, ZN => S_FWA_1_port);
   U39 : INV_X1 port map( A => n81, ZN => n80);
   U42 : INV_X1 port map( A => D3_i(1), ZN => n81);
   U43 : INV_X1 port map( A => n23, ZN => n76);
   U44 : INV_X1 port map( A => D3_i(2), ZN => n23);
   U45 : CLKBUF_X1 port map( A => D3_i(0), Z => n77);
   U46 : OR2_X1 port map( A1 => n61, A2 => n31, ZN => n8);
   U47 : INV_X1 port map( A => D2_i(0), ZN => n34);
   U48 : INV_X1 port map( A => D2_i(1), ZN => n38);
   U49 : INV_X1 port map( A => D2_i(3), ZN => n37);
   U50 : NAND2_X1 port map( A1 => S_mem_W, A2 => S_mem_LOAD_BAR, ZN => n31);
   U51 : INV_X1 port map( A => n74, ZN => n67);
   U52 : OAI22_X1 port map( A1 => n22, A2 => rB_i(0), B1 => n23, B2 => rB_i(2),
                           ZN => n16);
   U54 : NOR3_X1 port map( A1 => n33, A2 => n78, A3 => n32, ZN => n9);
   U56 : NAND3_X1 port map( A1 => n15, A2 => n14, A3 => n13, ZN => n12);
   U57 : NAND2_X1 port map( A1 => n47, A2 => rB_i(4), ZN => n46);
   U58 : NAND2_X1 port map( A1 => n20, A2 => rB_i(0), ZN => n19);
   U59 : NAND2_X1 port map( A1 => n27, A2 => rB_i(3), ZN => n26);
   U60 : OAI211_X1 port map( C1 => n29, C2 => rB_i(4), A => n46, B => S_wb_W, 
                           ZN => n28);
   U61 : NOR2_X1 port map( A1 => n17, A2 => n16, ZN => n15);
   U62 : NOR2_X1 port map( A1 => n33, A2 => n32, ZN => n10);
   U63 : OAI22_X1 port map( A1 => rB_i(1), A2 => n81, B1 => n79, B2 => rB_i(3),
                           ZN => n21);
   U64 : NOR2_X1 port map( A1 => n24, A2 => n21, ZN => n14);
   U65 : NAND3_X1 port map( A1 => n69, A2 => n67, A3 => n68, ZN => n48);
   U66 : NAND2_X1 port map( A1 => n37, A2 => rAdec_i(3), ZN => n72);
   U67 : NAND2_X1 port map( A1 => n72, A2 => n73, ZN => n70);
   U68 : OAI22_X1 port map( A1 => n1, A2 => rAdec_i(2), B1 => rAdec_i(0), B2 =>
                           n34, ZN => n74);
   U69 : NAND2_X1 port map( A1 => n38, A2 => rAdec_i(1), ZN => n73);
   U70 : OAI22_X1 port map( A1 => n37, A2 => rAdec_i(3), B1 => n6, B2 => 
                           rAdec_i(1), ZN => n71);
   U71 : NOR2_X1 port map( A1 => n70, A2 => n71, ZN => n69);
   U72 : NAND2_X1 port map( A1 => n50, A2 => n66, ZN => n49);
   U73 : XNOR2_X1 port map( A => rAdec_i(4), B => D2_i(4), ZN => n66);
   U74 : AOI22_X1 port map( A1 => n1, A2 => rAdec_i(2), B1 => rAdec_i(0), B2 =>
                           n34, ZN => n68);
   U75 : AOI22_X1 port map( A1 => n79, A2 => rAdec_i(3), B1 => rAdec_i(1), B2 
                           => n81, ZN => n44);
   U76 : AOI22_X1 port map( A1 => n22, A2 => rAdec_i(0), B1 => rAdec_i(2), B2 
                           => n23, ZN => n43);
   U77 : OAI221_X1 port map( B1 => n5, B2 => n45, C1 => n29, C2 => rAdec_i(4), 
                           A => S_wb_W, ZN => n40);
   U78 : OAI221_X1 port map( B1 => n79, B2 => rAdec_i(3), C1 => n81, C2 => 
                           rAdec_i(1), A => n44, ZN => n41);
   U79 : OAI221_X1 port map( B1 => n22, B2 => rAdec_i(0), C1 => n23, C2 => 
                           rAdec_i(2), A => n43, ZN => n42);
   U80 : OAI221_X1 port map( B1 => n37, B2 => rA_i(3), C1 => n6, C2 => rA_i(1),
                           A => n65, ZN => n62);
   U81 : AOI22_X1 port map( A1 => n54, A2 => n77, B1 => n76, B2 => n55, ZN => 
                           n56);
   U82 : OAI221_X1 port map( B1 => n34, B2 => rA_i(0), C1 => n1, C2 => rA_i(2),
                           A => n64, ZN => n63);
   U83 : AOI22_X1 port map( A1 => n57, A2 => n7, B1 => n80, B2 => n58, ZN => 
                           n59);
   U84 : AOI22_X1 port map( A1 => n37, A2 => rA_i(3), B1 => rA_i(1), B2 => n6, 
                           ZN => n65);
   U85 : NAND3_X1 port map( A1 => n36, A2 => n83, A3 => n82, ZN => n33);
   U86 : OAI221_X1 port map( B1 => rA_i(4), B2 => n29, C1 => n60, C2 => n5, A 
                           => S_wb_W, ZN => n51);
   U87 : OAI221_X1 port map( B1 => n57, B2 => n7, C1 => n58, C2 => n80, A => 
                           n59, ZN => n52);
   U88 : OAI221_X1 port map( B1 => n54, B2 => n77, C1 => n55, C2 => n76, A => 
                           n56, ZN => n53);
   U89 : AOI22_X1 port map( A1 => n34, A2 => rA_i(0), B1 => rA_i(2), B2 => n35,
                           ZN => n64);
   U90 : NAND3_X1 port map( A1 => n85, A2 => n86, A3 => n39, ZN => n32);
   U91 : AOI22_X1 port map( A1 => n34, A2 => rB_i(0), B1 => rB_i(2), B2 => n35,
                           ZN => n36);
   U92 : AOI22_X1 port map( A1 => n37, A2 => rB_i(3), B1 => n38, B2 => rB_i(1),
                           ZN => n39);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity mem_block is

   port( X_i, LOAD_i : in std_logic_vector (31 downto 0);  W_o : out 
         std_logic_vector (31 downto 0);  S_MUX_MEM_i_BAR : in std_logic);

end mem_block;

architecture SYN_struct of mem_block is

   component mux21_2
      port( IN0, IN1 : in std_logic_vector (31 downto 0);  OUT1 : out 
            std_logic_vector (31 downto 0);  CTRL_BAR : in std_logic);
   end component;

begin
   
   MUXMEM : mux21_2 port map( IN0(31) => X_i(31), IN0(30) => X_i(30), IN0(29) 
                           => X_i(29), IN0(28) => X_i(28), IN0(27) => X_i(27), 
                           IN0(26) => X_i(26), IN0(25) => X_i(25), IN0(24) => 
                           X_i(24), IN0(23) => X_i(23), IN0(22) => X_i(22), 
                           IN0(21) => X_i(21), IN0(20) => X_i(20), IN0(19) => 
                           X_i(19), IN0(18) => X_i(18), IN0(17) => X_i(17), 
                           IN0(16) => X_i(16), IN0(15) => X_i(15), IN0(14) => 
                           X_i(14), IN0(13) => X_i(13), IN0(12) => X_i(12), 
                           IN0(11) => X_i(11), IN0(10) => X_i(10), IN0(9) => 
                           X_i(9), IN0(8) => X_i(8), IN0(7) => X_i(7), IN0(6) 
                           => X_i(6), IN0(5) => X_i(5), IN0(4) => X_i(4), 
                           IN0(3) => X_i(3), IN0(2) => X_i(2), IN0(1) => X_i(1)
                           , IN0(0) => X_i(0), IN1(31) => LOAD_i(31), IN1(30) 
                           => LOAD_i(30), IN1(29) => LOAD_i(29), IN1(28) => 
                           LOAD_i(28), IN1(27) => LOAD_i(27), IN1(26) => 
                           LOAD_i(26), IN1(25) => LOAD_i(25), IN1(24) => 
                           LOAD_i(24), IN1(23) => LOAD_i(23), IN1(22) => 
                           LOAD_i(22), IN1(21) => LOAD_i(21), IN1(20) => 
                           LOAD_i(20), IN1(19) => LOAD_i(19), IN1(18) => 
                           LOAD_i(18), IN1(17) => LOAD_i(17), IN1(16) => 
                           LOAD_i(16), IN1(15) => LOAD_i(15), IN1(14) => 
                           LOAD_i(14), IN1(13) => LOAD_i(13), IN1(12) => 
                           LOAD_i(12), IN1(11) => LOAD_i(11), IN1(10) => 
                           LOAD_i(10), IN1(9) => LOAD_i(9), IN1(8) => LOAD_i(8)
                           , IN1(7) => LOAD_i(7), IN1(6) => LOAD_i(6), IN1(5) 
                           => LOAD_i(5), IN1(4) => LOAD_i(4), IN1(3) => 
                           LOAD_i(3), IN1(2) => LOAD_i(2), IN1(1) => LOAD_i(1),
                           IN1(0) => LOAD_i(0), OUT1(31) => W_o(31), OUT1(30) 
                           => W_o(30), OUT1(29) => W_o(29), OUT1(28) => W_o(28)
                           , OUT1(27) => W_o(27), OUT1(26) => W_o(26), OUT1(25)
                           => W_o(25), OUT1(24) => W_o(24), OUT1(23) => W_o(23)
                           , OUT1(22) => W_o(22), OUT1(21) => W_o(21), OUT1(20)
                           => W_o(20), OUT1(19) => W_o(19), OUT1(18) => W_o(18)
                           , OUT1(17) => W_o(17), OUT1(16) => W_o(16), OUT1(15)
                           => W_o(15), OUT1(14) => W_o(14), OUT1(13) => W_o(13)
                           , OUT1(12) => W_o(12), OUT1(11) => W_o(11), OUT1(10)
                           => W_o(10), OUT1(9) => W_o(9), OUT1(8) => W_o(8), 
                           OUT1(7) => W_o(7), OUT1(6) => W_o(6), OUT1(5) => 
                           W_o(5), OUT1(4) => W_o(4), OUT1(3) => W_o(3), 
                           OUT1(2) => W_o(2), OUT1(1) => W_o(1), OUT1(0) => 
                           W_o(0), CTRL_BAR => S_MUX_MEM_i_BAR);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity mem_regs is

   port( W_i : in std_logic_vector (31 downto 0);  D3_i : in std_logic_vector 
         (4 downto 0);  W_o : out std_logic_vector (31 downto 0);  D3_o : out 
         std_logic_vector (4 downto 0);  clk, rst : in std_logic);

end mem_regs;

architecture SYN_Struct of mem_regs is

   component ff32_SIZE5
      port( D : in std_logic_vector (4 downto 0);  clk, rst : in std_logic;  Q 
            : out std_logic_vector (4 downto 0));
   end component;
   
   component ff32_SIZE32
      port( D : in std_logic_vector (31 downto 0);  clk, rst : in std_logic;  Q
            : out std_logic_vector (31 downto 0));
   end component;

begin
   
   W : ff32_SIZE32 port map( D(31) => W_i(31), D(30) => W_i(30), D(29) => 
                           W_i(29), D(28) => W_i(28), D(27) => W_i(27), D(26) 
                           => W_i(26), D(25) => W_i(25), D(24) => W_i(24), 
                           D(23) => W_i(23), D(22) => W_i(22), D(21) => W_i(21)
                           , D(20) => W_i(20), D(19) => W_i(19), D(18) => 
                           W_i(18), D(17) => W_i(17), D(16) => W_i(16), D(15) 
                           => W_i(15), D(14) => W_i(14), D(13) => W_i(13), 
                           D(12) => W_i(12), D(11) => W_i(11), D(10) => W_i(10)
                           , D(9) => W_i(9), D(8) => W_i(8), D(7) => W_i(7), 
                           D(6) => W_i(6), D(5) => W_i(5), D(4) => W_i(4), D(3)
                           => W_i(3), D(2) => W_i(2), D(1) => W_i(1), D(0) => 
                           W_i(0), clk => clk, rst => rst, Q(31) => W_o(31), 
                           Q(30) => W_o(30), Q(29) => W_o(29), Q(28) => W_o(28)
                           , Q(27) => W_o(27), Q(26) => W_o(26), Q(25) => 
                           W_o(25), Q(24) => W_o(24), Q(23) => W_o(23), Q(22) 
                           => W_o(22), Q(21) => W_o(21), Q(20) => W_o(20), 
                           Q(19) => W_o(19), Q(18) => W_o(18), Q(17) => W_o(17)
                           , Q(16) => W_o(16), Q(15) => W_o(15), Q(14) => 
                           W_o(14), Q(13) => W_o(13), Q(12) => W_o(12), Q(11) 
                           => W_o(11), Q(10) => W_o(10), Q(9) => W_o(9), Q(8) 
                           => W_o(8), Q(7) => W_o(7), Q(6) => W_o(6), Q(5) => 
                           W_o(5), Q(4) => W_o(4), Q(3) => W_o(3), Q(2) => 
                           W_o(2), Q(1) => W_o(1), Q(0) => W_o(0));
   D3 : ff32_SIZE5 port map( D(4) => D3_i(4), D(3) => D3_i(3), D(2) => D3_i(2),
                           D(1) => D3_i(1), D(0) => D3_i(0), clk => clk, rst =>
                           rst, Q(4) => D3_o(4), Q(3) => D3_o(3), Q(2) => 
                           D3_o(2), Q(1) => D3_o(1), Q(0) => D3_o(0));

end SYN_Struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity execute_block is

   port( IMM_i, A_i : in std_logic_vector (31 downto 0);  rB_i, rC_i : in 
         std_logic_vector (4 downto 0);  MUXED_B_i : in std_logic_vector (31 
         downto 0);  S_MUX_ALUIN_i : in std_logic;  FW_X_i, FW_W_i : in 
         std_logic_vector (31 downto 0);  S_FW_A_i, S_FW_B_i : in 
         std_logic_vector (1 downto 0);  muxed_dest : out std_logic_vector (4 
         downto 0);  muxed_B : out std_logic_vector (31 downto 0);  
         S_MUX_DEST_i : in std_logic_vector (1 downto 0);  OP : in 
         std_logic_vector (0 to 4);  ALUW_i : in std_logic_vector (12 downto 0)
         ;  DOUT : out std_logic_vector (31 downto 0);  stall_o : out std_logic
         ;  Clock, Reset : in std_logic);

end execute_block;

architecture SYN_struct of execute_block is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component mux41_MUX_SIZE32_1
      port( IN0, IN1, IN2, IN3 : in std_logic_vector (31 downto 0);  CTRL : in 
            std_logic_vector (1 downto 0);  OUT1 : out std_logic_vector (31 
            downto 0));
   end component;
   
   component mux41_MUX_SIZE32_2
      port( IN0, IN1, IN2, IN3 : in std_logic_vector (31 downto 0);  CTRL : in 
            std_logic_vector (1 downto 0);  OUT1 : out std_logic_vector (31 
            downto 0));
   end component;
   
   component mux41_MUX_SIZE5
      port( IN0, IN1, IN2, IN3 : in std_logic_vector (4 downto 0);  CTRL : in 
            std_logic_vector (1 downto 0);  OUT1 : out std_logic_vector (4 
            downto 0));
   end component;
   
   component real_alu_DATA_SIZE32
      port( IN1, IN2 : in std_logic_vector (31 downto 0);  ALUW_i : in 
            std_logic_vector (12 downto 0);  DOUT : out std_logic_vector (31 
            downto 0);  stall_o : out std_logic;  Clock, Reset : in std_logic);
   end component;
   
   component mux21_3
      port( IN0, IN1 : in std_logic_vector (31 downto 0);  CTRL : in std_logic;
            OUT1 : out std_logic_vector (31 downto 0));
   end component;
   
   signal X_Logic1_port, X_Logic0_port, muxed_B_31_port, muxed_B_30_port, 
      muxed_B_29_port, muxed_B_28_port, muxed_B_27_port, muxed_B_26_port, 
      muxed_B_25_port, muxed_B_24_port, muxed_B_23_port, muxed_B_22_port, 
      muxed_B_21_port, muxed_B_20_port, muxed_B_19_port, muxed_B_18_port, 
      muxed_B_17_port, muxed_B_16_port, muxed_B_15_port, muxed_B_14_port, 
      muxed_B_13_port, muxed_B_12_port, muxed_B_11_port, muxed_B_10_port, 
      muxed_B_9_port, muxed_B_8_port, muxed_B_7_port, muxed_B_6_port, 
      muxed_B_5_port, muxed_B_4_port, muxed_B_3_port, muxed_B_2_port, n5, 
      FWB2alu_31_port, FWB2alu_30_port, FWB2alu_29_port, FWB2alu_28_port, 
      FWB2alu_27_port, FWB2alu_26_port, FWB2alu_25_port, FWB2alu_24_port, 
      FWB2alu_23_port, FWB2alu_22_port, FWB2alu_20_port, FWB2alu_19_port, 
      FWB2alu_18_port, FWB2alu_17_port, FWB2alu_16_port, FWB2alu_15_port, 
      FWB2alu_14_port, FWB2alu_13_port, FWB2alu_12_port, FWB2alu_11_port, 
      FWB2alu_10_port, FWB2alu_9_port, FWB2alu_8_port, FWB2alu_7_port, 
      FWB2alu_6_port, FWB2alu_5_port, FWB2alu_4_port, FWB2alu_3_port, 
      FWB2alu_2_port, FWB2alu_1_port, FWB2alu_0_port, FWA2alu_31_port, 
      FWA2alu_30_port, FWA2alu_29_port, FWA2alu_28_port, FWA2alu_27_port, 
      FWA2alu_26_port, FWA2alu_25_port, FWA2alu_24_port, FWA2alu_23_port, 
      FWA2alu_22_port, FWA2alu_21_port, FWA2alu_20_port, FWA2alu_19_port, 
      FWA2alu_18_port, FWA2alu_17_port, FWA2alu_16_port, FWA2alu_15_port, 
      FWA2alu_14_port, FWA2alu_13_port, FWA2alu_12_port, FWA2alu_11_port, 
      FWA2alu_10_port, FWA2alu_9_port, FWA2alu_8_port, FWA2alu_7_port, 
      FWA2alu_6_port, FWA2alu_5_port, FWA2alu_4_port, FWA2alu_3_port, 
      FWA2alu_2_port, FWA2alu_1_port, FWA2alu_0_port, n1, muxed_B_0_port, n3, 
      muxed_B_1_port : std_logic;

begin
   muxed_B <= ( muxed_B_31_port, muxed_B_30_port, muxed_B_29_port, 
      muxed_B_28_port, muxed_B_27_port, muxed_B_26_port, muxed_B_25_port, 
      muxed_B_24_port, muxed_B_23_port, muxed_B_22_port, muxed_B_21_port, 
      muxed_B_20_port, muxed_B_19_port, muxed_B_18_port, muxed_B_17_port, 
      muxed_B_16_port, muxed_B_15_port, muxed_B_14_port, muxed_B_13_port, 
      muxed_B_12_port, muxed_B_11_port, muxed_B_10_port, muxed_B_9_port, 
      muxed_B_8_port, muxed_B_7_port, muxed_B_6_port, muxed_B_5_port, 
      muxed_B_4_port, muxed_B_3_port, muxed_B_2_port, muxed_B_1_port, 
      muxed_B_0_port );
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   n1 <= '0';
   ALUIN_MUX : mux21_3 port map( IN0(31) => muxed_B_31_port, IN0(30) => 
                           muxed_B_30_port, IN0(29) => muxed_B_29_port, IN0(28)
                           => muxed_B_28_port, IN0(27) => muxed_B_27_port, 
                           IN0(26) => muxed_B_26_port, IN0(25) => 
                           muxed_B_25_port, IN0(24) => muxed_B_24_port, IN0(23)
                           => muxed_B_23_port, IN0(22) => muxed_B_22_port, 
                           IN0(21) => muxed_B_21_port, IN0(20) => 
                           muxed_B_20_port, IN0(19) => muxed_B_19_port, IN0(18)
                           => muxed_B_18_port, IN0(17) => muxed_B_17_port, 
                           IN0(16) => muxed_B_16_port, IN0(15) => 
                           muxed_B_15_port, IN0(14) => muxed_B_14_port, IN0(13)
                           => muxed_B_13_port, IN0(12) => muxed_B_12_port, 
                           IN0(11) => muxed_B_11_port, IN0(10) => 
                           muxed_B_10_port, IN0(9) => muxed_B_9_port, IN0(8) =>
                           muxed_B_8_port, IN0(7) => muxed_B_7_port, IN0(6) => 
                           muxed_B_6_port, IN0(5) => muxed_B_5_port, IN0(4) => 
                           muxed_B_4_port, IN0(3) => muxed_B_3_port, IN0(2) => 
                           muxed_B_2_port, IN0(1) => muxed_B_1_port, IN0(0) => 
                           n5, IN1(31) => IMM_i(31), IN1(30) => IMM_i(30), 
                           IN1(29) => IMM_i(29), IN1(28) => IMM_i(28), IN1(27) 
                           => IMM_i(27), IN1(26) => IMM_i(26), IN1(25) => 
                           IMM_i(25), IN1(24) => IMM_i(24), IN1(23) => 
                           IMM_i(23), IN1(22) => IMM_i(22), IN1(21) => 
                           IMM_i(21), IN1(20) => IMM_i(20), IN1(19) => 
                           IMM_i(19), IN1(18) => IMM_i(18), IN1(17) => 
                           IMM_i(17), IN1(16) => IMM_i(16), IN1(15) => 
                           IMM_i(15), IN1(14) => IMM_i(14), IN1(13) => 
                           IMM_i(13), IN1(12) => IMM_i(12), IN1(11) => 
                           IMM_i(11), IN1(10) => IMM_i(10), IN1(9) => IMM_i(9),
                           IN1(8) => IMM_i(8), IN1(7) => IMM_i(7), IN1(6) => 
                           IMM_i(6), IN1(5) => IMM_i(5), IN1(4) => IMM_i(4), 
                           IN1(3) => IMM_i(3), IN1(2) => IMM_i(2), IN1(1) => 
                           IMM_i(1), IN1(0) => IMM_i(0), CTRL => S_MUX_ALUIN_i,
                           OUT1(31) => FWB2alu_31_port, OUT1(30) => 
                           FWB2alu_30_port, OUT1(29) => FWB2alu_29_port, 
                           OUT1(28) => FWB2alu_28_port, OUT1(27) => 
                           FWB2alu_27_port, OUT1(26) => FWB2alu_26_port, 
                           OUT1(25) => FWB2alu_25_port, OUT1(24) => 
                           FWB2alu_24_port, OUT1(23) => FWB2alu_23_port, 
                           OUT1(22) => FWB2alu_22_port, OUT1(21) => n3, 
                           OUT1(20) => FWB2alu_20_port, OUT1(19) => 
                           FWB2alu_19_port, OUT1(18) => FWB2alu_18_port, 
                           OUT1(17) => FWB2alu_17_port, OUT1(16) => 
                           FWB2alu_16_port, OUT1(15) => FWB2alu_15_port, 
                           OUT1(14) => FWB2alu_14_port, OUT1(13) => 
                           FWB2alu_13_port, OUT1(12) => FWB2alu_12_port, 
                           OUT1(11) => FWB2alu_11_port, OUT1(10) => 
                           FWB2alu_10_port, OUT1(9) => FWB2alu_9_port, OUT1(8) 
                           => FWB2alu_8_port, OUT1(7) => FWB2alu_7_port, 
                           OUT1(6) => FWB2alu_6_port, OUT1(5) => FWB2alu_5_port
                           , OUT1(4) => FWB2alu_4_port, OUT1(3) => 
                           FWB2alu_3_port, OUT1(2) => FWB2alu_2_port, OUT1(1) 
                           => FWB2alu_1_port, OUT1(0) => FWB2alu_0_port);
   ALU : real_alu_DATA_SIZE32 port map( IN1(31) => FWA2alu_31_port, IN1(30) => 
                           FWA2alu_30_port, IN1(29) => FWA2alu_29_port, IN1(28)
                           => FWA2alu_28_port, IN1(27) => FWA2alu_27_port, 
                           IN1(26) => FWA2alu_26_port, IN1(25) => 
                           FWA2alu_25_port, IN1(24) => FWA2alu_24_port, IN1(23)
                           => FWA2alu_23_port, IN1(22) => FWA2alu_22_port, 
                           IN1(21) => FWA2alu_21_port, IN1(20) => 
                           FWA2alu_20_port, IN1(19) => FWA2alu_19_port, IN1(18)
                           => FWA2alu_18_port, IN1(17) => FWA2alu_17_port, 
                           IN1(16) => FWA2alu_16_port, IN1(15) => 
                           FWA2alu_15_port, IN1(14) => FWA2alu_14_port, IN1(13)
                           => FWA2alu_13_port, IN1(12) => FWA2alu_12_port, 
                           IN1(11) => FWA2alu_11_port, IN1(10) => 
                           FWA2alu_10_port, IN1(9) => FWA2alu_9_port, IN1(8) =>
                           FWA2alu_8_port, IN1(7) => FWA2alu_7_port, IN1(6) => 
                           FWA2alu_6_port, IN1(5) => FWA2alu_5_port, IN1(4) => 
                           FWA2alu_4_port, IN1(3) => FWA2alu_3_port, IN1(2) => 
                           FWA2alu_2_port, IN1(1) => FWA2alu_1_port, IN1(0) => 
                           FWA2alu_0_port, IN2(31) => FWB2alu_31_port, IN2(30) 
                           => FWB2alu_30_port, IN2(29) => FWB2alu_29_port, 
                           IN2(28) => FWB2alu_28_port, IN2(27) => 
                           FWB2alu_27_port, IN2(26) => FWB2alu_26_port, IN2(25)
                           => FWB2alu_25_port, IN2(24) => FWB2alu_24_port, 
                           IN2(23) => FWB2alu_23_port, IN2(22) => 
                           FWB2alu_22_port, IN2(21) => n3, IN2(20) => 
                           FWB2alu_20_port, IN2(19) => FWB2alu_19_port, IN2(18)
                           => FWB2alu_18_port, IN2(17) => FWB2alu_17_port, 
                           IN2(16) => FWB2alu_16_port, IN2(15) => 
                           FWB2alu_15_port, IN2(14) => FWB2alu_14_port, IN2(13)
                           => FWB2alu_13_port, IN2(12) => FWB2alu_12_port, 
                           IN2(11) => FWB2alu_11_port, IN2(10) => 
                           FWB2alu_10_port, IN2(9) => FWB2alu_9_port, IN2(8) =>
                           FWB2alu_8_port, IN2(7) => FWB2alu_7_port, IN2(6) => 
                           FWB2alu_6_port, IN2(5) => FWB2alu_5_port, IN2(4) => 
                           FWB2alu_4_port, IN2(3) => FWB2alu_3_port, IN2(2) => 
                           FWB2alu_2_port, IN2(1) => FWB2alu_1_port, IN2(0) => 
                           FWB2alu_0_port, ALUW_i(12) => ALUW_i(12), ALUW_i(11)
                           => ALUW_i(11), ALUW_i(10) => ALUW_i(10), ALUW_i(9) 
                           => ALUW_i(9), ALUW_i(8) => ALUW_i(8), ALUW_i(7) => 
                           ALUW_i(7), ALUW_i(6) => ALUW_i(6), ALUW_i(5) => 
                           ALUW_i(5), ALUW_i(4) => ALUW_i(4), ALUW_i(3) => 
                           ALUW_i(3), ALUW_i(2) => ALUW_i(2), ALUW_i(1) => 
                           ALUW_i(1), ALUW_i(0) => ALUW_i(0), DOUT(31) => 
                           DOUT(31), DOUT(30) => DOUT(30), DOUT(29) => DOUT(29)
                           , DOUT(28) => DOUT(28), DOUT(27) => DOUT(27), 
                           DOUT(26) => DOUT(26), DOUT(25) => DOUT(25), DOUT(24)
                           => DOUT(24), DOUT(23) => DOUT(23), DOUT(22) => 
                           DOUT(22), DOUT(21) => DOUT(21), DOUT(20) => DOUT(20)
                           , DOUT(19) => DOUT(19), DOUT(18) => DOUT(18), 
                           DOUT(17) => DOUT(17), DOUT(16) => DOUT(16), DOUT(15)
                           => DOUT(15), DOUT(14) => DOUT(14), DOUT(13) => 
                           DOUT(13), DOUT(12) => DOUT(12), DOUT(11) => DOUT(11)
                           , DOUT(10) => DOUT(10), DOUT(9) => DOUT(9), DOUT(8) 
                           => DOUT(8), DOUT(7) => DOUT(7), DOUT(6) => DOUT(6), 
                           DOUT(5) => DOUT(5), DOUT(4) => DOUT(4), DOUT(3) => 
                           DOUT(3), DOUT(2) => DOUT(2), DOUT(1) => DOUT(1), 
                           DOUT(0) => DOUT(0), stall_o => stall_o, Clock => 
                           Clock, Reset => Reset);
   MUXDEST : mux41_MUX_SIZE5 port map( IN0(4) => X_Logic0_port, IN0(3) => 
                           X_Logic0_port, IN0(2) => X_Logic0_port, IN0(1) => 
                           X_Logic0_port, IN0(0) => X_Logic0_port, IN1(4) => 
                           rC_i(4), IN1(3) => rC_i(3), IN1(2) => rC_i(2), 
                           IN1(1) => rC_i(1), IN1(0) => rC_i(0), IN2(4) => 
                           rB_i(4), IN2(3) => rB_i(3), IN2(2) => rB_i(2), 
                           IN2(1) => rB_i(1), IN2(0) => rB_i(0), IN3(4) => 
                           X_Logic1_port, IN3(3) => X_Logic1_port, IN3(2) => 
                           X_Logic1_port, IN3(1) => X_Logic1_port, IN3(0) => 
                           X_Logic1_port, CTRL(1) => S_MUX_DEST_i(1), CTRL(0) 
                           => S_MUX_DEST_i(0), OUT1(4) => muxed_dest(4), 
                           OUT1(3) => muxed_dest(3), OUT1(2) => muxed_dest(2), 
                           OUT1(1) => muxed_dest(1), OUT1(0) => muxed_dest(0));
   MUX_FWA : mux41_MUX_SIZE32_2 port map( IN0(31) => A_i(31), IN0(30) => 
                           A_i(30), IN0(29) => A_i(29), IN0(28) => A_i(28), 
                           IN0(27) => A_i(27), IN0(26) => A_i(26), IN0(25) => 
                           A_i(25), IN0(24) => A_i(24), IN0(23) => A_i(23), 
                           IN0(22) => A_i(22), IN0(21) => A_i(21), IN0(20) => 
                           A_i(20), IN0(19) => A_i(19), IN0(18) => A_i(18), 
                           IN0(17) => A_i(17), IN0(16) => A_i(16), IN0(15) => 
                           A_i(15), IN0(14) => A_i(14), IN0(13) => A_i(13), 
                           IN0(12) => A_i(12), IN0(11) => A_i(11), IN0(10) => 
                           A_i(10), IN0(9) => A_i(9), IN0(8) => A_i(8), IN0(7) 
                           => A_i(7), IN0(6) => A_i(6), IN0(5) => A_i(5), 
                           IN0(4) => A_i(4), IN0(3) => A_i(3), IN0(2) => A_i(2)
                           , IN0(1) => A_i(1), IN0(0) => A_i(0), IN1(31) => 
                           FW_X_i(31), IN1(30) => FW_X_i(30), IN1(29) => 
                           FW_X_i(29), IN1(28) => FW_X_i(28), IN1(27) => 
                           FW_X_i(27), IN1(26) => FW_X_i(26), IN1(25) => 
                           FW_X_i(25), IN1(24) => FW_X_i(24), IN1(23) => 
                           FW_X_i(23), IN1(22) => FW_X_i(22), IN1(21) => 
                           FW_X_i(21), IN1(20) => FW_X_i(20), IN1(19) => 
                           FW_X_i(19), IN1(18) => FW_X_i(18), IN1(17) => 
                           FW_X_i(17), IN1(16) => FW_X_i(16), IN1(15) => 
                           FW_X_i(15), IN1(14) => FW_X_i(14), IN1(13) => 
                           FW_X_i(13), IN1(12) => FW_X_i(12), IN1(11) => 
                           FW_X_i(11), IN1(10) => FW_X_i(10), IN1(9) => 
                           FW_X_i(9), IN1(8) => FW_X_i(8), IN1(7) => FW_X_i(7),
                           IN1(6) => FW_X_i(6), IN1(5) => FW_X_i(5), IN1(4) => 
                           FW_X_i(4), IN1(3) => FW_X_i(3), IN1(2) => FW_X_i(2),
                           IN1(1) => FW_X_i(1), IN1(0) => FW_X_i(0), IN2(31) =>
                           FW_W_i(31), IN2(30) => FW_W_i(30), IN2(29) => 
                           FW_W_i(29), IN2(28) => FW_W_i(28), IN2(27) => 
                           FW_W_i(27), IN2(26) => FW_W_i(26), IN2(25) => 
                           FW_W_i(25), IN2(24) => FW_W_i(24), IN2(23) => 
                           FW_W_i(23), IN2(22) => FW_W_i(22), IN2(21) => 
                           FW_W_i(21), IN2(20) => FW_W_i(20), IN2(19) => 
                           FW_W_i(19), IN2(18) => FW_W_i(18), IN2(17) => 
                           FW_W_i(17), IN2(16) => FW_W_i(16), IN2(15) => 
                           FW_W_i(15), IN2(14) => FW_W_i(14), IN2(13) => 
                           FW_W_i(13), IN2(12) => FW_W_i(12), IN2(11) => 
                           FW_W_i(11), IN2(10) => FW_W_i(10), IN2(9) => 
                           FW_W_i(9), IN2(8) => FW_W_i(8), IN2(7) => FW_W_i(7),
                           IN2(6) => FW_W_i(6), IN2(5) => FW_W_i(5), IN2(4) => 
                           FW_W_i(4), IN2(3) => FW_W_i(3), IN2(2) => FW_W_i(2),
                           IN2(1) => FW_W_i(1), IN2(0) => FW_W_i(0), IN3(31) =>
                           n1, IN3(30) => n1, IN3(29) => n1, IN3(28) => n1, 
                           IN3(27) => n1, IN3(26) => n1, IN3(25) => n1, IN3(24)
                           => n1, IN3(23) => n1, IN3(22) => n1, IN3(21) => n1, 
                           IN3(20) => n1, IN3(19) => n1, IN3(18) => n1, IN3(17)
                           => n1, IN3(16) => n1, IN3(15) => n1, IN3(14) => n1, 
                           IN3(13) => n1, IN3(12) => n1, IN3(11) => n1, IN3(10)
                           => n1, IN3(9) => n1, IN3(8) => n1, IN3(7) => n1, 
                           IN3(6) => n1, IN3(5) => n1, IN3(4) => n1, IN3(3) => 
                           n1, IN3(2) => n1, IN3(1) => n1, IN3(0) => n1, 
                           CTRL(1) => S_FW_A_i(1), CTRL(0) => S_FW_A_i(0), 
                           OUT1(31) => FWA2alu_31_port, OUT1(30) => 
                           FWA2alu_30_port, OUT1(29) => FWA2alu_29_port, 
                           OUT1(28) => FWA2alu_28_port, OUT1(27) => 
                           FWA2alu_27_port, OUT1(26) => FWA2alu_26_port, 
                           OUT1(25) => FWA2alu_25_port, OUT1(24) => 
                           FWA2alu_24_port, OUT1(23) => FWA2alu_23_port, 
                           OUT1(22) => FWA2alu_22_port, OUT1(21) => 
                           FWA2alu_21_port, OUT1(20) => FWA2alu_20_port, 
                           OUT1(19) => FWA2alu_19_port, OUT1(18) => 
                           FWA2alu_18_port, OUT1(17) => FWA2alu_17_port, 
                           OUT1(16) => FWA2alu_16_port, OUT1(15) => 
                           FWA2alu_15_port, OUT1(14) => FWA2alu_14_port, 
                           OUT1(13) => FWA2alu_13_port, OUT1(12) => 
                           FWA2alu_12_port, OUT1(11) => FWA2alu_11_port, 
                           OUT1(10) => FWA2alu_10_port, OUT1(9) => 
                           FWA2alu_9_port, OUT1(8) => FWA2alu_8_port, OUT1(7) 
                           => FWA2alu_7_port, OUT1(6) => FWA2alu_6_port, 
                           OUT1(5) => FWA2alu_5_port, OUT1(4) => FWA2alu_4_port
                           , OUT1(3) => FWA2alu_3_port, OUT1(2) => 
                           FWA2alu_2_port, OUT1(1) => FWA2alu_1_port, OUT1(0) 
                           => FWA2alu_0_port);
   MUX_FWB : mux41_MUX_SIZE32_1 port map( IN0(31) => MUXED_B_i(31), IN0(30) => 
                           MUXED_B_i(30), IN0(29) => MUXED_B_i(29), IN0(28) => 
                           MUXED_B_i(28), IN0(27) => MUXED_B_i(27), IN0(26) => 
                           MUXED_B_i(26), IN0(25) => MUXED_B_i(25), IN0(24) => 
                           MUXED_B_i(24), IN0(23) => MUXED_B_i(23), IN0(22) => 
                           MUXED_B_i(22), IN0(21) => MUXED_B_i(21), IN0(20) => 
                           MUXED_B_i(20), IN0(19) => MUXED_B_i(19), IN0(18) => 
                           MUXED_B_i(18), IN0(17) => MUXED_B_i(17), IN0(16) => 
                           MUXED_B_i(16), IN0(15) => MUXED_B_i(15), IN0(14) => 
                           MUXED_B_i(14), IN0(13) => MUXED_B_i(13), IN0(12) => 
                           MUXED_B_i(12), IN0(11) => MUXED_B_i(11), IN0(10) => 
                           MUXED_B_i(10), IN0(9) => MUXED_B_i(9), IN0(8) => 
                           MUXED_B_i(8), IN0(7) => MUXED_B_i(7), IN0(6) => 
                           MUXED_B_i(6), IN0(5) => MUXED_B_i(5), IN0(4) => 
                           MUXED_B_i(4), IN0(3) => MUXED_B_i(3), IN0(2) => 
                           MUXED_B_i(2), IN0(1) => MUXED_B_i(1), IN0(0) => 
                           MUXED_B_i(0), IN1(31) => FW_X_i(31), IN1(30) => 
                           FW_X_i(30), IN1(29) => FW_X_i(29), IN1(28) => 
                           FW_X_i(28), IN1(27) => FW_X_i(27), IN1(26) => 
                           FW_X_i(26), IN1(25) => FW_X_i(25), IN1(24) => 
                           FW_X_i(24), IN1(23) => FW_X_i(23), IN1(22) => 
                           FW_X_i(22), IN1(21) => FW_X_i(21), IN1(20) => 
                           FW_X_i(20), IN1(19) => FW_X_i(19), IN1(18) => 
                           FW_X_i(18), IN1(17) => FW_X_i(17), IN1(16) => 
                           FW_X_i(16), IN1(15) => FW_X_i(15), IN1(14) => 
                           FW_X_i(14), IN1(13) => FW_X_i(13), IN1(12) => 
                           FW_X_i(12), IN1(11) => FW_X_i(11), IN1(10) => 
                           FW_X_i(10), IN1(9) => FW_X_i(9), IN1(8) => FW_X_i(8)
                           , IN1(7) => FW_X_i(7), IN1(6) => FW_X_i(6), IN1(5) 
                           => FW_X_i(5), IN1(4) => FW_X_i(4), IN1(3) => 
                           FW_X_i(3), IN1(2) => FW_X_i(2), IN1(1) => FW_X_i(1),
                           IN1(0) => FW_X_i(0), IN2(31) => FW_W_i(31), IN2(30) 
                           => FW_W_i(30), IN2(29) => FW_W_i(29), IN2(28) => 
                           FW_W_i(28), IN2(27) => FW_W_i(27), IN2(26) => 
                           FW_W_i(26), IN2(25) => FW_W_i(25), IN2(24) => 
                           FW_W_i(24), IN2(23) => FW_W_i(23), IN2(22) => 
                           FW_W_i(22), IN2(21) => FW_W_i(21), IN2(20) => 
                           FW_W_i(20), IN2(19) => FW_W_i(19), IN2(18) => 
                           FW_W_i(18), IN2(17) => FW_W_i(17), IN2(16) => 
                           FW_W_i(16), IN2(15) => FW_W_i(15), IN2(14) => 
                           FW_W_i(14), IN2(13) => FW_W_i(13), IN2(12) => 
                           FW_W_i(12), IN2(11) => FW_W_i(11), IN2(10) => 
                           FW_W_i(10), IN2(9) => FW_W_i(9), IN2(8) => FW_W_i(8)
                           , IN2(7) => FW_W_i(7), IN2(6) => FW_W_i(6), IN2(5) 
                           => FW_W_i(5), IN2(4) => FW_W_i(4), IN2(3) => 
                           FW_W_i(3), IN2(2) => FW_W_i(2), IN2(1) => FW_W_i(1),
                           IN2(0) => FW_W_i(0), IN3(31) => n1, IN3(30) => n1, 
                           IN3(29) => n1, IN3(28) => n1, IN3(27) => n1, IN3(26)
                           => n1, IN3(25) => n1, IN3(24) => n1, IN3(23) => n1, 
                           IN3(22) => n1, IN3(21) => n1, IN3(20) => n1, IN3(19)
                           => n1, IN3(18) => n1, IN3(17) => n1, IN3(16) => n1, 
                           IN3(15) => n1, IN3(14) => n1, IN3(13) => n1, IN3(12)
                           => n1, IN3(11) => n1, IN3(10) => n1, IN3(9) => n1, 
                           IN3(8) => n1, IN3(7) => n1, IN3(6) => n1, IN3(5) => 
                           n1, IN3(4) => n1, IN3(3) => n1, IN3(2) => n1, IN3(1)
                           => n1, IN3(0) => n1, CTRL(1) => S_FW_B_i(1), CTRL(0)
                           => S_FW_B_i(0), OUT1(31) => muxed_B_31_port, 
                           OUT1(30) => muxed_B_30_port, OUT1(29) => 
                           muxed_B_29_port, OUT1(28) => muxed_B_28_port, 
                           OUT1(27) => muxed_B_27_port, OUT1(26) => 
                           muxed_B_26_port, OUT1(25) => muxed_B_25_port, 
                           OUT1(24) => muxed_B_24_port, OUT1(23) => 
                           muxed_B_23_port, OUT1(22) => muxed_B_22_port, 
                           OUT1(21) => muxed_B_21_port, OUT1(20) => 
                           muxed_B_20_port, OUT1(19) => muxed_B_19_port, 
                           OUT1(18) => muxed_B_18_port, OUT1(17) => 
                           muxed_B_17_port, OUT1(16) => muxed_B_16_port, 
                           OUT1(15) => muxed_B_15_port, OUT1(14) => 
                           muxed_B_14_port, OUT1(13) => muxed_B_13_port, 
                           OUT1(12) => muxed_B_12_port, OUT1(11) => 
                           muxed_B_11_port, OUT1(10) => muxed_B_10_port, 
                           OUT1(9) => muxed_B_9_port, OUT1(8) => muxed_B_8_port
                           , OUT1(7) => muxed_B_7_port, OUT1(6) => 
                           muxed_B_6_port, OUT1(5) => muxed_B_5_port, OUT1(4) 
                           => muxed_B_4_port, OUT1(3) => muxed_B_3_port, 
                           OUT1(2) => muxed_B_2_port, OUT1(1) => muxed_B_1_port
                           , OUT1(0) => n5);
   U5 : CLKBUF_X1 port map( A => n5, Z => muxed_B_0_port);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity execute_regs is

   port( X_i, S_i : in std_logic_vector (31 downto 0);  D2_i : in 
         std_logic_vector (4 downto 0);  X_o, S_o : out std_logic_vector (31 
         downto 0);  D2_o : out std_logic_vector (4 downto 0);  stall_i, clk, 
         rst : in std_logic);

end execute_regs;

architecture SYN_struct of execute_regs is

   component ff32_en_SIZE5_1
      port( D : in std_logic_vector (4 downto 0);  en, clk, rst : in std_logic;
            Q : out std_logic_vector (4 downto 0));
   end component;
   
   component ff32_en_SIZE32_2
      port( D : in std_logic_vector (31 downto 0);  en, clk, rst : in std_logic
            ;  Q : out std_logic_vector (31 downto 0));
   end component;
   
   component ff32_en_SIZE32_3
      port( D : in std_logic_vector (31 downto 0);  en, clk, rst : in std_logic
            ;  Q : out std_logic_vector (31 downto 0));
   end component;
   
   signal n3 : std_logic;

begin
   
   X : ff32_en_SIZE32_3 port map( D(31) => X_i(31), D(30) => X_i(30), D(29) => 
                           X_i(29), D(28) => X_i(28), D(27) => X_i(27), D(26) 
                           => X_i(26), D(25) => X_i(25), D(24) => X_i(24), 
                           D(23) => X_i(23), D(22) => X_i(22), D(21) => X_i(21)
                           , D(20) => X_i(20), D(19) => X_i(19), D(18) => 
                           X_i(18), D(17) => X_i(17), D(16) => X_i(16), D(15) 
                           => X_i(15), D(14) => X_i(14), D(13) => X_i(13), 
                           D(12) => X_i(12), D(11) => X_i(11), D(10) => X_i(10)
                           , D(9) => X_i(9), D(8) => X_i(8), D(7) => X_i(7), 
                           D(6) => X_i(6), D(5) => X_i(5), D(4) => X_i(4), D(3)
                           => X_i(3), D(2) => X_i(2), D(1) => X_i(1), D(0) => 
                           X_i(0), en => n3, clk => clk, rst => rst, Q(31) => 
                           X_o(31), Q(30) => X_o(30), Q(29) => X_o(29), Q(28) 
                           => X_o(28), Q(27) => X_o(27), Q(26) => X_o(26), 
                           Q(25) => X_o(25), Q(24) => X_o(24), Q(23) => X_o(23)
                           , Q(22) => X_o(22), Q(21) => X_o(21), Q(20) => 
                           X_o(20), Q(19) => X_o(19), Q(18) => X_o(18), Q(17) 
                           => X_o(17), Q(16) => X_o(16), Q(15) => X_o(15), 
                           Q(14) => X_o(14), Q(13) => X_o(13), Q(12) => X_o(12)
                           , Q(11) => X_o(11), Q(10) => X_o(10), Q(9) => X_o(9)
                           , Q(8) => X_o(8), Q(7) => X_o(7), Q(6) => X_o(6), 
                           Q(5) => X_o(5), Q(4) => X_o(4), Q(3) => X_o(3), Q(2)
                           => X_o(2), Q(1) => X_o(1), Q(0) => X_o(0));
   S : ff32_en_SIZE32_2 port map( D(31) => S_i(31), D(30) => S_i(30), D(29) => 
                           S_i(29), D(28) => S_i(28), D(27) => S_i(27), D(26) 
                           => S_i(26), D(25) => S_i(25), D(24) => S_i(24), 
                           D(23) => S_i(23), D(22) => S_i(22), D(21) => S_i(21)
                           , D(20) => S_i(20), D(19) => S_i(19), D(18) => 
                           S_i(18), D(17) => S_i(17), D(16) => S_i(16), D(15) 
                           => S_i(15), D(14) => S_i(14), D(13) => S_i(13), 
                           D(12) => S_i(12), D(11) => S_i(11), D(10) => S_i(10)
                           , D(9) => S_i(9), D(8) => S_i(8), D(7) => S_i(7), 
                           D(6) => S_i(6), D(5) => S_i(5), D(4) => S_i(4), D(3)
                           => S_i(3), D(2) => S_i(2), D(1) => S_i(1), D(0) => 
                           S_i(0), en => n3, clk => clk, rst => rst, Q(31) => 
                           S_o(31), Q(30) => S_o(30), Q(29) => S_o(29), Q(28) 
                           => S_o(28), Q(27) => S_o(27), Q(26) => S_o(26), 
                           Q(25) => S_o(25), Q(24) => S_o(24), Q(23) => S_o(23)
                           , Q(22) => S_o(22), Q(21) => S_o(21), Q(20) => 
                           S_o(20), Q(19) => S_o(19), Q(18) => S_o(18), Q(17) 
                           => S_o(17), Q(16) => S_o(16), Q(15) => S_o(15), 
                           Q(14) => S_o(14), Q(13) => S_o(13), Q(12) => S_o(12)
                           , Q(11) => S_o(11), Q(10) => S_o(10), Q(9) => S_o(9)
                           , Q(8) => S_o(8), Q(7) => S_o(7), Q(6) => S_o(6), 
                           Q(5) => S_o(5), Q(4) => S_o(4), Q(3) => S_o(3), Q(2)
                           => S_o(2), Q(1) => S_o(1), Q(0) => S_o(0));
   D2 : ff32_en_SIZE5_1 port map( D(4) => D2_i(4), D(3) => D2_i(3), D(2) => 
                           D2_i(2), D(1) => D2_i(1), D(0) => D2_i(0), en => n3,
                           clk => clk, rst => rst, Q(4) => D2_o(4), Q(3) => 
                           D2_o(3), Q(2) => D2_o(2), Q(1) => D2_o(1), Q(0) => 
                           D2_o(0));
   n3 <= '1';

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity decode_regs is

   port( A_i, B_i : in std_logic_vector (31 downto 0);  rA_i, rB_i, rC_i : in 
         std_logic_vector (4 downto 0);  IMM_i : in std_logic_vector (31 downto
         0);  ALUW_i : in std_logic_vector (12 downto 0);  A_o, B_o : out 
         std_logic_vector (31 downto 0);  rA_o, rB_o, rC_o : out 
         std_logic_vector (4 downto 0);  IMM_o : out std_logic_vector (31 
         downto 0);  ALUW_o : out std_logic_vector (12 downto 0);  stall_i, clk
         , rst : in std_logic);

end decode_regs;

architecture SYN_struct of decode_regs is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component ff32_en_SIZE13
      port( D : in std_logic_vector (12 downto 0);  en, clk, rst : in std_logic
            ;  Q : out std_logic_vector (12 downto 0));
   end component;
   
   component ff32_en_SIZE32_4
      port( D : in std_logic_vector (31 downto 0);  en, clk, rst : in std_logic
            ;  Q : out std_logic_vector (31 downto 0));
   end component;
   
   component ff32_en_SIZE5_2
      port( D : in std_logic_vector (4 downto 0);  en, clk, rst : in std_logic;
            Q : out std_logic_vector (4 downto 0));
   end component;
   
   component ff32_en_SIZE5_3
      port( D : in std_logic_vector (4 downto 0);  en, clk, rst : in std_logic;
            Q : out std_logic_vector (4 downto 0));
   end component;
   
   component ff32_en_SIZE5_0
      port( D : in std_logic_vector (4 downto 0);  en, clk, rst : in std_logic;
            Q : out std_logic_vector (4 downto 0));
   end component;
   
   component ff32_en_SIZE32_5
      port( D : in std_logic_vector (31 downto 0);  en, clk, rst : in std_logic
            ;  Q : out std_logic_vector (31 downto 0));
   end component;
   
   component ff32_en_SIZE32_0
      port( D : in std_logic_vector (31 downto 0);  en, clk, rst : in std_logic
            ;  Q : out std_logic_vector (31 downto 0));
   end component;
   
   signal enable : std_logic;

begin
   
   A : ff32_en_SIZE32_0 port map( D(31) => A_i(31), D(30) => A_i(30), D(29) => 
                           A_i(29), D(28) => A_i(28), D(27) => A_i(27), D(26) 
                           => A_i(26), D(25) => A_i(25), D(24) => A_i(24), 
                           D(23) => A_i(23), D(22) => A_i(22), D(21) => A_i(21)
                           , D(20) => A_i(20), D(19) => A_i(19), D(18) => 
                           A_i(18), D(17) => A_i(17), D(16) => A_i(16), D(15) 
                           => A_i(15), D(14) => A_i(14), D(13) => A_i(13), 
                           D(12) => A_i(12), D(11) => A_i(11), D(10) => A_i(10)
                           , D(9) => A_i(9), D(8) => A_i(8), D(7) => A_i(7), 
                           D(6) => A_i(6), D(5) => A_i(5), D(4) => A_i(4), D(3)
                           => A_i(3), D(2) => A_i(2), D(1) => A_i(1), D(0) => 
                           A_i(0), en => enable, clk => clk, rst => rst, Q(31) 
                           => A_o(31), Q(30) => A_o(30), Q(29) => A_o(29), 
                           Q(28) => A_o(28), Q(27) => A_o(27), Q(26) => A_o(26)
                           , Q(25) => A_o(25), Q(24) => A_o(24), Q(23) => 
                           A_o(23), Q(22) => A_o(22), Q(21) => A_o(21), Q(20) 
                           => A_o(20), Q(19) => A_o(19), Q(18) => A_o(18), 
                           Q(17) => A_o(17), Q(16) => A_o(16), Q(15) => A_o(15)
                           , Q(14) => A_o(14), Q(13) => A_o(13), Q(12) => 
                           A_o(12), Q(11) => A_o(11), Q(10) => A_o(10), Q(9) =>
                           A_o(9), Q(8) => A_o(8), Q(7) => A_o(7), Q(6) => 
                           A_o(6), Q(5) => A_o(5), Q(4) => A_o(4), Q(3) => 
                           A_o(3), Q(2) => A_o(2), Q(1) => A_o(1), Q(0) => 
                           A_o(0));
   B : ff32_en_SIZE32_5 port map( D(31) => B_i(31), D(30) => B_i(30), D(29) => 
                           B_i(29), D(28) => B_i(28), D(27) => B_i(27), D(26) 
                           => B_i(26), D(25) => B_i(25), D(24) => B_i(24), 
                           D(23) => B_i(23), D(22) => B_i(22), D(21) => B_i(21)
                           , D(20) => B_i(20), D(19) => B_i(19), D(18) => 
                           B_i(18), D(17) => B_i(17), D(16) => B_i(16), D(15) 
                           => B_i(15), D(14) => B_i(14), D(13) => B_i(13), 
                           D(12) => B_i(12), D(11) => B_i(11), D(10) => B_i(10)
                           , D(9) => B_i(9), D(8) => B_i(8), D(7) => B_i(7), 
                           D(6) => B_i(6), D(5) => B_i(5), D(4) => B_i(4), D(3)
                           => B_i(3), D(2) => B_i(2), D(1) => B_i(1), D(0) => 
                           B_i(0), en => enable, clk => clk, rst => rst, Q(31) 
                           => B_o(31), Q(30) => B_o(30), Q(29) => B_o(29), 
                           Q(28) => B_o(28), Q(27) => B_o(27), Q(26) => B_o(26)
                           , Q(25) => B_o(25), Q(24) => B_o(24), Q(23) => 
                           B_o(23), Q(22) => B_o(22), Q(21) => B_o(21), Q(20) 
                           => B_o(20), Q(19) => B_o(19), Q(18) => B_o(18), 
                           Q(17) => B_o(17), Q(16) => B_o(16), Q(15) => B_o(15)
                           , Q(14) => B_o(14), Q(13) => B_o(13), Q(12) => 
                           B_o(12), Q(11) => B_o(11), Q(10) => B_o(10), Q(9) =>
                           B_o(9), Q(8) => B_o(8), Q(7) => B_o(7), Q(6) => 
                           B_o(6), Q(5) => B_o(5), Q(4) => B_o(4), Q(3) => 
                           B_o(3), Q(2) => B_o(2), Q(1) => B_o(1), Q(0) => 
                           B_o(0));
   rA : ff32_en_SIZE5_0 port map( D(4) => rA_i(4), D(3) => rA_i(3), D(2) => 
                           rA_i(2), D(1) => rA_i(1), D(0) => rA_i(0), en => 
                           enable, clk => clk, rst => rst, Q(4) => rA_o(4), 
                           Q(3) => rA_o(3), Q(2) => rA_o(2), Q(1) => rA_o(1), 
                           Q(0) => rA_o(0));
   rB : ff32_en_SIZE5_3 port map( D(4) => rB_i(4), D(3) => rB_i(3), D(2) => 
                           rB_i(2), D(1) => rB_i(1), D(0) => rB_i(0), en => 
                           enable, clk => clk, rst => rst, Q(4) => rB_o(4), 
                           Q(3) => rB_o(3), Q(2) => rB_o(2), Q(1) => rB_o(1), 
                           Q(0) => rB_o(0));
   rC : ff32_en_SIZE5_2 port map( D(4) => rC_i(4), D(3) => rC_i(3), D(2) => 
                           rC_i(2), D(1) => rC_i(1), D(0) => rC_i(0), en => 
                           enable, clk => clk, rst => rst, Q(4) => rC_o(4), 
                           Q(3) => rC_o(3), Q(2) => rC_o(2), Q(1) => rC_o(1), 
                           Q(0) => rC_o(0));
   IMM : ff32_en_SIZE32_4 port map( D(31) => IMM_i(31), D(30) => IMM_i(30), 
                           D(29) => IMM_i(29), D(28) => IMM_i(28), D(27) => 
                           IMM_i(27), D(26) => IMM_i(26), D(25) => IMM_i(25), 
                           D(24) => IMM_i(24), D(23) => IMM_i(23), D(22) => 
                           IMM_i(22), D(21) => IMM_i(21), D(20) => IMM_i(20), 
                           D(19) => IMM_i(19), D(18) => IMM_i(18), D(17) => 
                           IMM_i(17), D(16) => IMM_i(16), D(15) => IMM_i(15), 
                           D(14) => IMM_i(14), D(13) => IMM_i(13), D(12) => 
                           IMM_i(12), D(11) => IMM_i(11), D(10) => IMM_i(10), 
                           D(9) => IMM_i(9), D(8) => IMM_i(8), D(7) => IMM_i(7)
                           , D(6) => IMM_i(6), D(5) => IMM_i(5), D(4) => 
                           IMM_i(4), D(3) => IMM_i(3), D(2) => IMM_i(2), D(1) 
                           => IMM_i(1), D(0) => IMM_i(0), en => enable, clk => 
                           clk, rst => rst, Q(31) => IMM_o(31), Q(30) => 
                           IMM_o(30), Q(29) => IMM_o(29), Q(28) => IMM_o(28), 
                           Q(27) => IMM_o(27), Q(26) => IMM_o(26), Q(25) => 
                           IMM_o(25), Q(24) => IMM_o(24), Q(23) => IMM_o(23), 
                           Q(22) => IMM_o(22), Q(21) => IMM_o(21), Q(20) => 
                           IMM_o(20), Q(19) => IMM_o(19), Q(18) => IMM_o(18), 
                           Q(17) => IMM_o(17), Q(16) => IMM_o(16), Q(15) => 
                           IMM_o(15), Q(14) => IMM_o(14), Q(13) => IMM_o(13), 
                           Q(12) => IMM_o(12), Q(11) => IMM_o(11), Q(10) => 
                           IMM_o(10), Q(9) => IMM_o(9), Q(8) => IMM_o(8), Q(7) 
                           => IMM_o(7), Q(6) => IMM_o(6), Q(5) => IMM_o(5), 
                           Q(4) => IMM_o(4), Q(3) => IMM_o(3), Q(2) => IMM_o(2)
                           , Q(1) => IMM_o(1), Q(0) => IMM_o(0));
   ALUW : ff32_en_SIZE13 port map( D(12) => ALUW_i(12), D(11) => ALUW_i(11), 
                           D(10) => ALUW_i(10), D(9) => ALUW_i(9), D(8) => 
                           ALUW_i(8), D(7) => ALUW_i(7), D(6) => ALUW_i(6), 
                           D(5) => ALUW_i(5), D(4) => ALUW_i(4), D(3) => 
                           ALUW_i(3), D(2) => ALUW_i(2), D(1) => ALUW_i(1), 
                           D(0) => ALUW_i(0), en => enable, clk => clk, rst => 
                           rst, Q(12) => ALUW_o(12), Q(11) => ALUW_o(11), Q(10)
                           => ALUW_o(10), Q(9) => ALUW_o(9), Q(8) => ALUW_o(8),
                           Q(7) => ALUW_o(7), Q(6) => ALUW_o(6), Q(5) => 
                           ALUW_o(5), Q(4) => ALUW_o(4), Q(3) => ALUW_o(3), 
                           Q(2) => ALUW_o(2), Q(1) => ALUW_o(1), Q(0) => 
                           ALUW_o(0));
   U1 : INV_X1 port map( A => stall_i, ZN => enable);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity dlx_regfile is

   port( Clk, Rst, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, 
         ADD_RD2 : in std_logic_vector (4 downto 0);  DATAIN : in 
         std_logic_vector (31 downto 0);  OUT1, OUT2 : out std_logic_vector (31
         downto 0));

end dlx_regfile;

architecture SYN_A of dlx_regfile is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_dlx_regfile_1
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_dlx_regfile_2
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_dlx_regfile_3
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_dlx_regfile_4
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_dlx_regfile_5
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_dlx_regfile_6
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_dlx_regfile_7
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_dlx_regfile_8
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_dlx_regfile_9
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_dlx_regfile_10
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_dlx_regfile_11
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_dlx_regfile_12
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_dlx_regfile_13
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_dlx_regfile_14
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_dlx_regfile_15
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_dlx_regfile_16
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_dlx_regfile_17
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_dlx_regfile_18
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_dlx_regfile_19
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_dlx_regfile_20
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_dlx_regfile_21
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_dlx_regfile_22
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_dlx_regfile_23
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_dlx_regfile_24
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_dlx_regfile_25
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_dlx_regfile_26
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_dlx_regfile_27
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_dlx_regfile_28
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_dlx_regfile_29
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_dlx_regfile_30
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_dlx_regfile_31
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_dlx_regfile_32
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_dlx_regfile_33
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_dlx_regfile_0
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal N2503, N2567, N2631, N2695, N2759, N2823, N2887, N2951, N3015, N3079,
      N3143, N3207, N3271, N3335, N3399, N3463, N3527, N3591, N3655, N3719, 
      N3783, N3847, N3911, N3975, N4039, N4103, N4167, N4231, N4295, N4359, 
      N4423, N4490, N4492, N4494, N4496, N4498, N4500, N4502, N4504, N4506, 
      N4508, N4510, N4512, N4514, N4516, N4518, N4520, N4522, N4524, N4526, 
      N4528, N4530, N4532, N4534, N4536, N4538, N4540, N4542, N4544, N4546, 
      N4548, N4550, N4552, N4554, N4556, N4558, N4560, N4562, N4564, N4566, 
      N4568, N4570, N4572, N4574, N4576, N4578, N4580, N4582, N4584, N4586, 
      N4588, N4590, N4592, N4594, N4596, N4598, N4600, N4602, N4604, N4606, 
      N4608, N4610, N4612, N4614, N4615, N4616, net3391, net3396, net3401, 
      net3406, net3411, net3416, net3421, net3426, net3431, net3436, net3441, 
      net3446, net3451, net3456, net3461, net3466, net3471, net3476, net3481, 
      net3486, net3491, net3496, net3501, net3506, net3511, net3516, net3521, 
      net3526, net3531, net3536, net3541, net3546, net3551, net3556, n4, n5, n6
      , n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
      n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36
      , n38, n40, n42, n44, n46, n48, n50, n52, n54, n56, n58, n60, n62, n64, 
      n66, n68, n70, n72, n74, n76, n78, n80, n82, n84, n86, n88, n90, n92, n94
      , n96, n98, n1094, n1150, n1172, n1194, n1216, n1238, n1260, n1282, n1304
      , n1326, n1348, n1370, n1392, n1414, n1436, n1458, n1480, n1502, n1524, 
      n1546, n1568, n1590, n1612, n1634, n1656, n1678, n1700, n1722, n1744, 
      n1766, n1788, n1810, n1, n2, n3, n37, n39, n41, n43, n45, n47, n49, n51, 
      n53, n55, n57, n59, n61, n63, n65, n67, n69, n71, n73, n75, n77, n79, n81
      , n83, n85, n87, n89, n91, n93, n95, n97, n99, n100, n101, n102, n103, 
      n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, 
      n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, 
      n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, 
      n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, 
      n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, 
      n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, 
      n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, 
      n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, 
      n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, 
      n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, 
      n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, 
      n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, 
      n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, 
      n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, 
      n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, 
      n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, 
      n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, 
      n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, 
      n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, 
      n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, 
      n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, 
      n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, 
      n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, 
      n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, 
      n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, 
      n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, 
      n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, 
      n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, 
      n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, 
      n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, 
      n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, 
      n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, 
      n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, 
      n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, 
      n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, 
      n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, 
      n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, 
      n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, 
      n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, 
      n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, 
      n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, 
      n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, 
      n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, 
      n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, 
      n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, 
      n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, 
      n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, 
      n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, 
      n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, 
      n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, 
      n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, 
      n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, 
      n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, 
      n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, 
      n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, 
      n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, 
      n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, 
      n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, 
      n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, 
      n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, 
      n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, 
      n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, 
      n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, 
      n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, 
      n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, 
      n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, 
      n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, 
      n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, 
      n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, 
      n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, 
      n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, 
      n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, 
      n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, 
      n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, 
      n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, 
      n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, 
      n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, 
      n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, 
      n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, 
      n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, 
      n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, 
      n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, 
      n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, 
      n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, 
      n1093, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, 
      n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, 
      n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, 
      n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, 
      n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, 
      n1144, n1145, n1146, n1147, n1148, n1149, n1151, n1152, n1153, n1154, 
      n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, 
      n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1173, n1174, n1175, 
      n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, 
      n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1195, n1196, 
      n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, 
      n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1217, 
      n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, 
      n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, 
      n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, 
      n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, 
      n1259, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, 
      n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, 
      n1280, n1281, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, 
      n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, 
      n1301, n1302, n1303, n1305, n1306, n1307, n1308, n1309, n1310, n1311, 
      n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, 
      n1322, n1323, n1324, n1325, n1327, n1328, n1329, n1330, n1331, n1332, 
      n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, 
      n1343, n1344, n1345, n1346, n1347, n1349, n1350, n1351, n1352, n1353, 
      n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, 
      n1364, n1365, n1366, n1367, n1368, n1369, n1371, n1372, n1373, n1374, 
      n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, 
      n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1393, n1394, n1395, 
      n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, 
      n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1415, n1416, 
      n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, 
      n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1437, 
      n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, 
      n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, 
      n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, 
      n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, 
      n1479, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, 
      n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, 
      n1500, n1501, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, 
      n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, 
      n1521, n1522, n1523, n1525, n1526, n1527, n1528, n1529, n1530, n1531, 
      n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, 
      n1542, n1543, n1544, n1545, n1547, n1548, n1549, n1550, n1551, n1552, 
      n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, 
      n1563, n1564, n1565, n1566, n1567, n1569, n1570, n1571, n1572, n1573, 
      n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, 
      n1584, n1585, n1586, n1587, n1588, n1589, n1591, n1592, n1593, n1594, 
      n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, 
      n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1613, n1614, n1615, 
      n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, 
      n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1635, n1636, 
      n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, 
      n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1657, 
      n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, 
      n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, 
      n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, 
      n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, 
      n1699, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, 
      n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, 
      n1720, n1721, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, 
      n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, 
      n1741, n1742, n1743, n1745, n1746, n1747, n1748, n1749, n1750, n1751, 
      n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, 
      n1762, n1763, n1764, n1765, n1767, n1768, n1769, n1770, n1771, n1772, 
      n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, 
      n1783, n1784, n1785, n1786, n1787, n1789, n1790, n1791, n1792, n1793, 
      n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, 
      n1804, n1805, n1806, n1807, n1808, n1809, n1811, n1812, n1813, n1814, 
      n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, 
      n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, 
      n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, 
      n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, 
      n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, 
      n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, 
      n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, 
      n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, 
      n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, 
      n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, 
      n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, 
      n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, 
      n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, 
      n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, 
      n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, 
      n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, 
      n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, 
      n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, 
      n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, 
      n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, 
      n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, 
      n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, 
      n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, 
      n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, 
      n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, 
      n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, 
      n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, 
      n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, 
      n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, 
      n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, 
      n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, 
      n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, 
      n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, 
      n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, 
      n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, 
      n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, 
      n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, 
      n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, 
      n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, 
      n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, 
      n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, 
      n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, 
      n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, 
      n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, 
      n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, 
      n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, 
      n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, 
      n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, 
      n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, 
      n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, 
      n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, 
      n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, 
      n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, 
      n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, 
      n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, 
      n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, 
      n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, 
      n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, 
      n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, 
      n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, 
      n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, 
      n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, 
      n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, 
      n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, 
      n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, 
      n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, 
      n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, 
      n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, 
      n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503_port, n2504
      , n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, 
      n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, 
      n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, 
      n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, 
      n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, 
      n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, 
      n2565, n2566, n2567_port, n2568, n2569, n2570, n2571, n2572, n2573, n2574
      , n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, 
      n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, 
      n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, 
      n2605, n2606, n2607, n2608, n2609, net47689, net47690, net47691, net47692
      , net47693, net47694, net47695, net47696, net47697, net47698, net47699, 
      net47700, net47701, net47702, net47703, net47704, net47705, net47706, 
      net47707, net47708, net47709, net47710, net47711, net47712, net47713, 
      net47714, net47715, net47716, net47717, net47718, net47719, net47720, 
      net47721, net47722, net47723, net47724, net47725, net47726, net47727, 
      net47728, net47729, net47730, net47731, net47732, net47733, net47734, 
      net47735, net47736, net47737, net47738, net47739, net47740, net47741, 
      net47742, net47743, net47744, net47745, net47746, net47747, net47748, 
      net47749, net47750, net47751, net47752, net47753, net47754, net47755, 
      net47756, net47757, net47758, net47759, net47760, net47761, net47762, 
      net47763, net47764, net47765, net47766, net47767, net47768, net47769, 
      net47770, net47771, net47772, net47773, net47774, net47775, net47776, 
      net47777, net47778, net47779, net47780, net47781, net47782, net47783, 
      net47784, net47785, net47786, net47787, net47788, net47789, net47790, 
      net47791, net47792, net47793, net47794, net47795, net47796, net47797, 
      net47798, net47799, net47800, net47801, net47802, net47803, net47804, 
      net47805, net47806, net47807, net47808, net47809, net47810, net47811, 
      net47812, net47813, net47814, net47815, net47816, net47817, net47818, 
      net47819, net47820, net47821, net47822, net47823, net47824, net47825, 
      net47826, net47827, net47828, net47829, net47830, net47831, net47832, 
      net47833, net47834, net47835, net47836, net47837, net47838, net47839, 
      net47840, net47841, net47842, net47843, net47844, net47845, net47846, 
      net47847, net47848, net47849, net47850, net47851, net47852, net47853, 
      net47854, net47855, net47856, net47857, net47858, net47859, net47860, 
      net47861, net47862, net47863, net47864, net47865, net47866, net47867, 
      net47868, net47869, net47870, net47871, net47872, net47873, net47874, 
      net47875, net47876, net47877, net47878, net47879, net47880, net47881, 
      net47882, net47883, net47884, net47885, net47886, net47887, net47888, 
      net47889, net47890, net47891, net47892, net47893, net47894, net47895, 
      net47896, net47897, net47898, net47899, net47900, net47901, net47902, 
      net47903, net47904, net47905, net47906, net47907, net47908, net47909, 
      net47910, net47911, net47912, net47913, net47914, net47915, net47916, 
      net47917, net47918, net47919, net47920, net47921, net47922, net47923, 
      net47924, net47925, net47926, net47927, net47928, net47929, net47930, 
      net47931, net47932, net47933, net47934, net47935, net47936, net47937, 
      net47938, net47939, net47940, net47941, net47942, net47943, net47944, 
      net47945, net47946, net47947, net47948, net47949, net47950, net47951, 
      net47952, net47953, net47954, net47955, net47956, net47957, net47958, 
      net47959, net47960, net47961, net47962, net47963, net47964, net47965, 
      net47966, net47967, net47968, net47969, net47970, net47971, net47972, 
      net47973, net47974, net47975, net47976, net47977, net47978, net47979, 
      net47980, net47981, net47982, net47983, net47984, net47985, net47986, 
      net47987, net47988, net47989, net47990, net47991, net47992, net47993, 
      net47994, net47995, net47996, net47997, net47998, net47999, net48000, 
      net48001, net48002, net48003, net48004, net48005, net48006, net48007, 
      net48008, net48009, net48010, net48011, net48012, net48013, net48014, 
      net48015, net48016, net48017, net48018, net48019, net48020, net48021, 
      net48022, net48023, net48024, net48025, net48026, net48027, net48028, 
      net48029, net48030, net48031, net48032, net48033, net48034, net48035, 
      net48036, net48037, net48038, net48039, net48040, net48041, net48042, 
      net48043, net48044, net48045, net48046, net48047, net48048, net48049, 
      net48050, net48051, net48052, net48053, net48054, net48055, net48056, 
      net48057, net48058, net48059, net48060, net48061, net48062, net48063, 
      net48064, net48065, net48066, net48067, net48068, net48069, net48070, 
      net48071, net48072, net48073, net48074, net48075, net48076, net48077, 
      net48078, net48079, net48080, net48081, net48082, net48083, net48084, 
      net48085, net48086, net48087, net48088, net48089, net48090, net48091, 
      net48092, net48093, net48094, net48095, net48096, net48097, net48098, 
      net48099, net48100, net48101, net48102, net48103, net48104, net48105, 
      net48106, net48107, net48108, net48109, net48110, net48111, net48112, 
      net48113, net48114, net48115, net48116, net48117, net48118, net48119, 
      net48120, net48121, net48122, net48123, net48124, net48125, net48126, 
      net48127, net48128, net48129, net48130, net48131, net48132, net48133, 
      net48134, net48135, net48136, net48137, net48138, net48139, net48140, 
      net48141, net48142, net48143, net48144, net48145, net48146, net48147, 
      net48148, net48149, net48150, net48151, net48152, net48153, net48154, 
      net48155, net48156, net48157, net48158, net48159, net48160, net48161, 
      net48162, net48163, net48164, net48165, net48166, net48167, net48168, 
      net48169, net48170, net48171, net48172, net48173, net48174, net48175, 
      net48176, net48177, net48178, net48179, net48180, net48181, net48182, 
      net48183, net48184, net48185, net48186, net48187, net48188, net48189, 
      net48190, net48191, net48192, net48193, net48194, net48195, net48196, 
      net48197, net48198, net48199, net48200, net48201, net48202, net48203, 
      net48204, net48205, net48206, net48207, net48208, net48209, net48210, 
      net48211, net48212, net48213, net48214, net48215, net48216, net48217, 
      net48218, net48219, net48220, net48221, net48222, net48223, net48224, 
      net48225, net48226, net48227, net48228, net48229, net48230, net48231, 
      net48232, net48233, net48234, net48235, net48236, net48237, net48238, 
      net48239, net48240, net48241, net48242, net48243, net48244, net48245, 
      net48246, net48247, net48248, net48249, net48250, net48251, net48252, 
      net48253, net48254, net48255, net48256, net48257, net48258, net48259, 
      net48260, net48261, net48262, net48263, net48264, net48265, net48266, 
      net48267, net48268, net48269, net48270, net48271, net48272, net48273, 
      net48274, net48275, net48276, net48277, net48278, net48279, net48280, 
      net48281, net48282, net48283, net48284, net48285, net48286, net48287, 
      net48288, net48289, net48290, net48291, net48292, net48293, net48294, 
      net48295, net48296, net48297, net48298, net48299, net48300, net48301, 
      net48302, net48303, net48304, net48305, net48306, net48307, net48308, 
      net48309, net48310, net48311, net48312, net48313, net48314, net48315, 
      net48316, net48317, net48318, net48319, net48320, net48321, net48322, 
      net48323, net48324, net48325, net48326, net48327, net48328, net48329, 
      net48330, net48331, net48332, net48333, net48334, net48335, net48336, 
      net48337, net48338, net48339, net48340, net48341, net48342, net48343, 
      net48344, net48345, net48346, net48347, net48348, net48349, net48350, 
      net48351, net48352, net48353, net48354, net48355, net48356, net48357, 
      net48358, net48359, net48360, net48361, net48362, net48363, net48364, 
      net48365, net48366, net48367, net48368, net48369, net48370, net48371, 
      net48372, net48373, net48374, net48375, net48376, net48377, net48378, 
      net48379, net48380, net48381, net48382, net48383, net48384, net48385, 
      net48386, net48387, net48388, net48389, net48390, net48391, net48392, 
      net48393, net48394, net48395, net48396, net48397, net48398, net48399, 
      net48400, net48401, net48402, net48403, net48404, net48405, net48406, 
      net48407, net48408, net48409, net48410, net48411, net48412, net48413, 
      net48414, net48415, net48416, net48417, net48418, net48419, net48420, 
      net48421, net48422, net48423, net48424, net48425, net48426, net48427, 
      net48428, net48429, net48430, net48431, net48432, net48433, net48434, 
      net48435, net48436, net48437, net48438, net48439, net48440, net48441, 
      net48442, net48443, net48444, net48445, net48446, net48447, net48448, 
      net48449, net48450, net48451, net48452, net48453, net48454, net48455, 
      net48456, net48457, net48458, net48459, net48460, net48461, net48462, 
      net48463, net48464, net48465, net48466, net48467, net48468, net48469, 
      net48470, net48471, net48472, net48473, net48474, net48475, net48476, 
      net48477, net48478, net48479, net48480, net48481, net48482, net48483, 
      net48484, net48485, net48486, net48487, net48488, net48489, net48490, 
      net48491, net48492, net48493, net48494, net48495, net48496, net48497, 
      net48498, net48499, net48500, net48501, net48502, net48503, net48504, 
      net48505, net48506, net48507, net48508, net48509, net48510, net48511, 
      net48512, net48513, net48514, net48515, net48516, net48517, net48518, 
      net48519, net48520, net48521, net48522, net48523, net48524, net48525, 
      net48526, net48527, net48528, net48529, net48530, net48531, net48532, 
      net48533, net48534, net48535, net48536, net48537, net48538, net48539, 
      net48540, net48541, net48542, net48543, net48544, net48545, net48546, 
      net48547, net48548, net48549, net48550, net48551, net48552, net48553, 
      net48554, net48555, net48556, net48557, net48558, net48559, net48560, 
      net48561, net48562, net48563, net48564, net48565, net48566, net48567, 
      net48568, net48569, net48570, net48571, net48572, net48573, net48574, 
      net48575, net48576, net48577, net48578, net48579, net48580, net48581, 
      net48582, net48583, net48584, net48585, net48586, net48587, net48588, 
      net48589, net48590, net48591, net48592, net48593, net48594, net48595, 
      net48596, net48597, net48598, net48599, net48600, net48601, net48602, 
      net48603, net48604, net48605, net48606, net48607, net48608, net48609, 
      net48610, net48611, net48612, net48613, net48614, net48615, net48616, 
      net48617, net48618, net48619, net48620, net48621, net48622, net48623, 
      net48624, net48625, net48626, net48627, net48628, net48629, net48630, 
      net48631, net48632, net48633, net48634, net48635, net48636, net48637, 
      net48638, net48639, net48640, net48641, net48642, net48643, net48644, 
      net48645, net48646, net48647, net48648, net48649, net48650, net48651, 
      net48652, net48653, net48654, net48655, net48656, net48657, net48658, 
      net48659, net48660, net48661, net48662, net48663, net48664, net48665, 
      net48666, net48667, net48668, net48669, net48670, net48671, net48672, 
      net48673, net48674, net48675, net48676, net48677, net48678, net48679, 
      net48680, net48681, net48682, net48683, net48684, net48685, net48686, 
      net48687, net48688, net48689, net48690, net48691, net48692, net48693, 
      net48694, net48695, net48696, net48697, net48698, net48699, net48700, 
      net48701, net48702, net48703, net48704, net48705, net48706, net48707, 
      net48708, net48709, net48710, net48711, net48712 : std_logic;

begin
   
   REGISTERS_reg_0_31_inst : DFF_X1 port map( D => n1094, CK => net3396, Q => 
                           n177, QN => net48712);
   REGISTERS_reg_0_30_inst : DFF_X1 port map( D => n1150, CK => net3396, Q => 
                           n176, QN => net48711);
   REGISTERS_reg_0_29_inst : DFF_X1 port map( D => n1172, CK => net3396, Q => 
                           n174, QN => net48710);
   REGISTERS_reg_0_28_inst : DFF_X1 port map( D => n1194, CK => net3396, Q => 
                           n173, QN => net48709);
   REGISTERS_reg_0_27_inst : DFF_X1 port map( D => n1216, CK => net3396, Q => 
                           n172, QN => net48708);
   REGISTERS_reg_0_26_inst : DFF_X1 port map( D => n1238, CK => net3396, Q => 
                           n171, QN => net48707);
   REGISTERS_reg_0_25_inst : DFF_X1 port map( D => n1260, CK => net3396, Q => 
                           n170, QN => net48706);
   REGISTERS_reg_0_24_inst : DFF_X1 port map( D => n1282, CK => net3396, Q => 
                           n169, QN => net48705);
   REGISTERS_reg_0_23_inst : DFF_X1 port map( D => n1304, CK => net3396, Q => 
                           n168, QN => net48704);
   REGISTERS_reg_0_22_inst : DFF_X1 port map( D => n1326, CK => net3396, Q => 
                           n167, QN => net48703);
   REGISTERS_reg_0_21_inst : DFF_X1 port map( D => n1348, CK => net3396, Q => 
                           n166, QN => net48702);
   REGISTERS_reg_0_20_inst : DFF_X1 port map( D => n1370, CK => net3396, Q => 
                           n165, QN => net48701);
   REGISTERS_reg_0_19_inst : DFF_X1 port map( D => n1392, CK => net3396, Q => 
                           n163, QN => net48700);
   REGISTERS_reg_0_18_inst : DFF_X1 port map( D => n1414, CK => net3396, Q => 
                           n162, QN => net48699);
   REGISTERS_reg_0_17_inst : DFF_X1 port map( D => n1436, CK => net3396, Q => 
                           n161, QN => net48698);
   REGISTERS_reg_0_16_inst : DFF_X1 port map( D => n1458, CK => net3396, Q => 
                           n160, QN => net48697);
   REGISTERS_reg_0_15_inst : DFF_X1 port map( D => n1480, CK => net3396, Q => 
                           n159, QN => net48696);
   REGISTERS_reg_0_14_inst : DFF_X1 port map( D => n1502, CK => net3396, Q => 
                           n158, QN => net48695);
   REGISTERS_reg_0_13_inst : DFF_X1 port map( D => n1524, CK => net3396, Q => 
                           n157, QN => net48694);
   REGISTERS_reg_0_12_inst : DFF_X1 port map( D => n1546, CK => net3396, Q => 
                           n156, QN => net48693);
   REGISTERS_reg_0_11_inst : DFF_X1 port map( D => n1568, CK => net3396, Q => 
                           n155, QN => net48692);
   REGISTERS_reg_0_10_inst : DFF_X1 port map( D => n1590, CK => net3396, Q => 
                           n154, QN => net48691);
   REGISTERS_reg_0_9_inst : DFF_X1 port map( D => n1612, CK => net3396, Q => 
                           n152, QN => net48690);
   REGISTERS_reg_0_8_inst : DFF_X1 port map( D => n1634, CK => net3396, Q => 
                           n151, QN => net48689);
   REGISTERS_reg_0_7_inst : DFF_X1 port map( D => n1656, CK => net3396, Q => 
                           n150, QN => net48688);
   REGISTERS_reg_0_6_inst : DFF_X1 port map( D => n1678, CK => net3396, Q => 
                           n149, QN => net48687);
   REGISTERS_reg_0_5_inst : DFF_X1 port map( D => n1700, CK => net3396, Q => 
                           n148, QN => net48686);
   REGISTERS_reg_0_4_inst : DFF_X1 port map( D => n1722, CK => net3396, Q => 
                           n147, QN => net48685);
   REGISTERS_reg_0_3_inst : DFF_X1 port map( D => n1744, CK => net3396, Q => 
                           n146, QN => net48684);
   REGISTERS_reg_0_2_inst : DFF_X1 port map( D => n1766, CK => net3396, Q => 
                           n145, QN => net48683);
   REGISTERS_reg_0_1_inst : DFF_X1 port map( D => n1788, CK => net3396, Q => 
                           n144, QN => net48682);
   REGISTERS_reg_0_0_inst : DFF_X1 port map( D => n1810, CK => net3396, Q => 
                           n143, QN => net48681);
   REGISTERS_reg_1_31_inst : DFF_X1 port map( D => n1094, CK => net3401, Q => 
                           n141, QN => net48680);
   REGISTERS_reg_1_30_inst : DFF_X1 port map( D => n1150, CK => net3401, Q => 
                           n140, QN => net48679);
   REGISTERS_reg_1_29_inst : DFF_X1 port map( D => n1172, CK => net3401, Q => 
                           n139, QN => net48678);
   REGISTERS_reg_1_28_inst : DFF_X1 port map( D => n1194, CK => net3401, Q => 
                           n138, QN => net48677);
   REGISTERS_reg_1_27_inst : DFF_X1 port map( D => n1216, CK => net3401, Q => 
                           n137, QN => net48676);
   REGISTERS_reg_1_26_inst : DFF_X1 port map( D => n1238, CK => net3401, Q => 
                           n136, QN => net48675);
   REGISTERS_reg_1_25_inst : DFF_X1 port map( D => n1260, CK => net3401, Q => 
                           n135, QN => net48674);
   REGISTERS_reg_1_24_inst : DFF_X1 port map( D => n1282, CK => net3401, Q => 
                           n134, QN => net48673);
   REGISTERS_reg_1_23_inst : DFF_X1 port map( D => n1304, CK => net3401, Q => 
                           n133, QN => net48672);
   REGISTERS_reg_1_22_inst : DFF_X1 port map( D => n1326, CK => net3401, Q => 
                           n132, QN => net48671);
   REGISTERS_reg_1_21_inst : DFF_X1 port map( D => n1348, CK => net3401, Q => 
                           n130, QN => net48670);
   REGISTERS_reg_1_20_inst : DFF_X1 port map( D => n1370, CK => net3401, Q => 
                           n129, QN => net48669);
   REGISTERS_reg_1_19_inst : DFF_X1 port map( D => n1392, CK => net3401, Q => 
                           n128, QN => net48668);
   REGISTERS_reg_1_18_inst : DFF_X1 port map( D => n1414, CK => net3401, Q => 
                           n127, QN => net48667);
   REGISTERS_reg_1_17_inst : DFF_X1 port map( D => n1436, CK => net3401, Q => 
                           n126, QN => net48666);
   REGISTERS_reg_1_16_inst : DFF_X1 port map( D => n1458, CK => net3401, Q => 
                           n125, QN => net48665);
   REGISTERS_reg_1_15_inst : DFF_X1 port map( D => n1480, CK => net3401, Q => 
                           n124, QN => net48664);
   REGISTERS_reg_1_14_inst : DFF_X1 port map( D => n1502, CK => net3401, Q => 
                           n123, QN => net48663);
   REGISTERS_reg_1_13_inst : DFF_X1 port map( D => n1524, CK => net3401, Q => 
                           n122, QN => net48662);
   REGISTERS_reg_1_12_inst : DFF_X1 port map( D => n1546, CK => net3401, Q => 
                           n121, QN => net48661);
   REGISTERS_reg_1_11_inst : DFF_X1 port map( D => n1568, CK => net3401, Q => 
                           n119, QN => net48660);
   REGISTERS_reg_1_10_inst : DFF_X1 port map( D => n1590, CK => net3401, Q => 
                           n118, QN => net48659);
   REGISTERS_reg_1_9_inst : DFF_X1 port map( D => n1612, CK => net3401, Q => 
                           n117, QN => net48658);
   REGISTERS_reg_1_8_inst : DFF_X1 port map( D => n1634, CK => net3401, Q => 
                           n116, QN => net48657);
   REGISTERS_reg_1_7_inst : DFF_X1 port map( D => n1656, CK => net3401, Q => 
                           n115, QN => net48656);
   REGISTERS_reg_1_6_inst : DFF_X1 port map( D => n1678, CK => net3401, Q => 
                           n114, QN => net48655);
   REGISTERS_reg_1_5_inst : DFF_X1 port map( D => n1700, CK => net3401, Q => 
                           n113, QN => net48654);
   REGISTERS_reg_1_4_inst : DFF_X1 port map( D => n1722, CK => net3401, Q => 
                           n112, QN => net48653);
   REGISTERS_reg_1_3_inst : DFF_X1 port map( D => n1744, CK => net3401, Q => 
                           n111, QN => net48652);
   REGISTERS_reg_1_2_inst : DFF_X1 port map( D => n1766, CK => net3401, Q => 
                           n110, QN => net48651);
   REGISTERS_reg_1_1_inst : DFF_X1 port map( D => n1788, CK => net3401, Q => 
                           n108, QN => net48650);
   REGISTERS_reg_1_0_inst : DFF_X1 port map( D => n1810, CK => net3401, Q => 
                           n107, QN => net48649);
   REGISTERS_reg_2_31_inst : DFF_X1 port map( D => n1094, CK => net3406, Q => 
                           n106, QN => net48648);
   REGISTERS_reg_2_30_inst : DFF_X1 port map( D => n1150, CK => net3406, Q => 
                           n105, QN => net48647);
   REGISTERS_reg_2_29_inst : DFF_X1 port map( D => n1172, CK => net3406, Q => 
                           n104, QN => net48646);
   REGISTERS_reg_2_28_inst : DFF_X1 port map( D => n1194, CK => net3406, Q => 
                           n103, QN => net48645);
   REGISTERS_reg_2_27_inst : DFF_X1 port map( D => n1216, CK => net3406, Q => 
                           n102, QN => net48644);
   REGISTERS_reg_2_26_inst : DFF_X1 port map( D => n1238, CK => net3406, Q => 
                           n101, QN => net48643);
   REGISTERS_reg_2_25_inst : DFF_X1 port map( D => n1260, CK => net3406, Q => 
                           n100, QN => net48642);
   REGISTERS_reg_2_24_inst : DFF_X1 port map( D => n1282, CK => net3406, Q => 
                           n99, QN => net48641);
   REGISTERS_reg_2_23_inst : DFF_X1 port map( D => n1304, CK => net3406, Q => 
                           n95, QN => net48640);
   REGISTERS_reg_2_22_inst : DFF_X1 port map( D => n1326, CK => net3406, Q => 
                           n93, QN => net48639);
   REGISTERS_reg_2_21_inst : DFF_X1 port map( D => n1348, CK => net3406, Q => 
                           n91, QN => net48638);
   REGISTERS_reg_2_20_inst : DFF_X1 port map( D => n1370, CK => net3406, Q => 
                           n89, QN => net48637);
   REGISTERS_reg_2_19_inst : DFF_X1 port map( D => n1392, CK => net3406, Q => 
                           n87, QN => net48636);
   REGISTERS_reg_2_18_inst : DFF_X1 port map( D => n1414, CK => net3406, Q => 
                           n85, QN => net48635);
   REGISTERS_reg_2_17_inst : DFF_X1 port map( D => n1436, CK => net3406, Q => 
                           n83, QN => net48634);
   REGISTERS_reg_2_16_inst : DFF_X1 port map( D => n1458, CK => net3406, Q => 
                           n81, QN => net48633);
   REGISTERS_reg_2_15_inst : DFF_X1 port map( D => n1480, CK => net3406, Q => 
                           n79, QN => net48632);
   REGISTERS_reg_2_14_inst : DFF_X1 port map( D => n1502, CK => net3406, Q => 
                           n77, QN => net48631);
   REGISTERS_reg_2_13_inst : DFF_X1 port map( D => n1524, CK => net3406, Q => 
                           n73, QN => net48630);
   REGISTERS_reg_2_12_inst : DFF_X1 port map( D => n1546, CK => net3406, Q => 
                           n71, QN => net48629);
   REGISTERS_reg_2_11_inst : DFF_X1 port map( D => n1568, CK => net3406, Q => 
                           n69, QN => net48628);
   REGISTERS_reg_2_10_inst : DFF_X1 port map( D => n1590, CK => net3406, Q => 
                           n67, QN => net48627);
   REGISTERS_reg_2_9_inst : DFF_X1 port map( D => n1612, CK => net3406, Q => 
                           n65, QN => net48626);
   REGISTERS_reg_2_8_inst : DFF_X1 port map( D => n1634, CK => net3406, Q => 
                           n63, QN => net48625);
   REGISTERS_reg_2_7_inst : DFF_X1 port map( D => n1656, CK => net3406, Q => 
                           n61, QN => net48624);
   REGISTERS_reg_2_6_inst : DFF_X1 port map( D => n1678, CK => net3406, Q => 
                           n59, QN => net48623);
   REGISTERS_reg_2_5_inst : DFF_X1 port map( D => n1700, CK => net3406, Q => 
                           n57, QN => net48622);
   REGISTERS_reg_2_4_inst : DFF_X1 port map( D => n1722, CK => net3406, Q => 
                           n55, QN => net48621);
   REGISTERS_reg_2_3_inst : DFF_X1 port map( D => n1744, CK => net3406, Q => 
                           n1100, QN => net48620);
   REGISTERS_reg_2_2_inst : DFF_X1 port map( D => n1766, CK => net3406, Q => 
                           n1099, QN => net48619);
   REGISTERS_reg_2_1_inst : DFF_X1 port map( D => n1788, CK => net3406, Q => 
                           n1098, QN => net48618);
   REGISTERS_reg_2_0_inst : DFF_X1 port map( D => n1810, CK => net3406, Q => 
                           n1097, QN => net48617);
   REGISTERS_reg_3_31_inst : DFF_X1 port map( D => n1094, CK => net3411, Q => 
                           n1096, QN => net48616);
   REGISTERS_reg_3_30_inst : DFF_X1 port map( D => n1150, CK => net3411, Q => 
                           n1095, QN => net48615);
   REGISTERS_reg_3_29_inst : DFF_X1 port map( D => n1172, CK => net3411, Q => 
                           n1093, QN => net48614);
   REGISTERS_reg_3_28_inst : DFF_X1 port map( D => n1194, CK => net3411, Q => 
                           n1092, QN => net48613);
   REGISTERS_reg_3_27_inst : DFF_X1 port map( D => n1216, CK => net3411, Q => 
                           n1091, QN => net48612);
   REGISTERS_reg_3_26_inst : DFF_X1 port map( D => n1238, CK => net3411, Q => 
                           n1090, QN => net48611);
   REGISTERS_reg_3_25_inst : DFF_X1 port map( D => n1260, CK => net3411, Q => 
                           n1088, QN => net48610);
   REGISTERS_reg_3_24_inst : DFF_X1 port map( D => n1282, CK => net3411, Q => 
                           n1087, QN => net48609);
   REGISTERS_reg_3_23_inst : DFF_X1 port map( D => n1304, CK => net3411, Q => 
                           n1086, QN => net48608);
   REGISTERS_reg_3_22_inst : DFF_X1 port map( D => n1326, CK => net3411, Q => 
                           n1085, QN => net48607);
   REGISTERS_reg_3_21_inst : DFF_X1 port map( D => n1348, CK => net3411, Q => 
                           n1084, QN => net48606);
   REGISTERS_reg_3_20_inst : DFF_X1 port map( D => n1370, CK => net3411, Q => 
                           n1083, QN => net48605);
   REGISTERS_reg_3_19_inst : DFF_X1 port map( D => n1392, CK => net3411, Q => 
                           n1082, QN => net48604);
   REGISTERS_reg_3_18_inst : DFF_X1 port map( D => n1414, CK => net3411, Q => 
                           n1081, QN => net48603);
   REGISTERS_reg_3_17_inst : DFF_X1 port map( D => n1436, CK => net3411, Q => 
                           n1080, QN => net48602);
   REGISTERS_reg_3_16_inst : DFF_X1 port map( D => n1458, CK => net3411, Q => 
                           n1079, QN => net48601);
   REGISTERS_reg_3_15_inst : DFF_X1 port map( D => n1480, CK => net3411, Q => 
                           n1078, QN => net48600);
   REGISTERS_reg_3_14_inst : DFF_X1 port map( D => n1502, CK => net3411, Q => 
                           n1077, QN => net48599);
   REGISTERS_reg_3_13_inst : DFF_X1 port map( D => n1524, CK => net3411, Q => 
                           n1076, QN => net48598);
   REGISTERS_reg_3_12_inst : DFF_X1 port map( D => n1546, CK => net3411, Q => 
                           n1075, QN => net48597);
   REGISTERS_reg_3_11_inst : DFF_X1 port map( D => n1568, CK => net3411, Q => 
                           n1074, QN => net48596);
   REGISTERS_reg_3_10_inst : DFF_X1 port map( D => n1590, CK => net3411, Q => 
                           n1073, QN => net48595);
   REGISTERS_reg_3_9_inst : DFF_X1 port map( D => n1612, CK => net3411, Q => 
                           n1072, QN => net48594);
   REGISTERS_reg_3_8_inst : DFF_X1 port map( D => n1634, CK => net3411, Q => 
                           n1071, QN => net48593);
   REGISTERS_reg_3_7_inst : DFF_X1 port map( D => n1656, CK => net3411, Q => 
                           n1070, QN => net48592);
   REGISTERS_reg_3_6_inst : DFF_X1 port map( D => n1678, CK => net3411, Q => 
                           n1069, QN => net48591);
   REGISTERS_reg_3_5_inst : DFF_X1 port map( D => n1700, CK => net3411, Q => 
                           n1067, QN => net48590);
   REGISTERS_reg_3_4_inst : DFF_X1 port map( D => n1722, CK => net3411, Q => 
                           n1066, QN => net48589);
   REGISTERS_reg_3_3_inst : DFF_X1 port map( D => n1744, CK => net3411, Q => 
                           n1065, QN => net48588);
   REGISTERS_reg_3_2_inst : DFF_X1 port map( D => n1766, CK => net3411, Q => 
                           n1064, QN => net48587);
   REGISTERS_reg_3_1_inst : DFF_X1 port map( D => n1788, CK => net3411, Q => 
                           n1063, QN => net48586);
   REGISTERS_reg_3_0_inst : DFF_X1 port map( D => n1810, CK => net3411, Q => 
                           n1062, QN => net48585);
   REGISTERS_reg_4_31_inst : DFF_X1 port map( D => n1094, CK => net3416, Q => 
                           n1061, QN => net48584);
   REGISTERS_reg_4_30_inst : DFF_X1 port map( D => n1150, CK => net3416, Q => 
                           n1060, QN => net48583);
   REGISTERS_reg_4_29_inst : DFF_X1 port map( D => n1172, CK => net3416, Q => 
                           n1059, QN => net48582);
   REGISTERS_reg_4_28_inst : DFF_X1 port map( D => n1194, CK => net3416, Q => 
                           n1058, QN => net48581);
   REGISTERS_reg_4_27_inst : DFF_X1 port map( D => n1216, CK => net3416, Q => 
                           n1057, QN => net48580);
   REGISTERS_reg_4_26_inst : DFF_X1 port map( D => n1238, CK => net3416, Q => 
                           n1056, QN => net48579);
   REGISTERS_reg_4_25_inst : DFF_X1 port map( D => n1260, CK => net3416, Q => 
                           n1055, QN => net48578);
   REGISTERS_reg_4_24_inst : DFF_X1 port map( D => n1282, CK => net3416, Q => 
                           n1054, QN => net48577);
   REGISTERS_reg_4_23_inst : DFF_X1 port map( D => n1304, CK => net3416, Q => 
                           n1053, QN => net48576);
   REGISTERS_reg_4_22_inst : DFF_X1 port map( D => n1326, CK => net3416, Q => 
                           n1052, QN => net48575);
   REGISTERS_reg_4_21_inst : DFF_X1 port map( D => n1348, CK => net3416, Q => 
                           n1051, QN => net48574);
   REGISTERS_reg_4_20_inst : DFF_X1 port map( D => n1370, CK => net3416, Q => 
                           n1050, QN => net48573);
   REGISTERS_reg_4_19_inst : DFF_X1 port map( D => n1392, CK => net3416, Q => 
                           n1049, QN => net48572);
   REGISTERS_reg_4_18_inst : DFF_X1 port map( D => n1414, CK => net3416, Q => 
                           n1048, QN => net48571);
   REGISTERS_reg_4_17_inst : DFF_X1 port map( D => n1436, CK => net3416, Q => 
                           n1046, QN => net48570);
   REGISTERS_reg_4_16_inst : DFF_X1 port map( D => n1458, CK => net3416, Q => 
                           n1045, QN => net48569);
   REGISTERS_reg_4_15_inst : DFF_X1 port map( D => n1480, CK => net3416, Q => 
                           n1044, QN => net48568);
   REGISTERS_reg_4_14_inst : DFF_X1 port map( D => n1502, CK => net3416, Q => 
                           n1043, QN => net48567);
   REGISTERS_reg_4_13_inst : DFF_X1 port map( D => n1524, CK => net3416, Q => 
                           n1042, QN => net48566);
   REGISTERS_reg_4_12_inst : DFF_X1 port map( D => n1546, CK => net3416, Q => 
                           n1041, QN => net48565);
   REGISTERS_reg_4_11_inst : DFF_X1 port map( D => n1568, CK => net3416, Q => 
                           n1040, QN => net48564);
   REGISTERS_reg_4_10_inst : DFF_X1 port map( D => n1590, CK => net3416, Q => 
                           n1039, QN => net48563);
   REGISTERS_reg_4_9_inst : DFF_X1 port map( D => n1612, CK => net3416, Q => 
                           n1038, QN => net48562);
   REGISTERS_reg_4_8_inst : DFF_X1 port map( D => n1634, CK => net3416, Q => 
                           n1037, QN => net48561);
   REGISTERS_reg_4_7_inst : DFF_X1 port map( D => n1656, CK => net3416, Q => 
                           n1036, QN => net48560);
   REGISTERS_reg_4_6_inst : DFF_X1 port map( D => n1678, CK => net3416, Q => 
                           n1035, QN => net48559);
   REGISTERS_reg_4_5_inst : DFF_X1 port map( D => n1700, CK => net3416, Q => 
                           n1034, QN => net48558);
   REGISTERS_reg_4_4_inst : DFF_X1 port map( D => n1722, CK => net3416, Q => 
                           n1033, QN => net48557);
   REGISTERS_reg_4_3_inst : DFF_X1 port map( D => n1744, CK => net3416, Q => 
                           n1032, QN => net48556);
   REGISTERS_reg_4_2_inst : DFF_X1 port map( D => n1766, CK => net3416, Q => 
                           n1031, QN => net48555);
   REGISTERS_reg_4_1_inst : DFF_X1 port map( D => n1788, CK => net3416, Q => 
                           n1030, QN => net48554);
   REGISTERS_reg_4_0_inst : DFF_X1 port map( D => n1810, CK => net3416, Q => 
                           n1029, QN => net48553);
   REGISTERS_reg_5_31_inst : DFF_X1 port map( D => n1094, CK => net3421, Q => 
                           n1028, QN => net48552);
   REGISTERS_reg_5_30_inst : DFF_X1 port map( D => n1150, CK => net3421, Q => 
                           n1027, QN => net48551);
   REGISTERS_reg_5_29_inst : DFF_X1 port map( D => n1172, CK => net3421, Q => 
                           n1025, QN => net48550);
   REGISTERS_reg_5_28_inst : DFF_X1 port map( D => n1194, CK => net3421, Q => 
                           n1024, QN => net48549);
   REGISTERS_reg_5_27_inst : DFF_X1 port map( D => n1216, CK => net3421, Q => 
                           n1023, QN => net48548);
   REGISTERS_reg_5_26_inst : DFF_X1 port map( D => n1238, CK => net3421, Q => 
                           n1022, QN => net48547);
   REGISTERS_reg_5_25_inst : DFF_X1 port map( D => n1260, CK => net3421, Q => 
                           n1021, QN => net48546);
   REGISTERS_reg_5_24_inst : DFF_X1 port map( D => n1282, CK => net3421, Q => 
                           n1020, QN => net48545);
   REGISTERS_reg_5_23_inst : DFF_X1 port map( D => n1304, CK => net3421, Q => 
                           n1019, QN => net48544);
   REGISTERS_reg_5_22_inst : DFF_X1 port map( D => n1326, CK => net3421, Q => 
                           n1018, QN => net48543);
   REGISTERS_reg_5_21_inst : DFF_X1 port map( D => n1348, CK => net3421, Q => 
                           n1017, QN => net48542);
   REGISTERS_reg_5_20_inst : DFF_X1 port map( D => n1370, CK => net3421, Q => 
                           n1016, QN => net48541);
   REGISTERS_reg_5_19_inst : DFF_X1 port map( D => n1392, CK => net3421, Q => 
                           n1015, QN => net48540);
   REGISTERS_reg_5_18_inst : DFF_X1 port map( D => n1414, CK => net3421, Q => 
                           n1014, QN => net48539);
   REGISTERS_reg_5_17_inst : DFF_X1 port map( D => n1436, CK => net3421, Q => 
                           n1013, QN => net48538);
   REGISTERS_reg_5_16_inst : DFF_X1 port map( D => n1458, CK => net3421, Q => 
                           n1012, QN => net48537);
   REGISTERS_reg_5_15_inst : DFF_X1 port map( D => n1480, CK => net3421, Q => 
                           n1011, QN => net48536);
   REGISTERS_reg_5_14_inst : DFF_X1 port map( D => n1502, CK => net3421, Q => 
                           n1010, QN => net48535);
   REGISTERS_reg_5_13_inst : DFF_X1 port map( D => n1524, CK => net3421, Q => 
                           n1009, QN => net48534);
   REGISTERS_reg_5_12_inst : DFF_X1 port map( D => n1546, CK => net3421, Q => 
                           n1008, QN => net48533);
   REGISTERS_reg_5_11_inst : DFF_X1 port map( D => n1568, CK => net3421, Q => 
                           n1007, QN => net48532);
   REGISTERS_reg_5_10_inst : DFF_X1 port map( D => n1590, CK => net3421, Q => 
                           n1006, QN => net48531);
   REGISTERS_reg_5_9_inst : DFF_X1 port map( D => n1612, CK => net3421, Q => 
                           n1004, QN => net48530);
   REGISTERS_reg_5_8_inst : DFF_X1 port map( D => n1634, CK => net3421, Q => 
                           n1003, QN => net48529);
   REGISTERS_reg_5_7_inst : DFF_X1 port map( D => n1656, CK => net3421, Q => 
                           n1002, QN => net48528);
   REGISTERS_reg_5_6_inst : DFF_X1 port map( D => n1678, CK => net3421, Q => 
                           n1001, QN => net48527);
   REGISTERS_reg_5_5_inst : DFF_X1 port map( D => n1700, CK => net3421, Q => 
                           n1000, QN => net48526);
   REGISTERS_reg_5_4_inst : DFF_X1 port map( D => n1722, CK => net3421, Q => 
                           n999, QN => net48525);
   REGISTERS_reg_5_3_inst : DFF_X1 port map( D => n1744, CK => net3421, Q => 
                           n998, QN => net48524);
   REGISTERS_reg_5_2_inst : DFF_X1 port map( D => n1766, CK => net3421, Q => 
                           n997, QN => net48523);
   REGISTERS_reg_5_1_inst : DFF_X1 port map( D => n1788, CK => net3421, Q => 
                           n996, QN => net48522);
   REGISTERS_reg_5_0_inst : DFF_X1 port map( D => n1810, CK => net3421, Q => 
                           n995, QN => net48521);
   REGISTERS_reg_6_31_inst : DFF_X1 port map( D => n1094, CK => net3426, Q => 
                           n994, QN => net48520);
   REGISTERS_reg_6_30_inst : DFF_X1 port map( D => n1150, CK => net3426, Q => 
                           n993, QN => net48519);
   REGISTERS_reg_6_29_inst : DFF_X1 port map( D => n1172, CK => net3426, Q => 
                           n992, QN => net48518);
   REGISTERS_reg_6_28_inst : DFF_X1 port map( D => n1194, CK => net3426, Q => 
                           n991, QN => net48517);
   REGISTERS_reg_6_27_inst : DFF_X1 port map( D => n1216, CK => net3426, Q => 
                           n990, QN => net48516);
   REGISTERS_reg_6_26_inst : DFF_X1 port map( D => n1238, CK => net3426, Q => 
                           n989, QN => net48515);
   REGISTERS_reg_6_25_inst : DFF_X1 port map( D => n1260, CK => net3426, Q => 
                           n988, QN => net48514);
   REGISTERS_reg_6_24_inst : DFF_X1 port map( D => n1282, CK => net3426, Q => 
                           n987, QN => net48513);
   REGISTERS_reg_6_23_inst : DFF_X1 port map( D => n1304, CK => net3426, Q => 
                           n986, QN => net48512);
   REGISTERS_reg_6_22_inst : DFF_X1 port map( D => n1326, CK => net3426, Q => 
                           n985, QN => net48511);
   REGISTERS_reg_6_21_inst : DFF_X1 port map( D => n1348, CK => net3426, Q => 
                           n983, QN => net48510);
   REGISTERS_reg_6_20_inst : DFF_X1 port map( D => n1370, CK => net3426, Q => 
                           n982, QN => net48509);
   REGISTERS_reg_6_19_inst : DFF_X1 port map( D => n1392, CK => net3426, Q => 
                           n981, QN => net48508);
   REGISTERS_reg_6_18_inst : DFF_X1 port map( D => n1414, CK => net3426, Q => 
                           n980, QN => net48507);
   REGISTERS_reg_6_17_inst : DFF_X1 port map( D => n1436, CK => net3426, Q => 
                           n979, QN => net48506);
   REGISTERS_reg_6_16_inst : DFF_X1 port map( D => n1458, CK => net3426, Q => 
                           n978, QN => net48505);
   REGISTERS_reg_6_15_inst : DFF_X1 port map( D => n1480, CK => net3426, Q => 
                           n977, QN => net48504);
   REGISTERS_reg_6_14_inst : DFF_X1 port map( D => n1502, CK => net3426, Q => 
                           n976, QN => net48503);
   REGISTERS_reg_6_13_inst : DFF_X1 port map( D => n1524, CK => net3426, Q => 
                           n975, QN => net48502);
   REGISTERS_reg_6_12_inst : DFF_X1 port map( D => n1546, CK => net3426, Q => 
                           n974, QN => net48501);
   REGISTERS_reg_6_11_inst : DFF_X1 port map( D => n1568, CK => net3426, Q => 
                           n973, QN => net48500);
   REGISTERS_reg_6_10_inst : DFF_X1 port map( D => n1590, CK => net3426, Q => 
                           n972, QN => net48499);
   REGISTERS_reg_6_9_inst : DFF_X1 port map( D => n1612, CK => net3426, Q => 
                           n971, QN => net48498);
   REGISTERS_reg_6_8_inst : DFF_X1 port map( D => n1634, CK => net3426, Q => 
                           n970, QN => net48497);
   REGISTERS_reg_6_7_inst : DFF_X1 port map( D => n1656, CK => net3426, Q => 
                           n969, QN => net48496);
   REGISTERS_reg_6_6_inst : DFF_X1 port map( D => n1678, CK => net3426, Q => 
                           n968, QN => net48495);
   REGISTERS_reg_6_5_inst : DFF_X1 port map( D => n1700, CK => net3426, Q => 
                           n967, QN => net48494);
   REGISTERS_reg_6_4_inst : DFF_X1 port map( D => n1722, CK => net3426, Q => 
                           n966, QN => net48493);
   REGISTERS_reg_6_3_inst : DFF_X1 port map( D => n1744, CK => net3426, Q => 
                           n965, QN => net48492);
   REGISTERS_reg_6_2_inst : DFF_X1 port map( D => n1766, CK => net3426, Q => 
                           n964, QN => net48491);
   REGISTERS_reg_6_1_inst : DFF_X1 port map( D => n1788, CK => net3426, Q => 
                           n962, QN => net48490);
   REGISTERS_reg_6_0_inst : DFF_X1 port map( D => n1810, CK => net3426, Q => 
                           n961, QN => net48489);
   REGISTERS_reg_7_31_inst : DFF_X1 port map( D => n1094, CK => net3431, Q => 
                           n960, QN => net48488);
   REGISTERS_reg_7_30_inst : DFF_X1 port map( D => n1150, CK => net3431, Q => 
                           n959, QN => net48487);
   REGISTERS_reg_7_29_inst : DFF_X1 port map( D => n1172, CK => net3431, Q => 
                           n958, QN => net48486);
   REGISTERS_reg_7_28_inst : DFF_X1 port map( D => n1194, CK => net3431, Q => 
                           n957, QN => net48485);
   REGISTERS_reg_7_27_inst : DFF_X1 port map( D => n1216, CK => net3431, Q => 
                           n956, QN => net48484);
   REGISTERS_reg_7_26_inst : DFF_X1 port map( D => n1238, CK => net3431, Q => 
                           n955, QN => net48483);
   REGISTERS_reg_7_25_inst : DFF_X1 port map( D => n1260, CK => net3431, Q => 
                           n954, QN => net48482);
   REGISTERS_reg_7_24_inst : DFF_X1 port map( D => n1282, CK => net3431, Q => 
                           n953, QN => net48481);
   REGISTERS_reg_7_23_inst : DFF_X1 port map( D => n1304, CK => net3431, Q => 
                           n952, QN => net48480);
   REGISTERS_reg_7_22_inst : DFF_X1 port map( D => n1326, CK => net3431, Q => 
                           n951, QN => net48479);
   REGISTERS_reg_7_21_inst : DFF_X1 port map( D => n1348, CK => net3431, Q => 
                           n950, QN => net48478);
   REGISTERS_reg_7_20_inst : DFF_X1 port map( D => n1370, CK => net3431, Q => 
                           n949, QN => net48477);
   REGISTERS_reg_7_19_inst : DFF_X1 port map( D => n1392, CK => net3431, Q => 
                           n948, QN => net48476);
   REGISTERS_reg_7_18_inst : DFF_X1 port map( D => n1414, CK => net3431, Q => 
                           n947, QN => net48475);
   REGISTERS_reg_7_17_inst : DFF_X1 port map( D => n1436, CK => net3431, Q => 
                           n946, QN => net48474);
   REGISTERS_reg_7_16_inst : DFF_X1 port map( D => n1458, CK => net3431, Q => 
                           n945, QN => net48473);
   REGISTERS_reg_7_15_inst : DFF_X1 port map( D => n1480, CK => net3431, Q => 
                           n944, QN => net48472);
   REGISTERS_reg_7_14_inst : DFF_X1 port map( D => n1502, CK => net3431, Q => 
                           n943, QN => net48471);
   REGISTERS_reg_7_13_inst : DFF_X1 port map( D => n1524, CK => net3431, Q => 
                           n941, QN => net48470);
   REGISTERS_reg_7_12_inst : DFF_X1 port map( D => n1546, CK => net3431, Q => 
                           n940, QN => net48469);
   REGISTERS_reg_7_11_inst : DFF_X1 port map( D => n1568, CK => net3431, Q => 
                           n939, QN => net48468);
   REGISTERS_reg_7_10_inst : DFF_X1 port map( D => n1590, CK => net3431, Q => 
                           n938, QN => net48467);
   REGISTERS_reg_7_9_inst : DFF_X1 port map( D => n1612, CK => net3431, Q => 
                           n937, QN => net48466);
   REGISTERS_reg_7_8_inst : DFF_X1 port map( D => n1634, CK => net3431, Q => 
                           n936, QN => net48465);
   REGISTERS_reg_7_7_inst : DFF_X1 port map( D => n1656, CK => net3431, Q => 
                           n935, QN => net48464);
   REGISTERS_reg_7_6_inst : DFF_X1 port map( D => n1678, CK => net3431, Q => 
                           n934, QN => net48463);
   REGISTERS_reg_7_5_inst : DFF_X1 port map( D => n1700, CK => net3431, Q => 
                           n933, QN => net48462);
   REGISTERS_reg_7_4_inst : DFF_X1 port map( D => n1722, CK => net3431, Q => 
                           n932, QN => net48461);
   REGISTERS_reg_7_3_inst : DFF_X1 port map( D => n1744, CK => net3431, Q => 
                           n931, QN => net48460);
   REGISTERS_reg_7_2_inst : DFF_X1 port map( D => n1766, CK => net3431, Q => 
                           n930, QN => net48459);
   REGISTERS_reg_7_1_inst : DFF_X1 port map( D => n1788, CK => net3431, Q => 
                           n929, QN => net48458);
   REGISTERS_reg_7_0_inst : DFF_X1 port map( D => n1810, CK => net3431, Q => 
                           n928, QN => net48457);
   REGISTERS_reg_8_31_inst : DFF_X1 port map( D => n1094, CK => net3436, Q => 
                           n927, QN => net48456);
   REGISTERS_reg_8_30_inst : DFF_X1 port map( D => n1150, CK => net3436, Q => 
                           n926, QN => net48455);
   REGISTERS_reg_8_29_inst : DFF_X1 port map( D => n1172, CK => net3436, Q => 
                           n925, QN => net48454);
   REGISTERS_reg_8_28_inst : DFF_X1 port map( D => n1194, CK => net3436, Q => 
                           n924, QN => net48453);
   REGISTERS_reg_8_27_inst : DFF_X1 port map( D => n1216, CK => net3436, Q => 
                           n923, QN => net48452);
   REGISTERS_reg_8_26_inst : DFF_X1 port map( D => n1238, CK => net3436, Q => 
                           n922, QN => net48451);
   REGISTERS_reg_8_25_inst : DFF_X1 port map( D => n1260, CK => net3436, Q => 
                           n920, QN => net48450);
   REGISTERS_reg_8_24_inst : DFF_X1 port map( D => n1282, CK => net3436, Q => 
                           n919, QN => net48449);
   REGISTERS_reg_8_23_inst : DFF_X1 port map( D => n1304, CK => net3436, Q => 
                           n918, QN => net48448);
   REGISTERS_reg_8_22_inst : DFF_X1 port map( D => n1326, CK => net3436, Q => 
                           n917, QN => net48447);
   REGISTERS_reg_8_21_inst : DFF_X1 port map( D => n1348, CK => net3436, Q => 
                           n916, QN => net48446);
   REGISTERS_reg_8_20_inst : DFF_X1 port map( D => n1370, CK => net3436, Q => 
                           n915, QN => net48445);
   REGISTERS_reg_8_19_inst : DFF_X1 port map( D => n1392, CK => net3436, Q => 
                           n914, QN => net48444);
   REGISTERS_reg_8_18_inst : DFF_X1 port map( D => n1414, CK => net3436, Q => 
                           n913, QN => net48443);
   REGISTERS_reg_8_17_inst : DFF_X1 port map( D => n1436, CK => net3436, Q => 
                           n912, QN => net48442);
   REGISTERS_reg_8_16_inst : DFF_X1 port map( D => n1458, CK => net3436, Q => 
                           n911, QN => net48441);
   REGISTERS_reg_8_15_inst : DFF_X1 port map( D => n1480, CK => net3436, Q => 
                           n910, QN => net48440);
   REGISTERS_reg_8_14_inst : DFF_X1 port map( D => n1502, CK => net3436, Q => 
                           n909, QN => net48439);
   REGISTERS_reg_8_13_inst : DFF_X1 port map( D => n1524, CK => net3436, Q => 
                           n908, QN => net48438);
   REGISTERS_reg_8_12_inst : DFF_X1 port map( D => n1546, CK => net3436, Q => 
                           n907, QN => net48437);
   REGISTERS_reg_8_11_inst : DFF_X1 port map( D => n1568, CK => net3436, Q => 
                           n906, QN => net48436);
   REGISTERS_reg_8_10_inst : DFF_X1 port map( D => n1590, CK => net3436, Q => 
                           n905, QN => net48435);
   REGISTERS_reg_8_9_inst : DFF_X1 port map( D => n1612, CK => net3436, Q => 
                           n904, QN => net48434);
   REGISTERS_reg_8_8_inst : DFF_X1 port map( D => n1634, CK => net3436, Q => 
                           n903, QN => net48433);
   REGISTERS_reg_8_7_inst : DFF_X1 port map( D => n1656, CK => net3436, Q => 
                           n902, QN => net48432);
   REGISTERS_reg_8_6_inst : DFF_X1 port map( D => n1678, CK => net3436, Q => 
                           n901, QN => net48431);
   REGISTERS_reg_8_5_inst : DFF_X1 port map( D => n1700, CK => net3436, Q => 
                           n899, QN => net48430);
   REGISTERS_reg_8_4_inst : DFF_X1 port map( D => n1722, CK => net3436, Q => 
                           n898, QN => net48429);
   REGISTERS_reg_8_3_inst : DFF_X1 port map( D => n1744, CK => net3436, Q => 
                           n897, QN => net48428);
   REGISTERS_reg_8_2_inst : DFF_X1 port map( D => n1766, CK => net3436, Q => 
                           n896, QN => net48427);
   REGISTERS_reg_8_1_inst : DFF_X1 port map( D => n1788, CK => net3436, Q => 
                           n895, QN => net48426);
   REGISTERS_reg_8_0_inst : DFF_X1 port map( D => n1810, CK => net3436, Q => 
                           n894, QN => net48425);
   REGISTERS_reg_9_31_inst : DFF_X1 port map( D => n1094, CK => net3441, Q => 
                           n893, QN => net48424);
   REGISTERS_reg_9_30_inst : DFF_X1 port map( D => n1150, CK => net3441, Q => 
                           n892, QN => net48423);
   REGISTERS_reg_9_29_inst : DFF_X1 port map( D => n1172, CK => net3441, Q => 
                           n891, QN => net48422);
   REGISTERS_reg_9_28_inst : DFF_X1 port map( D => n1194, CK => net3441, Q => 
                           n890, QN => net48421);
   REGISTERS_reg_9_27_inst : DFF_X1 port map( D => n1216, CK => net3441, Q => 
                           n889, QN => net48420);
   REGISTERS_reg_9_26_inst : DFF_X1 port map( D => n1238, CK => net3441, Q => 
                           n888, QN => net48419);
   REGISTERS_reg_9_25_inst : DFF_X1 port map( D => n1260, CK => net3441, Q => 
                           n887, QN => net48418);
   REGISTERS_reg_9_24_inst : DFF_X1 port map( D => n1282, CK => net3441, Q => 
                           n886, QN => net48417);
   REGISTERS_reg_9_23_inst : DFF_X1 port map( D => n1304, CK => net3441, Q => 
                           n885, QN => net48416);
   REGISTERS_reg_9_22_inst : DFF_X1 port map( D => n1326, CK => net3441, Q => 
                           n884, QN => net48415);
   REGISTERS_reg_9_21_inst : DFF_X1 port map( D => n1348, CK => net3441, Q => 
                           n883, QN => net48414);
   REGISTERS_reg_9_20_inst : DFF_X1 port map( D => n1370, CK => net3441, Q => 
                           n882, QN => net48413);
   REGISTERS_reg_9_19_inst : DFF_X1 port map( D => n1392, CK => net3441, Q => 
                           n881, QN => net48412);
   REGISTERS_reg_9_18_inst : DFF_X1 port map( D => n1414, CK => net3441, Q => 
                           n880, QN => net48411);
   REGISTERS_reg_9_17_inst : DFF_X1 port map( D => n1436, CK => net3441, Q => 
                           n878, QN => net48410);
   REGISTERS_reg_9_16_inst : DFF_X1 port map( D => n1458, CK => net3441, Q => 
                           n877, QN => net48409);
   REGISTERS_reg_9_15_inst : DFF_X1 port map( D => n1480, CK => net3441, Q => 
                           n876, QN => net48408);
   REGISTERS_reg_9_14_inst : DFF_X1 port map( D => n1502, CK => net3441, Q => 
                           n875, QN => net48407);
   REGISTERS_reg_9_13_inst : DFF_X1 port map( D => n1524, CK => net3441, Q => 
                           n874, QN => net48406);
   REGISTERS_reg_9_12_inst : DFF_X1 port map( D => n1546, CK => net3441, Q => 
                           n873, QN => net48405);
   REGISTERS_reg_9_11_inst : DFF_X1 port map( D => n1568, CK => net3441, Q => 
                           n872, QN => net48404);
   REGISTERS_reg_9_10_inst : DFF_X1 port map( D => n1590, CK => net3441, Q => 
                           n871, QN => net48403);
   REGISTERS_reg_9_9_inst : DFF_X1 port map( D => n1612, CK => net3441, Q => 
                           n870, QN => net48402);
   REGISTERS_reg_9_8_inst : DFF_X1 port map( D => n1634, CK => net3441, Q => 
                           n869, QN => net48401);
   REGISTERS_reg_9_7_inst : DFF_X1 port map( D => n1656, CK => net3441, Q => 
                           n868, QN => net48400);
   REGISTERS_reg_9_6_inst : DFF_X1 port map( D => n1678, CK => net3441, Q => 
                           n867, QN => net48399);
   REGISTERS_reg_9_5_inst : DFF_X1 port map( D => n1700, CK => net3441, Q => 
                           n866, QN => net48398);
   REGISTERS_reg_9_4_inst : DFF_X1 port map( D => n1722, CK => net3441, Q => 
                           n865, QN => net48397);
   REGISTERS_reg_9_3_inst : DFF_X1 port map( D => n1744, CK => net3441, Q => 
                           n864, QN => net48396);
   REGISTERS_reg_9_2_inst : DFF_X1 port map( D => n1766, CK => net3441, Q => 
                           n863, QN => net48395);
   REGISTERS_reg_9_1_inst : DFF_X1 port map( D => n1788, CK => net3441, Q => 
                           n862, QN => net48394);
   REGISTERS_reg_9_0_inst : DFF_X1 port map( D => n1810, CK => net3441, Q => 
                           n861, QN => net48393);
   REGISTERS_reg_10_31_inst : DFF_X1 port map( D => n1094, CK => net3446, Q => 
                           n860, QN => net48392);
   REGISTERS_reg_10_30_inst : DFF_X1 port map( D => n1150, CK => net3446, Q => 
                           n859, QN => net48391);
   REGISTERS_reg_10_29_inst : DFF_X1 port map( D => n1172, CK => net3446, Q => 
                           n857, QN => net48390);
   REGISTERS_reg_10_28_inst : DFF_X1 port map( D => n1194, CK => net3446, Q => 
                           n856, QN => net48389);
   REGISTERS_reg_10_27_inst : DFF_X1 port map( D => n1216, CK => net3446, Q => 
                           n855, QN => net48388);
   REGISTERS_reg_10_26_inst : DFF_X1 port map( D => n1238, CK => net3446, Q => 
                           n854, QN => net48387);
   REGISTERS_reg_10_25_inst : DFF_X1 port map( D => n1260, CK => net3446, Q => 
                           n853, QN => net48386);
   REGISTERS_reg_10_24_inst : DFF_X1 port map( D => n1282, CK => net3446, Q => 
                           n852, QN => net48385);
   REGISTERS_reg_10_23_inst : DFF_X1 port map( D => n1304, CK => net3446, Q => 
                           n851, QN => net48384);
   REGISTERS_reg_10_22_inst : DFF_X1 port map( D => n1326, CK => net3446, Q => 
                           n850, QN => net48383);
   REGISTERS_reg_10_21_inst : DFF_X1 port map( D => n1348, CK => net3446, Q => 
                           n849, QN => net48382);
   REGISTERS_reg_10_20_inst : DFF_X1 port map( D => n1370, CK => net3446, Q => 
                           n848, QN => net48381);
   REGISTERS_reg_10_19_inst : DFF_X1 port map( D => n1392, CK => net3446, Q => 
                           n847, QN => net48380);
   REGISTERS_reg_10_18_inst : DFF_X1 port map( D => n1414, CK => net3446, Q => 
                           n846, QN => net48379);
   REGISTERS_reg_10_17_inst : DFF_X1 port map( D => n1436, CK => net3446, Q => 
                           n845, QN => net48378);
   REGISTERS_reg_10_16_inst : DFF_X1 port map( D => n1458, CK => net3446, Q => 
                           n844, QN => net48377);
   REGISTERS_reg_10_15_inst : DFF_X1 port map( D => n1480, CK => net3446, Q => 
                           n843, QN => net48376);
   REGISTERS_reg_10_14_inst : DFF_X1 port map( D => n1502, CK => net3446, Q => 
                           n842, QN => net48375);
   REGISTERS_reg_10_13_inst : DFF_X1 port map( D => n1524, CK => net3446, Q => 
                           n841, QN => net48374);
   REGISTERS_reg_10_12_inst : DFF_X1 port map( D => n1546, CK => net3446, Q => 
                           n840, QN => net48373);
   REGISTERS_reg_10_11_inst : DFF_X1 port map( D => n1568, CK => net3446, Q => 
                           n839, QN => net48372);
   REGISTERS_reg_10_10_inst : DFF_X1 port map( D => n1590, CK => net3446, Q => 
                           n838, QN => net48371);
   REGISTERS_reg_10_9_inst : DFF_X1 port map( D => n1612, CK => net3446, Q => 
                           n836, QN => net48370);
   REGISTERS_reg_10_8_inst : DFF_X1 port map( D => n1634, CK => net3446, Q => 
                           n835, QN => net48369);
   REGISTERS_reg_10_7_inst : DFF_X1 port map( D => n1656, CK => net3446, Q => 
                           n834, QN => net48368);
   REGISTERS_reg_10_6_inst : DFF_X1 port map( D => n1678, CK => net3446, Q => 
                           n833, QN => net48367);
   REGISTERS_reg_10_5_inst : DFF_X1 port map( D => n1700, CK => net3446, Q => 
                           n832, QN => net48366);
   REGISTERS_reg_10_4_inst : DFF_X1 port map( D => n1722, CK => net3446, Q => 
                           n831, QN => net48365);
   REGISTERS_reg_10_3_inst : DFF_X1 port map( D => n1744, CK => net3446, Q => 
                           n830, QN => net48364);
   REGISTERS_reg_10_2_inst : DFF_X1 port map( D => n1766, CK => net3446, Q => 
                           n829, QN => net48363);
   REGISTERS_reg_10_1_inst : DFF_X1 port map( D => n1788, CK => net3446, Q => 
                           n828, QN => net48362);
   REGISTERS_reg_10_0_inst : DFF_X1 port map( D => n1810, CK => net3446, Q => 
                           n827, QN => net48361);
   REGISTERS_reg_11_31_inst : DFF_X1 port map( D => n1094, CK => net3451, Q => 
                           n826, QN => net48360);
   REGISTERS_reg_11_30_inst : DFF_X1 port map( D => n1150, CK => net3451, Q => 
                           n825, QN => net48359);
   REGISTERS_reg_11_29_inst : DFF_X1 port map( D => n1172, CK => net3451, Q => 
                           n824, QN => net48358);
   REGISTERS_reg_11_28_inst : DFF_X1 port map( D => n1194, CK => net3451, Q => 
                           n823, QN => net48357);
   REGISTERS_reg_11_27_inst : DFF_X1 port map( D => n1216, CK => net3451, Q => 
                           n822, QN => net48356);
   REGISTERS_reg_11_26_inst : DFF_X1 port map( D => n1238, CK => net3451, Q => 
                           n821, QN => net48355);
   REGISTERS_reg_11_25_inst : DFF_X1 port map( D => n1260, CK => net3451, Q => 
                           n820, QN => net48354);
   REGISTERS_reg_11_24_inst : DFF_X1 port map( D => n1282, CK => net3451, Q => 
                           n819, QN => net48353);
   REGISTERS_reg_11_23_inst : DFF_X1 port map( D => n1304, CK => net3451, Q => 
                           n818, QN => net48352);
   REGISTERS_reg_11_22_inst : DFF_X1 port map( D => n1326, CK => net3451, Q => 
                           n817, QN => net48351);
   REGISTERS_reg_11_21_inst : DFF_X1 port map( D => n1348, CK => net3451, Q => 
                           n815, QN => net48350);
   REGISTERS_reg_11_20_inst : DFF_X1 port map( D => n1370, CK => net3451, Q => 
                           n814, QN => net48349);
   REGISTERS_reg_11_19_inst : DFF_X1 port map( D => n1392, CK => net3451, Q => 
                           n813, QN => net48348);
   REGISTERS_reg_11_18_inst : DFF_X1 port map( D => n1414, CK => net3451, Q => 
                           n812, QN => net48347);
   REGISTERS_reg_11_17_inst : DFF_X1 port map( D => n1436, CK => net3451, Q => 
                           n811, QN => net48346);
   REGISTERS_reg_11_16_inst : DFF_X1 port map( D => n1458, CK => net3451, Q => 
                           n810, QN => net48345);
   REGISTERS_reg_11_15_inst : DFF_X1 port map( D => n1480, CK => net3451, Q => 
                           n809, QN => net48344);
   REGISTERS_reg_11_14_inst : DFF_X1 port map( D => n1502, CK => net3451, Q => 
                           n808, QN => net48343);
   REGISTERS_reg_11_13_inst : DFF_X1 port map( D => n1524, CK => net3451, Q => 
                           n807, QN => net48342);
   REGISTERS_reg_11_12_inst : DFF_X1 port map( D => n1546, CK => net3451, Q => 
                           n806, QN => net48341);
   REGISTERS_reg_11_11_inst : DFF_X1 port map( D => n1568, CK => net3451, Q => 
                           n805, QN => net48340);
   REGISTERS_reg_11_10_inst : DFF_X1 port map( D => n1590, CK => net3451, Q => 
                           n804, QN => net48339);
   REGISTERS_reg_11_9_inst : DFF_X1 port map( D => n1612, CK => net3451, Q => 
                           n803, QN => net48338);
   REGISTERS_reg_11_8_inst : DFF_X1 port map( D => n1634, CK => net3451, Q => 
                           n802, QN => net48337);
   REGISTERS_reg_11_7_inst : DFF_X1 port map( D => n1656, CK => net3451, Q => 
                           n801, QN => net48336);
   REGISTERS_reg_11_6_inst : DFF_X1 port map( D => n1678, CK => net3451, Q => 
                           n800, QN => net48335);
   REGISTERS_reg_11_5_inst : DFF_X1 port map( D => n1700, CK => net3451, Q => 
                           n799, QN => net48334);
   REGISTERS_reg_11_4_inst : DFF_X1 port map( D => n1722, CK => net3451, Q => 
                           n798, QN => net48333);
   REGISTERS_reg_11_3_inst : DFF_X1 port map( D => n1744, CK => net3451, Q => 
                           n797, QN => net48332);
   REGISTERS_reg_11_2_inst : DFF_X1 port map( D => n1766, CK => net3451, Q => 
                           n796, QN => net48331);
   REGISTERS_reg_11_1_inst : DFF_X1 port map( D => n1788, CK => net3451, Q => 
                           n794, QN => net48330);
   REGISTERS_reg_11_0_inst : DFF_X1 port map( D => n1810, CK => net3451, Q => 
                           n793, QN => net48329);
   REGISTERS_reg_12_31_inst : DFF_X1 port map( D => n1094, CK => net3456, Q => 
                           n792, QN => net48328);
   REGISTERS_reg_12_30_inst : DFF_X1 port map( D => n1150, CK => net3456, Q => 
                           n791, QN => net48327);
   REGISTERS_reg_12_29_inst : DFF_X1 port map( D => n1172, CK => net3456, Q => 
                           n790, QN => net48326);
   REGISTERS_reg_12_28_inst : DFF_X1 port map( D => n1194, CK => net3456, Q => 
                           n789, QN => net48325);
   REGISTERS_reg_12_27_inst : DFF_X1 port map( D => n1216, CK => net3456, Q => 
                           n788, QN => net48324);
   REGISTERS_reg_12_26_inst : DFF_X1 port map( D => n1238, CK => net3456, Q => 
                           n787, QN => net48323);
   REGISTERS_reg_12_25_inst : DFF_X1 port map( D => n1260, CK => net3456, Q => 
                           n786, QN => net48322);
   REGISTERS_reg_12_24_inst : DFF_X1 port map( D => n1282, CK => net3456, Q => 
                           n785, QN => net48321);
   REGISTERS_reg_12_23_inst : DFF_X1 port map( D => n1304, CK => net3456, Q => 
                           n784, QN => net48320);
   REGISTERS_reg_12_22_inst : DFF_X1 port map( D => n1326, CK => net3456, Q => 
                           n783, QN => net48319);
   REGISTERS_reg_12_21_inst : DFF_X1 port map( D => n1348, CK => net3456, Q => 
                           n782, QN => net48318);
   REGISTERS_reg_12_20_inst : DFF_X1 port map( D => n1370, CK => net3456, Q => 
                           n781, QN => net48317);
   REGISTERS_reg_12_19_inst : DFF_X1 port map( D => n1392, CK => net3456, Q => 
                           n780, QN => net48316);
   REGISTERS_reg_12_18_inst : DFF_X1 port map( D => n1414, CK => net3456, Q => 
                           n779, QN => net48315);
   REGISTERS_reg_12_17_inst : DFF_X1 port map( D => n1436, CK => net3456, Q => 
                           n778, QN => net48314);
   REGISTERS_reg_12_16_inst : DFF_X1 port map( D => n1458, CK => net3456, Q => 
                           n777, QN => net48313);
   REGISTERS_reg_12_15_inst : DFF_X1 port map( D => n1480, CK => net3456, Q => 
                           n776, QN => net48312);
   REGISTERS_reg_12_14_inst : DFF_X1 port map( D => n1502, CK => net3456, Q => 
                           n775, QN => net48311);
   REGISTERS_reg_12_13_inst : DFF_X1 port map( D => n1524, CK => net3456, Q => 
                           n773, QN => net48310);
   REGISTERS_reg_12_12_inst : DFF_X1 port map( D => n1546, CK => net3456, Q => 
                           n772, QN => net48309);
   REGISTERS_reg_12_11_inst : DFF_X1 port map( D => n1568, CK => net3456, Q => 
                           n771, QN => net48308);
   REGISTERS_reg_12_10_inst : DFF_X1 port map( D => n1590, CK => net3456, Q => 
                           n770, QN => net48307);
   REGISTERS_reg_12_9_inst : DFF_X1 port map( D => n1612, CK => net3456, Q => 
                           n769, QN => net48306);
   REGISTERS_reg_12_8_inst : DFF_X1 port map( D => n1634, CK => net3456, Q => 
                           n768, QN => net48305);
   REGISTERS_reg_12_7_inst : DFF_X1 port map( D => n1656, CK => net3456, Q => 
                           n767, QN => net48304);
   REGISTERS_reg_12_6_inst : DFF_X1 port map( D => n1678, CK => net3456, Q => 
                           n766, QN => net48303);
   REGISTERS_reg_12_5_inst : DFF_X1 port map( D => n1700, CK => net3456, Q => 
                           n765, QN => net48302);
   REGISTERS_reg_12_4_inst : DFF_X1 port map( D => n1722, CK => net3456, Q => 
                           n764, QN => net48301);
   REGISTERS_reg_12_3_inst : DFF_X1 port map( D => n1744, CK => net3456, Q => 
                           n763, QN => net48300);
   REGISTERS_reg_12_2_inst : DFF_X1 port map( D => n1766, CK => net3456, Q => 
                           n762, QN => net48299);
   REGISTERS_reg_12_1_inst : DFF_X1 port map( D => n1788, CK => net3456, Q => 
                           n761, QN => net48298);
   REGISTERS_reg_12_0_inst : DFF_X1 port map( D => n1810, CK => net3456, Q => 
                           n760, QN => net48297);
   REGISTERS_reg_13_31_inst : DFF_X1 port map( D => n1094, CK => net3461, Q => 
                           n759, QN => net48296);
   REGISTERS_reg_13_30_inst : DFF_X1 port map( D => n1150, CK => net3461, Q => 
                           n758, QN => net48295);
   REGISTERS_reg_13_29_inst : DFF_X1 port map( D => n1172, CK => net3461, Q => 
                           n757, QN => net48294);
   REGISTERS_reg_13_28_inst : DFF_X1 port map( D => n1194, CK => net3461, Q => 
                           n756, QN => net48293);
   REGISTERS_reg_13_27_inst : DFF_X1 port map( D => n1216, CK => net3461, Q => 
                           n755, QN => net48292);
   REGISTERS_reg_13_26_inst : DFF_X1 port map( D => n1238, CK => net3461, Q => 
                           n754, QN => net48291);
   REGISTERS_reg_13_25_inst : DFF_X1 port map( D => n1260, CK => net3461, Q => 
                           n752, QN => net48290);
   REGISTERS_reg_13_24_inst : DFF_X1 port map( D => n1282, CK => net3461, Q => 
                           n751, QN => net48289);
   REGISTERS_reg_13_23_inst : DFF_X1 port map( D => n1304, CK => net3461, Q => 
                           n750, QN => net48288);
   REGISTERS_reg_13_22_inst : DFF_X1 port map( D => n1326, CK => net3461, Q => 
                           n749, QN => net48287);
   REGISTERS_reg_13_21_inst : DFF_X1 port map( D => n1348, CK => net3461, Q => 
                           n748, QN => net48286);
   REGISTERS_reg_13_20_inst : DFF_X1 port map( D => n1370, CK => net3461, Q => 
                           n747, QN => net48285);
   REGISTERS_reg_13_19_inst : DFF_X1 port map( D => n1392, CK => net3461, Q => 
                           n746, QN => net48284);
   REGISTERS_reg_13_18_inst : DFF_X1 port map( D => n1414, CK => net3461, Q => 
                           n745, QN => net48283);
   REGISTERS_reg_13_17_inst : DFF_X1 port map( D => n1436, CK => net3461, Q => 
                           n744, QN => net48282);
   REGISTERS_reg_13_16_inst : DFF_X1 port map( D => n1458, CK => net3461, Q => 
                           n743, QN => net48281);
   REGISTERS_reg_13_15_inst : DFF_X1 port map( D => n1480, CK => net3461, Q => 
                           n742, QN => net48280);
   REGISTERS_reg_13_14_inst : DFF_X1 port map( D => n1502, CK => net3461, Q => 
                           n741, QN => net48279);
   REGISTERS_reg_13_13_inst : DFF_X1 port map( D => n1524, CK => net3461, Q => 
                           n740, QN => net48278);
   REGISTERS_reg_13_12_inst : DFF_X1 port map( D => n1546, CK => net3461, Q => 
                           n739, QN => net48277);
   REGISTERS_reg_13_11_inst : DFF_X1 port map( D => n1568, CK => net3461, Q => 
                           n738, QN => net48276);
   REGISTERS_reg_13_10_inst : DFF_X1 port map( D => n1590, CK => net3461, Q => 
                           n737, QN => net48275);
   REGISTERS_reg_13_9_inst : DFF_X1 port map( D => n1612, CK => net3461, Q => 
                           n736, QN => net48274);
   REGISTERS_reg_13_8_inst : DFF_X1 port map( D => n1634, CK => net3461, Q => 
                           n735, QN => net48273);
   REGISTERS_reg_13_7_inst : DFF_X1 port map( D => n1656, CK => net3461, Q => 
                           n734, QN => net48272);
   REGISTERS_reg_13_6_inst : DFF_X1 port map( D => n1678, CK => net3461, Q => 
                           n733, QN => net48271);
   REGISTERS_reg_13_5_inst : DFF_X1 port map( D => n1700, CK => net3461, Q => 
                           n731, QN => net48270);
   REGISTERS_reg_13_4_inst : DFF_X1 port map( D => n1722, CK => net3461, Q => 
                           n730, QN => net48269);
   REGISTERS_reg_13_3_inst : DFF_X1 port map( D => n1744, CK => net3461, Q => 
                           n729, QN => net48268);
   REGISTERS_reg_13_2_inst : DFF_X1 port map( D => n1766, CK => net3461, Q => 
                           n728, QN => net48267);
   REGISTERS_reg_13_1_inst : DFF_X1 port map( D => n1788, CK => net3461, Q => 
                           n727, QN => net48266);
   REGISTERS_reg_13_0_inst : DFF_X1 port map( D => n1810, CK => net3461, Q => 
                           n726, QN => net48265);
   REGISTERS_reg_14_31_inst : DFF_X1 port map( D => n1094, CK => net3466, Q => 
                           n725, QN => net48264);
   REGISTERS_reg_14_30_inst : DFF_X1 port map( D => n1150, CK => net3466, Q => 
                           n724, QN => net48263);
   REGISTERS_reg_14_29_inst : DFF_X1 port map( D => n1172, CK => net3466, Q => 
                           n723, QN => net48262);
   REGISTERS_reg_14_28_inst : DFF_X1 port map( D => n1194, CK => net3466, Q => 
                           n722, QN => net48261);
   REGISTERS_reg_14_27_inst : DFF_X1 port map( D => n1216, CK => net3466, Q => 
                           n721, QN => net48260);
   REGISTERS_reg_14_26_inst : DFF_X1 port map( D => n1238, CK => net3466, Q => 
                           n720, QN => net48259);
   REGISTERS_reg_14_25_inst : DFF_X1 port map( D => n1260, CK => net3466, Q => 
                           n719, QN => net48258);
   REGISTERS_reg_14_24_inst : DFF_X1 port map( D => n1282, CK => net3466, Q => 
                           n718, QN => net48257);
   REGISTERS_reg_14_23_inst : DFF_X1 port map( D => n1304, CK => net3466, Q => 
                           n717, QN => net48256);
   REGISTERS_reg_14_22_inst : DFF_X1 port map( D => n1326, CK => net3466, Q => 
                           n716, QN => net48255);
   REGISTERS_reg_14_21_inst : DFF_X1 port map( D => n1348, CK => net3466, Q => 
                           n715, QN => net48254);
   REGISTERS_reg_14_20_inst : DFF_X1 port map( D => n1370, CK => net3466, Q => 
                           n714, QN => net48253);
   REGISTERS_reg_14_19_inst : DFF_X1 port map( D => n1392, CK => net3466, Q => 
                           n713, QN => net48252);
   REGISTERS_reg_14_18_inst : DFF_X1 port map( D => n1414, CK => net3466, Q => 
                           n712, QN => net48251);
   REGISTERS_reg_14_17_inst : DFF_X1 port map( D => n1436, CK => net3466, Q => 
                           n710, QN => net48250);
   REGISTERS_reg_14_16_inst : DFF_X1 port map( D => n1458, CK => net3466, Q => 
                           n709, QN => net48249);
   REGISTERS_reg_14_15_inst : DFF_X1 port map( D => n1480, CK => net3466, Q => 
                           n708, QN => net48248);
   REGISTERS_reg_14_14_inst : DFF_X1 port map( D => n1502, CK => net3466, Q => 
                           n707, QN => net48247);
   REGISTERS_reg_14_13_inst : DFF_X1 port map( D => n1524, CK => net3466, Q => 
                           n706, QN => net48246);
   REGISTERS_reg_14_12_inst : DFF_X1 port map( D => n1546, CK => net3466, Q => 
                           n705, QN => net48245);
   REGISTERS_reg_14_11_inst : DFF_X1 port map( D => n1568, CK => net3466, Q => 
                           n704, QN => net48244);
   REGISTERS_reg_14_10_inst : DFF_X1 port map( D => n1590, CK => net3466, Q => 
                           n703, QN => net48243);
   REGISTERS_reg_14_9_inst : DFF_X1 port map( D => n1612, CK => net3466, Q => 
                           n702, QN => net48242);
   REGISTERS_reg_14_8_inst : DFF_X1 port map( D => n1634, CK => net3466, Q => 
                           n701, QN => net48241);
   REGISTERS_reg_14_7_inst : DFF_X1 port map( D => n1656, CK => net3466, Q => 
                           n700, QN => net48240);
   REGISTERS_reg_14_6_inst : DFF_X1 port map( D => n1678, CK => net3466, Q => 
                           n699, QN => net48239);
   REGISTERS_reg_14_5_inst : DFF_X1 port map( D => n1700, CK => net3466, Q => 
                           n698, QN => net48238);
   REGISTERS_reg_14_4_inst : DFF_X1 port map( D => n1722, CK => net3466, Q => 
                           n697, QN => net48237);
   REGISTERS_reg_14_3_inst : DFF_X1 port map( D => n1744, CK => net3466, Q => 
                           n696, QN => net48236);
   REGISTERS_reg_14_2_inst : DFF_X1 port map( D => n1766, CK => net3466, Q => 
                           n695, QN => net48235);
   REGISTERS_reg_14_1_inst : DFF_X1 port map( D => n1788, CK => net3466, Q => 
                           n694, QN => net48234);
   REGISTERS_reg_14_0_inst : DFF_X1 port map( D => n1810, CK => net3466, Q => 
                           n693, QN => net48233);
   REGISTERS_reg_15_31_inst : DFF_X1 port map( D => n1094, CK => net3471, Q => 
                           n692, QN => net48232);
   REGISTERS_reg_15_30_inst : DFF_X1 port map( D => n1150, CK => net3471, Q => 
                           n691, QN => net48231);
   REGISTERS_reg_15_29_inst : DFF_X1 port map( D => n1172, CK => net3471, Q => 
                           n689, QN => net48230);
   REGISTERS_reg_15_28_inst : DFF_X1 port map( D => n1194, CK => net3471, Q => 
                           n688, QN => net48229);
   REGISTERS_reg_15_27_inst : DFF_X1 port map( D => n1216, CK => net3471, Q => 
                           n687, QN => net48228);
   REGISTERS_reg_15_26_inst : DFF_X1 port map( D => n1238, CK => net3471, Q => 
                           n686, QN => net48227);
   REGISTERS_reg_15_25_inst : DFF_X1 port map( D => n1260, CK => net3471, Q => 
                           n685, QN => net48226);
   REGISTERS_reg_15_24_inst : DFF_X1 port map( D => n1282, CK => net3471, Q => 
                           n684, QN => net48225);
   REGISTERS_reg_15_23_inst : DFF_X1 port map( D => n1304, CK => net3471, Q => 
                           n683, QN => net48224);
   REGISTERS_reg_15_22_inst : DFF_X1 port map( D => n1326, CK => net3471, Q => 
                           n682, QN => net48223);
   REGISTERS_reg_15_21_inst : DFF_X1 port map( D => n1348, CK => net3471, Q => 
                           n681, QN => net48222);
   REGISTERS_reg_15_20_inst : DFF_X1 port map( D => n1370, CK => net3471, Q => 
                           n680, QN => net48221);
   REGISTERS_reg_15_19_inst : DFF_X1 port map( D => n1392, CK => net3471, Q => 
                           n679, QN => net48220);
   REGISTERS_reg_15_18_inst : DFF_X1 port map( D => n1414, CK => net3471, Q => 
                           n678, QN => net48219);
   REGISTERS_reg_15_17_inst : DFF_X1 port map( D => n1436, CK => net3471, Q => 
                           n677, QN => net48218);
   REGISTERS_reg_15_16_inst : DFF_X1 port map( D => n1458, CK => net3471, Q => 
                           n676, QN => net48217);
   REGISTERS_reg_15_15_inst : DFF_X1 port map( D => n1480, CK => net3471, Q => 
                           n675, QN => net48216);
   REGISTERS_reg_15_14_inst : DFF_X1 port map( D => n1502, CK => net3471, Q => 
                           n674, QN => net48215);
   REGISTERS_reg_15_13_inst : DFF_X1 port map( D => n1524, CK => net3471, Q => 
                           n673, QN => net48214);
   REGISTERS_reg_15_12_inst : DFF_X1 port map( D => n1546, CK => net3471, Q => 
                           n672, QN => net48213);
   REGISTERS_reg_15_11_inst : DFF_X1 port map( D => n1568, CK => net3471, Q => 
                           n671, QN => net48212);
   REGISTERS_reg_15_10_inst : DFF_X1 port map( D => n1590, CK => net3471, Q => 
                           n670, QN => net48211);
   REGISTERS_reg_15_9_inst : DFF_X1 port map( D => n1612, CK => net3471, Q => 
                           n668, QN => net48210);
   REGISTERS_reg_15_8_inst : DFF_X1 port map( D => n1634, CK => net3471, Q => 
                           n667, QN => net48209);
   REGISTERS_reg_15_7_inst : DFF_X1 port map( D => n1656, CK => net3471, Q => 
                           n666, QN => net48208);
   REGISTERS_reg_15_6_inst : DFF_X1 port map( D => n1678, CK => net3471, Q => 
                           n665, QN => net48207);
   REGISTERS_reg_15_5_inst : DFF_X1 port map( D => n1700, CK => net3471, Q => 
                           n664, QN => net48206);
   REGISTERS_reg_15_4_inst : DFF_X1 port map( D => n1722, CK => net3471, Q => 
                           n663, QN => net48205);
   REGISTERS_reg_15_3_inst : DFF_X1 port map( D => n1744, CK => net3471, Q => 
                           n662, QN => net48204);
   REGISTERS_reg_15_2_inst : DFF_X1 port map( D => n1766, CK => net3471, Q => 
                           n661, QN => net48203);
   REGISTERS_reg_15_1_inst : DFF_X1 port map( D => n1788, CK => net3471, Q => 
                           n660, QN => net48202);
   REGISTERS_reg_15_0_inst : DFF_X1 port map( D => n1810, CK => net3471, Q => 
                           n659, QN => net48201);
   REGISTERS_reg_16_31_inst : DFF_X1 port map( D => n1094, CK => net3476, Q => 
                           n658, QN => net48200);
   REGISTERS_reg_16_30_inst : DFF_X1 port map( D => n1150, CK => net3476, Q => 
                           n657, QN => net48199);
   REGISTERS_reg_16_29_inst : DFF_X1 port map( D => n1172, CK => net3476, Q => 
                           n656, QN => net48198);
   REGISTERS_reg_16_28_inst : DFF_X1 port map( D => n1194, CK => net3476, Q => 
                           n655, QN => net48197);
   REGISTERS_reg_16_27_inst : DFF_X1 port map( D => n1216, CK => net3476, Q => 
                           n654, QN => net48196);
   REGISTERS_reg_16_26_inst : DFF_X1 port map( D => n1238, CK => net3476, Q => 
                           n653, QN => net48195);
   REGISTERS_reg_16_25_inst : DFF_X1 port map( D => n1260, CK => net3476, Q => 
                           n652, QN => net48194);
   REGISTERS_reg_16_24_inst : DFF_X1 port map( D => n1282, CK => net3476, Q => 
                           n651, QN => net48193);
   REGISTERS_reg_16_23_inst : DFF_X1 port map( D => n1304, CK => net3476, Q => 
                           n650, QN => net48192);
   REGISTERS_reg_16_22_inst : DFF_X1 port map( D => n1326, CK => net3476, Q => 
                           n649, QN => net48191);
   REGISTERS_reg_16_21_inst : DFF_X1 port map( D => n1348, CK => net3476, Q => 
                           n647, QN => net48190);
   REGISTERS_reg_16_20_inst : DFF_X1 port map( D => n1370, CK => net3476, Q => 
                           n646, QN => net48189);
   REGISTERS_reg_16_19_inst : DFF_X1 port map( D => n1392, CK => net3476, Q => 
                           n645, QN => net48188);
   REGISTERS_reg_16_18_inst : DFF_X1 port map( D => n1414, CK => net3476, Q => 
                           n644, QN => net48187);
   REGISTERS_reg_16_17_inst : DFF_X1 port map( D => n1436, CK => net3476, Q => 
                           n643, QN => net48186);
   REGISTERS_reg_16_16_inst : DFF_X1 port map( D => n1458, CK => net3476, Q => 
                           n642, QN => net48185);
   REGISTERS_reg_16_15_inst : DFF_X1 port map( D => n1480, CK => net3476, Q => 
                           n641, QN => net48184);
   REGISTERS_reg_16_14_inst : DFF_X1 port map( D => n1502, CK => net3476, Q => 
                           n640, QN => net48183);
   REGISTERS_reg_16_13_inst : DFF_X1 port map( D => n1524, CK => net3476, Q => 
                           n639, QN => net48182);
   REGISTERS_reg_16_12_inst : DFF_X1 port map( D => n1546, CK => net3476, Q => 
                           n638, QN => net48181);
   REGISTERS_reg_16_11_inst : DFF_X1 port map( D => n1568, CK => net3476, Q => 
                           n637, QN => net48180);
   REGISTERS_reg_16_10_inst : DFF_X1 port map( D => n1590, CK => net3476, Q => 
                           n636, QN => net48179);
   REGISTERS_reg_16_9_inst : DFF_X1 port map( D => n1612, CK => net3476, Q => 
                           n635, QN => net48178);
   REGISTERS_reg_16_8_inst : DFF_X1 port map( D => n1634, CK => net3476, Q => 
                           n634, QN => net48177);
   REGISTERS_reg_16_7_inst : DFF_X1 port map( D => n1656, CK => net3476, Q => 
                           n633, QN => net48176);
   REGISTERS_reg_16_6_inst : DFF_X1 port map( D => n1678, CK => net3476, Q => 
                           n632, QN => net48175);
   REGISTERS_reg_16_5_inst : DFF_X1 port map( D => n1700, CK => net3476, Q => 
                           n631, QN => net48174);
   REGISTERS_reg_16_4_inst : DFF_X1 port map( D => n1722, CK => net3476, Q => 
                           n630, QN => net48173);
   REGISTERS_reg_16_3_inst : DFF_X1 port map( D => n1744, CK => net3476, Q => 
                           n629, QN => net48172);
   REGISTERS_reg_16_2_inst : DFF_X1 port map( D => n1766, CK => net3476, Q => 
                           n628, QN => net48171);
   REGISTERS_reg_16_1_inst : DFF_X1 port map( D => n1788, CK => net3476, Q => 
                           n626, QN => net48170);
   REGISTERS_reg_16_0_inst : DFF_X1 port map( D => n1810, CK => net3476, Q => 
                           n625, QN => net48169);
   REGISTERS_reg_17_31_inst : DFF_X1 port map( D => n1094, CK => net3481, Q => 
                           n624, QN => net48168);
   REGISTERS_reg_17_30_inst : DFF_X1 port map( D => n1150, CK => net3481, Q => 
                           n623, QN => net48167);
   REGISTERS_reg_17_29_inst : DFF_X1 port map( D => n1172, CK => net3481, Q => 
                           n622, QN => net48166);
   REGISTERS_reg_17_28_inst : DFF_X1 port map( D => n1194, CK => net3481, Q => 
                           n621, QN => net48165);
   REGISTERS_reg_17_27_inst : DFF_X1 port map( D => n1216, CK => net3481, Q => 
                           n620, QN => net48164);
   REGISTERS_reg_17_26_inst : DFF_X1 port map( D => n1238, CK => net3481, Q => 
                           n619, QN => net48163);
   REGISTERS_reg_17_25_inst : DFF_X1 port map( D => n1260, CK => net3481, Q => 
                           n618, QN => net48162);
   REGISTERS_reg_17_24_inst : DFF_X1 port map( D => n1282, CK => net3481, Q => 
                           n617, QN => net48161);
   REGISTERS_reg_17_23_inst : DFF_X1 port map( D => n1304, CK => net3481, Q => 
                           n616, QN => net48160);
   REGISTERS_reg_17_22_inst : DFF_X1 port map( D => n1326, CK => net3481, Q => 
                           n615, QN => net48159);
   REGISTERS_reg_17_21_inst : DFF_X1 port map( D => n1348, CK => net3481, Q => 
                           n614, QN => net48158);
   REGISTERS_reg_17_20_inst : DFF_X1 port map( D => n1370, CK => net3481, Q => 
                           n613, QN => net48157);
   REGISTERS_reg_17_19_inst : DFF_X1 port map( D => n1392, CK => net3481, Q => 
                           n612, QN => net48156);
   REGISTERS_reg_17_18_inst : DFF_X1 port map( D => n1414, CK => net3481, Q => 
                           n611, QN => net48155);
   REGISTERS_reg_17_17_inst : DFF_X1 port map( D => n1436, CK => net3481, Q => 
                           n610, QN => net48154);
   REGISTERS_reg_17_16_inst : DFF_X1 port map( D => n1458, CK => net3481, Q => 
                           n609, QN => net48153);
   REGISTERS_reg_17_15_inst : DFF_X1 port map( D => n1480, CK => net3481, Q => 
                           n608, QN => net48152);
   REGISTERS_reg_17_14_inst : DFF_X1 port map( D => n1502, CK => net3481, Q => 
                           n607, QN => net48151);
   REGISTERS_reg_17_13_inst : DFF_X1 port map( D => n1524, CK => net3481, Q => 
                           n605, QN => net48150);
   REGISTERS_reg_17_12_inst : DFF_X1 port map( D => n1546, CK => net3481, Q => 
                           n604, QN => net48149);
   REGISTERS_reg_17_11_inst : DFF_X1 port map( D => n1568, CK => net3481, Q => 
                           n603, QN => net48148);
   REGISTERS_reg_17_10_inst : DFF_X1 port map( D => n1590, CK => net3481, Q => 
                           n602, QN => net48147);
   REGISTERS_reg_17_9_inst : DFF_X1 port map( D => n1612, CK => net3481, Q => 
                           n601, QN => net48146);
   REGISTERS_reg_17_8_inst : DFF_X1 port map( D => n1634, CK => net3481, Q => 
                           n600, QN => net48145);
   REGISTERS_reg_17_7_inst : DFF_X1 port map( D => n1656, CK => net3481, Q => 
                           n599, QN => net48144);
   REGISTERS_reg_17_6_inst : DFF_X1 port map( D => n1678, CK => net3481, Q => 
                           n598, QN => net48143);
   REGISTERS_reg_17_5_inst : DFF_X1 port map( D => n1700, CK => net3481, Q => 
                           n597, QN => net48142);
   REGISTERS_reg_17_4_inst : DFF_X1 port map( D => n1722, CK => net3481, Q => 
                           n596, QN => net48141);
   REGISTERS_reg_17_3_inst : DFF_X1 port map( D => n1744, CK => net3481, Q => 
                           n595, QN => net48140);
   REGISTERS_reg_17_2_inst : DFF_X1 port map( D => n1766, CK => net3481, Q => 
                           n594, QN => net48139);
   REGISTERS_reg_17_1_inst : DFF_X1 port map( D => n1788, CK => net3481, Q => 
                           n593, QN => net48138);
   REGISTERS_reg_17_0_inst : DFF_X1 port map( D => n1810, CK => net3481, Q => 
                           n592, QN => net48137);
   REGISTERS_reg_18_31_inst : DFF_X1 port map( D => n1094, CK => net3486, Q => 
                           n591, QN => net48136);
   REGISTERS_reg_18_30_inst : DFF_X1 port map( D => n1150, CK => net3486, Q => 
                           n590, QN => net48135);
   REGISTERS_reg_18_29_inst : DFF_X1 port map( D => n1172, CK => net3486, Q => 
                           n589, QN => net48134);
   REGISTERS_reg_18_28_inst : DFF_X1 port map( D => n1194, CK => net3486, Q => 
                           n588, QN => net48133);
   REGISTERS_reg_18_27_inst : DFF_X1 port map( D => n1216, CK => net3486, Q => 
                           n587, QN => net48132);
   REGISTERS_reg_18_26_inst : DFF_X1 port map( D => n1238, CK => net3486, Q => 
                           n586, QN => net48131);
   REGISTERS_reg_18_25_inst : DFF_X1 port map( D => n1260, CK => net3486, Q => 
                           n584, QN => net48130);
   REGISTERS_reg_18_24_inst : DFF_X1 port map( D => n1282, CK => net3486, Q => 
                           n583, QN => net48129);
   REGISTERS_reg_18_23_inst : DFF_X1 port map( D => n1304, CK => net3486, Q => 
                           n582, QN => net48128);
   REGISTERS_reg_18_22_inst : DFF_X1 port map( D => n1326, CK => net3486, Q => 
                           n581, QN => net48127);
   REGISTERS_reg_18_21_inst : DFF_X1 port map( D => n1348, CK => net3486, Q => 
                           n580, QN => net48126);
   REGISTERS_reg_18_20_inst : DFF_X1 port map( D => n1370, CK => net3486, Q => 
                           n579, QN => net48125);
   REGISTERS_reg_18_19_inst : DFF_X1 port map( D => n1392, CK => net3486, Q => 
                           n578, QN => net48124);
   REGISTERS_reg_18_18_inst : DFF_X1 port map( D => n1414, CK => net3486, Q => 
                           n577, QN => net48123);
   REGISTERS_reg_18_17_inst : DFF_X1 port map( D => n1436, CK => net3486, Q => 
                           n576, QN => net48122);
   REGISTERS_reg_18_16_inst : DFF_X1 port map( D => n1458, CK => net3486, Q => 
                           n575, QN => net48121);
   REGISTERS_reg_18_15_inst : DFF_X1 port map( D => n1480, CK => net3486, Q => 
                           n574, QN => net48120);
   REGISTERS_reg_18_14_inst : DFF_X1 port map( D => n1502, CK => net3486, Q => 
                           n573, QN => net48119);
   REGISTERS_reg_18_13_inst : DFF_X1 port map( D => n1524, CK => net3486, Q => 
                           n572, QN => net48118);
   REGISTERS_reg_18_12_inst : DFF_X1 port map( D => n1546, CK => net3486, Q => 
                           n571, QN => net48117);
   REGISTERS_reg_18_11_inst : DFF_X1 port map( D => n1568, CK => net3486, Q => 
                           n570, QN => net48116);
   REGISTERS_reg_18_10_inst : DFF_X1 port map( D => n1590, CK => net3486, Q => 
                           n569, QN => net48115);
   REGISTERS_reg_18_9_inst : DFF_X1 port map( D => n1612, CK => net3486, Q => 
                           n568, QN => net48114);
   REGISTERS_reg_18_8_inst : DFF_X1 port map( D => n1634, CK => net3486, Q => 
                           n567, QN => net48113);
   REGISTERS_reg_18_7_inst : DFF_X1 port map( D => n1656, CK => net3486, Q => 
                           n566, QN => net48112);
   REGISTERS_reg_18_6_inst : DFF_X1 port map( D => n1678, CK => net3486, Q => 
                           n565, QN => net48111);
   REGISTERS_reg_18_5_inst : DFF_X1 port map( D => n1700, CK => net3486, Q => 
                           n563, QN => net48110);
   REGISTERS_reg_18_4_inst : DFF_X1 port map( D => n1722, CK => net3486, Q => 
                           n562, QN => net48109);
   REGISTERS_reg_18_3_inst : DFF_X1 port map( D => n1744, CK => net3486, Q => 
                           n561, QN => net48108);
   REGISTERS_reg_18_2_inst : DFF_X1 port map( D => n1766, CK => net3486, Q => 
                           n560, QN => net48107);
   REGISTERS_reg_18_1_inst : DFF_X1 port map( D => n1788, CK => net3486, Q => 
                           n559, QN => net48106);
   REGISTERS_reg_18_0_inst : DFF_X1 port map( D => n1810, CK => net3486, Q => 
                           n558, QN => net48105);
   REGISTERS_reg_19_31_inst : DFF_X1 port map( D => n1094, CK => net3491, Q => 
                           n557, QN => net48104);
   REGISTERS_reg_19_30_inst : DFF_X1 port map( D => n1150, CK => net3491, Q => 
                           n556, QN => net48103);
   REGISTERS_reg_19_29_inst : DFF_X1 port map( D => n1172, CK => net3491, Q => 
                           n555, QN => net48102);
   REGISTERS_reg_19_28_inst : DFF_X1 port map( D => n1194, CK => net3491, Q => 
                           n554, QN => net48101);
   REGISTERS_reg_19_27_inst : DFF_X1 port map( D => n1216, CK => net3491, Q => 
                           n553, QN => net48100);
   REGISTERS_reg_19_26_inst : DFF_X1 port map( D => n1238, CK => net3491, Q => 
                           n552, QN => net48099);
   REGISTERS_reg_19_25_inst : DFF_X1 port map( D => n1260, CK => net3491, Q => 
                           n551, QN => net48098);
   REGISTERS_reg_19_24_inst : DFF_X1 port map( D => n1282, CK => net3491, Q => 
                           n550, QN => net48097);
   REGISTERS_reg_19_23_inst : DFF_X1 port map( D => n1304, CK => net3491, Q => 
                           n549, QN => net48096);
   REGISTERS_reg_19_22_inst : DFF_X1 port map( D => n1326, CK => net3491, Q => 
                           n548, QN => net48095);
   REGISTERS_reg_19_21_inst : DFF_X1 port map( D => n1348, CK => net3491, Q => 
                           n547, QN => net48094);
   REGISTERS_reg_19_20_inst : DFF_X1 port map( D => n1370, CK => net3491, Q => 
                           n546, QN => net48093);
   REGISTERS_reg_19_19_inst : DFF_X1 port map( D => n1392, CK => net3491, Q => 
                           n545, QN => net48092);
   REGISTERS_reg_19_18_inst : DFF_X1 port map( D => n1414, CK => net3491, Q => 
                           n544, QN => net48091);
   REGISTERS_reg_19_17_inst : DFF_X1 port map( D => n1436, CK => net3491, Q => 
                           n542, QN => net48090);
   REGISTERS_reg_19_16_inst : DFF_X1 port map( D => n1458, CK => net3491, Q => 
                           n541, QN => net48089);
   REGISTERS_reg_19_15_inst : DFF_X1 port map( D => n1480, CK => net3491, Q => 
                           n540, QN => net48088);
   REGISTERS_reg_19_14_inst : DFF_X1 port map( D => n1502, CK => net3491, Q => 
                           n539, QN => net48087);
   REGISTERS_reg_19_13_inst : DFF_X1 port map( D => n1524, CK => net3491, Q => 
                           n538, QN => net48086);
   REGISTERS_reg_19_12_inst : DFF_X1 port map( D => n1546, CK => net3491, Q => 
                           n537, QN => net48085);
   REGISTERS_reg_19_11_inst : DFF_X1 port map( D => n1568, CK => net3491, Q => 
                           n536, QN => net48084);
   REGISTERS_reg_19_10_inst : DFF_X1 port map( D => n1590, CK => net3491, Q => 
                           n535, QN => net48083);
   REGISTERS_reg_19_9_inst : DFF_X1 port map( D => n1612, CK => net3491, Q => 
                           n534, QN => net48082);
   REGISTERS_reg_19_8_inst : DFF_X1 port map( D => n1634, CK => net3491, Q => 
                           n533, QN => net48081);
   REGISTERS_reg_19_7_inst : DFF_X1 port map( D => n1656, CK => net3491, Q => 
                           n532, QN => net48080);
   REGISTERS_reg_19_6_inst : DFF_X1 port map( D => n1678, CK => net3491, Q => 
                           n531, QN => net48079);
   REGISTERS_reg_19_5_inst : DFF_X1 port map( D => n1700, CK => net3491, Q => 
                           n530, QN => net48078);
   REGISTERS_reg_19_4_inst : DFF_X1 port map( D => n1722, CK => net3491, Q => 
                           n529, QN => net48077);
   REGISTERS_reg_19_3_inst : DFF_X1 port map( D => n1744, CK => net3491, Q => 
                           n528, QN => net48076);
   REGISTERS_reg_19_2_inst : DFF_X1 port map( D => n1766, CK => net3491, Q => 
                           n527, QN => net48075);
   REGISTERS_reg_19_1_inst : DFF_X1 port map( D => n1788, CK => net3491, Q => 
                           n526, QN => net48074);
   REGISTERS_reg_19_0_inst : DFF_X1 port map( D => n1810, CK => net3491, Q => 
                           n525, QN => net48073);
   REGISTERS_reg_20_31_inst : DFF_X1 port map( D => n1094, CK => net3496, Q => 
                           n524, QN => net48072);
   REGISTERS_reg_20_30_inst : DFF_X1 port map( D => n1150, CK => net3496, Q => 
                           n523, QN => net48071);
   REGISTERS_reg_20_29_inst : DFF_X1 port map( D => n1172, CK => net3496, Q => 
                           n521, QN => net48070);
   REGISTERS_reg_20_28_inst : DFF_X1 port map( D => n1194, CK => net3496, Q => 
                           n520, QN => net48069);
   REGISTERS_reg_20_27_inst : DFF_X1 port map( D => n1216, CK => net3496, Q => 
                           n519, QN => net48068);
   REGISTERS_reg_20_26_inst : DFF_X1 port map( D => n1238, CK => net3496, Q => 
                           n518, QN => net48067);
   REGISTERS_reg_20_25_inst : DFF_X1 port map( D => n1260, CK => net3496, Q => 
                           n517, QN => net48066);
   REGISTERS_reg_20_24_inst : DFF_X1 port map( D => n1282, CK => net3496, Q => 
                           n516, QN => net48065);
   REGISTERS_reg_20_23_inst : DFF_X1 port map( D => n1304, CK => net3496, Q => 
                           n515, QN => net48064);
   REGISTERS_reg_20_22_inst : DFF_X1 port map( D => n1326, CK => net3496, Q => 
                           n514, QN => net48063);
   REGISTERS_reg_20_21_inst : DFF_X1 port map( D => n1348, CK => net3496, Q => 
                           n513, QN => net48062);
   REGISTERS_reg_20_20_inst : DFF_X1 port map( D => n1370, CK => net3496, Q => 
                           n512, QN => net48061);
   REGISTERS_reg_20_19_inst : DFF_X1 port map( D => n1392, CK => net3496, Q => 
                           n511, QN => net48060);
   REGISTERS_reg_20_18_inst : DFF_X1 port map( D => n1414, CK => net3496, Q => 
                           n510, QN => net48059);
   REGISTERS_reg_20_17_inst : DFF_X1 port map( D => n1436, CK => net3496, Q => 
                           n509, QN => net48058);
   REGISTERS_reg_20_16_inst : DFF_X1 port map( D => n1458, CK => net3496, Q => 
                           n508, QN => net48057);
   REGISTERS_reg_20_15_inst : DFF_X1 port map( D => n1480, CK => net3496, Q => 
                           n507, QN => net48056);
   REGISTERS_reg_20_14_inst : DFF_X1 port map( D => n1502, CK => net3496, Q => 
                           n506, QN => net48055);
   REGISTERS_reg_20_13_inst : DFF_X1 port map( D => n1524, CK => net3496, Q => 
                           n505, QN => net48054);
   REGISTERS_reg_20_12_inst : DFF_X1 port map( D => n1546, CK => net3496, Q => 
                           n504, QN => net48053);
   REGISTERS_reg_20_11_inst : DFF_X1 port map( D => n1568, CK => net3496, Q => 
                           n503, QN => net48052);
   REGISTERS_reg_20_10_inst : DFF_X1 port map( D => n1590, CK => net3496, Q => 
                           n502, QN => net48051);
   REGISTERS_reg_20_9_inst : DFF_X1 port map( D => n1612, CK => net3496, Q => 
                           n500, QN => net48050);
   REGISTERS_reg_20_8_inst : DFF_X1 port map( D => n1634, CK => net3496, Q => 
                           n499, QN => net48049);
   REGISTERS_reg_20_7_inst : DFF_X1 port map( D => n1656, CK => net3496, Q => 
                           n498, QN => net48048);
   REGISTERS_reg_20_6_inst : DFF_X1 port map( D => n1678, CK => net3496, Q => 
                           n497, QN => net48047);
   REGISTERS_reg_20_5_inst : DFF_X1 port map( D => n1700, CK => net3496, Q => 
                           n496, QN => net48046);
   REGISTERS_reg_20_4_inst : DFF_X1 port map( D => n1722, CK => net3496, Q => 
                           n495, QN => net48045);
   REGISTERS_reg_20_3_inst : DFF_X1 port map( D => n1744, CK => net3496, Q => 
                           n494, QN => net48044);
   REGISTERS_reg_20_2_inst : DFF_X1 port map( D => n1766, CK => net3496, Q => 
                           n493, QN => net48043);
   REGISTERS_reg_20_1_inst : DFF_X1 port map( D => n1788, CK => net3496, Q => 
                           n492, QN => net48042);
   REGISTERS_reg_20_0_inst : DFF_X1 port map( D => n1810, CK => net3496, Q => 
                           n491, QN => net48041);
   REGISTERS_reg_21_31_inst : DFF_X1 port map( D => n1094, CK => net3501, Q => 
                           n490, QN => net48040);
   REGISTERS_reg_21_30_inst : DFF_X1 port map( D => n1150, CK => net3501, Q => 
                           n489, QN => net48039);
   REGISTERS_reg_21_29_inst : DFF_X1 port map( D => n1172, CK => net3501, Q => 
                           n488, QN => net48038);
   REGISTERS_reg_21_28_inst : DFF_X1 port map( D => n1194, CK => net3501, Q => 
                           n487, QN => net48037);
   REGISTERS_reg_21_27_inst : DFF_X1 port map( D => n1216, CK => net3501, Q => 
                           n486, QN => net48036);
   REGISTERS_reg_21_26_inst : DFF_X1 port map( D => n1238, CK => net3501, Q => 
                           n485, QN => net48035);
   REGISTERS_reg_21_25_inst : DFF_X1 port map( D => n1260, CK => net3501, Q => 
                           n484, QN => net48034);
   REGISTERS_reg_21_24_inst : DFF_X1 port map( D => n1282, CK => net3501, Q => 
                           n483, QN => net48033);
   REGISTERS_reg_21_23_inst : DFF_X1 port map( D => n1304, CK => net3501, Q => 
                           n482, QN => net48032);
   REGISTERS_reg_21_22_inst : DFF_X1 port map( D => n1326, CK => net3501, Q => 
                           n481, QN => net48031);
   REGISTERS_reg_21_21_inst : DFF_X1 port map( D => n1348, CK => net3501, Q => 
                           n479, QN => net48030);
   REGISTERS_reg_21_20_inst : DFF_X1 port map( D => n1370, CK => net3501, Q => 
                           n478, QN => net48029);
   REGISTERS_reg_21_19_inst : DFF_X1 port map( D => n1392, CK => net3501, Q => 
                           n477, QN => net48028);
   REGISTERS_reg_21_18_inst : DFF_X1 port map( D => n1414, CK => net3501, Q => 
                           n476, QN => net48027);
   REGISTERS_reg_21_17_inst : DFF_X1 port map( D => n1436, CK => net3501, Q => 
                           n475, QN => net48026);
   REGISTERS_reg_21_16_inst : DFF_X1 port map( D => n1458, CK => net3501, Q => 
                           n474, QN => net48025);
   REGISTERS_reg_21_15_inst : DFF_X1 port map( D => n1480, CK => net3501, Q => 
                           n473, QN => net48024);
   REGISTERS_reg_21_14_inst : DFF_X1 port map( D => n1502, CK => net3501, Q => 
                           n472, QN => net48023);
   REGISTERS_reg_21_13_inst : DFF_X1 port map( D => n1524, CK => net3501, Q => 
                           n471, QN => net48022);
   REGISTERS_reg_21_12_inst : DFF_X1 port map( D => n1546, CK => net3501, Q => 
                           n470, QN => net48021);
   REGISTERS_reg_21_11_inst : DFF_X1 port map( D => n1568, CK => net3501, Q => 
                           n469, QN => net48020);
   REGISTERS_reg_21_10_inst : DFF_X1 port map( D => n1590, CK => net3501, Q => 
                           n468, QN => net48019);
   REGISTERS_reg_21_9_inst : DFF_X1 port map( D => n1612, CK => net3501, Q => 
                           n467, QN => net48018);
   REGISTERS_reg_21_8_inst : DFF_X1 port map( D => n1634, CK => net3501, Q => 
                           n466, QN => net48017);
   REGISTERS_reg_21_7_inst : DFF_X1 port map( D => n1656, CK => net3501, Q => 
                           n465, QN => net48016);
   REGISTERS_reg_21_6_inst : DFF_X1 port map( D => n1678, CK => net3501, Q => 
                           n464, QN => net48015);
   REGISTERS_reg_21_5_inst : DFF_X1 port map( D => n1700, CK => net3501, Q => 
                           n463, QN => net48014);
   REGISTERS_reg_21_4_inst : DFF_X1 port map( D => n1722, CK => net3501, Q => 
                           n462, QN => net48013);
   REGISTERS_reg_21_3_inst : DFF_X1 port map( D => n1744, CK => net3501, Q => 
                           n461, QN => net48012);
   REGISTERS_reg_21_2_inst : DFF_X1 port map( D => n1766, CK => net3501, Q => 
                           n460, QN => net48011);
   REGISTERS_reg_21_1_inst : DFF_X1 port map( D => n1788, CK => net3501, Q => 
                           n458, QN => net48010);
   REGISTERS_reg_21_0_inst : DFF_X1 port map( D => n1810, CK => net3501, Q => 
                           n457, QN => net48009);
   REGISTERS_reg_22_31_inst : DFF_X1 port map( D => n1094, CK => net3506, Q => 
                           n456, QN => net48008);
   REGISTERS_reg_22_30_inst : DFF_X1 port map( D => n1150, CK => net3506, Q => 
                           n455, QN => net48007);
   REGISTERS_reg_22_29_inst : DFF_X1 port map( D => n1172, CK => net3506, Q => 
                           n454, QN => net48006);
   REGISTERS_reg_22_28_inst : DFF_X1 port map( D => n1194, CK => net3506, Q => 
                           n453, QN => net48005);
   REGISTERS_reg_22_27_inst : DFF_X1 port map( D => n1216, CK => net3506, Q => 
                           n452, QN => net48004);
   REGISTERS_reg_22_26_inst : DFF_X1 port map( D => n1238, CK => net3506, Q => 
                           n451, QN => net48003);
   REGISTERS_reg_22_25_inst : DFF_X1 port map( D => n1260, CK => net3506, Q => 
                           n450, QN => net48002);
   REGISTERS_reg_22_24_inst : DFF_X1 port map( D => n1282, CK => net3506, Q => 
                           n449, QN => net48001);
   REGISTERS_reg_22_23_inst : DFF_X1 port map( D => n1304, CK => net3506, Q => 
                           n448, QN => net48000);
   REGISTERS_reg_22_22_inst : DFF_X1 port map( D => n1326, CK => net3506, Q => 
                           n447, QN => net47999);
   REGISTERS_reg_22_21_inst : DFF_X1 port map( D => n1348, CK => net3506, Q => 
                           n446, QN => net47998);
   REGISTERS_reg_22_20_inst : DFF_X1 port map( D => n1370, CK => net3506, Q => 
                           n445, QN => net47997);
   REGISTERS_reg_22_19_inst : DFF_X1 port map( D => n1392, CK => net3506, Q => 
                           n444, QN => net47996);
   REGISTERS_reg_22_18_inst : DFF_X1 port map( D => n1414, CK => net3506, Q => 
                           n443, QN => net47995);
   REGISTERS_reg_22_17_inst : DFF_X1 port map( D => n1436, CK => net3506, Q => 
                           n442, QN => net47994);
   REGISTERS_reg_22_16_inst : DFF_X1 port map( D => n1458, CK => net3506, Q => 
                           n441, QN => net47993);
   REGISTERS_reg_22_15_inst : DFF_X1 port map( D => n1480, CK => net3506, Q => 
                           n440, QN => net47992);
   REGISTERS_reg_22_14_inst : DFF_X1 port map( D => n1502, CK => net3506, Q => 
                           n439, QN => net47991);
   REGISTERS_reg_22_13_inst : DFF_X1 port map( D => n1524, CK => net3506, Q => 
                           n437, QN => net47990);
   REGISTERS_reg_22_12_inst : DFF_X1 port map( D => n1546, CK => net3506, Q => 
                           n436, QN => net47989);
   REGISTERS_reg_22_11_inst : DFF_X1 port map( D => n1568, CK => net3506, Q => 
                           n435, QN => net47988);
   REGISTERS_reg_22_10_inst : DFF_X1 port map( D => n1590, CK => net3506, Q => 
                           n434, QN => net47987);
   REGISTERS_reg_22_9_inst : DFF_X1 port map( D => n1612, CK => net3506, Q => 
                           n433, QN => net47986);
   REGISTERS_reg_22_8_inst : DFF_X1 port map( D => n1634, CK => net3506, Q => 
                           n432, QN => net47985);
   REGISTERS_reg_22_7_inst : DFF_X1 port map( D => n1656, CK => net3506, Q => 
                           n431, QN => net47984);
   REGISTERS_reg_22_6_inst : DFF_X1 port map( D => n1678, CK => net3506, Q => 
                           n430, QN => net47983);
   REGISTERS_reg_22_5_inst : DFF_X1 port map( D => n1700, CK => net3506, Q => 
                           n429, QN => net47982);
   REGISTERS_reg_22_4_inst : DFF_X1 port map( D => n1722, CK => net3506, Q => 
                           n428, QN => net47981);
   REGISTERS_reg_22_3_inst : DFF_X1 port map( D => n1744, CK => net3506, Q => 
                           n427, QN => net47980);
   REGISTERS_reg_22_2_inst : DFF_X1 port map( D => n1766, CK => net3506, Q => 
                           n426, QN => net47979);
   REGISTERS_reg_22_1_inst : DFF_X1 port map( D => n1788, CK => net3506, Q => 
                           n425, QN => net47978);
   REGISTERS_reg_22_0_inst : DFF_X1 port map( D => n1810, CK => net3506, Q => 
                           n424, QN => net47977);
   REGISTERS_reg_23_31_inst : DFF_X1 port map( D => n1094, CK => net3511, Q => 
                           n423, QN => net47976);
   REGISTERS_reg_23_30_inst : DFF_X1 port map( D => n1150, CK => net3511, Q => 
                           n422, QN => net47975);
   REGISTERS_reg_23_29_inst : DFF_X1 port map( D => n1172, CK => net3511, Q => 
                           n421, QN => net47974);
   REGISTERS_reg_23_28_inst : DFF_X1 port map( D => n1194, CK => net3511, Q => 
                           n420, QN => net47973);
   REGISTERS_reg_23_27_inst : DFF_X1 port map( D => n1216, CK => net3511, Q => 
                           n419, QN => net47972);
   REGISTERS_reg_23_26_inst : DFF_X1 port map( D => n1238, CK => net3511, Q => 
                           n418, QN => net47971);
   REGISTERS_reg_23_25_inst : DFF_X1 port map( D => n1260, CK => net3511, Q => 
                           n417, QN => net47970);
   REGISTERS_reg_23_24_inst : DFF_X1 port map( D => n1282, CK => net3511, Q => 
                           n416, QN => net47969);
   REGISTERS_reg_23_23_inst : DFF_X1 port map( D => n1304, CK => net3511, Q => 
                           n415, QN => net47968);
   REGISTERS_reg_23_22_inst : DFF_X1 port map( D => n1326, CK => net3511, Q => 
                           n414, QN => net47967);
   REGISTERS_reg_23_21_inst : DFF_X1 port map( D => n1348, CK => net3511, Q => 
                           n413, QN => net47966);
   REGISTERS_reg_23_20_inst : DFF_X1 port map( D => n1370, CK => net3511, Q => 
                           n412, QN => net47965);
   REGISTERS_reg_23_19_inst : DFF_X1 port map( D => n1392, CK => net3511, Q => 
                           n411, QN => net47964);
   REGISTERS_reg_23_18_inst : DFF_X1 port map( D => n1414, CK => net3511, Q => 
                           n410, QN => net47963);
   REGISTERS_reg_23_17_inst : DFF_X1 port map( D => n1436, CK => net3511, Q => 
                           n409, QN => net47962);
   REGISTERS_reg_23_16_inst : DFF_X1 port map( D => n1458, CK => net3511, Q => 
                           n408, QN => net47961);
   REGISTERS_reg_23_15_inst : DFF_X1 port map( D => n1480, CK => net3511, Q => 
                           n407, QN => net47960);
   REGISTERS_reg_23_14_inst : DFF_X1 port map( D => n1502, CK => net3511, Q => 
                           n406, QN => net47959);
   REGISTERS_reg_23_13_inst : DFF_X1 port map( D => n1524, CK => net3511, Q => 
                           n405, QN => net47958);
   REGISTERS_reg_23_12_inst : DFF_X1 port map( D => n1546, CK => net3511, Q => 
                           n404, QN => net47957);
   REGISTERS_reg_23_11_inst : DFF_X1 port map( D => n1568, CK => net3511, Q => 
                           n403, QN => net47956);
   REGISTERS_reg_23_10_inst : DFF_X1 port map( D => n1590, CK => net3511, Q => 
                           n402, QN => net47955);
   REGISTERS_reg_23_9_inst : DFF_X1 port map( D => n1612, CK => net3511, Q => 
                           n401, QN => net47954);
   REGISTERS_reg_23_8_inst : DFF_X1 port map( D => n1634, CK => net3511, Q => 
                           n400, QN => net47953);
   REGISTERS_reg_23_7_inst : DFF_X1 port map( D => n1656, CK => net3511, Q => 
                           n399, QN => net47952);
   REGISTERS_reg_23_6_inst : DFF_X1 port map( D => n1678, CK => net3511, Q => 
                           n398, QN => net47951);
   REGISTERS_reg_23_5_inst : DFF_X1 port map( D => n1700, CK => net3511, Q => 
                           n397, QN => net47950);
   REGISTERS_reg_23_4_inst : DFF_X1 port map( D => n1722, CK => net3511, Q => 
                           n396, QN => net47949);
   REGISTERS_reg_23_3_inst : DFF_X1 port map( D => n1744, CK => net3511, Q => 
                           n395, QN => net47948);
   REGISTERS_reg_23_2_inst : DFF_X1 port map( D => n1766, CK => net3511, Q => 
                           n394, QN => net47947);
   REGISTERS_reg_23_1_inst : DFF_X1 port map( D => n1788, CK => net3511, Q => 
                           n393, QN => net47946);
   REGISTERS_reg_23_0_inst : DFF_X1 port map( D => n1810, CK => net3511, Q => 
                           n392, QN => net47945);
   REGISTERS_reg_24_31_inst : DFF_X1 port map( D => n1094, CK => net3516, Q => 
                           n391, QN => net47944);
   REGISTERS_reg_24_30_inst : DFF_X1 port map( D => n1150, CK => net3516, Q => 
                           n390, QN => net47943);
   REGISTERS_reg_24_29_inst : DFF_X1 port map( D => n1172, CK => net3516, Q => 
                           n389, QN => net47942);
   REGISTERS_reg_24_28_inst : DFF_X1 port map( D => n1194, CK => net3516, Q => 
                           n388, QN => net47941);
   REGISTERS_reg_24_27_inst : DFF_X1 port map( D => n1216, CK => net3516, Q => 
                           n387, QN => net47940);
   REGISTERS_reg_24_26_inst : DFF_X1 port map( D => n1238, CK => net3516, Q => 
                           n386, QN => net47939);
   REGISTERS_reg_24_25_inst : DFF_X1 port map( D => n1260, CK => net3516, Q => 
                           n385, QN => net47938);
   REGISTERS_reg_24_24_inst : DFF_X1 port map( D => n1282, CK => net3516, Q => 
                           n384, QN => net47937);
   REGISTERS_reg_24_23_inst : DFF_X1 port map( D => n1304, CK => net3516, Q => 
                           n383, QN => net47936);
   REGISTERS_reg_24_22_inst : DFF_X1 port map( D => n1326, CK => net3516, Q => 
                           n382, QN => net47935);
   REGISTERS_reg_24_21_inst : DFF_X1 port map( D => n1348, CK => net3516, Q => 
                           n381, QN => net47934);
   REGISTERS_reg_24_20_inst : DFF_X1 port map( D => n1370, CK => net3516, Q => 
                           n380, QN => net47933);
   REGISTERS_reg_24_19_inst : DFF_X1 port map( D => n1392, CK => net3516, Q => 
                           n379, QN => net47932);
   REGISTERS_reg_24_18_inst : DFF_X1 port map( D => n1414, CK => net3516, Q => 
                           n378, QN => net47931);
   REGISTERS_reg_24_17_inst : DFF_X1 port map( D => n1436, CK => net3516, Q => 
                           n377, QN => net47930);
   REGISTERS_reg_24_16_inst : DFF_X1 port map( D => n1458, CK => net3516, Q => 
                           n376, QN => net47929);
   REGISTERS_reg_24_15_inst : DFF_X1 port map( D => n1480, CK => net3516, Q => 
                           n375, QN => net47928);
   REGISTERS_reg_24_14_inst : DFF_X1 port map( D => n1502, CK => net3516, Q => 
                           n374, QN => net47927);
   REGISTERS_reg_24_13_inst : DFF_X1 port map( D => n1524, CK => net3516, Q => 
                           n373, QN => net47926);
   REGISTERS_reg_24_12_inst : DFF_X1 port map( D => n1546, CK => net3516, Q => 
                           n372, QN => net47925);
   REGISTERS_reg_24_11_inst : DFF_X1 port map( D => n1568, CK => net3516, Q => 
                           n371, QN => net47924);
   REGISTERS_reg_24_10_inst : DFF_X1 port map( D => n1590, CK => net3516, Q => 
                           n370, QN => net47923);
   REGISTERS_reg_24_9_inst : DFF_X1 port map( D => n1612, CK => net3516, Q => 
                           n369, QN => net47922);
   REGISTERS_reg_24_8_inst : DFF_X1 port map( D => n1634, CK => net3516, Q => 
                           n368, QN => net47921);
   REGISTERS_reg_24_7_inst : DFF_X1 port map( D => n1656, CK => net3516, Q => 
                           n367, QN => net47920);
   REGISTERS_reg_24_6_inst : DFF_X1 port map( D => n1678, CK => net3516, Q => 
                           n366, QN => net47919);
   REGISTERS_reg_24_5_inst : DFF_X1 port map( D => n1700, CK => net3516, Q => 
                           n365, QN => net47918);
   REGISTERS_reg_24_4_inst : DFF_X1 port map( D => n1722, CK => net3516, Q => 
                           n364, QN => net47917);
   REGISTERS_reg_24_3_inst : DFF_X1 port map( D => n1744, CK => net3516, Q => 
                           n363, QN => net47916);
   REGISTERS_reg_24_2_inst : DFF_X1 port map( D => n1766, CK => net3516, Q => 
                           n362, QN => net47915);
   REGISTERS_reg_24_1_inst : DFF_X1 port map( D => n1788, CK => net3516, Q => 
                           n361, QN => net47914);
   REGISTERS_reg_24_0_inst : DFF_X1 port map( D => n1810, CK => net3516, Q => 
                           n360, QN => net47913);
   REGISTERS_reg_25_31_inst : DFF_X1 port map( D => n1094, CK => net3521, Q => 
                           n359, QN => net47912);
   REGISTERS_reg_25_30_inst : DFF_X1 port map( D => n1150, CK => net3521, Q => 
                           n358, QN => net47911);
   REGISTERS_reg_25_29_inst : DFF_X1 port map( D => n1172, CK => net3521, Q => 
                           n357, QN => net47910);
   REGISTERS_reg_25_28_inst : DFF_X1 port map( D => n1194, CK => net3521, Q => 
                           n356, QN => net47909);
   REGISTERS_reg_25_27_inst : DFF_X1 port map( D => n1216, CK => net3521, Q => 
                           n355, QN => net47908);
   REGISTERS_reg_25_26_inst : DFF_X1 port map( D => n1238, CK => net3521, Q => 
                           n354, QN => net47907);
   REGISTERS_reg_25_25_inst : DFF_X1 port map( D => n1260, CK => net3521, Q => 
                           n353, QN => net47906);
   REGISTERS_reg_25_24_inst : DFF_X1 port map( D => n1282, CK => net3521, Q => 
                           n352, QN => net47905);
   REGISTERS_reg_25_23_inst : DFF_X1 port map( D => n1304, CK => net3521, Q => 
                           n351, QN => net47904);
   REGISTERS_reg_25_22_inst : DFF_X1 port map( D => n1326, CK => net3521, Q => 
                           n350, QN => net47903);
   REGISTERS_reg_25_21_inst : DFF_X1 port map( D => n1348, CK => net3521, Q => 
                           n349, QN => net47902);
   REGISTERS_reg_25_20_inst : DFF_X1 port map( D => n1370, CK => net3521, Q => 
                           n348, QN => net47901);
   REGISTERS_reg_25_19_inst : DFF_X1 port map( D => n1392, CK => net3521, Q => 
                           n347, QN => net47900);
   REGISTERS_reg_25_18_inst : DFF_X1 port map( D => n1414, CK => net3521, Q => 
                           n346, QN => net47899);
   REGISTERS_reg_25_17_inst : DFF_X1 port map( D => n1436, CK => net3521, Q => 
                           n345, QN => net47898);
   REGISTERS_reg_25_16_inst : DFF_X1 port map( D => n1458, CK => net3521, Q => 
                           n344, QN => net47897);
   REGISTERS_reg_25_15_inst : DFF_X1 port map( D => n1480, CK => net3521, Q => 
                           n343, QN => net47896);
   REGISTERS_reg_25_14_inst : DFF_X1 port map( D => n1502, CK => net3521, Q => 
                           n342, QN => net47895);
   REGISTERS_reg_25_13_inst : DFF_X1 port map( D => n1524, CK => net3521, Q => 
                           n341, QN => net47894);
   REGISTERS_reg_25_12_inst : DFF_X1 port map( D => n1546, CK => net3521, Q => 
                           n340, QN => net47893);
   REGISTERS_reg_25_11_inst : DFF_X1 port map( D => n1568, CK => net3521, Q => 
                           n339, QN => net47892);
   REGISTERS_reg_25_10_inst : DFF_X1 port map( D => n1590, CK => net3521, Q => 
                           n338, QN => net47891);
   REGISTERS_reg_25_9_inst : DFF_X1 port map( D => n1612, CK => net3521, Q => 
                           n337, QN => net47890);
   REGISTERS_reg_25_8_inst : DFF_X1 port map( D => n1634, CK => net3521, Q => 
                           n336, QN => net47889);
   REGISTERS_reg_25_7_inst : DFF_X1 port map( D => n1656, CK => net3521, Q => 
                           n335, QN => net47888);
   REGISTERS_reg_25_6_inst : DFF_X1 port map( D => n1678, CK => net3521, Q => 
                           n334, QN => net47887);
   REGISTERS_reg_25_5_inst : DFF_X1 port map( D => n1700, CK => net3521, Q => 
                           n333, QN => net47886);
   REGISTERS_reg_25_4_inst : DFF_X1 port map( D => n1722, CK => net3521, Q => 
                           n332, QN => net47885);
   REGISTERS_reg_25_3_inst : DFF_X1 port map( D => n1744, CK => net3521, Q => 
                           n331, QN => net47884);
   REGISTERS_reg_25_2_inst : DFF_X1 port map( D => n1766, CK => net3521, Q => 
                           n330, QN => net47883);
   REGISTERS_reg_25_1_inst : DFF_X1 port map( D => n1788, CK => net3521, Q => 
                           n329, QN => net47882);
   REGISTERS_reg_25_0_inst : DFF_X1 port map( D => n1810, CK => net3521, Q => 
                           n328, QN => net47881);
   REGISTERS_reg_26_31_inst : DFF_X1 port map( D => n1094, CK => net3526, Q => 
                           n327, QN => net47880);
   REGISTERS_reg_26_30_inst : DFF_X1 port map( D => n1150, CK => net3526, Q => 
                           n326, QN => net47879);
   REGISTERS_reg_26_29_inst : DFF_X1 port map( D => n1172, CK => net3526, Q => 
                           n325, QN => net47878);
   REGISTERS_reg_26_28_inst : DFF_X1 port map( D => n1194, CK => net3526, Q => 
                           n324, QN => net47877);
   REGISTERS_reg_26_27_inst : DFF_X1 port map( D => n1216, CK => net3526, Q => 
                           n323, QN => net47876);
   REGISTERS_reg_26_26_inst : DFF_X1 port map( D => n1238, CK => net3526, Q => 
                           n322, QN => net47875);
   REGISTERS_reg_26_25_inst : DFF_X1 port map( D => n1260, CK => net3526, Q => 
                           n321, QN => net47874);
   REGISTERS_reg_26_24_inst : DFF_X1 port map( D => n1282, CK => net3526, Q => 
                           n320, QN => net47873);
   REGISTERS_reg_26_23_inst : DFF_X1 port map( D => n1304, CK => net3526, Q => 
                           n319, QN => net47872);
   REGISTERS_reg_26_22_inst : DFF_X1 port map( D => n1326, CK => net3526, Q => 
                           n318, QN => net47871);
   REGISTERS_reg_26_21_inst : DFF_X1 port map( D => n1348, CK => net3526, Q => 
                           n317, QN => net47870);
   REGISTERS_reg_26_20_inst : DFF_X1 port map( D => n1370, CK => net3526, Q => 
                           n316, QN => net47869);
   REGISTERS_reg_26_19_inst : DFF_X1 port map( D => n1392, CK => net3526, Q => 
                           n315, QN => net47868);
   REGISTERS_reg_26_18_inst : DFF_X1 port map( D => n1414, CK => net3526, Q => 
                           n314, QN => net47867);
   REGISTERS_reg_26_17_inst : DFF_X1 port map( D => n1436, CK => net3526, Q => 
                           n313, QN => net47866);
   REGISTERS_reg_26_16_inst : DFF_X1 port map( D => n1458, CK => net3526, Q => 
                           n312, QN => net47865);
   REGISTERS_reg_26_15_inst : DFF_X1 port map( D => n1480, CK => net3526, Q => 
                           n311, QN => net47864);
   REGISTERS_reg_26_14_inst : DFF_X1 port map( D => n1502, CK => net3526, Q => 
                           n310, QN => net47863);
   REGISTERS_reg_26_13_inst : DFF_X1 port map( D => n1524, CK => net3526, Q => 
                           n309, QN => net47862);
   REGISTERS_reg_26_12_inst : DFF_X1 port map( D => n1546, CK => net3526, Q => 
                           n308, QN => net47861);
   REGISTERS_reg_26_11_inst : DFF_X1 port map( D => n1568, CK => net3526, Q => 
                           n307, QN => net47860);
   REGISTERS_reg_26_10_inst : DFF_X1 port map( D => n1590, CK => net3526, Q => 
                           n306, QN => net47859);
   REGISTERS_reg_26_9_inst : DFF_X1 port map( D => n1612, CK => net3526, Q => 
                           n305, QN => net47858);
   REGISTERS_reg_26_8_inst : DFF_X1 port map( D => n1634, CK => net3526, Q => 
                           n304, QN => net47857);
   REGISTERS_reg_26_7_inst : DFF_X1 port map( D => n1656, CK => net3526, Q => 
                           n303, QN => net47856);
   REGISTERS_reg_26_6_inst : DFF_X1 port map( D => n1678, CK => net3526, Q => 
                           n302, QN => net47855);
   REGISTERS_reg_26_5_inst : DFF_X1 port map( D => n1700, CK => net3526, Q => 
                           n301, QN => net47854);
   REGISTERS_reg_26_4_inst : DFF_X1 port map( D => n1722, CK => net3526, Q => 
                           n300, QN => net47853);
   REGISTERS_reg_26_3_inst : DFF_X1 port map( D => n1744, CK => net3526, Q => 
                           n299, QN => net47852);
   REGISTERS_reg_26_2_inst : DFF_X1 port map( D => n1766, CK => net3526, Q => 
                           n298, QN => net47851);
   REGISTERS_reg_26_1_inst : DFF_X1 port map( D => n1788, CK => net3526, Q => 
                           n297, QN => net47850);
   REGISTERS_reg_26_0_inst : DFF_X1 port map( D => n1810, CK => net3526, Q => 
                           n296, QN => net47849);
   REGISTERS_reg_27_31_inst : DFF_X1 port map( D => n1094, CK => net3531, Q => 
                           n295, QN => net47848);
   REGISTERS_reg_27_30_inst : DFF_X1 port map( D => n1150, CK => net3531, Q => 
                           n294, QN => net47847);
   REGISTERS_reg_27_29_inst : DFF_X1 port map( D => n1172, CK => net3531, Q => 
                           n293, QN => net47846);
   REGISTERS_reg_27_28_inst : DFF_X1 port map( D => n1194, CK => net3531, Q => 
                           n292, QN => net47845);
   REGISTERS_reg_27_27_inst : DFF_X1 port map( D => n1216, CK => net3531, Q => 
                           n291, QN => net47844);
   REGISTERS_reg_27_26_inst : DFF_X1 port map( D => n1238, CK => net3531, Q => 
                           n290, QN => net47843);
   REGISTERS_reg_27_25_inst : DFF_X1 port map( D => n1260, CK => net3531, Q => 
                           n289, QN => net47842);
   REGISTERS_reg_27_24_inst : DFF_X1 port map( D => n1282, CK => net3531, Q => 
                           n288, QN => net47841);
   REGISTERS_reg_27_23_inst : DFF_X1 port map( D => n1304, CK => net3531, Q => 
                           n287, QN => net47840);
   REGISTERS_reg_27_22_inst : DFF_X1 port map( D => n1326, CK => net3531, Q => 
                           n286, QN => net47839);
   REGISTERS_reg_27_21_inst : DFF_X1 port map( D => n1348, CK => net3531, Q => 
                           n285, QN => net47838);
   REGISTERS_reg_27_20_inst : DFF_X1 port map( D => n1370, CK => net3531, Q => 
                           n284, QN => net47837);
   REGISTERS_reg_27_19_inst : DFF_X1 port map( D => n1392, CK => net3531, Q => 
                           n283, QN => net47836);
   REGISTERS_reg_27_18_inst : DFF_X1 port map( D => n1414, CK => net3531, Q => 
                           n282, QN => net47835);
   REGISTERS_reg_27_17_inst : DFF_X1 port map( D => n1436, CK => net3531, Q => 
                           n281, QN => net47834);
   REGISTERS_reg_27_16_inst : DFF_X1 port map( D => n1458, CK => net3531, Q => 
                           n280, QN => net47833);
   REGISTERS_reg_27_15_inst : DFF_X1 port map( D => n1480, CK => net3531, Q => 
                           n279, QN => net47832);
   REGISTERS_reg_27_14_inst : DFF_X1 port map( D => n1502, CK => net3531, Q => 
                           n278, QN => net47831);
   REGISTERS_reg_27_13_inst : DFF_X1 port map( D => n1524, CK => net3531, Q => 
                           n277, QN => net47830);
   REGISTERS_reg_27_12_inst : DFF_X1 port map( D => n1546, CK => net3531, Q => 
                           n276, QN => net47829);
   REGISTERS_reg_27_11_inst : DFF_X1 port map( D => n1568, CK => net3531, Q => 
                           n275, QN => net47828);
   REGISTERS_reg_27_10_inst : DFF_X1 port map( D => n1590, CK => net3531, Q => 
                           n274, QN => net47827);
   REGISTERS_reg_27_9_inst : DFF_X1 port map( D => n1612, CK => net3531, Q => 
                           n273, QN => net47826);
   REGISTERS_reg_27_8_inst : DFF_X1 port map( D => n1634, CK => net3531, Q => 
                           n272, QN => net47825);
   REGISTERS_reg_27_7_inst : DFF_X1 port map( D => n1656, CK => net3531, Q => 
                           n271, QN => net47824);
   REGISTERS_reg_27_6_inst : DFF_X1 port map( D => n1678, CK => net3531, Q => 
                           n270, QN => net47823);
   REGISTERS_reg_27_5_inst : DFF_X1 port map( D => n1700, CK => net3531, Q => 
                           n269, QN => net47822);
   REGISTERS_reg_27_4_inst : DFF_X1 port map( D => n1722, CK => net3531, Q => 
                           n268, QN => net47821);
   REGISTERS_reg_27_3_inst : DFF_X1 port map( D => n1744, CK => net3531, Q => 
                           n267, QN => net47820);
   REGISTERS_reg_27_2_inst : DFF_X1 port map( D => n1766, CK => net3531, Q => 
                           n266, QN => net47819);
   REGISTERS_reg_27_1_inst : DFF_X1 port map( D => n1788, CK => net3531, Q => 
                           n265, QN => net47818);
   REGISTERS_reg_27_0_inst : DFF_X1 port map( D => n1810, CK => net3531, Q => 
                           n264, QN => net47817);
   REGISTERS_reg_28_31_inst : DFF_X1 port map( D => n1094, CK => net3536, Q => 
                           n263, QN => net47816);
   REGISTERS_reg_28_30_inst : DFF_X1 port map( D => n1150, CK => net3536, Q => 
                           n262, QN => net47815);
   REGISTERS_reg_28_29_inst : DFF_X1 port map( D => n1172, CK => net3536, Q => 
                           n261, QN => net47814);
   REGISTERS_reg_28_28_inst : DFF_X1 port map( D => n1194, CK => net3536, Q => 
                           n260, QN => net47813);
   REGISTERS_reg_28_27_inst : DFF_X1 port map( D => n1216, CK => net3536, Q => 
                           n259, QN => net47812);
   REGISTERS_reg_28_26_inst : DFF_X1 port map( D => n1238, CK => net3536, Q => 
                           n258, QN => net47811);
   REGISTERS_reg_28_25_inst : DFF_X1 port map( D => n1260, CK => net3536, Q => 
                           n257, QN => net47810);
   REGISTERS_reg_28_24_inst : DFF_X1 port map( D => n1282, CK => net3536, Q => 
                           n256, QN => net47809);
   REGISTERS_reg_28_23_inst : DFF_X1 port map( D => n1304, CK => net3536, Q => 
                           n255, QN => net47808);
   REGISTERS_reg_28_22_inst : DFF_X1 port map( D => n1326, CK => net3536, Q => 
                           n254, QN => net47807);
   REGISTERS_reg_28_21_inst : DFF_X1 port map( D => n1348, CK => net3536, Q => 
                           n253, QN => net47806);
   REGISTERS_reg_28_20_inst : DFF_X1 port map( D => n1370, CK => net3536, Q => 
                           n252, QN => net47805);
   REGISTERS_reg_28_19_inst : DFF_X1 port map( D => n1392, CK => net3536, Q => 
                           n251, QN => net47804);
   REGISTERS_reg_28_18_inst : DFF_X1 port map( D => n1414, CK => net3536, Q => 
                           n250, QN => net47803);
   REGISTERS_reg_28_17_inst : DFF_X1 port map( D => n1436, CK => net3536, Q => 
                           n249, QN => net47802);
   REGISTERS_reg_28_16_inst : DFF_X1 port map( D => n1458, CK => net3536, Q => 
                           n248, QN => net47801);
   REGISTERS_reg_28_15_inst : DFF_X1 port map( D => n1480, CK => net3536, Q => 
                           n247, QN => net47800);
   REGISTERS_reg_28_14_inst : DFF_X1 port map( D => n1502, CK => net3536, Q => 
                           n246, QN => net47799);
   REGISTERS_reg_28_13_inst : DFF_X1 port map( D => n1524, CK => net3536, Q => 
                           n245, QN => net47798);
   REGISTERS_reg_28_12_inst : DFF_X1 port map( D => n1546, CK => net3536, Q => 
                           n244, QN => net47797);
   REGISTERS_reg_28_11_inst : DFF_X1 port map( D => n1568, CK => net3536, Q => 
                           n243, QN => net47796);
   REGISTERS_reg_28_10_inst : DFF_X1 port map( D => n1590, CK => net3536, Q => 
                           n242, QN => net47795);
   REGISTERS_reg_28_9_inst : DFF_X1 port map( D => n1612, CK => net3536, Q => 
                           n241, QN => net47794);
   REGISTERS_reg_28_8_inst : DFF_X1 port map( D => n1634, CK => net3536, Q => 
                           n240, QN => net47793);
   REGISTERS_reg_28_7_inst : DFF_X1 port map( D => n1656, CK => net3536, Q => 
                           n239, QN => net47792);
   REGISTERS_reg_28_6_inst : DFF_X1 port map( D => n1678, CK => net3536, Q => 
                           n238, QN => net47791);
   REGISTERS_reg_28_5_inst : DFF_X1 port map( D => n1700, CK => net3536, Q => 
                           n237, QN => net47790);
   REGISTERS_reg_28_4_inst : DFF_X1 port map( D => n1722, CK => net3536, Q => 
                           n236, QN => net47789);
   REGISTERS_reg_28_3_inst : DFF_X1 port map( D => n1744, CK => net3536, Q => 
                           n235, QN => net47788);
   REGISTERS_reg_28_2_inst : DFF_X1 port map( D => n1766, CK => net3536, Q => 
                           n234, QN => net47787);
   REGISTERS_reg_28_1_inst : DFF_X1 port map( D => n1788, CK => net3536, Q => 
                           n233, QN => net47786);
   REGISTERS_reg_28_0_inst : DFF_X1 port map( D => n1810, CK => net3536, Q => 
                           n232, QN => net47785);
   REGISTERS_reg_29_31_inst : DFF_X1 port map( D => n1094, CK => net3541, Q => 
                           n231, QN => net47784);
   REGISTERS_reg_29_30_inst : DFF_X1 port map( D => n1150, CK => net3541, Q => 
                           n230, QN => net47783);
   REGISTERS_reg_29_29_inst : DFF_X1 port map( D => n1172, CK => net3541, Q => 
                           n229, QN => net47782);
   REGISTERS_reg_29_28_inst : DFF_X1 port map( D => n1194, CK => net3541, Q => 
                           n228, QN => net47781);
   REGISTERS_reg_29_27_inst : DFF_X1 port map( D => n1216, CK => net3541, Q => 
                           n227, QN => net47780);
   REGISTERS_reg_29_26_inst : DFF_X1 port map( D => n1238, CK => net3541, Q => 
                           n226, QN => net47779);
   REGISTERS_reg_29_25_inst : DFF_X1 port map( D => n1260, CK => net3541, Q => 
                           n225, QN => net47778);
   REGISTERS_reg_29_24_inst : DFF_X1 port map( D => n1282, CK => net3541, Q => 
                           n224, QN => net47777);
   REGISTERS_reg_29_23_inst : DFF_X1 port map( D => n1304, CK => net3541, Q => 
                           n223, QN => net47776);
   REGISTERS_reg_29_22_inst : DFF_X1 port map( D => n1326, CK => net3541, Q => 
                           n222, QN => net47775);
   REGISTERS_reg_29_21_inst : DFF_X1 port map( D => n1348, CK => net3541, Q => 
                           n221, QN => net47774);
   REGISTERS_reg_29_20_inst : DFF_X1 port map( D => n1370, CK => net3541, Q => 
                           n220, QN => net47773);
   REGISTERS_reg_29_19_inst : DFF_X1 port map( D => n1392, CK => net3541, Q => 
                           n219, QN => net47772);
   REGISTERS_reg_29_18_inst : DFF_X1 port map( D => n1414, CK => net3541, Q => 
                           n218, QN => net47771);
   REGISTERS_reg_29_17_inst : DFF_X1 port map( D => n1436, CK => net3541, Q => 
                           n217, QN => net47770);
   REGISTERS_reg_29_16_inst : DFF_X1 port map( D => n1458, CK => net3541, Q => 
                           n216, QN => net47769);
   REGISTERS_reg_29_15_inst : DFF_X1 port map( D => n1480, CK => net3541, Q => 
                           n215, QN => net47768);
   REGISTERS_reg_29_14_inst : DFF_X1 port map( D => n1502, CK => net3541, Q => 
                           n214, QN => net47767);
   REGISTERS_reg_29_13_inst : DFF_X1 port map( D => n1524, CK => net3541, Q => 
                           n213, QN => net47766);
   REGISTERS_reg_29_12_inst : DFF_X1 port map( D => n1546, CK => net3541, Q => 
                           n212, QN => net47765);
   REGISTERS_reg_29_11_inst : DFF_X1 port map( D => n1568, CK => net3541, Q => 
                           n211, QN => net47764);
   REGISTERS_reg_29_10_inst : DFF_X1 port map( D => n1590, CK => net3541, Q => 
                           n210, QN => net47763);
   REGISTERS_reg_29_9_inst : DFF_X1 port map( D => n1612, CK => net3541, Q => 
                           n209, QN => net47762);
   REGISTERS_reg_29_8_inst : DFF_X1 port map( D => n1634, CK => net3541, Q => 
                           n208, QN => net47761);
   REGISTERS_reg_29_7_inst : DFF_X1 port map( D => n1656, CK => net3541, Q => 
                           n207, QN => net47760);
   REGISTERS_reg_29_6_inst : DFF_X1 port map( D => n1678, CK => net3541, Q => 
                           n206, QN => net47759);
   REGISTERS_reg_29_5_inst : DFF_X1 port map( D => n1700, CK => net3541, Q => 
                           n205, QN => net47758);
   REGISTERS_reg_29_4_inst : DFF_X1 port map( D => n1722, CK => net3541, Q => 
                           n204, QN => net47757);
   REGISTERS_reg_29_3_inst : DFF_X1 port map( D => n1744, CK => net3541, Q => 
                           n203, QN => net47756);
   REGISTERS_reg_29_2_inst : DFF_X1 port map( D => n1766, CK => net3541, Q => 
                           n202, QN => net47755);
   REGISTERS_reg_29_1_inst : DFF_X1 port map( D => n1788, CK => net3541, Q => 
                           n201, QN => net47754);
   REGISTERS_reg_29_0_inst : DFF_X1 port map( D => n1810, CK => net3541, Q => 
                           n200, QN => net47753);
   REGISTERS_reg_30_31_inst : DFF_X1 port map( D => n1094, CK => net3546, Q => 
                           n199, QN => net47752);
   REGISTERS_reg_30_30_inst : DFF_X1 port map( D => n1150, CK => net3546, Q => 
                           n198, QN => net47751);
   REGISTERS_reg_30_29_inst : DFF_X1 port map( D => n1172, CK => net3546, Q => 
                           n197, QN => net47750);
   REGISTERS_reg_30_28_inst : DFF_X1 port map( D => n1194, CK => net3546, Q => 
                           n196, QN => net47749);
   REGISTERS_reg_30_27_inst : DFF_X1 port map( D => n1216, CK => net3546, Q => 
                           n195, QN => net47748);
   REGISTERS_reg_30_26_inst : DFF_X1 port map( D => n1238, CK => net3546, Q => 
                           n194, QN => net47747);
   REGISTERS_reg_30_25_inst : DFF_X1 port map( D => n1260, CK => net3546, Q => 
                           n193, QN => net47746);
   REGISTERS_reg_30_24_inst : DFF_X1 port map( D => n1282, CK => net3546, Q => 
                           n192, QN => net47745);
   REGISTERS_reg_30_23_inst : DFF_X1 port map( D => n1304, CK => net3546, Q => 
                           n191, QN => net47744);
   REGISTERS_reg_30_22_inst : DFF_X1 port map( D => n1326, CK => net3546, Q => 
                           n190, QN => net47743);
   REGISTERS_reg_30_21_inst : DFF_X1 port map( D => n1348, CK => net3546, Q => 
                           n189, QN => net47742);
   REGISTERS_reg_30_20_inst : DFF_X1 port map( D => n1370, CK => net3546, Q => 
                           n188, QN => net47741);
   REGISTERS_reg_30_19_inst : DFF_X1 port map( D => n1392, CK => net3546, Q => 
                           n187, QN => net47740);
   REGISTERS_reg_30_18_inst : DFF_X1 port map( D => n1414, CK => net3546, Q => 
                           n186, QN => net47739);
   REGISTERS_reg_30_17_inst : DFF_X1 port map( D => n1436, CK => net3546, Q => 
                           n185, QN => net47738);
   REGISTERS_reg_30_16_inst : DFF_X1 port map( D => n1458, CK => net3546, Q => 
                           n184, QN => net47737);
   REGISTERS_reg_30_15_inst : DFF_X1 port map( D => n1480, CK => net3546, Q => 
                           n183, QN => net47736);
   REGISTERS_reg_30_14_inst : DFF_X1 port map( D => n1502, CK => net3546, Q => 
                           n182, QN => net47735);
   REGISTERS_reg_30_13_inst : DFF_X1 port map( D => n1524, CK => net3546, Q => 
                           n181, QN => net47734);
   REGISTERS_reg_30_12_inst : DFF_X1 port map( D => n1546, CK => net3546, Q => 
                           n180, QN => net47733);
   REGISTERS_reg_30_11_inst : DFF_X1 port map( D => n1568, CK => net3546, Q => 
                           n179, QN => net47732);
   REGISTERS_reg_30_10_inst : DFF_X1 port map( D => n1590, CK => net3546, Q => 
                           n178, QN => net47731);
   REGISTERS_reg_30_9_inst : DFF_X1 port map( D => n1612, CK => net3546, Q => 
                           n175, QN => net47730);
   REGISTERS_reg_30_8_inst : DFF_X1 port map( D => n1634, CK => net3546, Q => 
                           n164, QN => net47729);
   REGISTERS_reg_30_7_inst : DFF_X1 port map( D => n1656, CK => net3546, Q => 
                           n153, QN => net47728);
   REGISTERS_reg_30_6_inst : DFF_X1 port map( D => n1678, CK => net3546, Q => 
                           n142, QN => net47727);
   REGISTERS_reg_30_5_inst : DFF_X1 port map( D => n1700, CK => net3546, Q => 
                           n131, QN => net47726);
   REGISTERS_reg_30_4_inst : DFF_X1 port map( D => n1722, CK => net3546, Q => 
                           n120, QN => net47725);
   REGISTERS_reg_30_3_inst : DFF_X1 port map( D => n1744, CK => net3546, Q => 
                           n109, QN => net47724);
   REGISTERS_reg_30_2_inst : DFF_X1 port map( D => n1766, CK => net3546, Q => 
                           n97, QN => net47723);
   REGISTERS_reg_30_1_inst : DFF_X1 port map( D => n1788, CK => net3546, Q => 
                           n75, QN => net47722);
   REGISTERS_reg_30_0_inst : DFF_X1 port map( D => n1810, CK => net3546, Q => 
                           n53, QN => net47721);
   REGISTERS_reg_31_31_inst : DFF_X1 port map( D => n1094, CK => net3551, Q => 
                           n1089, QN => net47720);
   OUT2_reg_31_inst : DFF_X1 port map( D => N4616, CK => net3391, Q => OUT2(31)
                           , QN => n98);
   REGISTERS_reg_31_30_inst : DFF_X1 port map( D => n1150, CK => net3551, Q => 
                           n1068, QN => net47719);
   OUT2_reg_30_inst : DFF_X1 port map( D => N4614, CK => net3391, Q => OUT2(30)
                           , QN => n96);
   REGISTERS_reg_31_29_inst : DFF_X1 port map( D => n1172, CK => net3551, Q => 
                           n1047, QN => net47718);
   OUT2_reg_29_inst : DFF_X1 port map( D => N4612, CK => net3391, Q => OUT2(29)
                           , QN => n94);
   REGISTERS_reg_31_28_inst : DFF_X1 port map( D => n1194, CK => net3551, Q => 
                           n1026, QN => net47717);
   OUT2_reg_28_inst : DFF_X1 port map( D => N4610, CK => net3391, Q => OUT2(28)
                           , QN => n92);
   REGISTERS_reg_31_27_inst : DFF_X1 port map( D => n1216, CK => net3551, Q => 
                           n1005, QN => net47716);
   OUT2_reg_27_inst : DFF_X1 port map( D => N4608, CK => net3391, Q => OUT2(27)
                           , QN => n90);
   REGISTERS_reg_31_26_inst : DFF_X1 port map( D => n1238, CK => net3551, Q => 
                           n984, QN => net47715);
   OUT2_reg_26_inst : DFF_X1 port map( D => N4606, CK => net3391, Q => OUT2(26)
                           , QN => n88);
   REGISTERS_reg_31_25_inst : DFF_X1 port map( D => n1260, CK => net3551, Q => 
                           n963, QN => net47714);
   OUT2_reg_25_inst : DFF_X1 port map( D => N4604, CK => net3391, Q => OUT2(25)
                           , QN => n86);
   REGISTERS_reg_31_24_inst : DFF_X1 port map( D => n1282, CK => net3551, Q => 
                           n942, QN => net47713);
   OUT2_reg_24_inst : DFF_X1 port map( D => N4602, CK => net3391, Q => OUT2(24)
                           , QN => n84);
   REGISTERS_reg_31_23_inst : DFF_X1 port map( D => n1304, CK => net3551, Q => 
                           n921, QN => net47712);
   OUT2_reg_23_inst : DFF_X1 port map( D => N4600, CK => net3391, Q => OUT2(23)
                           , QN => n82);
   REGISTERS_reg_31_22_inst : DFF_X1 port map( D => n1326, CK => net3551, Q => 
                           n900, QN => net47711);
   OUT2_reg_22_inst : DFF_X1 port map( D => N4598, CK => net3391, Q => OUT2(22)
                           , QN => n80);
   REGISTERS_reg_31_21_inst : DFF_X1 port map( D => n1348, CK => net3551, Q => 
                           n879, QN => net47710);
   OUT2_reg_21_inst : DFF_X1 port map( D => N4596, CK => net3391, Q => OUT2(21)
                           , QN => n78);
   REGISTERS_reg_31_20_inst : DFF_X1 port map( D => n1370, CK => net3551, Q => 
                           n858, QN => net47709);
   OUT2_reg_20_inst : DFF_X1 port map( D => N4594, CK => net3391, Q => OUT2(20)
                           , QN => n76);
   REGISTERS_reg_31_19_inst : DFF_X1 port map( D => n1392, CK => net3551, Q => 
                           n837, QN => net47708);
   OUT2_reg_19_inst : DFF_X1 port map( D => N4592, CK => net3391, Q => OUT2(19)
                           , QN => n74);
   REGISTERS_reg_31_18_inst : DFF_X1 port map( D => n1414, CK => net3551, Q => 
                           n816, QN => net47707);
   OUT2_reg_18_inst : DFF_X1 port map( D => N4590, CK => net3391, Q => OUT2(18)
                           , QN => n72);
   REGISTERS_reg_31_17_inst : DFF_X1 port map( D => n1436, CK => net3551, Q => 
                           n795, QN => net47706);
   OUT2_reg_17_inst : DFF_X1 port map( D => N4588, CK => net3391, Q => OUT2(17)
                           , QN => n70);
   REGISTERS_reg_31_16_inst : DFF_X1 port map( D => n1458, CK => net3551, Q => 
                           n774, QN => net47705);
   OUT2_reg_16_inst : DFF_X1 port map( D => N4586, CK => net3391, Q => OUT2(16)
                           , QN => n68);
   REGISTERS_reg_31_15_inst : DFF_X1 port map( D => n1480, CK => net3551, Q => 
                           n753, QN => net47704);
   OUT2_reg_15_inst : DFF_X1 port map( D => N4584, CK => net3391, Q => OUT2(15)
                           , QN => n66);
   REGISTERS_reg_31_14_inst : DFF_X1 port map( D => n1502, CK => net3551, Q => 
                           n732, QN => net47703);
   OUT2_reg_14_inst : DFF_X1 port map( D => N4582, CK => net3391, Q => OUT2(14)
                           , QN => n64);
   REGISTERS_reg_31_13_inst : DFF_X1 port map( D => n1524, CK => net3551, Q => 
                           n711, QN => net47702);
   OUT2_reg_13_inst : DFF_X1 port map( D => N4580, CK => net3391, Q => OUT2(13)
                           , QN => n62);
   REGISTERS_reg_31_12_inst : DFF_X1 port map( D => n1546, CK => net3551, Q => 
                           n690, QN => net47701);
   OUT2_reg_12_inst : DFF_X1 port map( D => N4578, CK => net3391, Q => OUT2(12)
                           , QN => n60);
   REGISTERS_reg_31_11_inst : DFF_X1 port map( D => n1568, CK => net3551, Q => 
                           n669, QN => net47700);
   OUT2_reg_11_inst : DFF_X1 port map( D => N4576, CK => net3391, Q => OUT2(11)
                           , QN => n58);
   REGISTERS_reg_31_10_inst : DFF_X1 port map( D => n1590, CK => net3551, Q => 
                           n648, QN => net47699);
   OUT2_reg_10_inst : DFF_X1 port map( D => N4574, CK => net3391, Q => OUT2(10)
                           , QN => n56);
   REGISTERS_reg_31_9_inst : DFF_X1 port map( D => n1612, CK => net3551, Q => 
                           n627, QN => net47698);
   OUT2_reg_9_inst : DFF_X1 port map( D => N4572, CK => net3391, Q => OUT2(9), 
                           QN => n54);
   REGISTERS_reg_31_8_inst : DFF_X1 port map( D => n1634, CK => net3551, Q => 
                           n606, QN => net47697);
   OUT2_reg_8_inst : DFF_X1 port map( D => N4570, CK => net3391, Q => OUT2(8), 
                           QN => n52);
   REGISTERS_reg_31_7_inst : DFF_X1 port map( D => n1656, CK => net3551, Q => 
                           n585, QN => net47696);
   OUT2_reg_7_inst : DFF_X1 port map( D => N4568, CK => net3391, Q => OUT2(7), 
                           QN => n50);
   REGISTERS_reg_31_6_inst : DFF_X1 port map( D => n1678, CK => net3551, Q => 
                           n564, QN => net47695);
   OUT2_reg_6_inst : DFF_X1 port map( D => N4566, CK => net3391, Q => OUT2(6), 
                           QN => n48);
   REGISTERS_reg_31_5_inst : DFF_X1 port map( D => n1700, CK => net3551, Q => 
                           n543, QN => net47694);
   OUT2_reg_5_inst : DFF_X1 port map( D => N4564, CK => net3391, Q => OUT2(5), 
                           QN => n46);
   REGISTERS_reg_31_4_inst : DFF_X1 port map( D => n1722, CK => net3551, Q => 
                           n522, QN => net47693);
   OUT2_reg_4_inst : DFF_X1 port map( D => N4562, CK => net3391, Q => OUT2(4), 
                           QN => n44);
   REGISTERS_reg_31_3_inst : DFF_X1 port map( D => n1744, CK => net3551, Q => 
                           n501, QN => net47692);
   OUT2_reg_3_inst : DFF_X1 port map( D => N4560, CK => net3391, Q => OUT2(3), 
                           QN => n42);
   REGISTERS_reg_31_2_inst : DFF_X1 port map( D => n1766, CK => net3551, Q => 
                           n480, QN => net47691);
   OUT2_reg_2_inst : DFF_X1 port map( D => N4558, CK => net3391, Q => OUT2(2), 
                           QN => n40);
   REGISTERS_reg_31_1_inst : DFF_X1 port map( D => n1788, CK => net3551, Q => 
                           n459, QN => net47690);
   OUT2_reg_1_inst : DFF_X1 port map( D => N4556, CK => net3391, Q => OUT2(1), 
                           QN => n38);
   REGISTERS_reg_31_0_inst : DFF_X1 port map( D => n1810, CK => net3551, Q => 
                           n438, QN => net47689);
   OUT2_reg_0_inst : DFF_X1 port map( D => N4554, CK => net3391, Q => OUT2(0), 
                           QN => n36);
   OUT1_reg_31_inst : DFF_X1 port map( D => N4552, CK => net3556, Q => OUT1(31)
                           , QN => n35);
   OUT1_reg_30_inst : DFF_X1 port map( D => N4550, CK => net3556, Q => OUT1(30)
                           , QN => n34);
   OUT1_reg_29_inst : DFF_X1 port map( D => N4548, CK => net3556, Q => OUT1(29)
                           , QN => n33);
   OUT1_reg_28_inst : DFF_X1 port map( D => N4546, CK => net3556, Q => OUT1(28)
                           , QN => n32);
   OUT1_reg_27_inst : DFF_X1 port map( D => N4544, CK => net3556, Q => OUT1(27)
                           , QN => n31);
   OUT1_reg_26_inst : DFF_X1 port map( D => N4542, CK => net3556, Q => OUT1(26)
                           , QN => n30);
   OUT1_reg_25_inst : DFF_X1 port map( D => N4540, CK => net3556, Q => OUT1(25)
                           , QN => n29);
   OUT1_reg_24_inst : DFF_X1 port map( D => N4538, CK => net3556, Q => OUT1(24)
                           , QN => n28);
   OUT1_reg_23_inst : DFF_X1 port map( D => N4536, CK => net3556, Q => OUT1(23)
                           , QN => n27);
   OUT1_reg_22_inst : DFF_X1 port map( D => N4534, CK => net3556, Q => OUT1(22)
                           , QN => n26);
   OUT1_reg_21_inst : DFF_X1 port map( D => N4532, CK => net3556, Q => OUT1(21)
                           , QN => n25);
   OUT1_reg_20_inst : DFF_X1 port map( D => N4530, CK => net3556, Q => OUT1(20)
                           , QN => n24);
   OUT1_reg_19_inst : DFF_X1 port map( D => N4528, CK => net3556, Q => OUT1(19)
                           , QN => n23);
   OUT1_reg_18_inst : DFF_X1 port map( D => N4526, CK => net3556, Q => OUT1(18)
                           , QN => n22);
   OUT1_reg_17_inst : DFF_X1 port map( D => N4524, CK => net3556, Q => OUT1(17)
                           , QN => n21);
   OUT1_reg_16_inst : DFF_X1 port map( D => N4522, CK => net3556, Q => OUT1(16)
                           , QN => n20);
   OUT1_reg_15_inst : DFF_X1 port map( D => N4520, CK => net3556, Q => OUT1(15)
                           , QN => n19);
   OUT1_reg_14_inst : DFF_X1 port map( D => N4518, CK => net3556, Q => OUT1(14)
                           , QN => n18);
   OUT1_reg_13_inst : DFF_X1 port map( D => N4516, CK => net3556, Q => OUT1(13)
                           , QN => n17);
   OUT1_reg_12_inst : DFF_X1 port map( D => N4514, CK => net3556, Q => OUT1(12)
                           , QN => n16);
   OUT1_reg_11_inst : DFF_X1 port map( D => N4512, CK => net3556, Q => OUT1(11)
                           , QN => n15);
   OUT1_reg_10_inst : DFF_X1 port map( D => N4510, CK => net3556, Q => OUT1(10)
                           , QN => n14);
   OUT1_reg_9_inst : DFF_X1 port map( D => N4508, CK => net3556, Q => OUT1(9), 
                           QN => n13);
   OUT1_reg_8_inst : DFF_X1 port map( D => N4506, CK => net3556, Q => OUT1(8), 
                           QN => n12);
   OUT1_reg_7_inst : DFF_X1 port map( D => N4504, CK => net3556, Q => OUT1(7), 
                           QN => n11);
   OUT1_reg_6_inst : DFF_X1 port map( D => N4502, CK => net3556, Q => OUT1(6), 
                           QN => n10);
   OUT1_reg_5_inst : DFF_X1 port map( D => N4500, CK => net3556, Q => OUT1(5), 
                           QN => n9);
   OUT1_reg_4_inst : DFF_X1 port map( D => N4498, CK => net3556, Q => OUT1(4), 
                           QN => n8);
   OUT1_reg_3_inst : DFF_X1 port map( D => N4496, CK => net3556, Q => OUT1(3), 
                           QN => n7);
   OUT1_reg_2_inst : DFF_X1 port map( D => N4494, CK => net3556, Q => OUT1(2), 
                           QN => n6);
   OUT1_reg_1_inst : DFF_X1 port map( D => N4492, CK => net3556, Q => OUT1(1), 
                           QN => n5);
   OUT1_reg_0_inst : DFF_X1 port map( D => N4490, CK => net3556, Q => OUT1(0), 
                           QN => n4);
   clk_gate_OUT2_reg : SNPS_CLOCK_GATE_HIGH_dlx_regfile_0 port map( CLK => Clk,
                           EN => N4615, ENCLK => net3391);
   clk_gate_REGISTERS_reg_0_inst : SNPS_CLOCK_GATE_HIGH_dlx_regfile_33 port 
                           map( CLK => Clk, EN => Rst, ENCLK => net3396);
   clk_gate_REGISTERS_reg_1_inst : SNPS_CLOCK_GATE_HIGH_dlx_regfile_32 port 
                           map( CLK => Clk, EN => N4423, ENCLK => net3401);
   clk_gate_REGISTERS_reg_2_inst : SNPS_CLOCK_GATE_HIGH_dlx_regfile_31 port 
                           map( CLK => Clk, EN => N4359, ENCLK => net3406);
   clk_gate_REGISTERS_reg_3_inst : SNPS_CLOCK_GATE_HIGH_dlx_regfile_30 port 
                           map( CLK => Clk, EN => N4295, ENCLK => net3411);
   clk_gate_REGISTERS_reg_4_inst : SNPS_CLOCK_GATE_HIGH_dlx_regfile_29 port 
                           map( CLK => Clk, EN => N4231, ENCLK => net3416);
   clk_gate_REGISTERS_reg_5_inst : SNPS_CLOCK_GATE_HIGH_dlx_regfile_28 port 
                           map( CLK => Clk, EN => N4167, ENCLK => net3421);
   clk_gate_REGISTERS_reg_6_inst : SNPS_CLOCK_GATE_HIGH_dlx_regfile_27 port 
                           map( CLK => Clk, EN => N4103, ENCLK => net3426);
   clk_gate_REGISTERS_reg_7_inst : SNPS_CLOCK_GATE_HIGH_dlx_regfile_26 port 
                           map( CLK => Clk, EN => N4039, ENCLK => net3431);
   clk_gate_REGISTERS_reg_8_inst : SNPS_CLOCK_GATE_HIGH_dlx_regfile_25 port 
                           map( CLK => Clk, EN => N3975, ENCLK => net3436);
   clk_gate_REGISTERS_reg_9_inst : SNPS_CLOCK_GATE_HIGH_dlx_regfile_24 port 
                           map( CLK => Clk, EN => N3911, ENCLK => net3441);
   clk_gate_REGISTERS_reg_10_inst : SNPS_CLOCK_GATE_HIGH_dlx_regfile_23 port 
                           map( CLK => Clk, EN => N3847, ENCLK => net3446);
   clk_gate_REGISTERS_reg_11_inst : SNPS_CLOCK_GATE_HIGH_dlx_regfile_22 port 
                           map( CLK => Clk, EN => N3783, ENCLK => net3451);
   clk_gate_REGISTERS_reg_12_inst : SNPS_CLOCK_GATE_HIGH_dlx_regfile_21 port 
                           map( CLK => Clk, EN => N3719, ENCLK => net3456);
   clk_gate_REGISTERS_reg_13_inst : SNPS_CLOCK_GATE_HIGH_dlx_regfile_20 port 
                           map( CLK => Clk, EN => N3655, ENCLK => net3461);
   clk_gate_REGISTERS_reg_14_inst : SNPS_CLOCK_GATE_HIGH_dlx_regfile_19 port 
                           map( CLK => Clk, EN => N3591, ENCLK => net3466);
   clk_gate_REGISTERS_reg_15_inst : SNPS_CLOCK_GATE_HIGH_dlx_regfile_18 port 
                           map( CLK => Clk, EN => N3527, ENCLK => net3471);
   clk_gate_REGISTERS_reg_16_inst : SNPS_CLOCK_GATE_HIGH_dlx_regfile_17 port 
                           map( CLK => Clk, EN => N3463, ENCLK => net3476);
   clk_gate_REGISTERS_reg_17_inst : SNPS_CLOCK_GATE_HIGH_dlx_regfile_16 port 
                           map( CLK => Clk, EN => N3399, ENCLK => net3481);
   clk_gate_REGISTERS_reg_18_inst : SNPS_CLOCK_GATE_HIGH_dlx_regfile_15 port 
                           map( CLK => Clk, EN => N3335, ENCLK => net3486);
   clk_gate_REGISTERS_reg_19_inst : SNPS_CLOCK_GATE_HIGH_dlx_regfile_14 port 
                           map( CLK => Clk, EN => N3271, ENCLK => net3491);
   clk_gate_REGISTERS_reg_20_inst : SNPS_CLOCK_GATE_HIGH_dlx_regfile_13 port 
                           map( CLK => Clk, EN => N3207, ENCLK => net3496);
   clk_gate_REGISTERS_reg_21_inst : SNPS_CLOCK_GATE_HIGH_dlx_regfile_12 port 
                           map( CLK => Clk, EN => N3143, ENCLK => net3501);
   clk_gate_REGISTERS_reg_22_inst : SNPS_CLOCK_GATE_HIGH_dlx_regfile_11 port 
                           map( CLK => Clk, EN => N3079, ENCLK => net3506);
   clk_gate_REGISTERS_reg_23_inst : SNPS_CLOCK_GATE_HIGH_dlx_regfile_10 port 
                           map( CLK => Clk, EN => N3015, ENCLK => net3511);
   clk_gate_REGISTERS_reg_24_inst : SNPS_CLOCK_GATE_HIGH_dlx_regfile_9 port 
                           map( CLK => Clk, EN => N2951, ENCLK => net3516);
   clk_gate_REGISTERS_reg_25_inst : SNPS_CLOCK_GATE_HIGH_dlx_regfile_8 port 
                           map( CLK => Clk, EN => N2887, ENCLK => net3521);
   clk_gate_REGISTERS_reg_26_inst : SNPS_CLOCK_GATE_HIGH_dlx_regfile_7 port 
                           map( CLK => Clk, EN => N2823, ENCLK => net3526);
   clk_gate_REGISTERS_reg_27_inst : SNPS_CLOCK_GATE_HIGH_dlx_regfile_6 port 
                           map( CLK => Clk, EN => N2759, ENCLK => net3531);
   clk_gate_REGISTERS_reg_28_inst : SNPS_CLOCK_GATE_HIGH_dlx_regfile_5 port 
                           map( CLK => Clk, EN => N2695, ENCLK => net3536);
   clk_gate_REGISTERS_reg_29_inst : SNPS_CLOCK_GATE_HIGH_dlx_regfile_4 port 
                           map( CLK => Clk, EN => N2631, ENCLK => net3541);
   clk_gate_REGISTERS_reg_30_inst : SNPS_CLOCK_GATE_HIGH_dlx_regfile_3 port 
                           map( CLK => Clk, EN => N2567, ENCLK => net3546);
   clk_gate_REGISTERS_reg_31_inst : SNPS_CLOCK_GATE_HIGH_dlx_regfile_2 port 
                           map( CLK => Clk, EN => N2503, ENCLK => net3551);
   clk_gate_OUT1_reg : SNPS_CLOCK_GATE_HIGH_dlx_regfile_1 port map( CLK => Clk,
                           EN => N4615, ENCLK => net3556);
   U3 : INV_X1 port map( A => Rst, ZN => n51);
   U4 : INV_X1 port map( A => Rst, ZN => n47);
   U5 : INV_X2 port map( A => Rst, ZN => n49);
   U6 : NAND2_X2 port map( A1 => n49, A2 => n1868, ZN => n1867);
   U7 : NAND2_X2 port map( A1 => n47, A2 => n1103, ZN => n1102);
   U8 : NAND3_X2 port map( A1 => n1819, A2 => n1820, A3 => n1821, ZN => n1103);
   U9 : NAND3_X2 port map( A1 => n1819, A2 => n2553, A3 => n2554, ZN => n1868);
   U10 : NAND2_X2 port map( A1 => DATAIN(1), A2 => n49, ZN => n1788);
   U11 : NAND2_X2 port map( A1 => DATAIN(31), A2 => n47, ZN => n1094);
   U12 : NAND2_X2 port map( A1 => DATAIN(2), A2 => n49, ZN => n1766);
   U13 : NAND2_X2 port map( A1 => DATAIN(3), A2 => n51, ZN => n1744);
   U14 : NAND2_X2 port map( A1 => DATAIN(30), A2 => n47, ZN => n1150);
   U15 : NAND2_X2 port map( A1 => DATAIN(4), A2 => n51, ZN => n1722);
   U16 : NAND2_X2 port map( A1 => DATAIN(5), A2 => n51, ZN => n1700);
   U17 : NAND2_X2 port map( A1 => DATAIN(29), A2 => n47, ZN => n1172);
   U18 : NAND2_X2 port map( A1 => DATAIN(6), A2 => n51, ZN => n1678);
   U19 : NAND2_X2 port map( A1 => DATAIN(7), A2 => n51, ZN => n1656);
   U20 : NAND2_X2 port map( A1 => DATAIN(28), A2 => n47, ZN => n1194);
   U21 : NAND2_X2 port map( A1 => DATAIN(8), A2 => n51, ZN => n1634);
   U22 : NAND2_X2 port map( A1 => DATAIN(0), A2 => n47, ZN => n1810);
   U23 : NAND2_X2 port map( A1 => DATAIN(16), A2 => n49, ZN => n1458);
   U24 : NAND2_X2 port map( A1 => DATAIN(17), A2 => n49, ZN => n1436);
   U25 : NAND2_X2 port map( A1 => DATAIN(23), A2 => n49, ZN => n1304);
   U26 : NAND2_X2 port map( A1 => DATAIN(18), A2 => n49, ZN => n1414);
   U27 : NAND2_X2 port map( A1 => DATAIN(19), A2 => n49, ZN => n1392);
   U28 : NAND2_X2 port map( A1 => DATAIN(22), A2 => n49, ZN => n1326);
   U29 : NAND2_X2 port map( A1 => DATAIN(20), A2 => n49, ZN => n1370);
   U30 : NAND2_X2 port map( A1 => DATAIN(21), A2 => n49, ZN => n1348);
   U31 : NAND2_X2 port map( A1 => DATAIN(9), A2 => n51, ZN => n1612);
   U32 : NAND2_X2 port map( A1 => DATAIN(27), A2 => n47, ZN => n1216);
   U33 : NAND2_X2 port map( A1 => DATAIN(10), A2 => n51, ZN => n1590);
   U34 : NAND2_X2 port map( A1 => DATAIN(11), A2 => n51, ZN => n1568);
   U35 : NAND2_X2 port map( A1 => DATAIN(26), A2 => n49, ZN => n1238);
   U36 : NAND2_X2 port map( A1 => DATAIN(12), A2 => n51, ZN => n1546);
   U37 : NAND2_X2 port map( A1 => DATAIN(13), A2 => n51, ZN => n1524);
   U38 : NAND2_X2 port map( A1 => DATAIN(25), A2 => n49, ZN => n1260);
   U39 : NAND2_X2 port map( A1 => DATAIN(14), A2 => n51, ZN => n1502);
   U40 : NAND2_X2 port map( A1 => DATAIN(15), A2 => n49, ZN => n1480);
   U41 : NAND2_X2 port map( A1 => DATAIN(24), A2 => n49, ZN => n1282);
   U42 : BUF_X1 port map( A => n1154, Z => n3);
   U43 : BUF_X1 port map( A => n1153, Z => n2);
   U44 : BUF_X1 port map( A => n1142, Z => n1);
   U45 : BUF_X1 port map( A => n1156, Z => n37);
   U46 : BUF_X1 port map( A => n1918, Z => n43);
   U47 : BUF_X1 port map( A => n1907, Z => n39);
   U48 : BUF_X1 port map( A => n1917, Z => n41);
   U49 : BUF_X1 port map( A => n1920, Z => n45);
   U50 : NAND2_X2 port map( A1 => n2572, A2 => n2597, ZN => n1914);
   U51 : NAND2_X2 port map( A1 => n2575, A2 => n2597, ZN => n1916);
   U52 : NAND2_X2 port map( A1 => n2598, A2 => n2575, ZN => n1915);
   U53 : NAND2_X2 port map( A1 => n2591, A2 => n2577, ZN => n1908);
   U54 : NAND2_X2 port map( A1 => n2572, A2 => n2573, ZN => n1878);
   U55 : NAND2_X2 port map( A1 => n2572, A2 => n2574, ZN => n1877);
   U56 : NAND2_X2 port map( A1 => n2575, A2 => n2573, ZN => n1880);
   U57 : NAND2_X2 port map( A1 => n2575, A2 => n2574, ZN => n1879);
   U58 : NAND2_X2 port map( A1 => n2576, A2 => n2573, ZN => n1882);
   U59 : NAND2_X2 port map( A1 => n2576, A2 => n2574, ZN => n1881);
   U60 : NAND2_X2 port map( A1 => n2577, A2 => n2573, ZN => n1884);
   U61 : NAND2_X2 port map( A1 => n2577, A2 => n2574, ZN => n1883);
   U62 : NAND2_X2 port map( A1 => n2572, A2 => n2585, ZN => n1890);
   U63 : NAND2_X2 port map( A1 => n2572, A2 => n2586, ZN => n1889);
   U64 : NAND2_X2 port map( A1 => n2585, A2 => n2575, ZN => n1892);
   U65 : NAND2_X2 port map( A1 => n2586, A2 => n2575, ZN => n1891);
   U66 : NAND2_X2 port map( A1 => n2576, A2 => n2585, ZN => n1894);
   U67 : NAND2_X2 port map( A1 => n2576, A2 => n2586, ZN => n1893);
   U68 : NAND2_X2 port map( A1 => n2577, A2 => n2585, ZN => n1896);
   U69 : NAND2_X2 port map( A1 => n2577, A2 => n2586, ZN => n1895);
   U70 : NAND2_X2 port map( A1 => n2572, A2 => n2591, ZN => n1902);
   U71 : NAND2_X2 port map( A1 => n2572, A2 => n2592, ZN => n1901);
   U72 : NAND2_X2 port map( A1 => n2591, A2 => n2575, ZN => n1904);
   U73 : NAND2_X2 port map( A1 => n2575, A2 => n2592, ZN => n1903);
   U74 : NAND2_X2 port map( A1 => n2576, A2 => n2591, ZN => n1906);
   U75 : NAND2_X2 port map( A1 => n2576, A2 => n2592, ZN => n1905);
   U76 : NAND2_X2 port map( A1 => n1865, A2 => n1842, ZN => n1151);
   U77 : NAND2_X2 port map( A1 => n1842, A2 => n1864, ZN => n1152);
   U78 : NAND2_X2 port map( A1 => n1839, A2 => n1864, ZN => n1149);
   U79 : NAND2_X2 port map( A1 => n1858, A2 => n1844, ZN => n1143);
   U80 : NAND2_X2 port map( A1 => n1843, A2 => n1859, ZN => n1140);
   U81 : NAND2_X2 port map( A1 => n1843, A2 => n1858, ZN => n1141);
   U82 : NAND2_X2 port map( A1 => n1842, A2 => n1859, ZN => n1138);
   U83 : NAND2_X2 port map( A1 => n1858, A2 => n1842, ZN => n1139);
   U84 : NAND2_X2 port map( A1 => n1839, A2 => n1859, ZN => n1136);
   U85 : NAND2_X2 port map( A1 => n1839, A2 => n1858, ZN => n1137);
   U86 : NAND2_X2 port map( A1 => n1844, A2 => n1853, ZN => n1130);
   U87 : NAND2_X2 port map( A1 => n1844, A2 => n1852, ZN => n1131);
   U88 : NAND2_X2 port map( A1 => n1843, A2 => n1853, ZN => n1128);
   U89 : NAND2_X2 port map( A1 => n1843, A2 => n1852, ZN => n1129);
   U90 : NAND2_X2 port map( A1 => n1853, A2 => n1842, ZN => n1126);
   U91 : NAND2_X2 port map( A1 => n1852, A2 => n1842, ZN => n1127);
   U92 : NAND2_X2 port map( A1 => n1839, A2 => n1853, ZN => n1124);
   U93 : NAND2_X2 port map( A1 => n1839, A2 => n1852, ZN => n1125);
   U94 : NAND2_X2 port map( A1 => n1844, A2 => n1841, ZN => n1118);
   U95 : NAND2_X2 port map( A1 => n1844, A2 => n1840, ZN => n1119);
   U96 : NAND2_X2 port map( A1 => n1843, A2 => n1841, ZN => n1116);
   U97 : NAND2_X2 port map( A1 => n1843, A2 => n1840, ZN => n1117);
   U98 : NAND2_X2 port map( A1 => n1842, A2 => n1841, ZN => n1114);
   U99 : NAND2_X2 port map( A1 => n1842, A2 => n1840, ZN => n1115);
   U100 : NAND2_X2 port map( A1 => n1839, A2 => n1841, ZN => n1112);
   U101 : NAND2_X2 port map( A1 => n1839, A2 => n1840, ZN => n1113);
   U102 : NAND2_X2 port map( A1 => n1865, A2 => n1844, ZN => n1155);
   U103 : NAND2_X2 port map( A1 => n1865, A2 => n1839, ZN => n1148);
   U104 : NAND2_X2 port map( A1 => n2598, A2 => n2577, ZN => n1919);
   U105 : NAND2_X2 port map( A1 => n2598, A2 => n2572, ZN => n1913);
   U106 : AND4_X1 port map( A1 => n1334, A2 => n1335, A3 => n1336, A4 => n1337,
                           ZN => n1333);
   U107 : AND4_X1 port map( A1 => n1202, A2 => n1203, A3 => n1204, A4 => n1205,
                           ZN => n1201);
   U108 : AND4_X1 port map( A1 => n1268, A2 => n1269, A3 => n1270, A4 => n1271,
                           ZN => n1267);
   U109 : AND4_X1 port map( A1 => n1554, A2 => n1555, A3 => n1556, A4 => n1557,
                           ZN => n1553);
   U110 : AND4_X1 port map( A1 => n1180, A2 => n1181, A3 => n1182, A4 => n1183,
                           ZN => n1179);
   U111 : AND4_X1 port map( A1 => n1356, A2 => n1357, A3 => n1358, A4 => n1359,
                           ZN => n1355);
   U112 : AND4_X1 port map( A1 => n1224, A2 => n1225, A3 => n1226, A4 => n1227,
                           ZN => n1223);
   U113 : AND4_X1 port map( A1 => n1532, A2 => n1533, A3 => n1534, A4 => n1535,
                           ZN => n1531);
   U114 : AND4_X1 port map( A1 => n1312, A2 => n1313, A3 => n1314, A4 => n1315,
                           ZN => n1311);
   U115 : AND4_X1 port map( A1 => n1422, A2 => n1423, A3 => n1424, A4 => n1425,
                           ZN => n1421);
   U116 : AND4_X1 port map( A1 => n1444, A2 => n1445, A3 => n1446, A4 => n1447,
                           ZN => n1443);
   U117 : AND4_X1 port map( A1 => n1510, A2 => n1511, A3 => n1512, A4 => n1513,
                           ZN => n1509);
   U118 : AND4_X1 port map( A1 => n1158, A2 => n1159, A3 => n1160, A4 => n1161,
                           ZN => n1157);
   U119 : AND4_X1 port map( A1 => n1400, A2 => n1401, A3 => n1402, A4 => n1403,
                           ZN => n1399);
   U120 : AND4_X1 port map( A1 => n1378, A2 => n1379, A3 => n1380, A4 => n1381,
                           ZN => n1377);
   U121 : AND4_X1 port map( A1 => n1488, A2 => n1489, A3 => n1490, A4 => n1491,
                           ZN => n1487);
   U122 : AND4_X1 port map( A1 => n1104, A2 => n1105, A3 => n1106, A4 => n1107,
                           ZN => n1101);
   U123 : AND4_X1 port map( A1 => n1466, A2 => n1467, A3 => n1468, A4 => n1469,
                           ZN => n1465);
   U124 : AND4_X1 port map( A1 => n1290, A2 => n1291, A3 => n1292, A4 => n1293,
                           ZN => n1289);
   U125 : AND4_X1 port map( A1 => n2279, A2 => n2280, A3 => n2281, A4 => n2282,
                           ZN => n2278);
   U126 : AND4_X1 port map( A1 => n2300, A2 => n2301, A3 => n2302, A4 => n2303,
                           ZN => n2299);
   U127 : AND4_X1 port map( A1 => n2174, A2 => n2175, A3 => n2176, A4 => n2177,
                           ZN => n2173);
   U128 : AND4_X1 port map( A1 => n2258, A2 => n2259, A3 => n2260, A4 => n2261,
                           ZN => n2257);
   U129 : AND4_X1 port map( A1 => n2027, A2 => n2028, A3 => n2029, A4 => n2030,
                           ZN => n2026);
   U130 : AND4_X1 port map( A1 => n1964, A2 => n1965, A3 => n1966, A4 => n1967,
                           ZN => n1963);
   U131 : AND4_X1 port map( A1 => n1985, A2 => n1986, A3 => n1987, A4 => n1988,
                           ZN => n1984);
   U132 : AND4_X1 port map( A1 => n2237, A2 => n2238, A3 => n2239, A4 => n2240,
                           ZN => n2236);
   U133 : AND4_X1 port map( A1 => n1943, A2 => n1944, A3 => n1945, A4 => n1946,
                           ZN => n1942);
   U134 : AND4_X1 port map( A1 => n2216, A2 => n2217, A3 => n2218, A4 => n2219,
                           ZN => n2215);
   U135 : AND4_X1 port map( A1 => n2153, A2 => n2154, A3 => n2155, A4 => n2156,
                           ZN => n2152);
   U136 : AND4_X1 port map( A1 => n2195, A2 => n2196, A3 => n2197, A4 => n2198,
                           ZN => n2194);
   U137 : AND4_X1 port map( A1 => n2090, A2 => n2091, A3 => n2092, A4 => n2093,
                           ZN => n2089);
   U138 : AND4_X1 port map( A1 => n1922, A2 => n1923, A3 => n1924, A4 => n1925,
                           ZN => n1921);
   U139 : AND4_X1 port map( A1 => n2069, A2 => n2070, A3 => n2071, A4 => n2072,
                           ZN => n2068);
   U140 : AND4_X1 port map( A1 => n1869, A2 => n1870, A3 => n1871, A4 => n1872,
                           ZN => n1866);
   U141 : AND4_X1 port map( A1 => n2048, A2 => n2049, A3 => n2050, A4 => n2051,
                           ZN => n2047);
   U142 : AND4_X1 port map( A1 => n2132, A2 => n2133, A3 => n2134, A4 => n2135,
                           ZN => n2131);
   U143 : AND4_X1 port map( A1 => n2111, A2 => n2112, A3 => n2113, A4 => n2114,
                           ZN => n2110);
   U144 : INV_X1 port map( A => n1773, ZN => n1767);
   U145 : AND4_X1 port map( A1 => n1730, A2 => n1731, A3 => n1732, A4 => n1733,
                           ZN => n1729);
   U146 : AND4_X1 port map( A1 => n1664, A2 => n1665, A3 => n1666, A4 => n1667,
                           ZN => n1663);
   U147 : AND4_X1 port map( A1 => n1686, A2 => n1687, A3 => n1688, A4 => n1689,
                           ZN => n1685);
   U148 : AND4_X1 port map( A1 => n1775, A2 => n1776, A3 => n1777, A4 => n1778,
                           ZN => n1774);
   U149 : AND4_X1 port map( A1 => n1831, A2 => n1832, A3 => n1833, A4 => n1834,
                           ZN => n1818);
   U150 : AND4_X1 port map( A1 => n1797, A2 => n1798, A3 => n1799, A4 => n1800,
                           ZN => n1796);
   U151 : AND4_X1 port map( A1 => n1708, A2 => n1709, A3 => n1710, A4 => n1711,
                           ZN => n1707);
   U152 : AND4_X1 port map( A1 => n2447, A2 => n2448, A3 => n2449, A4 => n2450,
                           ZN => n2446);
   U153 : AND4_X1 port map( A1 => n2532, A2 => n2533, A3 => n2534, A4 => n2535,
                           ZN => n2531);
   U154 : AND4_X1 port map( A1 => n2511, A2 => n2512, A3 => n2513, A4 => n2514,
                           ZN => n2510);
   U155 : AND4_X1 port map( A1 => n2564, A2 => n2565, A3 => n2566, A4 => 
                           n2567_port, ZN => n2552);
   U156 : AND4_X1 port map( A1 => n2405, A2 => n2406, A3 => n2407, A4 => n2408,
                           ZN => n2404);
   U157 : AND4_X1 port map( A1 => n2468, A2 => n2469, A3 => n2470, A4 => n2471,
                           ZN => n2467);
   U158 : INV_X1 port map( A => n2509, ZN => n2503_port);
   U159 : AND4_X1 port map( A1 => n2426, A2 => n2427, A3 => n2428, A4 => n2429,
                           ZN => n2425);
   U160 : AND4_X1 port map( A1 => n1598, A2 => n1599, A3 => n1600, A4 => n1601,
                           ZN => n1597);
   U161 : AND4_X1 port map( A1 => n1642, A2 => n1643, A3 => n1644, A4 => n1645,
                           ZN => n1641);
   U162 : AND4_X1 port map( A1 => n1576, A2 => n1577, A3 => n1578, A4 => n1579,
                           ZN => n1575);
   U163 : AND4_X1 port map( A1 => n1620, A2 => n1621, A3 => n1622, A4 => n1623,
                           ZN => n1619);
   U164 : AND4_X1 port map( A1 => n1246, A2 => n1247, A3 => n1248, A4 => n1249,
                           ZN => n1245);
   U165 : INV_X1 port map( A => ADD_RD2(4), ZN => n1828);
   U166 : INV_X1 port map( A => ADD_RD2(3), ZN => n1845);
   U167 : AND2_X1 port map( A1 => ADD_RD2(1), A2 => ADD_RD2(2), ZN => n1839);
   U168 : AND2_X1 port map( A1 => n1822, A2 => ADD_RD2(2), ZN => n1842);
   U169 : INV_X1 port map( A => ADD_RD2(1), ZN => n1822);
   U170 : INV_X1 port map( A => ADD_RD2(0), ZN => n1846);
   U171 : AND4_X1 port map( A1 => n2384, A2 => n2385, A3 => n2386, A4 => n2387,
                           ZN => n2383);
   U172 : AND4_X1 port map( A1 => n2363, A2 => n2364, A3 => n2365, A4 => n2366,
                           ZN => n2362);
   U173 : AND4_X1 port map( A1 => n2321, A2 => n2322, A3 => n2323, A4 => n2324,
                           ZN => n2320);
   U174 : AND4_X1 port map( A1 => n2006, A2 => n2007, A3 => n2008, A4 => n2009,
                           ZN => n2005);
   U175 : INV_X1 port map( A => n2563, ZN => n2560);
   U176 : AND4_X1 port map( A1 => n2342, A2 => n2343, A3 => n2344, A4 => n2345,
                           ZN => n2341);
   U177 : INV_X1 port map( A => ADD_RD1(4), ZN => n2558);
   U178 : INV_X1 port map( A => ADD_RD1(3), ZN => n2578);
   U179 : AND2_X1 port map( A1 => ADD_RD1(1), A2 => ADD_RD1(2), ZN => n2572);
   U180 : AND2_X1 port map( A1 => n2555, A2 => ADD_RD1(2), ZN => n2575);
   U181 : INV_X1 port map( A => ADD_RD1(1), ZN => n2555);
   U182 : INV_X1 port map( A => ADD_RD1(0), ZN => n2579);
   U183 : INV_X1 port map( A => ADD_WR(0), ZN => n1826);
   U184 : OR3_X1 port map( A1 => n1829, A2 => n2562, A3 => ADD_WR(4), ZN => 
                           n2607);
   U185 : INV_X1 port map( A => ADD_WR(3), ZN => n1829);
   U186 : INV_X1 port map( A => ADD_WR(1), ZN => n1823);
   U187 : OR2_X1 port map( A1 => Rst, A2 => ENABLE, ZN => N4615);
   U188 : INV_X1 port map( A => ADD_WR(2), ZN => n1825);
   U189 : NOR2_X1 port map( A1 => ADD_RD2(2), A2 => n1822, ZN => n1843);
   U190 : AOI21_X1 port map( B1 => n2560, B2 => n2561, A => n2562, ZN => n1819)
                           ;
   U191 : NOR2_X1 port map( A1 => ADD_RD1(2), A2 => n2555, ZN => n2576);
   U192 : NOR2_X1 port map( A1 => ADD_RD2(1), A2 => ADD_RD2(2), ZN => n1844);
   U193 : NOR2_X1 port map( A1 => ADD_RD1(1), A2 => ADD_RD1(2), ZN => n2577);
   U194 : NOR2_X1 port map( A1 => ADD_WR(4), A2 => ADD_WR(3), ZN => n2561);
   U195 : AOI221_X1 port map( B1 => ADD_WR(1), B2 => n1822, C1 => n1823, C2 => 
                           ADD_RD2(1), A => n1824, ZN => n1821);
   U196 : NOR2_X1 port map( A1 => ADD_RD2(0), A2 => n1847, ZN => n1841);
   U197 : AOI221_X1 port map( B1 => ADD_WR(1), B2 => n2555, C1 => n1823, C2 => 
                           ADD_RD1(1), A => n2556, ZN => n2554);
   U198 : NOR2_X1 port map( A1 => ADD_RD1(0), A2 => n2580, ZN => n2574);
   U199 : NAND3_X1 port map( A1 => n1826, A2 => n1825, A3 => n1823, ZN => n2563
                           );
   U200 : OAI22_X1 port map( A1 => n1101, A2 => n1102, B1 => n1103, B2 => n1094
                           , ZN => N4616);
   U201 : NOR4_X1 port map( A1 => n1108, A2 => n1109, A3 => n1110, A4 => n1111,
                           ZN => n1107);
   U202 : OAI22_X1 port map( A1 => n199, A2 => n1112, B1 => n1089, B2 => n1113,
                           ZN => n1111);
   U203 : OAI22_X1 port map( A1 => n263, A2 => n1114, B1 => n231, B2 => n1115, 
                           ZN => n1110);
   U204 : OAI22_X1 port map( A1 => n327, A2 => n1116, B1 => n295, B2 => n1117, 
                           ZN => n1109);
   U205 : OAI22_X1 port map( A1 => n391, A2 => n1118, B1 => n359, B2 => n1119, 
                           ZN => n1108);
   U206 : NOR4_X1 port map( A1 => n1120, A2 => n1121, A3 => n1122, A4 => n1123,
                           ZN => n1106);
   U207 : OAI22_X1 port map( A1 => n456, A2 => n1124, B1 => n423, B2 => n1125, 
                           ZN => n1123);
   U208 : OAI22_X1 port map( A1 => n524, A2 => n1126, B1 => n490, B2 => n1127, 
                           ZN => n1122);
   U209 : OAI22_X1 port map( A1 => n591, A2 => n1128, B1 => n557, B2 => n1129, 
                           ZN => n1121);
   U210 : OAI22_X1 port map( A1 => n658, A2 => n1130, B1 => n624, B2 => n1131, 
                           ZN => n1120);
   U211 : NOR4_X1 port map( A1 => n1132, A2 => n1133, A3 => n1134, A4 => n1135,
                           ZN => n1105);
   U212 : OAI22_X1 port map( A1 => n725, A2 => n1136, B1 => n692, B2 => n1137, 
                           ZN => n1135);
   U213 : OAI22_X1 port map( A1 => n792, A2 => n1138, B1 => n759, B2 => n1139, 
                           ZN => n1134);
   U214 : OAI22_X1 port map( A1 => n860, A2 => n1140, B1 => n826, B2 => n1141, 
                           ZN => n1133);
   U215 : OAI22_X1 port map( A1 => n927, A2 => n1142, B1 => n893, B2 => n1143, 
                           ZN => n1132);
   U216 : NOR4_X1 port map( A1 => n1144, A2 => n1145, A3 => n1146, A4 => n1147,
                           ZN => n1104);
   U217 : OAI22_X1 port map( A1 => n994, A2 => n1148, B1 => n960, B2 => n1149, 
                           ZN => n1147);
   U218 : OAI22_X1 port map( A1 => n1061, A2 => n1151, B1 => n1028, B2 => n1152
                           , ZN => n1146);
   U219 : OAI22_X1 port map( A1 => n106, A2 => n2, B1 => n1096, B2 => n1154, ZN
                           => n1145);
   U220 : OAI22_X1 port map( A1 => n177, A2 => n1155, B1 => n141, B2 => n1156, 
                           ZN => n1144);
   U221 : OAI22_X1 port map( A1 => n1157, A2 => n1102, B1 => n1103, B2 => n1150
                           , ZN => N4614);
   U222 : NOR4_X1 port map( A1 => n1162, A2 => n1163, A3 => n1164, A4 => n1165,
                           ZN => n1161);
   U223 : OAI22_X1 port map( A1 => n198, A2 => n1112, B1 => n1068, B2 => n1113,
                           ZN => n1165);
   U224 : OAI22_X1 port map( A1 => n262, A2 => n1114, B1 => n230, B2 => n1115, 
                           ZN => n1164);
   U225 : OAI22_X1 port map( A1 => n326, A2 => n1116, B1 => n294, B2 => n1117, 
                           ZN => n1163);
   U226 : OAI22_X1 port map( A1 => n390, A2 => n1118, B1 => n358, B2 => n1119, 
                           ZN => n1162);
   U227 : NOR4_X1 port map( A1 => n1166, A2 => n1167, A3 => n1168, A4 => n1169,
                           ZN => n1160);
   U228 : OAI22_X1 port map( A1 => n455, A2 => n1124, B1 => n422, B2 => n1125, 
                           ZN => n1169);
   U229 : OAI22_X1 port map( A1 => n523, A2 => n1126, B1 => n489, B2 => n1127, 
                           ZN => n1168);
   U230 : OAI22_X1 port map( A1 => n590, A2 => n1128, B1 => n556, B2 => n1129, 
                           ZN => n1167);
   U231 : OAI22_X1 port map( A1 => n657, A2 => n1130, B1 => n623, B2 => n1131, 
                           ZN => n1166);
   U232 : NOR4_X1 port map( A1 => n1170, A2 => n1171, A3 => n1173, A4 => n1174,
                           ZN => n1159);
   U233 : OAI22_X1 port map( A1 => n724, A2 => n1136, B1 => n691, B2 => n1137, 
                           ZN => n1174);
   U234 : OAI22_X1 port map( A1 => n791, A2 => n1138, B1 => n758, B2 => n1139, 
                           ZN => n1173);
   U235 : OAI22_X1 port map( A1 => n859, A2 => n1140, B1 => n825, B2 => n1141, 
                           ZN => n1171);
   U236 : OAI22_X1 port map( A1 => n926, A2 => n1, B1 => n892, B2 => n1143, ZN 
                           => n1170);
   U237 : NOR4_X1 port map( A1 => n1175, A2 => n1176, A3 => n1177, A4 => n1178,
                           ZN => n1158);
   U238 : OAI22_X1 port map( A1 => n993, A2 => n1148, B1 => n959, B2 => n1149, 
                           ZN => n1178);
   U239 : OAI22_X1 port map( A1 => n1060, A2 => n1151, B1 => n1027, B2 => n1152
                           , ZN => n1177);
   U240 : OAI22_X1 port map( A1 => n105, A2 => n1153, B1 => n1095, B2 => n1154,
                           ZN => n1176);
   U241 : OAI22_X1 port map( A1 => n176, A2 => n1155, B1 => n140, B2 => n37, ZN
                           => n1175);
   U242 : OAI22_X1 port map( A1 => n1179, A2 => n1102, B1 => n1103, B2 => n1172
                           , ZN => N4612);
   U243 : NOR4_X1 port map( A1 => n1184, A2 => n1185, A3 => n1186, A4 => n1187,
                           ZN => n1183);
   U244 : OAI22_X1 port map( A1 => n197, A2 => n1112, B1 => n1047, B2 => n1113,
                           ZN => n1187);
   U245 : OAI22_X1 port map( A1 => n261, A2 => n1114, B1 => n229, B2 => n1115, 
                           ZN => n1186);
   U246 : OAI22_X1 port map( A1 => n325, A2 => n1116, B1 => n293, B2 => n1117, 
                           ZN => n1185);
   U247 : OAI22_X1 port map( A1 => n389, A2 => n1118, B1 => n357, B2 => n1119, 
                           ZN => n1184);
   U248 : NOR4_X1 port map( A1 => n1188, A2 => n1189, A3 => n1190, A4 => n1191,
                           ZN => n1182);
   U249 : OAI22_X1 port map( A1 => n454, A2 => n1124, B1 => n421, B2 => n1125, 
                           ZN => n1191);
   U250 : OAI22_X1 port map( A1 => n521, A2 => n1126, B1 => n488, B2 => n1127, 
                           ZN => n1190);
   U251 : OAI22_X1 port map( A1 => n589, A2 => n1128, B1 => n555, B2 => n1129, 
                           ZN => n1189);
   U252 : OAI22_X1 port map( A1 => n656, A2 => n1130, B1 => n622, B2 => n1131, 
                           ZN => n1188);
   U253 : NOR4_X1 port map( A1 => n1192, A2 => n1193, A3 => n1195, A4 => n1196,
                           ZN => n1181);
   U254 : OAI22_X1 port map( A1 => n723, A2 => n1136, B1 => n689, B2 => n1137, 
                           ZN => n1196);
   U255 : OAI22_X1 port map( A1 => n790, A2 => n1138, B1 => n757, B2 => n1139, 
                           ZN => n1195);
   U256 : OAI22_X1 port map( A1 => n857, A2 => n1140, B1 => n824, B2 => n1141, 
                           ZN => n1193);
   U257 : OAI22_X1 port map( A1 => n925, A2 => n1142, B1 => n891, B2 => n1143, 
                           ZN => n1192);
   U258 : NOR4_X1 port map( A1 => n1197, A2 => n1198, A3 => n1199, A4 => n1200,
                           ZN => n1180);
   U259 : OAI22_X1 port map( A1 => n992, A2 => n1148, B1 => n958, B2 => n1149, 
                           ZN => n1200);
   U260 : OAI22_X1 port map( A1 => n1059, A2 => n1151, B1 => n1025, B2 => n1152
                           , ZN => n1199);
   U261 : OAI22_X1 port map( A1 => n104, A2 => n1153, B1 => n1093, B2 => n1154,
                           ZN => n1198);
   U262 : OAI22_X1 port map( A1 => n174, A2 => n1155, B1 => n139, B2 => n37, ZN
                           => n1197);
   U263 : OAI22_X1 port map( A1 => n1201, A2 => n1102, B1 => n1103, B2 => n1194
                           , ZN => N4610);
   U264 : NOR4_X1 port map( A1 => n1206, A2 => n1207, A3 => n1208, A4 => n1209,
                           ZN => n1205);
   U265 : OAI22_X1 port map( A1 => n196, A2 => n1112, B1 => n1026, B2 => n1113,
                           ZN => n1209);
   U266 : OAI22_X1 port map( A1 => n260, A2 => n1114, B1 => n228, B2 => n1115, 
                           ZN => n1208);
   U267 : OAI22_X1 port map( A1 => n324, A2 => n1116, B1 => n292, B2 => n1117, 
                           ZN => n1207);
   U268 : OAI22_X1 port map( A1 => n388, A2 => n1118, B1 => n356, B2 => n1119, 
                           ZN => n1206);
   U269 : NOR4_X1 port map( A1 => n1210, A2 => n1211, A3 => n1212, A4 => n1213,
                           ZN => n1204);
   U270 : OAI22_X1 port map( A1 => n453, A2 => n1124, B1 => n420, B2 => n1125, 
                           ZN => n1213);
   U271 : OAI22_X1 port map( A1 => n520, A2 => n1126, B1 => n487, B2 => n1127, 
                           ZN => n1212);
   U272 : OAI22_X1 port map( A1 => n588, A2 => n1128, B1 => n554, B2 => n1129, 
                           ZN => n1211);
   U273 : OAI22_X1 port map( A1 => n655, A2 => n1130, B1 => n621, B2 => n1131, 
                           ZN => n1210);
   U274 : NOR4_X1 port map( A1 => n1214, A2 => n1215, A3 => n1217, A4 => n1218,
                           ZN => n1203);
   U275 : OAI22_X1 port map( A1 => n722, A2 => n1136, B1 => n688, B2 => n1137, 
                           ZN => n1218);
   U276 : OAI22_X1 port map( A1 => n789, A2 => n1138, B1 => n756, B2 => n1139, 
                           ZN => n1217);
   U277 : OAI22_X1 port map( A1 => n856, A2 => n1140, B1 => n823, B2 => n1141, 
                           ZN => n1215);
   U278 : OAI22_X1 port map( A1 => n924, A2 => n1142, B1 => n890, B2 => n1143, 
                           ZN => n1214);
   U279 : NOR4_X1 port map( A1 => n1219, A2 => n1220, A3 => n1221, A4 => n1222,
                           ZN => n1202);
   U280 : OAI22_X1 port map( A1 => n991, A2 => n1148, B1 => n957, B2 => n1149, 
                           ZN => n1222);
   U281 : OAI22_X1 port map( A1 => n1058, A2 => n1151, B1 => n1024, B2 => n1152
                           , ZN => n1221);
   U282 : OAI22_X1 port map( A1 => n103, A2 => n1153, B1 => n1092, B2 => n3, ZN
                           => n1220);
   U283 : OAI22_X1 port map( A1 => n173, A2 => n1155, B1 => n138, B2 => n37, ZN
                           => n1219);
   U284 : OAI22_X1 port map( A1 => n1223, A2 => n1102, B1 => n1103, B2 => n1216
                           , ZN => N4608);
   U285 : NOR4_X1 port map( A1 => n1228, A2 => n1229, A3 => n1230, A4 => n1231,
                           ZN => n1227);
   U286 : OAI22_X1 port map( A1 => n195, A2 => n1112, B1 => n1005, B2 => n1113,
                           ZN => n1231);
   U287 : OAI22_X1 port map( A1 => n259, A2 => n1114, B1 => n227, B2 => n1115, 
                           ZN => n1230);
   U288 : OAI22_X1 port map( A1 => n323, A2 => n1116, B1 => n291, B2 => n1117, 
                           ZN => n1229);
   U289 : OAI22_X1 port map( A1 => n387, A2 => n1118, B1 => n355, B2 => n1119, 
                           ZN => n1228);
   U290 : NOR4_X1 port map( A1 => n1232, A2 => n1233, A3 => n1234, A4 => n1235,
                           ZN => n1226);
   U291 : OAI22_X1 port map( A1 => n452, A2 => n1124, B1 => n419, B2 => n1125, 
                           ZN => n1235);
   U292 : OAI22_X1 port map( A1 => n519, A2 => n1126, B1 => n486, B2 => n1127, 
                           ZN => n1234);
   U293 : OAI22_X1 port map( A1 => n587, A2 => n1128, B1 => n553, B2 => n1129, 
                           ZN => n1233);
   U294 : OAI22_X1 port map( A1 => n654, A2 => n1130, B1 => n620, B2 => n1131, 
                           ZN => n1232);
   U295 : NOR4_X1 port map( A1 => n1236, A2 => n1237, A3 => n1239, A4 => n1240,
                           ZN => n1225);
   U296 : OAI22_X1 port map( A1 => n721, A2 => n1136, B1 => n687, B2 => n1137, 
                           ZN => n1240);
   U297 : OAI22_X1 port map( A1 => n788, A2 => n1138, B1 => n755, B2 => n1139, 
                           ZN => n1239);
   U298 : OAI22_X1 port map( A1 => n855, A2 => n1140, B1 => n822, B2 => n1141, 
                           ZN => n1237);
   U299 : OAI22_X1 port map( A1 => n923, A2 => n1142, B1 => n889, B2 => n1143, 
                           ZN => n1236);
   U300 : NOR4_X1 port map( A1 => n1241, A2 => n1242, A3 => n1243, A4 => n1244,
                           ZN => n1224);
   U301 : OAI22_X1 port map( A1 => n990, A2 => n1148, B1 => n956, B2 => n1149, 
                           ZN => n1244);
   U302 : OAI22_X1 port map( A1 => n1057, A2 => n1151, B1 => n1023, B2 => n1152
                           , ZN => n1243);
   U303 : OAI22_X1 port map( A1 => n102, A2 => n1153, B1 => n1091, B2 => n3, ZN
                           => n1242);
   U304 : OAI22_X1 port map( A1 => n172, A2 => n1155, B1 => n137, B2 => n37, ZN
                           => n1241);
   U305 : OAI22_X1 port map( A1 => n1245, A2 => n1102, B1 => n1103, B2 => n1238
                           , ZN => N4606);
   U306 : NOR4_X1 port map( A1 => n1250, A2 => n1251, A3 => n1252, A4 => n1253,
                           ZN => n1249);
   U307 : OAI22_X1 port map( A1 => n194, A2 => n1112, B1 => n984, B2 => n1113, 
                           ZN => n1253);
   U308 : OAI22_X1 port map( A1 => n258, A2 => n1114, B1 => n226, B2 => n1115, 
                           ZN => n1252);
   U309 : OAI22_X1 port map( A1 => n322, A2 => n1116, B1 => n290, B2 => n1117, 
                           ZN => n1251);
   U310 : OAI22_X1 port map( A1 => n386, A2 => n1118, B1 => n354, B2 => n1119, 
                           ZN => n1250);
   U311 : NOR4_X1 port map( A1 => n1254, A2 => n1255, A3 => n1256, A4 => n1257,
                           ZN => n1248);
   U312 : OAI22_X1 port map( A1 => n451, A2 => n1124, B1 => n418, B2 => n1125, 
                           ZN => n1257);
   U313 : OAI22_X1 port map( A1 => n518, A2 => n1126, B1 => n485, B2 => n1127, 
                           ZN => n1256);
   U314 : OAI22_X1 port map( A1 => n586, A2 => n1128, B1 => n552, B2 => n1129, 
                           ZN => n1255);
   U315 : OAI22_X1 port map( A1 => n653, A2 => n1130, B1 => n619, B2 => n1131, 
                           ZN => n1254);
   U316 : NOR4_X1 port map( A1 => n1258, A2 => n1259, A3 => n1261, A4 => n1262,
                           ZN => n1247);
   U317 : OAI22_X1 port map( A1 => n720, A2 => n1136, B1 => n686, B2 => n1137, 
                           ZN => n1262);
   U318 : OAI22_X1 port map( A1 => n787, A2 => n1138, B1 => n754, B2 => n1139, 
                           ZN => n1261);
   U319 : OAI22_X1 port map( A1 => n854, A2 => n1140, B1 => n821, B2 => n1141, 
                           ZN => n1259);
   U320 : OAI22_X1 port map( A1 => n922, A2 => n1142, B1 => n888, B2 => n1143, 
                           ZN => n1258);
   U321 : NOR4_X1 port map( A1 => n1263, A2 => n1264, A3 => n1265, A4 => n1266,
                           ZN => n1246);
   U322 : OAI22_X1 port map( A1 => n989, A2 => n1148, B1 => n955, B2 => n1149, 
                           ZN => n1266);
   U323 : OAI22_X1 port map( A1 => n1056, A2 => n1151, B1 => n1022, B2 => n1152
                           , ZN => n1265);
   U324 : OAI22_X1 port map( A1 => n101, A2 => n1153, B1 => n1090, B2 => n1154,
                           ZN => n1264);
   U325 : OAI22_X1 port map( A1 => n171, A2 => n1155, B1 => n136, B2 => n37, ZN
                           => n1263);
   U326 : OAI22_X1 port map( A1 => n1267, A2 => n1102, B1 => n1103, B2 => n1260
                           , ZN => N4604);
   U327 : NOR4_X1 port map( A1 => n1272, A2 => n1273, A3 => n1274, A4 => n1275,
                           ZN => n1271);
   U328 : OAI22_X1 port map( A1 => n193, A2 => n1112, B1 => n963, B2 => n1113, 
                           ZN => n1275);
   U329 : OAI22_X1 port map( A1 => n257, A2 => n1114, B1 => n225, B2 => n1115, 
                           ZN => n1274);
   U330 : OAI22_X1 port map( A1 => n321, A2 => n1116, B1 => n289, B2 => n1117, 
                           ZN => n1273);
   U331 : OAI22_X1 port map( A1 => n385, A2 => n1118, B1 => n353, B2 => n1119, 
                           ZN => n1272);
   U332 : NOR4_X1 port map( A1 => n1276, A2 => n1277, A3 => n1278, A4 => n1279,
                           ZN => n1270);
   U333 : OAI22_X1 port map( A1 => n450, A2 => n1124, B1 => n417, B2 => n1125, 
                           ZN => n1279);
   U334 : OAI22_X1 port map( A1 => n517, A2 => n1126, B1 => n484, B2 => n1127, 
                           ZN => n1278);
   U335 : OAI22_X1 port map( A1 => n584, A2 => n1128, B1 => n551, B2 => n1129, 
                           ZN => n1277);
   U336 : OAI22_X1 port map( A1 => n652, A2 => n1130, B1 => n618, B2 => n1131, 
                           ZN => n1276);
   U337 : NOR4_X1 port map( A1 => n1280, A2 => n1281, A3 => n1283, A4 => n1284,
                           ZN => n1269);
   U338 : OAI22_X1 port map( A1 => n719, A2 => n1136, B1 => n685, B2 => n1137, 
                           ZN => n1284);
   U339 : OAI22_X1 port map( A1 => n786, A2 => n1138, B1 => n752, B2 => n1139, 
                           ZN => n1283);
   U340 : OAI22_X1 port map( A1 => n853, A2 => n1140, B1 => n820, B2 => n1141, 
                           ZN => n1281);
   U341 : OAI22_X1 port map( A1 => n920, A2 => n1142, B1 => n887, B2 => n1143, 
                           ZN => n1280);
   U342 : NOR4_X1 port map( A1 => n1285, A2 => n1286, A3 => n1287, A4 => n1288,
                           ZN => n1268);
   U343 : OAI22_X1 port map( A1 => n988, A2 => n1148, B1 => n954, B2 => n1149, 
                           ZN => n1288);
   U344 : OAI22_X1 port map( A1 => n1055, A2 => n1151, B1 => n1021, B2 => n1152
                           , ZN => n1287);
   U345 : OAI22_X1 port map( A1 => n100, A2 => n1153, B1 => n1088, B2 => n3, ZN
                           => n1286);
   U346 : OAI22_X1 port map( A1 => n170, A2 => n1155, B1 => n135, B2 => n37, ZN
                           => n1285);
   U347 : OAI22_X1 port map( A1 => n1289, A2 => n1102, B1 => n1103, B2 => n1282
                           , ZN => N4602);
   U348 : NOR4_X1 port map( A1 => n1294, A2 => n1295, A3 => n1296, A4 => n1297,
                           ZN => n1293);
   U349 : OAI22_X1 port map( A1 => n192, A2 => n1112, B1 => n942, B2 => n1113, 
                           ZN => n1297);
   U350 : OAI22_X1 port map( A1 => n256, A2 => n1114, B1 => n224, B2 => n1115, 
                           ZN => n1296);
   U351 : OAI22_X1 port map( A1 => n320, A2 => n1116, B1 => n288, B2 => n1117, 
                           ZN => n1295);
   U352 : OAI22_X1 port map( A1 => n384, A2 => n1118, B1 => n352, B2 => n1119, 
                           ZN => n1294);
   U353 : NOR4_X1 port map( A1 => n1298, A2 => n1299, A3 => n1300, A4 => n1301,
                           ZN => n1292);
   U354 : OAI22_X1 port map( A1 => n449, A2 => n1124, B1 => n416, B2 => n1125, 
                           ZN => n1301);
   U355 : OAI22_X1 port map( A1 => n516, A2 => n1126, B1 => n483, B2 => n1127, 
                           ZN => n1300);
   U356 : OAI22_X1 port map( A1 => n583, A2 => n1128, B1 => n550, B2 => n1129, 
                           ZN => n1299);
   U357 : OAI22_X1 port map( A1 => n651, A2 => n1130, B1 => n617, B2 => n1131, 
                           ZN => n1298);
   U358 : NOR4_X1 port map( A1 => n1302, A2 => n1303, A3 => n1305, A4 => n1306,
                           ZN => n1291);
   U359 : OAI22_X1 port map( A1 => n718, A2 => n1136, B1 => n684, B2 => n1137, 
                           ZN => n1306);
   U360 : OAI22_X1 port map( A1 => n785, A2 => n1138, B1 => n751, B2 => n1139, 
                           ZN => n1305);
   U361 : OAI22_X1 port map( A1 => n852, A2 => n1140, B1 => n819, B2 => n1141, 
                           ZN => n1303);
   U362 : OAI22_X1 port map( A1 => n919, A2 => n1142, B1 => n886, B2 => n1143, 
                           ZN => n1302);
   U363 : NOR4_X1 port map( A1 => n1307, A2 => n1308, A3 => n1309, A4 => n1310,
                           ZN => n1290);
   U364 : OAI22_X1 port map( A1 => n987, A2 => n1148, B1 => n953, B2 => n1149, 
                           ZN => n1310);
   U365 : OAI22_X1 port map( A1 => n1054, A2 => n1151, B1 => n1020, B2 => n1152
                           , ZN => n1309);
   U366 : OAI22_X1 port map( A1 => n99, A2 => n1153, B1 => n1087, B2 => n1154, 
                           ZN => n1308);
   U367 : OAI22_X1 port map( A1 => n169, A2 => n1155, B1 => n134, B2 => n37, ZN
                           => n1307);
   U368 : OAI22_X1 port map( A1 => n1311, A2 => n1102, B1 => n1103, B2 => n1304
                           , ZN => N4600);
   U369 : NOR4_X1 port map( A1 => n1316, A2 => n1317, A3 => n1318, A4 => n1319,
                           ZN => n1315);
   U370 : OAI22_X1 port map( A1 => n191, A2 => n1112, B1 => n921, B2 => n1113, 
                           ZN => n1319);
   U371 : OAI22_X1 port map( A1 => n255, A2 => n1114, B1 => n223, B2 => n1115, 
                           ZN => n1318);
   U372 : OAI22_X1 port map( A1 => n319, A2 => n1116, B1 => n287, B2 => n1117, 
                           ZN => n1317);
   U373 : OAI22_X1 port map( A1 => n383, A2 => n1118, B1 => n351, B2 => n1119, 
                           ZN => n1316);
   U374 : NOR4_X1 port map( A1 => n1320, A2 => n1321, A3 => n1322, A4 => n1323,
                           ZN => n1314);
   U375 : OAI22_X1 port map( A1 => n448, A2 => n1124, B1 => n415, B2 => n1125, 
                           ZN => n1323);
   U376 : OAI22_X1 port map( A1 => n515, A2 => n1126, B1 => n482, B2 => n1127, 
                           ZN => n1322);
   U377 : OAI22_X1 port map( A1 => n582, A2 => n1128, B1 => n549, B2 => n1129, 
                           ZN => n1321);
   U378 : OAI22_X1 port map( A1 => n650, A2 => n1130, B1 => n616, B2 => n1131, 
                           ZN => n1320);
   U379 : NOR4_X1 port map( A1 => n1324, A2 => n1325, A3 => n1327, A4 => n1328,
                           ZN => n1313);
   U380 : OAI22_X1 port map( A1 => n717, A2 => n1136, B1 => n683, B2 => n1137, 
                           ZN => n1328);
   U381 : OAI22_X1 port map( A1 => n784, A2 => n1138, B1 => n750, B2 => n1139, 
                           ZN => n1327);
   U382 : OAI22_X1 port map( A1 => n851, A2 => n1140, B1 => n818, B2 => n1141, 
                           ZN => n1325);
   U383 : OAI22_X1 port map( A1 => n918, A2 => n1142, B1 => n885, B2 => n1143, 
                           ZN => n1324);
   U384 : NOR4_X1 port map( A1 => n1329, A2 => n1330, A3 => n1331, A4 => n1332,
                           ZN => n1312);
   U385 : OAI22_X1 port map( A1 => n986, A2 => n1148, B1 => n952, B2 => n1149, 
                           ZN => n1332);
   U386 : OAI22_X1 port map( A1 => n1053, A2 => n1151, B1 => n1019, B2 => n1152
                           , ZN => n1331);
   U387 : OAI22_X1 port map( A1 => n95, A2 => n1153, B1 => n1086, B2 => n3, ZN 
                           => n1330);
   U388 : OAI22_X1 port map( A1 => n168, A2 => n1155, B1 => n133, B2 => n37, ZN
                           => n1329);
   U389 : OAI22_X1 port map( A1 => n1333, A2 => n1102, B1 => n1103, B2 => n1326
                           , ZN => N4598);
   U390 : NOR4_X1 port map( A1 => n1338, A2 => n1339, A3 => n1340, A4 => n1341,
                           ZN => n1337);
   U391 : OAI22_X1 port map( A1 => n190, A2 => n1112, B1 => n900, B2 => n1113, 
                           ZN => n1341);
   U392 : OAI22_X1 port map( A1 => n254, A2 => n1114, B1 => n222, B2 => n1115, 
                           ZN => n1340);
   U393 : OAI22_X1 port map( A1 => n318, A2 => n1116, B1 => n286, B2 => n1117, 
                           ZN => n1339);
   U394 : OAI22_X1 port map( A1 => n382, A2 => n1118, B1 => n350, B2 => n1119, 
                           ZN => n1338);
   U395 : NOR4_X1 port map( A1 => n1342, A2 => n1343, A3 => n1344, A4 => n1345,
                           ZN => n1336);
   U396 : OAI22_X1 port map( A1 => n447, A2 => n1124, B1 => n414, B2 => n1125, 
                           ZN => n1345);
   U397 : OAI22_X1 port map( A1 => n514, A2 => n1126, B1 => n481, B2 => n1127, 
                           ZN => n1344);
   U398 : OAI22_X1 port map( A1 => n581, A2 => n1128, B1 => n548, B2 => n1129, 
                           ZN => n1343);
   U399 : OAI22_X1 port map( A1 => n649, A2 => n1130, B1 => n615, B2 => n1131, 
                           ZN => n1342);
   U400 : NOR4_X1 port map( A1 => n1346, A2 => n1347, A3 => n1349, A4 => n1350,
                           ZN => n1335);
   U401 : OAI22_X1 port map( A1 => n716, A2 => n1136, B1 => n682, B2 => n1137, 
                           ZN => n1350);
   U402 : OAI22_X1 port map( A1 => n783, A2 => n1138, B1 => n749, B2 => n1139, 
                           ZN => n1349);
   U403 : OAI22_X1 port map( A1 => n850, A2 => n1140, B1 => n817, B2 => n1141, 
                           ZN => n1347);
   U404 : OAI22_X1 port map( A1 => n917, A2 => n1142, B1 => n884, B2 => n1143, 
                           ZN => n1346);
   U405 : NOR4_X1 port map( A1 => n1351, A2 => n1352, A3 => n1353, A4 => n1354,
                           ZN => n1334);
   U406 : OAI22_X1 port map( A1 => n985, A2 => n1148, B1 => n951, B2 => n1149, 
                           ZN => n1354);
   U407 : OAI22_X1 port map( A1 => n1052, A2 => n1151, B1 => n1018, B2 => n1152
                           , ZN => n1353);
   U408 : OAI22_X1 port map( A1 => n93, A2 => n1153, B1 => n1085, B2 => n3, ZN 
                           => n1352);
   U409 : OAI22_X1 port map( A1 => n167, A2 => n1155, B1 => n132, B2 => n37, ZN
                           => n1351);
   U410 : OAI22_X1 port map( A1 => n1355, A2 => n1102, B1 => n1103, B2 => n1348
                           , ZN => N4596);
   U411 : NOR4_X1 port map( A1 => n1360, A2 => n1361, A3 => n1362, A4 => n1363,
                           ZN => n1359);
   U412 : OAI22_X1 port map( A1 => n189, A2 => n1112, B1 => n879, B2 => n1113, 
                           ZN => n1363);
   U413 : OAI22_X1 port map( A1 => n253, A2 => n1114, B1 => n221, B2 => n1115, 
                           ZN => n1362);
   U414 : OAI22_X1 port map( A1 => n317, A2 => n1116, B1 => n285, B2 => n1117, 
                           ZN => n1361);
   U415 : OAI22_X1 port map( A1 => n381, A2 => n1118, B1 => n349, B2 => n1119, 
                           ZN => n1360);
   U416 : NOR4_X1 port map( A1 => n1364, A2 => n1365, A3 => n1366, A4 => n1367,
                           ZN => n1358);
   U417 : OAI22_X1 port map( A1 => n446, A2 => n1124, B1 => n413, B2 => n1125, 
                           ZN => n1367);
   U418 : OAI22_X1 port map( A1 => n513, A2 => n1126, B1 => n479, B2 => n1127, 
                           ZN => n1366);
   U419 : OAI22_X1 port map( A1 => n580, A2 => n1128, B1 => n547, B2 => n1129, 
                           ZN => n1365);
   U420 : OAI22_X1 port map( A1 => n647, A2 => n1130, B1 => n614, B2 => n1131, 
                           ZN => n1364);
   U421 : NOR4_X1 port map( A1 => n1368, A2 => n1369, A3 => n1371, A4 => n1372,
                           ZN => n1357);
   U422 : OAI22_X1 port map( A1 => n715, A2 => n1136, B1 => n681, B2 => n1137, 
                           ZN => n1372);
   U423 : OAI22_X1 port map( A1 => n782, A2 => n1138, B1 => n748, B2 => n1139, 
                           ZN => n1371);
   U424 : OAI22_X1 port map( A1 => n849, A2 => n1140, B1 => n815, B2 => n1141, 
                           ZN => n1369);
   U425 : OAI22_X1 port map( A1 => n916, A2 => n1142, B1 => n883, B2 => n1143, 
                           ZN => n1368);
   U426 : NOR4_X1 port map( A1 => n1373, A2 => n1374, A3 => n1375, A4 => n1376,
                           ZN => n1356);
   U427 : OAI22_X1 port map( A1 => n983, A2 => n1148, B1 => n950, B2 => n1149, 
                           ZN => n1376);
   U428 : OAI22_X1 port map( A1 => n1051, A2 => n1151, B1 => n1017, B2 => n1152
                           , ZN => n1375);
   U429 : OAI22_X1 port map( A1 => n91, A2 => n1153, B1 => n1084, B2 => n3, ZN 
                           => n1374);
   U430 : OAI22_X1 port map( A1 => n166, A2 => n1155, B1 => n130, B2 => n37, ZN
                           => n1373);
   U431 : OAI22_X1 port map( A1 => n1377, A2 => n1102, B1 => n1103, B2 => n1370
                           , ZN => N4594);
   U432 : NOR4_X1 port map( A1 => n1382, A2 => n1383, A3 => n1384, A4 => n1385,
                           ZN => n1381);
   U433 : OAI22_X1 port map( A1 => n188, A2 => n1112, B1 => n858, B2 => n1113, 
                           ZN => n1385);
   U434 : OAI22_X1 port map( A1 => n252, A2 => n1114, B1 => n220, B2 => n1115, 
                           ZN => n1384);
   U435 : OAI22_X1 port map( A1 => n316, A2 => n1116, B1 => n284, B2 => n1117, 
                           ZN => n1383);
   U436 : OAI22_X1 port map( A1 => n380, A2 => n1118, B1 => n348, B2 => n1119, 
                           ZN => n1382);
   U437 : NOR4_X1 port map( A1 => n1386, A2 => n1387, A3 => n1388, A4 => n1389,
                           ZN => n1380);
   U438 : OAI22_X1 port map( A1 => n445, A2 => n1124, B1 => n412, B2 => n1125, 
                           ZN => n1389);
   U439 : OAI22_X1 port map( A1 => n512, A2 => n1126, B1 => n478, B2 => n1127, 
                           ZN => n1388);
   U440 : OAI22_X1 port map( A1 => n579, A2 => n1128, B1 => n546, B2 => n1129, 
                           ZN => n1387);
   U441 : OAI22_X1 port map( A1 => n646, A2 => n1130, B1 => n613, B2 => n1131, 
                           ZN => n1386);
   U442 : NOR4_X1 port map( A1 => n1390, A2 => n1391, A3 => n1393, A4 => n1394,
                           ZN => n1379);
   U443 : OAI22_X1 port map( A1 => n714, A2 => n1136, B1 => n680, B2 => n1137, 
                           ZN => n1394);
   U444 : OAI22_X1 port map( A1 => n781, A2 => n1138, B1 => n747, B2 => n1139, 
                           ZN => n1393);
   U445 : OAI22_X1 port map( A1 => n848, A2 => n1140, B1 => n814, B2 => n1141, 
                           ZN => n1391);
   U446 : OAI22_X1 port map( A1 => n915, A2 => n1142, B1 => n882, B2 => n1143, 
                           ZN => n1390);
   U447 : NOR4_X1 port map( A1 => n1395, A2 => n1396, A3 => n1397, A4 => n1398,
                           ZN => n1378);
   U448 : OAI22_X1 port map( A1 => n982, A2 => n1148, B1 => n949, B2 => n1149, 
                           ZN => n1398);
   U449 : OAI22_X1 port map( A1 => n1050, A2 => n1151, B1 => n1016, B2 => n1152
                           , ZN => n1397);
   U450 : OAI22_X1 port map( A1 => n89, A2 => n1153, B1 => n1083, B2 => n3, ZN 
                           => n1396);
   U451 : OAI22_X1 port map( A1 => n165, A2 => n1155, B1 => n129, B2 => n1156, 
                           ZN => n1395);
   U452 : OAI22_X1 port map( A1 => n1399, A2 => n1102, B1 => n1103, B2 => n1392
                           , ZN => N4592);
   U453 : NOR4_X1 port map( A1 => n1404, A2 => n1405, A3 => n1406, A4 => n1407,
                           ZN => n1403);
   U454 : OAI22_X1 port map( A1 => n187, A2 => n1112, B1 => n837, B2 => n1113, 
                           ZN => n1407);
   U455 : OAI22_X1 port map( A1 => n251, A2 => n1114, B1 => n219, B2 => n1115, 
                           ZN => n1406);
   U456 : OAI22_X1 port map( A1 => n315, A2 => n1116, B1 => n283, B2 => n1117, 
                           ZN => n1405);
   U457 : OAI22_X1 port map( A1 => n379, A2 => n1118, B1 => n347, B2 => n1119, 
                           ZN => n1404);
   U458 : NOR4_X1 port map( A1 => n1408, A2 => n1409, A3 => n1410, A4 => n1411,
                           ZN => n1402);
   U459 : OAI22_X1 port map( A1 => n444, A2 => n1124, B1 => n411, B2 => n1125, 
                           ZN => n1411);
   U460 : OAI22_X1 port map( A1 => n511, A2 => n1126, B1 => n477, B2 => n1127, 
                           ZN => n1410);
   U461 : OAI22_X1 port map( A1 => n578, A2 => n1128, B1 => n545, B2 => n1129, 
                           ZN => n1409);
   U462 : OAI22_X1 port map( A1 => n645, A2 => n1130, B1 => n612, B2 => n1131, 
                           ZN => n1408);
   U463 : NOR4_X1 port map( A1 => n1412, A2 => n1413, A3 => n1415, A4 => n1416,
                           ZN => n1401);
   U464 : OAI22_X1 port map( A1 => n713, A2 => n1136, B1 => n679, B2 => n1137, 
                           ZN => n1416);
   U465 : OAI22_X1 port map( A1 => n780, A2 => n1138, B1 => n746, B2 => n1139, 
                           ZN => n1415);
   U466 : OAI22_X1 port map( A1 => n847, A2 => n1140, B1 => n813, B2 => n1141, 
                           ZN => n1413);
   U467 : OAI22_X1 port map( A1 => n914, A2 => n1142, B1 => n881, B2 => n1143, 
                           ZN => n1412);
   U468 : NOR4_X1 port map( A1 => n1417, A2 => n1418, A3 => n1419, A4 => n1420,
                           ZN => n1400);
   U469 : OAI22_X1 port map( A1 => n981, A2 => n1148, B1 => n948, B2 => n1149, 
                           ZN => n1420);
   U470 : OAI22_X1 port map( A1 => n1049, A2 => n1151, B1 => n1015, B2 => n1152
                           , ZN => n1419);
   U471 : OAI22_X1 port map( A1 => n87, A2 => n2, B1 => n1082, B2 => n3, ZN => 
                           n1418);
   U472 : OAI22_X1 port map( A1 => n163, A2 => n1155, B1 => n128, B2 => n1156, 
                           ZN => n1417);
   U473 : OAI22_X1 port map( A1 => n1421, A2 => n1102, B1 => n1103, B2 => n1414
                           , ZN => N4590);
   U474 : NOR4_X1 port map( A1 => n1426, A2 => n1427, A3 => n1428, A4 => n1429,
                           ZN => n1425);
   U475 : OAI22_X1 port map( A1 => n186, A2 => n1112, B1 => n816, B2 => n1113, 
                           ZN => n1429);
   U476 : OAI22_X1 port map( A1 => n250, A2 => n1114, B1 => n218, B2 => n1115, 
                           ZN => n1428);
   U477 : OAI22_X1 port map( A1 => n314, A2 => n1116, B1 => n282, B2 => n1117, 
                           ZN => n1427);
   U478 : OAI22_X1 port map( A1 => n378, A2 => n1118, B1 => n346, B2 => n1119, 
                           ZN => n1426);
   U479 : NOR4_X1 port map( A1 => n1430, A2 => n1431, A3 => n1432, A4 => n1433,
                           ZN => n1424);
   U480 : OAI22_X1 port map( A1 => n443, A2 => n1124, B1 => n410, B2 => n1125, 
                           ZN => n1433);
   U481 : OAI22_X1 port map( A1 => n510, A2 => n1126, B1 => n476, B2 => n1127, 
                           ZN => n1432);
   U482 : OAI22_X1 port map( A1 => n577, A2 => n1128, B1 => n544, B2 => n1129, 
                           ZN => n1431);
   U483 : OAI22_X1 port map( A1 => n644, A2 => n1130, B1 => n611, B2 => n1131, 
                           ZN => n1430);
   U484 : NOR4_X1 port map( A1 => n1434, A2 => n1435, A3 => n1437, A4 => n1438,
                           ZN => n1423);
   U485 : OAI22_X1 port map( A1 => n712, A2 => n1136, B1 => n678, B2 => n1137, 
                           ZN => n1438);
   U486 : OAI22_X1 port map( A1 => n779, A2 => n1138, B1 => n745, B2 => n1139, 
                           ZN => n1437);
   U487 : OAI22_X1 port map( A1 => n846, A2 => n1140, B1 => n812, B2 => n1141, 
                           ZN => n1435);
   U488 : OAI22_X1 port map( A1 => n913, A2 => n1142, B1 => n880, B2 => n1143, 
                           ZN => n1434);
   U489 : NOR4_X1 port map( A1 => n1439, A2 => n1440, A3 => n1441, A4 => n1442,
                           ZN => n1422);
   U490 : OAI22_X1 port map( A1 => n980, A2 => n1148, B1 => n947, B2 => n1149, 
                           ZN => n1442);
   U491 : OAI22_X1 port map( A1 => n1048, A2 => n1151, B1 => n1014, B2 => n1152
                           , ZN => n1441);
   U492 : OAI22_X1 port map( A1 => n85, A2 => n2, B1 => n1081, B2 => n3, ZN => 
                           n1440);
   U493 : OAI22_X1 port map( A1 => n162, A2 => n1155, B1 => n127, B2 => n1156, 
                           ZN => n1439);
   U494 : OAI22_X1 port map( A1 => n1443, A2 => n1102, B1 => n1103, B2 => n1436
                           , ZN => N4588);
   U495 : NOR4_X1 port map( A1 => n1448, A2 => n1449, A3 => n1450, A4 => n1451,
                           ZN => n1447);
   U496 : OAI22_X1 port map( A1 => n185, A2 => n1112, B1 => n795, B2 => n1113, 
                           ZN => n1451);
   U497 : OAI22_X1 port map( A1 => n249, A2 => n1114, B1 => n217, B2 => n1115, 
                           ZN => n1450);
   U498 : OAI22_X1 port map( A1 => n313, A2 => n1116, B1 => n281, B2 => n1117, 
                           ZN => n1449);
   U499 : OAI22_X1 port map( A1 => n377, A2 => n1118, B1 => n345, B2 => n1119, 
                           ZN => n1448);
   U500 : NOR4_X1 port map( A1 => n1452, A2 => n1453, A3 => n1454, A4 => n1455,
                           ZN => n1446);
   U501 : OAI22_X1 port map( A1 => n442, A2 => n1124, B1 => n409, B2 => n1125, 
                           ZN => n1455);
   U502 : OAI22_X1 port map( A1 => n509, A2 => n1126, B1 => n475, B2 => n1127, 
                           ZN => n1454);
   U503 : OAI22_X1 port map( A1 => n576, A2 => n1128, B1 => n542, B2 => n1129, 
                           ZN => n1453);
   U504 : OAI22_X1 port map( A1 => n643, A2 => n1130, B1 => n610, B2 => n1131, 
                           ZN => n1452);
   U505 : NOR4_X1 port map( A1 => n1456, A2 => n1457, A3 => n1459, A4 => n1460,
                           ZN => n1445);
   U506 : OAI22_X1 port map( A1 => n710, A2 => n1136, B1 => n677, B2 => n1137, 
                           ZN => n1460);
   U507 : OAI22_X1 port map( A1 => n778, A2 => n1138, B1 => n744, B2 => n1139, 
                           ZN => n1459);
   U508 : OAI22_X1 port map( A1 => n845, A2 => n1140, B1 => n811, B2 => n1141, 
                           ZN => n1457);
   U509 : OAI22_X1 port map( A1 => n912, A2 => n1142, B1 => n878, B2 => n1143, 
                           ZN => n1456);
   U510 : NOR4_X1 port map( A1 => n1461, A2 => n1462, A3 => n1463, A4 => n1464,
                           ZN => n1444);
   U511 : OAI22_X1 port map( A1 => n979, A2 => n1148, B1 => n946, B2 => n1149, 
                           ZN => n1464);
   U512 : OAI22_X1 port map( A1 => n1046, A2 => n1151, B1 => n1013, B2 => n1152
                           , ZN => n1463);
   U513 : OAI22_X1 port map( A1 => n83, A2 => n2, B1 => n1080, B2 => n3, ZN => 
                           n1462);
   U514 : OAI22_X1 port map( A1 => n161, A2 => n1155, B1 => n126, B2 => n1156, 
                           ZN => n1461);
   U515 : OAI22_X1 port map( A1 => n1465, A2 => n1102, B1 => n1103, B2 => n1458
                           , ZN => N4586);
   U516 : NOR4_X1 port map( A1 => n1470, A2 => n1471, A3 => n1472, A4 => n1473,
                           ZN => n1469);
   U517 : OAI22_X1 port map( A1 => n184, A2 => n1112, B1 => n774, B2 => n1113, 
                           ZN => n1473);
   U518 : OAI22_X1 port map( A1 => n248, A2 => n1114, B1 => n216, B2 => n1115, 
                           ZN => n1472);
   U519 : OAI22_X1 port map( A1 => n312, A2 => n1116, B1 => n280, B2 => n1117, 
                           ZN => n1471);
   U520 : OAI22_X1 port map( A1 => n376, A2 => n1118, B1 => n344, B2 => n1119, 
                           ZN => n1470);
   U521 : NOR4_X1 port map( A1 => n1474, A2 => n1475, A3 => n1476, A4 => n1477,
                           ZN => n1468);
   U522 : OAI22_X1 port map( A1 => n441, A2 => n1124, B1 => n408, B2 => n1125, 
                           ZN => n1477);
   U523 : OAI22_X1 port map( A1 => n508, A2 => n1126, B1 => n474, B2 => n1127, 
                           ZN => n1476);
   U524 : OAI22_X1 port map( A1 => n575, A2 => n1128, B1 => n541, B2 => n1129, 
                           ZN => n1475);
   U525 : OAI22_X1 port map( A1 => n642, A2 => n1130, B1 => n609, B2 => n1131, 
                           ZN => n1474);
   U526 : NOR4_X1 port map( A1 => n1478, A2 => n1479, A3 => n1481, A4 => n1482,
                           ZN => n1467);
   U527 : OAI22_X1 port map( A1 => n709, A2 => n1136, B1 => n676, B2 => n1137, 
                           ZN => n1482);
   U528 : OAI22_X1 port map( A1 => n777, A2 => n1138, B1 => n743, B2 => n1139, 
                           ZN => n1481);
   U529 : OAI22_X1 port map( A1 => n844, A2 => n1140, B1 => n810, B2 => n1141, 
                           ZN => n1479);
   U530 : OAI22_X1 port map( A1 => n911, A2 => n1142, B1 => n877, B2 => n1143, 
                           ZN => n1478);
   U531 : NOR4_X1 port map( A1 => n1483, A2 => n1484, A3 => n1485, A4 => n1486,
                           ZN => n1466);
   U532 : OAI22_X1 port map( A1 => n978, A2 => n1148, B1 => n945, B2 => n1149, 
                           ZN => n1486);
   U533 : OAI22_X1 port map( A1 => n1045, A2 => n1151, B1 => n1012, B2 => n1152
                           , ZN => n1485);
   U534 : OAI22_X1 port map( A1 => n81, A2 => n2, B1 => n1079, B2 => n3, ZN => 
                           n1484);
   U535 : OAI22_X1 port map( A1 => n160, A2 => n1155, B1 => n125, B2 => n1156, 
                           ZN => n1483);
   U536 : OAI22_X1 port map( A1 => n1487, A2 => n1102, B1 => n1103, B2 => n1480
                           , ZN => N4584);
   U537 : NOR4_X1 port map( A1 => n1492, A2 => n1493, A3 => n1494, A4 => n1495,
                           ZN => n1491);
   U538 : OAI22_X1 port map( A1 => n183, A2 => n1112, B1 => n753, B2 => n1113, 
                           ZN => n1495);
   U539 : OAI22_X1 port map( A1 => n247, A2 => n1114, B1 => n215, B2 => n1115, 
                           ZN => n1494);
   U540 : OAI22_X1 port map( A1 => n311, A2 => n1116, B1 => n279, B2 => n1117, 
                           ZN => n1493);
   U541 : OAI22_X1 port map( A1 => n375, A2 => n1118, B1 => n343, B2 => n1119, 
                           ZN => n1492);
   U542 : NOR4_X1 port map( A1 => n1496, A2 => n1497, A3 => n1498, A4 => n1499,
                           ZN => n1490);
   U543 : OAI22_X1 port map( A1 => n440, A2 => n1124, B1 => n407, B2 => n1125, 
                           ZN => n1499);
   U544 : OAI22_X1 port map( A1 => n507, A2 => n1126, B1 => n473, B2 => n1127, 
                           ZN => n1498);
   U545 : OAI22_X1 port map( A1 => n574, A2 => n1128, B1 => n540, B2 => n1129, 
                           ZN => n1497);
   U546 : OAI22_X1 port map( A1 => n641, A2 => n1130, B1 => n608, B2 => n1131, 
                           ZN => n1496);
   U547 : NOR4_X1 port map( A1 => n1500, A2 => n1501, A3 => n1503, A4 => n1504,
                           ZN => n1489);
   U548 : OAI22_X1 port map( A1 => n708, A2 => n1136, B1 => n675, B2 => n1137, 
                           ZN => n1504);
   U549 : OAI22_X1 port map( A1 => n776, A2 => n1138, B1 => n742, B2 => n1139, 
                           ZN => n1503);
   U550 : OAI22_X1 port map( A1 => n843, A2 => n1140, B1 => n809, B2 => n1141, 
                           ZN => n1501);
   U551 : OAI22_X1 port map( A1 => n910, A2 => n1142, B1 => n876, B2 => n1143, 
                           ZN => n1500);
   U552 : NOR4_X1 port map( A1 => n1505, A2 => n1506, A3 => n1507, A4 => n1508,
                           ZN => n1488);
   U553 : OAI22_X1 port map( A1 => n977, A2 => n1148, B1 => n944, B2 => n1149, 
                           ZN => n1508);
   U554 : OAI22_X1 port map( A1 => n1044, A2 => n1151, B1 => n1011, B2 => n1152
                           , ZN => n1507);
   U555 : OAI22_X1 port map( A1 => n79, A2 => n2, B1 => n1078, B2 => n3, ZN => 
                           n1506);
   U556 : OAI22_X1 port map( A1 => n159, A2 => n1155, B1 => n124, B2 => n1156, 
                           ZN => n1505);
   U557 : OAI22_X1 port map( A1 => n1509, A2 => n1102, B1 => n1103, B2 => n1502
                           , ZN => N4582);
   U558 : NOR4_X1 port map( A1 => n1514, A2 => n1515, A3 => n1516, A4 => n1517,
                           ZN => n1513);
   U559 : OAI22_X1 port map( A1 => n182, A2 => n1112, B1 => n732, B2 => n1113, 
                           ZN => n1517);
   U560 : OAI22_X1 port map( A1 => n246, A2 => n1114, B1 => n214, B2 => n1115, 
                           ZN => n1516);
   U561 : OAI22_X1 port map( A1 => n310, A2 => n1116, B1 => n278, B2 => n1117, 
                           ZN => n1515);
   U562 : OAI22_X1 port map( A1 => n374, A2 => n1118, B1 => n342, B2 => n1119, 
                           ZN => n1514);
   U563 : NOR4_X1 port map( A1 => n1518, A2 => n1519, A3 => n1520, A4 => n1521,
                           ZN => n1512);
   U564 : OAI22_X1 port map( A1 => n439, A2 => n1124, B1 => n406, B2 => n1125, 
                           ZN => n1521);
   U565 : OAI22_X1 port map( A1 => n506, A2 => n1126, B1 => n472, B2 => n1127, 
                           ZN => n1520);
   U566 : OAI22_X1 port map( A1 => n573, A2 => n1128, B1 => n539, B2 => n1129, 
                           ZN => n1519);
   U567 : OAI22_X1 port map( A1 => n640, A2 => n1130, B1 => n607, B2 => n1131, 
                           ZN => n1518);
   U568 : NOR4_X1 port map( A1 => n1522, A2 => n1523, A3 => n1525, A4 => n1526,
                           ZN => n1511);
   U569 : OAI22_X1 port map( A1 => n707, A2 => n1136, B1 => n674, B2 => n1137, 
                           ZN => n1526);
   U570 : OAI22_X1 port map( A1 => n775, A2 => n1138, B1 => n741, B2 => n1139, 
                           ZN => n1525);
   U571 : OAI22_X1 port map( A1 => n842, A2 => n1140, B1 => n808, B2 => n1141, 
                           ZN => n1523);
   U572 : OAI22_X1 port map( A1 => n909, A2 => n1142, B1 => n875, B2 => n1143, 
                           ZN => n1522);
   U573 : NOR4_X1 port map( A1 => n1527, A2 => n1528, A3 => n1529, A4 => n1530,
                           ZN => n1510);
   U574 : OAI22_X1 port map( A1 => n976, A2 => n1148, B1 => n943, B2 => n1149, 
                           ZN => n1530);
   U575 : OAI22_X1 port map( A1 => n1043, A2 => n1151, B1 => n1010, B2 => n1152
                           , ZN => n1529);
   U576 : OAI22_X1 port map( A1 => n77, A2 => n2, B1 => n1077, B2 => n3, ZN => 
                           n1528);
   U577 : OAI22_X1 port map( A1 => n158, A2 => n1155, B1 => n123, B2 => n1156, 
                           ZN => n1527);
   U578 : OAI22_X1 port map( A1 => n1531, A2 => n1102, B1 => n1103, B2 => n1524
                           , ZN => N4580);
   U579 : NOR4_X1 port map( A1 => n1536, A2 => n1537, A3 => n1538, A4 => n1539,
                           ZN => n1535);
   U580 : OAI22_X1 port map( A1 => n181, A2 => n1112, B1 => n711, B2 => n1113, 
                           ZN => n1539);
   U581 : OAI22_X1 port map( A1 => n245, A2 => n1114, B1 => n213, B2 => n1115, 
                           ZN => n1538);
   U582 : OAI22_X1 port map( A1 => n309, A2 => n1116, B1 => n277, B2 => n1117, 
                           ZN => n1537);
   U583 : OAI22_X1 port map( A1 => n373, A2 => n1118, B1 => n341, B2 => n1119, 
                           ZN => n1536);
   U584 : NOR4_X1 port map( A1 => n1540, A2 => n1541, A3 => n1542, A4 => n1543,
                           ZN => n1534);
   U585 : OAI22_X1 port map( A1 => n437, A2 => n1124, B1 => n405, B2 => n1125, 
                           ZN => n1543);
   U586 : OAI22_X1 port map( A1 => n505, A2 => n1126, B1 => n471, B2 => n1127, 
                           ZN => n1542);
   U587 : OAI22_X1 port map( A1 => n572, A2 => n1128, B1 => n538, B2 => n1129, 
                           ZN => n1541);
   U588 : OAI22_X1 port map( A1 => n639, A2 => n1130, B1 => n605, B2 => n1131, 
                           ZN => n1540);
   U589 : NOR4_X1 port map( A1 => n1544, A2 => n1545, A3 => n1547, A4 => n1548,
                           ZN => n1533);
   U590 : OAI22_X1 port map( A1 => n706, A2 => n1136, B1 => n673, B2 => n1137, 
                           ZN => n1548);
   U591 : OAI22_X1 port map( A1 => n773, A2 => n1138, B1 => n740, B2 => n1139, 
                           ZN => n1547);
   U592 : OAI22_X1 port map( A1 => n841, A2 => n1140, B1 => n807, B2 => n1141, 
                           ZN => n1545);
   U593 : OAI22_X1 port map( A1 => n908, A2 => n1142, B1 => n874, B2 => n1143, 
                           ZN => n1544);
   U594 : NOR4_X1 port map( A1 => n1549, A2 => n1550, A3 => n1551, A4 => n1552,
                           ZN => n1532);
   U595 : OAI22_X1 port map( A1 => n975, A2 => n1148, B1 => n941, B2 => n1149, 
                           ZN => n1552);
   U596 : OAI22_X1 port map( A1 => n1042, A2 => n1151, B1 => n1009, B2 => n1152
                           , ZN => n1551);
   U597 : OAI22_X1 port map( A1 => n73, A2 => n2, B1 => n1076, B2 => n3, ZN => 
                           n1550);
   U598 : OAI22_X1 port map( A1 => n157, A2 => n1155, B1 => n122, B2 => n1156, 
                           ZN => n1549);
   U599 : OAI22_X1 port map( A1 => n1553, A2 => n1102, B1 => n1103, B2 => n1546
                           , ZN => N4578);
   U600 : NOR4_X1 port map( A1 => n1558, A2 => n1559, A3 => n1560, A4 => n1561,
                           ZN => n1557);
   U601 : OAI22_X1 port map( A1 => n180, A2 => n1112, B1 => n690, B2 => n1113, 
                           ZN => n1561);
   U602 : OAI22_X1 port map( A1 => n244, A2 => n1114, B1 => n212, B2 => n1115, 
                           ZN => n1560);
   U603 : OAI22_X1 port map( A1 => n308, A2 => n1116, B1 => n276, B2 => n1117, 
                           ZN => n1559);
   U604 : OAI22_X1 port map( A1 => n372, A2 => n1118, B1 => n340, B2 => n1119, 
                           ZN => n1558);
   U605 : NOR4_X1 port map( A1 => n1562, A2 => n1563, A3 => n1564, A4 => n1565,
                           ZN => n1556);
   U606 : OAI22_X1 port map( A1 => n436, A2 => n1124, B1 => n404, B2 => n1125, 
                           ZN => n1565);
   U607 : OAI22_X1 port map( A1 => n504, A2 => n1126, B1 => n470, B2 => n1127, 
                           ZN => n1564);
   U608 : OAI22_X1 port map( A1 => n571, A2 => n1128, B1 => n537, B2 => n1129, 
                           ZN => n1563);
   U609 : OAI22_X1 port map( A1 => n638, A2 => n1130, B1 => n604, B2 => n1131, 
                           ZN => n1562);
   U610 : NOR4_X1 port map( A1 => n1566, A2 => n1567, A3 => n1569, A4 => n1570,
                           ZN => n1555);
   U611 : OAI22_X1 port map( A1 => n705, A2 => n1136, B1 => n672, B2 => n1137, 
                           ZN => n1570);
   U612 : OAI22_X1 port map( A1 => n772, A2 => n1138, B1 => n739, B2 => n1139, 
                           ZN => n1569);
   U613 : OAI22_X1 port map( A1 => n840, A2 => n1140, B1 => n806, B2 => n1141, 
                           ZN => n1567);
   U614 : OAI22_X1 port map( A1 => n907, A2 => n1142, B1 => n873, B2 => n1143, 
                           ZN => n1566);
   U615 : NOR4_X1 port map( A1 => n1571, A2 => n1572, A3 => n1573, A4 => n1574,
                           ZN => n1554);
   U616 : OAI22_X1 port map( A1 => n974, A2 => n1148, B1 => n940, B2 => n1149, 
                           ZN => n1574);
   U617 : OAI22_X1 port map( A1 => n1041, A2 => n1151, B1 => n1008, B2 => n1152
                           , ZN => n1573);
   U618 : OAI22_X1 port map( A1 => n71, A2 => n2, B1 => n1075, B2 => n3, ZN => 
                           n1572);
   U619 : OAI22_X1 port map( A1 => n156, A2 => n1155, B1 => n121, B2 => n1156, 
                           ZN => n1571);
   U620 : OAI22_X1 port map( A1 => n1575, A2 => n1102, B1 => n1103, B2 => n1568
                           , ZN => N4576);
   U621 : NOR4_X1 port map( A1 => n1580, A2 => n1581, A3 => n1582, A4 => n1583,
                           ZN => n1579);
   U622 : OAI22_X1 port map( A1 => n179, A2 => n1112, B1 => n669, B2 => n1113, 
                           ZN => n1583);
   U623 : OAI22_X1 port map( A1 => n243, A2 => n1114, B1 => n211, B2 => n1115, 
                           ZN => n1582);
   U624 : OAI22_X1 port map( A1 => n307, A2 => n1116, B1 => n275, B2 => n1117, 
                           ZN => n1581);
   U625 : OAI22_X1 port map( A1 => n371, A2 => n1118, B1 => n339, B2 => n1119, 
                           ZN => n1580);
   U626 : NOR4_X1 port map( A1 => n1584, A2 => n1585, A3 => n1586, A4 => n1587,
                           ZN => n1578);
   U627 : OAI22_X1 port map( A1 => n435, A2 => n1124, B1 => n403, B2 => n1125, 
                           ZN => n1587);
   U628 : OAI22_X1 port map( A1 => n503, A2 => n1126, B1 => n469, B2 => n1127, 
                           ZN => n1586);
   U629 : OAI22_X1 port map( A1 => n570, A2 => n1128, B1 => n536, B2 => n1129, 
                           ZN => n1585);
   U630 : OAI22_X1 port map( A1 => n637, A2 => n1130, B1 => n603, B2 => n1131, 
                           ZN => n1584);
   U631 : NOR4_X1 port map( A1 => n1588, A2 => n1589, A3 => n1591, A4 => n1592,
                           ZN => n1577);
   U632 : OAI22_X1 port map( A1 => n704, A2 => n1136, B1 => n671, B2 => n1137, 
                           ZN => n1592);
   U633 : OAI22_X1 port map( A1 => n771, A2 => n1138, B1 => n738, B2 => n1139, 
                           ZN => n1591);
   U634 : OAI22_X1 port map( A1 => n839, A2 => n1140, B1 => n805, B2 => n1141, 
                           ZN => n1589);
   U635 : OAI22_X1 port map( A1 => n906, A2 => n1, B1 => n872, B2 => n1143, ZN 
                           => n1588);
   U636 : NOR4_X1 port map( A1 => n1593, A2 => n1594, A3 => n1595, A4 => n1596,
                           ZN => n1576);
   U637 : OAI22_X1 port map( A1 => n973, A2 => n1148, B1 => n939, B2 => n1149, 
                           ZN => n1596);
   U638 : OAI22_X1 port map( A1 => n1040, A2 => n1151, B1 => n1007, B2 => n1152
                           , ZN => n1595);
   U639 : OAI22_X1 port map( A1 => n69, A2 => n2, B1 => n1074, B2 => n1154, ZN 
                           => n1594);
   U640 : OAI22_X1 port map( A1 => n155, A2 => n1155, B1 => n119, B2 => n1156, 
                           ZN => n1593);
   U641 : OAI22_X1 port map( A1 => n1597, A2 => n1102, B1 => n1103, B2 => n1590
                           , ZN => N4574);
   U642 : NOR4_X1 port map( A1 => n1602, A2 => n1603, A3 => n1604, A4 => n1605,
                           ZN => n1601);
   U643 : OAI22_X1 port map( A1 => n178, A2 => n1112, B1 => n648, B2 => n1113, 
                           ZN => n1605);
   U644 : OAI22_X1 port map( A1 => n242, A2 => n1114, B1 => n210, B2 => n1115, 
                           ZN => n1604);
   U645 : OAI22_X1 port map( A1 => n306, A2 => n1116, B1 => n274, B2 => n1117, 
                           ZN => n1603);
   U646 : OAI22_X1 port map( A1 => n370, A2 => n1118, B1 => n338, B2 => n1119, 
                           ZN => n1602);
   U647 : NOR4_X1 port map( A1 => n1606, A2 => n1607, A3 => n1608, A4 => n1609,
                           ZN => n1600);
   U648 : OAI22_X1 port map( A1 => n434, A2 => n1124, B1 => n402, B2 => n1125, 
                           ZN => n1609);
   U649 : OAI22_X1 port map( A1 => n502, A2 => n1126, B1 => n468, B2 => n1127, 
                           ZN => n1608);
   U650 : OAI22_X1 port map( A1 => n569, A2 => n1128, B1 => n535, B2 => n1129, 
                           ZN => n1607);
   U651 : OAI22_X1 port map( A1 => n636, A2 => n1130, B1 => n602, B2 => n1131, 
                           ZN => n1606);
   U652 : NOR4_X1 port map( A1 => n1610, A2 => n1611, A3 => n1613, A4 => n1614,
                           ZN => n1599);
   U653 : OAI22_X1 port map( A1 => n703, A2 => n1136, B1 => n670, B2 => n1137, 
                           ZN => n1614);
   U654 : OAI22_X1 port map( A1 => n770, A2 => n1138, B1 => n737, B2 => n1139, 
                           ZN => n1613);
   U655 : OAI22_X1 port map( A1 => n838, A2 => n1140, B1 => n804, B2 => n1141, 
                           ZN => n1611);
   U656 : OAI22_X1 port map( A1 => n905, A2 => n1, B1 => n871, B2 => n1143, ZN 
                           => n1610);
   U657 : NOR4_X1 port map( A1 => n1615, A2 => n1616, A3 => n1617, A4 => n1618,
                           ZN => n1598);
   U658 : OAI22_X1 port map( A1 => n972, A2 => n1148, B1 => n938, B2 => n1149, 
                           ZN => n1618);
   U659 : OAI22_X1 port map( A1 => n1039, A2 => n1151, B1 => n1006, B2 => n1152
                           , ZN => n1617);
   U660 : OAI22_X1 port map( A1 => n67, A2 => n2, B1 => n1073, B2 => n1154, ZN 
                           => n1616);
   U661 : OAI22_X1 port map( A1 => n154, A2 => n1155, B1 => n118, B2 => n1156, 
                           ZN => n1615);
   U662 : OAI22_X1 port map( A1 => n1619, A2 => n1102, B1 => n1103, B2 => n1612
                           , ZN => N4572);
   U663 : NOR4_X1 port map( A1 => n1624, A2 => n1625, A3 => n1626, A4 => n1627,
                           ZN => n1623);
   U664 : OAI22_X1 port map( A1 => n175, A2 => n1112, B1 => n627, B2 => n1113, 
                           ZN => n1627);
   U665 : OAI22_X1 port map( A1 => n241, A2 => n1114, B1 => n209, B2 => n1115, 
                           ZN => n1626);
   U666 : OAI22_X1 port map( A1 => n305, A2 => n1116, B1 => n273, B2 => n1117, 
                           ZN => n1625);
   U667 : OAI22_X1 port map( A1 => n369, A2 => n1118, B1 => n337, B2 => n1119, 
                           ZN => n1624);
   U668 : NOR4_X1 port map( A1 => n1628, A2 => n1629, A3 => n1630, A4 => n1631,
                           ZN => n1622);
   U669 : OAI22_X1 port map( A1 => n433, A2 => n1124, B1 => n401, B2 => n1125, 
                           ZN => n1631);
   U670 : OAI22_X1 port map( A1 => n500, A2 => n1126, B1 => n467, B2 => n1127, 
                           ZN => n1630);
   U671 : OAI22_X1 port map( A1 => n568, A2 => n1128, B1 => n534, B2 => n1129, 
                           ZN => n1629);
   U672 : OAI22_X1 port map( A1 => n635, A2 => n1130, B1 => n601, B2 => n1131, 
                           ZN => n1628);
   U673 : NOR4_X1 port map( A1 => n1632, A2 => n1633, A3 => n1635, A4 => n1636,
                           ZN => n1621);
   U674 : OAI22_X1 port map( A1 => n702, A2 => n1136, B1 => n668, B2 => n1137, 
                           ZN => n1636);
   U675 : OAI22_X1 port map( A1 => n769, A2 => n1138, B1 => n736, B2 => n1139, 
                           ZN => n1635);
   U676 : OAI22_X1 port map( A1 => n836, A2 => n1140, B1 => n803, B2 => n1141, 
                           ZN => n1633);
   U677 : OAI22_X1 port map( A1 => n904, A2 => n1, B1 => n870, B2 => n1143, ZN 
                           => n1632);
   U678 : NOR4_X1 port map( A1 => n1637, A2 => n1638, A3 => n1639, A4 => n1640,
                           ZN => n1620);
   U679 : OAI22_X1 port map( A1 => n971, A2 => n1148, B1 => n937, B2 => n1149, 
                           ZN => n1640);
   U680 : OAI22_X1 port map( A1 => n1038, A2 => n1151, B1 => n1004, B2 => n1152
                           , ZN => n1639);
   U681 : OAI22_X1 port map( A1 => n65, A2 => n2, B1 => n1072, B2 => n1154, ZN 
                           => n1638);
   U682 : OAI22_X1 port map( A1 => n152, A2 => n1155, B1 => n117, B2 => n1156, 
                           ZN => n1637);
   U683 : OAI22_X1 port map( A1 => n1641, A2 => n1102, B1 => n1103, B2 => n1634
                           , ZN => N4570);
   U684 : NOR4_X1 port map( A1 => n1646, A2 => n1647, A3 => n1648, A4 => n1649,
                           ZN => n1645);
   U685 : OAI22_X1 port map( A1 => n164, A2 => n1112, B1 => n606, B2 => n1113, 
                           ZN => n1649);
   U686 : OAI22_X1 port map( A1 => n240, A2 => n1114, B1 => n208, B2 => n1115, 
                           ZN => n1648);
   U687 : OAI22_X1 port map( A1 => n304, A2 => n1116, B1 => n272, B2 => n1117, 
                           ZN => n1647);
   U688 : OAI22_X1 port map( A1 => n368, A2 => n1118, B1 => n336, B2 => n1119, 
                           ZN => n1646);
   U689 : NOR4_X1 port map( A1 => n1650, A2 => n1651, A3 => n1652, A4 => n1653,
                           ZN => n1644);
   U690 : OAI22_X1 port map( A1 => n432, A2 => n1124, B1 => n400, B2 => n1125, 
                           ZN => n1653);
   U691 : OAI22_X1 port map( A1 => n499, A2 => n1126, B1 => n466, B2 => n1127, 
                           ZN => n1652);
   U692 : OAI22_X1 port map( A1 => n567, A2 => n1128, B1 => n533, B2 => n1129, 
                           ZN => n1651);
   U693 : OAI22_X1 port map( A1 => n634, A2 => n1130, B1 => n600, B2 => n1131, 
                           ZN => n1650);
   U694 : NOR4_X1 port map( A1 => n1654, A2 => n1655, A3 => n1657, A4 => n1658,
                           ZN => n1643);
   U695 : OAI22_X1 port map( A1 => n701, A2 => n1136, B1 => n667, B2 => n1137, 
                           ZN => n1658);
   U696 : OAI22_X1 port map( A1 => n768, A2 => n1138, B1 => n735, B2 => n1139, 
                           ZN => n1657);
   U697 : OAI22_X1 port map( A1 => n835, A2 => n1140, B1 => n802, B2 => n1141, 
                           ZN => n1655);
   U698 : OAI22_X1 port map( A1 => n903, A2 => n1, B1 => n869, B2 => n1143, ZN 
                           => n1654);
   U699 : NOR4_X1 port map( A1 => n1659, A2 => n1660, A3 => n1661, A4 => n1662,
                           ZN => n1642);
   U700 : OAI22_X1 port map( A1 => n970, A2 => n1148, B1 => n936, B2 => n1149, 
                           ZN => n1662);
   U701 : OAI22_X1 port map( A1 => n1037, A2 => n1151, B1 => n1003, B2 => n1152
                           , ZN => n1661);
   U702 : OAI22_X1 port map( A1 => n63, A2 => n2, B1 => n1071, B2 => n1154, ZN 
                           => n1660);
   U703 : OAI22_X1 port map( A1 => n151, A2 => n1155, B1 => n116, B2 => n37, ZN
                           => n1659);
   U704 : OAI22_X1 port map( A1 => n1663, A2 => n1102, B1 => n1103, B2 => n1656
                           , ZN => N4568);
   U705 : NOR4_X1 port map( A1 => n1668, A2 => n1669, A3 => n1670, A4 => n1671,
                           ZN => n1667);
   U706 : OAI22_X1 port map( A1 => n153, A2 => n1112, B1 => n585, B2 => n1113, 
                           ZN => n1671);
   U707 : OAI22_X1 port map( A1 => n239, A2 => n1114, B1 => n207, B2 => n1115, 
                           ZN => n1670);
   U708 : OAI22_X1 port map( A1 => n303, A2 => n1116, B1 => n271, B2 => n1117, 
                           ZN => n1669);
   U709 : OAI22_X1 port map( A1 => n367, A2 => n1118, B1 => n335, B2 => n1119, 
                           ZN => n1668);
   U710 : NOR4_X1 port map( A1 => n1672, A2 => n1673, A3 => n1674, A4 => n1675,
                           ZN => n1666);
   U711 : OAI22_X1 port map( A1 => n431, A2 => n1124, B1 => n399, B2 => n1125, 
                           ZN => n1675);
   U712 : OAI22_X1 port map( A1 => n498, A2 => n1126, B1 => n465, B2 => n1127, 
                           ZN => n1674);
   U713 : OAI22_X1 port map( A1 => n566, A2 => n1128, B1 => n532, B2 => n1129, 
                           ZN => n1673);
   U714 : OAI22_X1 port map( A1 => n633, A2 => n1130, B1 => n599, B2 => n1131, 
                           ZN => n1672);
   U715 : NOR4_X1 port map( A1 => n1676, A2 => n1677, A3 => n1679, A4 => n1680,
                           ZN => n1665);
   U716 : OAI22_X1 port map( A1 => n700, A2 => n1136, B1 => n666, B2 => n1137, 
                           ZN => n1680);
   U717 : OAI22_X1 port map( A1 => n767, A2 => n1138, B1 => n734, B2 => n1139, 
                           ZN => n1679);
   U718 : OAI22_X1 port map( A1 => n834, A2 => n1140, B1 => n801, B2 => n1141, 
                           ZN => n1677);
   U719 : OAI22_X1 port map( A1 => n902, A2 => n1, B1 => n868, B2 => n1143, ZN 
                           => n1676);
   U720 : NOR4_X1 port map( A1 => n1681, A2 => n1682, A3 => n1683, A4 => n1684,
                           ZN => n1664);
   U721 : OAI22_X1 port map( A1 => n969, A2 => n1148, B1 => n935, B2 => n1149, 
                           ZN => n1684);
   U722 : OAI22_X1 port map( A1 => n1036, A2 => n1151, B1 => n1002, B2 => n1152
                           , ZN => n1683);
   U723 : OAI22_X1 port map( A1 => n61, A2 => n2, B1 => n1070, B2 => n1154, ZN 
                           => n1682);
   U724 : OAI22_X1 port map( A1 => n150, A2 => n1155, B1 => n115, B2 => n1156, 
                           ZN => n1681);
   U725 : OAI22_X1 port map( A1 => n1685, A2 => n1102, B1 => n1103, B2 => n1678
                           , ZN => N4566);
   U726 : NOR4_X1 port map( A1 => n1690, A2 => n1691, A3 => n1692, A4 => n1693,
                           ZN => n1689);
   U727 : OAI22_X1 port map( A1 => n142, A2 => n1112, B1 => n564, B2 => n1113, 
                           ZN => n1693);
   U728 : OAI22_X1 port map( A1 => n238, A2 => n1114, B1 => n206, B2 => n1115, 
                           ZN => n1692);
   U729 : OAI22_X1 port map( A1 => n302, A2 => n1116, B1 => n270, B2 => n1117, 
                           ZN => n1691);
   U730 : OAI22_X1 port map( A1 => n366, A2 => n1118, B1 => n334, B2 => n1119, 
                           ZN => n1690);
   U731 : NOR4_X1 port map( A1 => n1694, A2 => n1695, A3 => n1696, A4 => n1697,
                           ZN => n1688);
   U732 : OAI22_X1 port map( A1 => n430, A2 => n1124, B1 => n398, B2 => n1125, 
                           ZN => n1697);
   U733 : OAI22_X1 port map( A1 => n497, A2 => n1126, B1 => n464, B2 => n1127, 
                           ZN => n1696);
   U734 : OAI22_X1 port map( A1 => n565, A2 => n1128, B1 => n531, B2 => n1129, 
                           ZN => n1695);
   U735 : OAI22_X1 port map( A1 => n632, A2 => n1130, B1 => n598, B2 => n1131, 
                           ZN => n1694);
   U736 : NOR4_X1 port map( A1 => n1698, A2 => n1699, A3 => n1701, A4 => n1702,
                           ZN => n1687);
   U737 : OAI22_X1 port map( A1 => n699, A2 => n1136, B1 => n665, B2 => n1137, 
                           ZN => n1702);
   U738 : OAI22_X1 port map( A1 => n766, A2 => n1138, B1 => n733, B2 => n1139, 
                           ZN => n1701);
   U739 : OAI22_X1 port map( A1 => n833, A2 => n1140, B1 => n800, B2 => n1141, 
                           ZN => n1699);
   U740 : OAI22_X1 port map( A1 => n901, A2 => n1, B1 => n867, B2 => n1143, ZN 
                           => n1698);
   U741 : NOR4_X1 port map( A1 => n1703, A2 => n1704, A3 => n1705, A4 => n1706,
                           ZN => n1686);
   U742 : OAI22_X1 port map( A1 => n968, A2 => n1148, B1 => n934, B2 => n1149, 
                           ZN => n1706);
   U743 : OAI22_X1 port map( A1 => n1035, A2 => n1151, B1 => n1001, B2 => n1152
                           , ZN => n1705);
   U744 : OAI22_X1 port map( A1 => n59, A2 => n1153, B1 => n1069, B2 => n1154, 
                           ZN => n1704);
   U745 : OAI22_X1 port map( A1 => n149, A2 => n1155, B1 => n114, B2 => n37, ZN
                           => n1703);
   U746 : OAI22_X1 port map( A1 => n1707, A2 => n1102, B1 => n1103, B2 => n1700
                           , ZN => N4564);
   U747 : NOR4_X1 port map( A1 => n1712, A2 => n1713, A3 => n1714, A4 => n1715,
                           ZN => n1711);
   U748 : OAI22_X1 port map( A1 => n131, A2 => n1112, B1 => n543, B2 => n1113, 
                           ZN => n1715);
   U749 : OAI22_X1 port map( A1 => n237, A2 => n1114, B1 => n205, B2 => n1115, 
                           ZN => n1714);
   U750 : OAI22_X1 port map( A1 => n301, A2 => n1116, B1 => n269, B2 => n1117, 
                           ZN => n1713);
   U751 : OAI22_X1 port map( A1 => n365, A2 => n1118, B1 => n333, B2 => n1119, 
                           ZN => n1712);
   U752 : NOR4_X1 port map( A1 => n1716, A2 => n1717, A3 => n1718, A4 => n1719,
                           ZN => n1710);
   U753 : OAI22_X1 port map( A1 => n429, A2 => n1124, B1 => n397, B2 => n1125, 
                           ZN => n1719);
   U754 : OAI22_X1 port map( A1 => n496, A2 => n1126, B1 => n463, B2 => n1127, 
                           ZN => n1718);
   U755 : OAI22_X1 port map( A1 => n563, A2 => n1128, B1 => n530, B2 => n1129, 
                           ZN => n1717);
   U756 : OAI22_X1 port map( A1 => n631, A2 => n1130, B1 => n597, B2 => n1131, 
                           ZN => n1716);
   U757 : NOR4_X1 port map( A1 => n1720, A2 => n1721, A3 => n1723, A4 => n1724,
                           ZN => n1709);
   U758 : OAI22_X1 port map( A1 => n698, A2 => n1136, B1 => n664, B2 => n1137, 
                           ZN => n1724);
   U759 : OAI22_X1 port map( A1 => n765, A2 => n1138, B1 => n731, B2 => n1139, 
                           ZN => n1723);
   U760 : OAI22_X1 port map( A1 => n832, A2 => n1140, B1 => n799, B2 => n1141, 
                           ZN => n1721);
   U761 : OAI22_X1 port map( A1 => n899, A2 => n1, B1 => n866, B2 => n1143, ZN 
                           => n1720);
   U762 : NOR4_X1 port map( A1 => n1725, A2 => n1726, A3 => n1727, A4 => n1728,
                           ZN => n1708);
   U763 : OAI22_X1 port map( A1 => n967, A2 => n1148, B1 => n933, B2 => n1149, 
                           ZN => n1728);
   U764 : OAI22_X1 port map( A1 => n1034, A2 => n1151, B1 => n1000, B2 => n1152
                           , ZN => n1727);
   U765 : OAI22_X1 port map( A1 => n57, A2 => n1153, B1 => n1067, B2 => n1154, 
                           ZN => n1726);
   U766 : OAI22_X1 port map( A1 => n148, A2 => n1155, B1 => n113, B2 => n1156, 
                           ZN => n1725);
   U767 : OAI22_X1 port map( A1 => n1729, A2 => n1102, B1 => n1103, B2 => n1722
                           , ZN => N4562);
   U768 : NOR4_X1 port map( A1 => n1734, A2 => n1735, A3 => n1736, A4 => n1737,
                           ZN => n1733);
   U769 : OAI22_X1 port map( A1 => n120, A2 => n1112, B1 => n522, B2 => n1113, 
                           ZN => n1737);
   U770 : OAI22_X1 port map( A1 => n236, A2 => n1114, B1 => n204, B2 => n1115, 
                           ZN => n1736);
   U771 : OAI22_X1 port map( A1 => n300, A2 => n1116, B1 => n268, B2 => n1117, 
                           ZN => n1735);
   U772 : OAI22_X1 port map( A1 => n364, A2 => n1118, B1 => n332, B2 => n1119, 
                           ZN => n1734);
   U773 : NOR4_X1 port map( A1 => n1738, A2 => n1739, A3 => n1740, A4 => n1741,
                           ZN => n1732);
   U774 : OAI22_X1 port map( A1 => n428, A2 => n1124, B1 => n396, B2 => n1125, 
                           ZN => n1741);
   U775 : OAI22_X1 port map( A1 => n495, A2 => n1126, B1 => n462, B2 => n1127, 
                           ZN => n1740);
   U776 : OAI22_X1 port map( A1 => n562, A2 => n1128, B1 => n529, B2 => n1129, 
                           ZN => n1739);
   U777 : OAI22_X1 port map( A1 => n630, A2 => n1130, B1 => n596, B2 => n1131, 
                           ZN => n1738);
   U778 : NOR4_X1 port map( A1 => n1742, A2 => n1743, A3 => n1745, A4 => n1746,
                           ZN => n1731);
   U779 : OAI22_X1 port map( A1 => n697, A2 => n1136, B1 => n663, B2 => n1137, 
                           ZN => n1746);
   U780 : OAI22_X1 port map( A1 => n764, A2 => n1138, B1 => n730, B2 => n1139, 
                           ZN => n1745);
   U781 : OAI22_X1 port map( A1 => n831, A2 => n1140, B1 => n798, B2 => n1141, 
                           ZN => n1743);
   U782 : OAI22_X1 port map( A1 => n898, A2 => n1, B1 => n865, B2 => n1143, ZN 
                           => n1742);
   U783 : NOR4_X1 port map( A1 => n1747, A2 => n1748, A3 => n1749, A4 => n1750,
                           ZN => n1730);
   U784 : OAI22_X1 port map( A1 => n966, A2 => n1148, B1 => n932, B2 => n1149, 
                           ZN => n1750);
   U785 : OAI22_X1 port map( A1 => n1033, A2 => n1151, B1 => n999, B2 => n1152,
                           ZN => n1749);
   U786 : OAI22_X1 port map( A1 => n55, A2 => n1153, B1 => n1066, B2 => n1154, 
                           ZN => n1748);
   U787 : OAI22_X1 port map( A1 => n147, A2 => n1155, B1 => n112, B2 => n1156, 
                           ZN => n1747);
   U788 : OAI22_X1 port map( A1 => n1751, A2 => n1102, B1 => n1744, B2 => n1103
                           , ZN => N4560);
   U789 : NOR4_X1 port map( A1 => n1752, A2 => n1753, A3 => n1754, A4 => n1755,
                           ZN => n1751);
   U790 : OAI211_X1 port map( C1 => n1100, C2 => n1153, A => n1756, B => n1757,
                           ZN => n1755);
   U791 : NOR4_X1 port map( A1 => n1758, A2 => n1759, A3 => n1760, A4 => n1761,
                           ZN => n1757);
   U792 : OAI22_X1 port map( A1 => n109, A2 => n1112, B1 => n203, B2 => n1115, 
                           ZN => n1761);
   U793 : OAI22_X1 port map( A1 => n235, A2 => n1114, B1 => n267, B2 => n1117, 
                           ZN => n1760);
   U794 : OAI22_X1 port map( A1 => n299, A2 => n1116, B1 => n331, B2 => n1119, 
                           ZN => n1759);
   U795 : OAI22_X1 port map( A1 => n363, A2 => n1118, B1 => n395, B2 => n1125, 
                           ZN => n1758);
   U796 : NOR4_X1 port map( A1 => n1762, A2 => n1763, A3 => n1764, A4 => n1765,
                           ZN => n1756);
   U797 : OAI22_X1 port map( A1 => n427, A2 => n1124, B1 => n461, B2 => n1127, 
                           ZN => n1765);
   U798 : OAI22_X1 port map( A1 => n494, A2 => n1126, B1 => n528, B2 => n1129, 
                           ZN => n1764);
   U799 : OAI22_X1 port map( A1 => n561, A2 => n1128, B1 => n595, B2 => n1131, 
                           ZN => n1763);
   U800 : OAI22_X1 port map( A1 => n629, A2 => n1130, B1 => n662, B2 => n1137, 
                           ZN => n1762);
   U801 : OAI211_X1 port map( C1 => n146, C2 => n1155, A => n1767, B => n1768, 
                           ZN => n1754);
   U802 : NOR4_X1 port map( A1 => n1769, A2 => n1770, A3 => n1771, A4 => n1772,
                           ZN => n1768);
   U803 : OAI22_X1 port map( A1 => n763, A2 => n1138, B1 => n797, B2 => n1141, 
                           ZN => n1772);
   U804 : OAI22_X1 port map( A1 => n696, A2 => n1136, B1 => n729, B2 => n1139, 
                           ZN => n1771);
   U805 : OAI22_X1 port map( A1 => n897, A2 => n1, B1 => n931, B2 => n1149, ZN 
                           => n1770);
   U806 : OAI22_X1 port map( A1 => n830, A2 => n1140, B1 => n864, B2 => n1143, 
                           ZN => n1769);
   U807 : OAI22_X1 port map( A1 => n1113, A2 => n501, B1 => n37, B2 => n111, ZN
                           => n1773);
   U808 : OAI22_X1 port map( A1 => n1032, A2 => n1151, B1 => n1065, B2 => n1154
                           , ZN => n1753);
   U809 : OAI22_X1 port map( A1 => n965, A2 => n1148, B1 => n998, B2 => n1152, 
                           ZN => n1752);
   U810 : OAI22_X1 port map( A1 => n1774, A2 => n1102, B1 => n1103, B2 => n1766
                           , ZN => N4558);
   U811 : NOR4_X1 port map( A1 => n1779, A2 => n1780, A3 => n1781, A4 => n1782,
                           ZN => n1778);
   U812 : OAI22_X1 port map( A1 => n97, A2 => n1112, B1 => n480, B2 => n1113, 
                           ZN => n1782);
   U813 : OAI22_X1 port map( A1 => n234, A2 => n1114, B1 => n202, B2 => n1115, 
                           ZN => n1781);
   U814 : OAI22_X1 port map( A1 => n298, A2 => n1116, B1 => n266, B2 => n1117, 
                           ZN => n1780);
   U815 : OAI22_X1 port map( A1 => n362, A2 => n1118, B1 => n330, B2 => n1119, 
                           ZN => n1779);
   U816 : NOR4_X1 port map( A1 => n1783, A2 => n1784, A3 => n1785, A4 => n1786,
                           ZN => n1777);
   U817 : OAI22_X1 port map( A1 => n426, A2 => n1124, B1 => n394, B2 => n1125, 
                           ZN => n1786);
   U818 : OAI22_X1 port map( A1 => n493, A2 => n1126, B1 => n460, B2 => n1127, 
                           ZN => n1785);
   U819 : OAI22_X1 port map( A1 => n560, A2 => n1128, B1 => n527, B2 => n1129, 
                           ZN => n1784);
   U820 : OAI22_X1 port map( A1 => n628, A2 => n1130, B1 => n594, B2 => n1131, 
                           ZN => n1783);
   U821 : NOR4_X1 port map( A1 => n1787, A2 => n1789, A3 => n1790, A4 => n1791,
                           ZN => n1776);
   U822 : OAI22_X1 port map( A1 => n695, A2 => n1136, B1 => n661, B2 => n1137, 
                           ZN => n1791);
   U823 : OAI22_X1 port map( A1 => n762, A2 => n1138, B1 => n728, B2 => n1139, 
                           ZN => n1790);
   U824 : OAI22_X1 port map( A1 => n829, A2 => n1140, B1 => n796, B2 => n1141, 
                           ZN => n1789);
   U825 : OAI22_X1 port map( A1 => n896, A2 => n1, B1 => n863, B2 => n1143, ZN 
                           => n1787);
   U826 : NOR4_X1 port map( A1 => n1792, A2 => n1793, A3 => n1794, A4 => n1795,
                           ZN => n1775);
   U827 : OAI22_X1 port map( A1 => n964, A2 => n1148, B1 => n930, B2 => n1149, 
                           ZN => n1795);
   U828 : OAI22_X1 port map( A1 => n1031, A2 => n1151, B1 => n997, B2 => n1152,
                           ZN => n1794);
   U829 : OAI22_X1 port map( A1 => n1099, A2 => n1153, B1 => n1064, B2 => n1154
                           , ZN => n1793);
   U830 : OAI22_X1 port map( A1 => n145, A2 => n1155, B1 => n110, B2 => n1156, 
                           ZN => n1792);
   U831 : OAI22_X1 port map( A1 => n1796, A2 => n1102, B1 => n1103, B2 => n1788
                           , ZN => N4556);
   U832 : NOR4_X1 port map( A1 => n1801, A2 => n1802, A3 => n1803, A4 => n1804,
                           ZN => n1800);
   U833 : OAI22_X1 port map( A1 => n75, A2 => n1112, B1 => n459, B2 => n1113, 
                           ZN => n1804);
   U834 : OAI22_X1 port map( A1 => n233, A2 => n1114, B1 => n201, B2 => n1115, 
                           ZN => n1803);
   U835 : OAI22_X1 port map( A1 => n297, A2 => n1116, B1 => n265, B2 => n1117, 
                           ZN => n1802);
   U836 : OAI22_X1 port map( A1 => n361, A2 => n1118, B1 => n329, B2 => n1119, 
                           ZN => n1801);
   U837 : NOR4_X1 port map( A1 => n1805, A2 => n1806, A3 => n1807, A4 => n1808,
                           ZN => n1799);
   U838 : OAI22_X1 port map( A1 => n425, A2 => n1124, B1 => n393, B2 => n1125, 
                           ZN => n1808);
   U839 : OAI22_X1 port map( A1 => n492, A2 => n1126, B1 => n458, B2 => n1127, 
                           ZN => n1807);
   U840 : OAI22_X1 port map( A1 => n559, A2 => n1128, B1 => n526, B2 => n1129, 
                           ZN => n1806);
   U841 : OAI22_X1 port map( A1 => n626, A2 => n1130, B1 => n593, B2 => n1131, 
                           ZN => n1805);
   U842 : NOR4_X1 port map( A1 => n1809, A2 => n1811, A3 => n1812, A4 => n1813,
                           ZN => n1798);
   U843 : OAI22_X1 port map( A1 => n694, A2 => n1136, B1 => n660, B2 => n1137, 
                           ZN => n1813);
   U844 : OAI22_X1 port map( A1 => n761, A2 => n1138, B1 => n727, B2 => n1139, 
                           ZN => n1812);
   U845 : OAI22_X1 port map( A1 => n828, A2 => n1140, B1 => n794, B2 => n1141, 
                           ZN => n1811);
   U846 : OAI22_X1 port map( A1 => n895, A2 => n1, B1 => n862, B2 => n1143, ZN 
                           => n1809);
   U847 : NOR4_X1 port map( A1 => n1814, A2 => n1815, A3 => n1816, A4 => n1817,
                           ZN => n1797);
   U848 : OAI22_X1 port map( A1 => n962, A2 => n1148, B1 => n929, B2 => n1149, 
                           ZN => n1817);
   U849 : OAI22_X1 port map( A1 => n1030, A2 => n1151, B1 => n996, B2 => n1152,
                           ZN => n1816);
   U850 : OAI22_X1 port map( A1 => n1098, A2 => n1153, B1 => n1063, B2 => n1154
                           , ZN => n1815);
   U851 : OAI22_X1 port map( A1 => n144, A2 => n1155, B1 => n108, B2 => n1156, 
                           ZN => n1814);
   U852 : OAI22_X1 port map( A1 => n1818, A2 => n1102, B1 => n1103, B2 => n1810
                           , ZN => N4554);
   U853 : OAI221_X1 port map( B1 => n1825, B2 => ADD_RD2(2), C1 => n1826, C2 =>
                           ADD_RD2(0), A => n1827, ZN => n1824);
   U854 : AOI22_X1 port map( A1 => n1825, A2 => ADD_RD2(2), B1 => n1826, B2 => 
                           ADD_RD2(0), ZN => n1827);
   U855 : AOI221_X1 port map( B1 => n1828, B2 => ADD_WR(4), C1 => n1829, C2 => 
                           ADD_RD2(3), A => n1830, ZN => n1820);
   U856 : OAI22_X1 port map( A1 => ADD_WR(4), A2 => n1828, B1 => n1829, B2 => 
                           ADD_RD2(3), ZN => n1830);
   U857 : NOR4_X1 port map( A1 => n1835, A2 => n1836, A3 => n1837, A4 => n1838,
                           ZN => n1834);
   U858 : OAI22_X1 port map( A1 => n53, A2 => n1112, B1 => n438, B2 => n1113, 
                           ZN => n1838);
   U859 : OAI22_X1 port map( A1 => n232, A2 => n1114, B1 => n200, B2 => n1115, 
                           ZN => n1837);
   U860 : OAI22_X1 port map( A1 => n296, A2 => n1116, B1 => n264, B2 => n1117, 
                           ZN => n1836);
   U861 : OAI22_X1 port map( A1 => n360, A2 => n1118, B1 => n328, B2 => n1119, 
                           ZN => n1835);
   U862 : NOR3_X1 port map( A1 => n1828, A2 => n1845, A3 => n1846, ZN => n1840)
                           ;
   U863 : NAND2_X1 port map( A1 => ADD_RD2(4), A2 => ADD_RD2(3), ZN => n1847);
   U864 : NOR4_X1 port map( A1 => n1848, A2 => n1849, A3 => n1850, A4 => n1851,
                           ZN => n1833);
   U865 : OAI22_X1 port map( A1 => n424, A2 => n1124, B1 => n392, B2 => n1125, 
                           ZN => n1851);
   U866 : OAI22_X1 port map( A1 => n491, A2 => n1126, B1 => n457, B2 => n1127, 
                           ZN => n1850);
   U867 : OAI22_X1 port map( A1 => n558, A2 => n1128, B1 => n525, B2 => n1129, 
                           ZN => n1849);
   U868 : OAI22_X1 port map( A1 => n625, A2 => n1130, B1 => n592, B2 => n1131, 
                           ZN => n1848);
   U869 : NOR3_X1 port map( A1 => ADD_RD2(3), A2 => n1828, A3 => n1846, ZN => 
                           n1852);
   U870 : NOR3_X1 port map( A1 => ADD_RD2(3), A2 => ADD_RD2(0), A3 => n1828, ZN
                           => n1853);
   U871 : NOR4_X1 port map( A1 => n1854, A2 => n1855, A3 => n1856, A4 => n1857,
                           ZN => n1832);
   U872 : OAI22_X1 port map( A1 => n693, A2 => n1136, B1 => n659, B2 => n1137, 
                           ZN => n1857);
   U873 : OAI22_X1 port map( A1 => n760, A2 => n1138, B1 => n726, B2 => n1139, 
                           ZN => n1856);
   U874 : OAI22_X1 port map( A1 => n827, A2 => n1140, B1 => n793, B2 => n1141, 
                           ZN => n1855);
   U875 : OAI22_X1 port map( A1 => n894, A2 => n1, B1 => n861, B2 => n1143, ZN 
                           => n1854);
   U876 : NOR3_X1 port map( A1 => ADD_RD2(4), A2 => n1845, A3 => n1846, ZN => 
                           n1858);
   U877 : NAND2_X1 port map( A1 => n1844, A2 => n1859, ZN => n1142);
   U878 : NOR3_X1 port map( A1 => ADD_RD2(4), A2 => ADD_RD2(0), A3 => n1845, ZN
                           => n1859);
   U879 : NOR4_X1 port map( A1 => n1860, A2 => n1861, A3 => n1862, A4 => n1863,
                           ZN => n1831);
   U880 : OAI22_X1 port map( A1 => n961, A2 => n1148, B1 => n928, B2 => n1149, 
                           ZN => n1863);
   U881 : OAI22_X1 port map( A1 => n1029, A2 => n1151, B1 => n995, B2 => n1152,
                           ZN => n1862);
   U882 : OAI22_X1 port map( A1 => n1097, A2 => n1153, B1 => n1062, B2 => n1154
                           , ZN => n1861);
   U883 : NAND2_X1 port map( A1 => n1843, A2 => n1864, ZN => n1154);
   U884 : NAND2_X1 port map( A1 => n1865, A2 => n1843, ZN => n1153);
   U885 : OAI22_X1 port map( A1 => n143, A2 => n1155, B1 => n107, B2 => n37, ZN
                           => n1860);
   U886 : NAND2_X1 port map( A1 => n1844, A2 => n1864, ZN => n1156);
   U887 : NOR3_X1 port map( A1 => ADD_RD2(4), A2 => ADD_RD2(3), A3 => n1846, ZN
                           => n1864);
   U888 : NOR3_X1 port map( A1 => ADD_RD2(4), A2 => ADD_RD2(3), A3 => 
                           ADD_RD2(0), ZN => n1865);
   U889 : OAI22_X1 port map( A1 => n1866, A2 => n1867, B1 => n1868, B2 => n1094
                           , ZN => N4552);
   U890 : NOR4_X1 port map( A1 => n1873, A2 => n1874, A3 => n1875, A4 => n1876,
                           ZN => n1872);
   U891 : OAI22_X1 port map( A1 => n199, A2 => n1877, B1 => n1089, B2 => n1878,
                           ZN => n1876);
   U892 : OAI22_X1 port map( A1 => n263, A2 => n1879, B1 => n231, B2 => n1880, 
                           ZN => n1875);
   U893 : OAI22_X1 port map( A1 => n327, A2 => n1881, B1 => n295, B2 => n1882, 
                           ZN => n1874);
   U894 : OAI22_X1 port map( A1 => n391, A2 => n1883, B1 => n359, B2 => n1884, 
                           ZN => n1873);
   U895 : NOR4_X1 port map( A1 => n1885, A2 => n1886, A3 => n1887, A4 => n1888,
                           ZN => n1871);
   U896 : OAI22_X1 port map( A1 => n456, A2 => n1889, B1 => n423, B2 => n1890, 
                           ZN => n1888);
   U897 : OAI22_X1 port map( A1 => n524, A2 => n1891, B1 => n490, B2 => n1892, 
                           ZN => n1887);
   U898 : OAI22_X1 port map( A1 => n591, A2 => n1893, B1 => n557, B2 => n1894, 
                           ZN => n1886);
   U899 : OAI22_X1 port map( A1 => n658, A2 => n1895, B1 => n624, B2 => n1896, 
                           ZN => n1885);
   U900 : NOR4_X1 port map( A1 => n1897, A2 => n1898, A3 => n1899, A4 => n1900,
                           ZN => n1870);
   U901 : OAI22_X1 port map( A1 => n725, A2 => n1901, B1 => n692, B2 => n1902, 
                           ZN => n1900);
   U902 : OAI22_X1 port map( A1 => n792, A2 => n1903, B1 => n759, B2 => n1904, 
                           ZN => n1899);
   U903 : OAI22_X1 port map( A1 => n860, A2 => n1905, B1 => n826, B2 => n1906, 
                           ZN => n1898);
   U904 : OAI22_X1 port map( A1 => n927, A2 => n1907, B1 => n893, B2 => n1908, 
                           ZN => n1897);
   U905 : NOR4_X1 port map( A1 => n1909, A2 => n1910, A3 => n1911, A4 => n1912,
                           ZN => n1869);
   U906 : OAI22_X1 port map( A1 => n994, A2 => n1913, B1 => n960, B2 => n1914, 
                           ZN => n1912);
   U907 : OAI22_X1 port map( A1 => n1061, A2 => n1915, B1 => n1028, B2 => n1916
                           , ZN => n1911);
   U908 : OAI22_X1 port map( A1 => n106, A2 => n41, B1 => n1096, B2 => n1918, 
                           ZN => n1910);
   U909 : OAI22_X1 port map( A1 => n177, A2 => n1919, B1 => n141, B2 => n1920, 
                           ZN => n1909);
   U910 : OAI22_X1 port map( A1 => n1921, A2 => n1867, B1 => n1868, B2 => n1150
                           , ZN => N4550);
   U911 : NOR4_X1 port map( A1 => n1926, A2 => n1927, A3 => n1928, A4 => n1929,
                           ZN => n1925);
   U912 : OAI22_X1 port map( A1 => n198, A2 => n1877, B1 => n1068, B2 => n1878,
                           ZN => n1929);
   U913 : OAI22_X1 port map( A1 => n262, A2 => n1879, B1 => n230, B2 => n1880, 
                           ZN => n1928);
   U914 : OAI22_X1 port map( A1 => n326, A2 => n1881, B1 => n294, B2 => n1882, 
                           ZN => n1927);
   U915 : OAI22_X1 port map( A1 => n390, A2 => n1883, B1 => n358, B2 => n1884, 
                           ZN => n1926);
   U916 : NOR4_X1 port map( A1 => n1930, A2 => n1931, A3 => n1932, A4 => n1933,
                           ZN => n1924);
   U917 : OAI22_X1 port map( A1 => n455, A2 => n1889, B1 => n422, B2 => n1890, 
                           ZN => n1933);
   U918 : OAI22_X1 port map( A1 => n523, A2 => n1891, B1 => n489, B2 => n1892, 
                           ZN => n1932);
   U919 : OAI22_X1 port map( A1 => n590, A2 => n1893, B1 => n556, B2 => n1894, 
                           ZN => n1931);
   U920 : OAI22_X1 port map( A1 => n657, A2 => n1895, B1 => n623, B2 => n1896, 
                           ZN => n1930);
   U921 : NOR4_X1 port map( A1 => n1934, A2 => n1935, A3 => n1936, A4 => n1937,
                           ZN => n1923);
   U922 : OAI22_X1 port map( A1 => n724, A2 => n1901, B1 => n691, B2 => n1902, 
                           ZN => n1937);
   U923 : OAI22_X1 port map( A1 => n791, A2 => n1903, B1 => n758, B2 => n1904, 
                           ZN => n1936);
   U924 : OAI22_X1 port map( A1 => n859, A2 => n1905, B1 => n825, B2 => n1906, 
                           ZN => n1935);
   U925 : OAI22_X1 port map( A1 => n926, A2 => n39, B1 => n892, B2 => n1908, ZN
                           => n1934);
   U926 : NOR4_X1 port map( A1 => n1938, A2 => n1939, A3 => n1940, A4 => n1941,
                           ZN => n1922);
   U927 : OAI22_X1 port map( A1 => n993, A2 => n1913, B1 => n959, B2 => n1914, 
                           ZN => n1941);
   U928 : OAI22_X1 port map( A1 => n1060, A2 => n1915, B1 => n1027, B2 => n1916
                           , ZN => n1940);
   U929 : OAI22_X1 port map( A1 => n105, A2 => n1917, B1 => n1095, B2 => n1918,
                           ZN => n1939);
   U930 : OAI22_X1 port map( A1 => n176, A2 => n1919, B1 => n140, B2 => n45, ZN
                           => n1938);
   U931 : OAI22_X1 port map( A1 => n1942, A2 => n1867, B1 => n1868, B2 => n1172
                           , ZN => N4548);
   U932 : NOR4_X1 port map( A1 => n1947, A2 => n1948, A3 => n1949, A4 => n1950,
                           ZN => n1946);
   U933 : OAI22_X1 port map( A1 => n197, A2 => n1877, B1 => n1047, B2 => n1878,
                           ZN => n1950);
   U934 : OAI22_X1 port map( A1 => n261, A2 => n1879, B1 => n229, B2 => n1880, 
                           ZN => n1949);
   U935 : OAI22_X1 port map( A1 => n325, A2 => n1881, B1 => n293, B2 => n1882, 
                           ZN => n1948);
   U936 : OAI22_X1 port map( A1 => n389, A2 => n1883, B1 => n357, B2 => n1884, 
                           ZN => n1947);
   U937 : NOR4_X1 port map( A1 => n1951, A2 => n1952, A3 => n1953, A4 => n1954,
                           ZN => n1945);
   U938 : OAI22_X1 port map( A1 => n454, A2 => n1889, B1 => n421, B2 => n1890, 
                           ZN => n1954);
   U939 : OAI22_X1 port map( A1 => n521, A2 => n1891, B1 => n488, B2 => n1892, 
                           ZN => n1953);
   U940 : OAI22_X1 port map( A1 => n589, A2 => n1893, B1 => n555, B2 => n1894, 
                           ZN => n1952);
   U941 : OAI22_X1 port map( A1 => n656, A2 => n1895, B1 => n622, B2 => n1896, 
                           ZN => n1951);
   U942 : NOR4_X1 port map( A1 => n1955, A2 => n1956, A3 => n1957, A4 => n1958,
                           ZN => n1944);
   U943 : OAI22_X1 port map( A1 => n723, A2 => n1901, B1 => n689, B2 => n1902, 
                           ZN => n1958);
   U944 : OAI22_X1 port map( A1 => n790, A2 => n1903, B1 => n757, B2 => n1904, 
                           ZN => n1957);
   U945 : OAI22_X1 port map( A1 => n857, A2 => n1905, B1 => n824, B2 => n1906, 
                           ZN => n1956);
   U946 : OAI22_X1 port map( A1 => n925, A2 => n1907, B1 => n891, B2 => n1908, 
                           ZN => n1955);
   U947 : NOR4_X1 port map( A1 => n1959, A2 => n1960, A3 => n1961, A4 => n1962,
                           ZN => n1943);
   U948 : OAI22_X1 port map( A1 => n992, A2 => n1913, B1 => n958, B2 => n1914, 
                           ZN => n1962);
   U949 : OAI22_X1 port map( A1 => n1059, A2 => n1915, B1 => n1025, B2 => n1916
                           , ZN => n1961);
   U950 : OAI22_X1 port map( A1 => n104, A2 => n1917, B1 => n1093, B2 => n1918,
                           ZN => n1960);
   U951 : OAI22_X1 port map( A1 => n174, A2 => n1919, B1 => n139, B2 => n45, ZN
                           => n1959);
   U952 : OAI22_X1 port map( A1 => n1963, A2 => n1867, B1 => n1868, B2 => n1194
                           , ZN => N4546);
   U953 : NOR4_X1 port map( A1 => n1968, A2 => n1969, A3 => n1970, A4 => n1971,
                           ZN => n1967);
   U954 : OAI22_X1 port map( A1 => n196, A2 => n1877, B1 => n1026, B2 => n1878,
                           ZN => n1971);
   U955 : OAI22_X1 port map( A1 => n260, A2 => n1879, B1 => n228, B2 => n1880, 
                           ZN => n1970);
   U956 : OAI22_X1 port map( A1 => n324, A2 => n1881, B1 => n292, B2 => n1882, 
                           ZN => n1969);
   U957 : OAI22_X1 port map( A1 => n388, A2 => n1883, B1 => n356, B2 => n1884, 
                           ZN => n1968);
   U958 : NOR4_X1 port map( A1 => n1972, A2 => n1973, A3 => n1974, A4 => n1975,
                           ZN => n1966);
   U959 : OAI22_X1 port map( A1 => n453, A2 => n1889, B1 => n420, B2 => n1890, 
                           ZN => n1975);
   U960 : OAI22_X1 port map( A1 => n520, A2 => n1891, B1 => n487, B2 => n1892, 
                           ZN => n1974);
   U961 : OAI22_X1 port map( A1 => n588, A2 => n1893, B1 => n554, B2 => n1894, 
                           ZN => n1973);
   U962 : OAI22_X1 port map( A1 => n655, A2 => n1895, B1 => n621, B2 => n1896, 
                           ZN => n1972);
   U963 : NOR4_X1 port map( A1 => n1976, A2 => n1977, A3 => n1978, A4 => n1979,
                           ZN => n1965);
   U964 : OAI22_X1 port map( A1 => n722, A2 => n1901, B1 => n688, B2 => n1902, 
                           ZN => n1979);
   U965 : OAI22_X1 port map( A1 => n789, A2 => n1903, B1 => n756, B2 => n1904, 
                           ZN => n1978);
   U966 : OAI22_X1 port map( A1 => n856, A2 => n1905, B1 => n823, B2 => n1906, 
                           ZN => n1977);
   U967 : OAI22_X1 port map( A1 => n924, A2 => n1907, B1 => n890, B2 => n1908, 
                           ZN => n1976);
   U968 : NOR4_X1 port map( A1 => n1980, A2 => n1981, A3 => n1982, A4 => n1983,
                           ZN => n1964);
   U969 : OAI22_X1 port map( A1 => n991, A2 => n1913, B1 => n957, B2 => n1914, 
                           ZN => n1983);
   U970 : OAI22_X1 port map( A1 => n1058, A2 => n1915, B1 => n1024, B2 => n1916
                           , ZN => n1982);
   U971 : OAI22_X1 port map( A1 => n103, A2 => n1917, B1 => n1092, B2 => n43, 
                           ZN => n1981);
   U972 : OAI22_X1 port map( A1 => n173, A2 => n1919, B1 => n138, B2 => n45, ZN
                           => n1980);
   U973 : OAI22_X1 port map( A1 => n1984, A2 => n1867, B1 => n1868, B2 => n1216
                           , ZN => N4544);
   U974 : NOR4_X1 port map( A1 => n1989, A2 => n1990, A3 => n1991, A4 => n1992,
                           ZN => n1988);
   U975 : OAI22_X1 port map( A1 => n195, A2 => n1877, B1 => n1005, B2 => n1878,
                           ZN => n1992);
   U976 : OAI22_X1 port map( A1 => n259, A2 => n1879, B1 => n227, B2 => n1880, 
                           ZN => n1991);
   U977 : OAI22_X1 port map( A1 => n323, A2 => n1881, B1 => n291, B2 => n1882, 
                           ZN => n1990);
   U978 : OAI22_X1 port map( A1 => n387, A2 => n1883, B1 => n355, B2 => n1884, 
                           ZN => n1989);
   U979 : NOR4_X1 port map( A1 => n1993, A2 => n1994, A3 => n1995, A4 => n1996,
                           ZN => n1987);
   U980 : OAI22_X1 port map( A1 => n452, A2 => n1889, B1 => n419, B2 => n1890, 
                           ZN => n1996);
   U981 : OAI22_X1 port map( A1 => n519, A2 => n1891, B1 => n486, B2 => n1892, 
                           ZN => n1995);
   U982 : OAI22_X1 port map( A1 => n587, A2 => n1893, B1 => n553, B2 => n1894, 
                           ZN => n1994);
   U983 : OAI22_X1 port map( A1 => n654, A2 => n1895, B1 => n620, B2 => n1896, 
                           ZN => n1993);
   U984 : NOR4_X1 port map( A1 => n1997, A2 => n1998, A3 => n1999, A4 => n2000,
                           ZN => n1986);
   U985 : OAI22_X1 port map( A1 => n721, A2 => n1901, B1 => n687, B2 => n1902, 
                           ZN => n2000);
   U986 : OAI22_X1 port map( A1 => n788, A2 => n1903, B1 => n755, B2 => n1904, 
                           ZN => n1999);
   U987 : OAI22_X1 port map( A1 => n855, A2 => n1905, B1 => n822, B2 => n1906, 
                           ZN => n1998);
   U988 : OAI22_X1 port map( A1 => n923, A2 => n1907, B1 => n889, B2 => n1908, 
                           ZN => n1997);
   U989 : NOR4_X1 port map( A1 => n2001, A2 => n2002, A3 => n2003, A4 => n2004,
                           ZN => n1985);
   U990 : OAI22_X1 port map( A1 => n990, A2 => n1913, B1 => n956, B2 => n1914, 
                           ZN => n2004);
   U991 : OAI22_X1 port map( A1 => n1057, A2 => n1915, B1 => n1023, B2 => n1916
                           , ZN => n2003);
   U992 : OAI22_X1 port map( A1 => n102, A2 => n1917, B1 => n1091, B2 => n43, 
                           ZN => n2002);
   U993 : OAI22_X1 port map( A1 => n172, A2 => n1919, B1 => n137, B2 => n45, ZN
                           => n2001);
   U994 : OAI22_X1 port map( A1 => n2005, A2 => n1867, B1 => n1868, B2 => n1238
                           , ZN => N4542);
   U995 : NOR4_X1 port map( A1 => n2010, A2 => n2011, A3 => n2012, A4 => n2013,
                           ZN => n2009);
   U996 : OAI22_X1 port map( A1 => n194, A2 => n1877, B1 => n984, B2 => n1878, 
                           ZN => n2013);
   U997 : OAI22_X1 port map( A1 => n258, A2 => n1879, B1 => n226, B2 => n1880, 
                           ZN => n2012);
   U998 : OAI22_X1 port map( A1 => n322, A2 => n1881, B1 => n290, B2 => n1882, 
                           ZN => n2011);
   U999 : OAI22_X1 port map( A1 => n386, A2 => n1883, B1 => n354, B2 => n1884, 
                           ZN => n2010);
   U1000 : NOR4_X1 port map( A1 => n2014, A2 => n2015, A3 => n2016, A4 => n2017
                           , ZN => n2008);
   U1001 : OAI22_X1 port map( A1 => n451, A2 => n1889, B1 => n418, B2 => n1890,
                           ZN => n2017);
   U1002 : OAI22_X1 port map( A1 => n518, A2 => n1891, B1 => n485, B2 => n1892,
                           ZN => n2016);
   U1003 : OAI22_X1 port map( A1 => n586, A2 => n1893, B1 => n552, B2 => n1894,
                           ZN => n2015);
   U1004 : OAI22_X1 port map( A1 => n653, A2 => n1895, B1 => n619, B2 => n1896,
                           ZN => n2014);
   U1005 : NOR4_X1 port map( A1 => n2018, A2 => n2019, A3 => n2020, A4 => n2021
                           , ZN => n2007);
   U1006 : OAI22_X1 port map( A1 => n720, A2 => n1901, B1 => n686, B2 => n1902,
                           ZN => n2021);
   U1007 : OAI22_X1 port map( A1 => n787, A2 => n1903, B1 => n754, B2 => n1904,
                           ZN => n2020);
   U1008 : OAI22_X1 port map( A1 => n854, A2 => n1905, B1 => n821, B2 => n1906,
                           ZN => n2019);
   U1009 : OAI22_X1 port map( A1 => n922, A2 => n1907, B1 => n888, B2 => n1908,
                           ZN => n2018);
   U1010 : NOR4_X1 port map( A1 => n2022, A2 => n2023, A3 => n2024, A4 => n2025
                           , ZN => n2006);
   U1011 : OAI22_X1 port map( A1 => n989, A2 => n1913, B1 => n955, B2 => n1914,
                           ZN => n2025);
   U1012 : OAI22_X1 port map( A1 => n1056, A2 => n1915, B1 => n1022, B2 => 
                           n1916, ZN => n2024);
   U1013 : OAI22_X1 port map( A1 => n101, A2 => n1917, B1 => n1090, B2 => n1918
                           , ZN => n2023);
   U1014 : OAI22_X1 port map( A1 => n171, A2 => n1919, B1 => n136, B2 => n45, 
                           ZN => n2022);
   U1015 : OAI22_X1 port map( A1 => n2026, A2 => n1867, B1 => n1868, B2 => 
                           n1260, ZN => N4540);
   U1016 : NOR4_X1 port map( A1 => n2031, A2 => n2032, A3 => n2033, A4 => n2034
                           , ZN => n2030);
   U1017 : OAI22_X1 port map( A1 => n193, A2 => n1877, B1 => n963, B2 => n1878,
                           ZN => n2034);
   U1018 : OAI22_X1 port map( A1 => n257, A2 => n1879, B1 => n225, B2 => n1880,
                           ZN => n2033);
   U1019 : OAI22_X1 port map( A1 => n321, A2 => n1881, B1 => n289, B2 => n1882,
                           ZN => n2032);
   U1020 : OAI22_X1 port map( A1 => n385, A2 => n1883, B1 => n353, B2 => n1884,
                           ZN => n2031);
   U1021 : NOR4_X1 port map( A1 => n2035, A2 => n2036, A3 => n2037, A4 => n2038
                           , ZN => n2029);
   U1022 : OAI22_X1 port map( A1 => n450, A2 => n1889, B1 => n417, B2 => n1890,
                           ZN => n2038);
   U1023 : OAI22_X1 port map( A1 => n517, A2 => n1891, B1 => n484, B2 => n1892,
                           ZN => n2037);
   U1024 : OAI22_X1 port map( A1 => n584, A2 => n1893, B1 => n551, B2 => n1894,
                           ZN => n2036);
   U1025 : OAI22_X1 port map( A1 => n652, A2 => n1895, B1 => n618, B2 => n1896,
                           ZN => n2035);
   U1026 : NOR4_X1 port map( A1 => n2039, A2 => n2040, A3 => n2041, A4 => n2042
                           , ZN => n2028);
   U1027 : OAI22_X1 port map( A1 => n719, A2 => n1901, B1 => n685, B2 => n1902,
                           ZN => n2042);
   U1028 : OAI22_X1 port map( A1 => n786, A2 => n1903, B1 => n752, B2 => n1904,
                           ZN => n2041);
   U1029 : OAI22_X1 port map( A1 => n853, A2 => n1905, B1 => n820, B2 => n1906,
                           ZN => n2040);
   U1030 : OAI22_X1 port map( A1 => n920, A2 => n1907, B1 => n887, B2 => n1908,
                           ZN => n2039);
   U1031 : NOR4_X1 port map( A1 => n2043, A2 => n2044, A3 => n2045, A4 => n2046
                           , ZN => n2027);
   U1032 : OAI22_X1 port map( A1 => n988, A2 => n1913, B1 => n954, B2 => n1914,
                           ZN => n2046);
   U1033 : OAI22_X1 port map( A1 => n1055, A2 => n1915, B1 => n1021, B2 => 
                           n1916, ZN => n2045);
   U1034 : OAI22_X1 port map( A1 => n100, A2 => n1917, B1 => n1088, B2 => n43, 
                           ZN => n2044);
   U1035 : OAI22_X1 port map( A1 => n170, A2 => n1919, B1 => n135, B2 => n45, 
                           ZN => n2043);
   U1036 : OAI22_X1 port map( A1 => n2047, A2 => n1867, B1 => n1868, B2 => 
                           n1282, ZN => N4538);
   U1037 : NOR4_X1 port map( A1 => n2052, A2 => n2053, A3 => n2054, A4 => n2055
                           , ZN => n2051);
   U1038 : OAI22_X1 port map( A1 => n192, A2 => n1877, B1 => n942, B2 => n1878,
                           ZN => n2055);
   U1039 : OAI22_X1 port map( A1 => n256, A2 => n1879, B1 => n224, B2 => n1880,
                           ZN => n2054);
   U1040 : OAI22_X1 port map( A1 => n320, A2 => n1881, B1 => n288, B2 => n1882,
                           ZN => n2053);
   U1041 : OAI22_X1 port map( A1 => n384, A2 => n1883, B1 => n352, B2 => n1884,
                           ZN => n2052);
   U1042 : NOR4_X1 port map( A1 => n2056, A2 => n2057, A3 => n2058, A4 => n2059
                           , ZN => n2050);
   U1043 : OAI22_X1 port map( A1 => n449, A2 => n1889, B1 => n416, B2 => n1890,
                           ZN => n2059);
   U1044 : OAI22_X1 port map( A1 => n516, A2 => n1891, B1 => n483, B2 => n1892,
                           ZN => n2058);
   U1045 : OAI22_X1 port map( A1 => n583, A2 => n1893, B1 => n550, B2 => n1894,
                           ZN => n2057);
   U1046 : OAI22_X1 port map( A1 => n651, A2 => n1895, B1 => n617, B2 => n1896,
                           ZN => n2056);
   U1047 : NOR4_X1 port map( A1 => n2060, A2 => n2061, A3 => n2062, A4 => n2063
                           , ZN => n2049);
   U1048 : OAI22_X1 port map( A1 => n718, A2 => n1901, B1 => n684, B2 => n1902,
                           ZN => n2063);
   U1049 : OAI22_X1 port map( A1 => n785, A2 => n1903, B1 => n751, B2 => n1904,
                           ZN => n2062);
   U1050 : OAI22_X1 port map( A1 => n852, A2 => n1905, B1 => n819, B2 => n1906,
                           ZN => n2061);
   U1051 : OAI22_X1 port map( A1 => n919, A2 => n1907, B1 => n886, B2 => n1908,
                           ZN => n2060);
   U1052 : NOR4_X1 port map( A1 => n2064, A2 => n2065, A3 => n2066, A4 => n2067
                           , ZN => n2048);
   U1053 : OAI22_X1 port map( A1 => n987, A2 => n1913, B1 => n953, B2 => n1914,
                           ZN => n2067);
   U1054 : OAI22_X1 port map( A1 => n1054, A2 => n1915, B1 => n1020, B2 => 
                           n1916, ZN => n2066);
   U1055 : OAI22_X1 port map( A1 => n99, A2 => n1917, B1 => n1087, B2 => n1918,
                           ZN => n2065);
   U1056 : OAI22_X1 port map( A1 => n169, A2 => n1919, B1 => n134, B2 => n45, 
                           ZN => n2064);
   U1057 : OAI22_X1 port map( A1 => n2068, A2 => n1867, B1 => n1868, B2 => 
                           n1304, ZN => N4536);
   U1058 : NOR4_X1 port map( A1 => n2073, A2 => n2074, A3 => n2075, A4 => n2076
                           , ZN => n2072);
   U1059 : OAI22_X1 port map( A1 => n191, A2 => n1877, B1 => n921, B2 => n1878,
                           ZN => n2076);
   U1060 : OAI22_X1 port map( A1 => n255, A2 => n1879, B1 => n223, B2 => n1880,
                           ZN => n2075);
   U1061 : OAI22_X1 port map( A1 => n319, A2 => n1881, B1 => n287, B2 => n1882,
                           ZN => n2074);
   U1062 : OAI22_X1 port map( A1 => n383, A2 => n1883, B1 => n351, B2 => n1884,
                           ZN => n2073);
   U1063 : NOR4_X1 port map( A1 => n2077, A2 => n2078, A3 => n2079, A4 => n2080
                           , ZN => n2071);
   U1064 : OAI22_X1 port map( A1 => n448, A2 => n1889, B1 => n415, B2 => n1890,
                           ZN => n2080);
   U1065 : OAI22_X1 port map( A1 => n515, A2 => n1891, B1 => n482, B2 => n1892,
                           ZN => n2079);
   U1066 : OAI22_X1 port map( A1 => n582, A2 => n1893, B1 => n549, B2 => n1894,
                           ZN => n2078);
   U1067 : OAI22_X1 port map( A1 => n650, A2 => n1895, B1 => n616, B2 => n1896,
                           ZN => n2077);
   U1068 : NOR4_X1 port map( A1 => n2081, A2 => n2082, A3 => n2083, A4 => n2084
                           , ZN => n2070);
   U1069 : OAI22_X1 port map( A1 => n717, A2 => n1901, B1 => n683, B2 => n1902,
                           ZN => n2084);
   U1070 : OAI22_X1 port map( A1 => n784, A2 => n1903, B1 => n750, B2 => n1904,
                           ZN => n2083);
   U1071 : OAI22_X1 port map( A1 => n851, A2 => n1905, B1 => n818, B2 => n1906,
                           ZN => n2082);
   U1072 : OAI22_X1 port map( A1 => n918, A2 => n1907, B1 => n885, B2 => n1908,
                           ZN => n2081);
   U1073 : NOR4_X1 port map( A1 => n2085, A2 => n2086, A3 => n2087, A4 => n2088
                           , ZN => n2069);
   U1074 : OAI22_X1 port map( A1 => n986, A2 => n1913, B1 => n952, B2 => n1914,
                           ZN => n2088);
   U1075 : OAI22_X1 port map( A1 => n1053, A2 => n1915, B1 => n1019, B2 => 
                           n1916, ZN => n2087);
   U1076 : OAI22_X1 port map( A1 => n95, A2 => n1917, B1 => n1086, B2 => n43, 
                           ZN => n2086);
   U1077 : OAI22_X1 port map( A1 => n168, A2 => n1919, B1 => n133, B2 => n45, 
                           ZN => n2085);
   U1078 : OAI22_X1 port map( A1 => n2089, A2 => n1867, B1 => n1868, B2 => 
                           n1326, ZN => N4534);
   U1079 : NOR4_X1 port map( A1 => n2094, A2 => n2095, A3 => n2096, A4 => n2097
                           , ZN => n2093);
   U1080 : OAI22_X1 port map( A1 => n190, A2 => n1877, B1 => n900, B2 => n1878,
                           ZN => n2097);
   U1081 : OAI22_X1 port map( A1 => n254, A2 => n1879, B1 => n222, B2 => n1880,
                           ZN => n2096);
   U1082 : OAI22_X1 port map( A1 => n318, A2 => n1881, B1 => n286, B2 => n1882,
                           ZN => n2095);
   U1083 : OAI22_X1 port map( A1 => n382, A2 => n1883, B1 => n350, B2 => n1884,
                           ZN => n2094);
   U1084 : NOR4_X1 port map( A1 => n2098, A2 => n2099, A3 => n2100, A4 => n2101
                           , ZN => n2092);
   U1085 : OAI22_X1 port map( A1 => n447, A2 => n1889, B1 => n414, B2 => n1890,
                           ZN => n2101);
   U1086 : OAI22_X1 port map( A1 => n514, A2 => n1891, B1 => n481, B2 => n1892,
                           ZN => n2100);
   U1087 : OAI22_X1 port map( A1 => n581, A2 => n1893, B1 => n548, B2 => n1894,
                           ZN => n2099);
   U1088 : OAI22_X1 port map( A1 => n649, A2 => n1895, B1 => n615, B2 => n1896,
                           ZN => n2098);
   U1089 : NOR4_X1 port map( A1 => n2102, A2 => n2103, A3 => n2104, A4 => n2105
                           , ZN => n2091);
   U1090 : OAI22_X1 port map( A1 => n716, A2 => n1901, B1 => n682, B2 => n1902,
                           ZN => n2105);
   U1091 : OAI22_X1 port map( A1 => n783, A2 => n1903, B1 => n749, B2 => n1904,
                           ZN => n2104);
   U1092 : OAI22_X1 port map( A1 => n850, A2 => n1905, B1 => n817, B2 => n1906,
                           ZN => n2103);
   U1093 : OAI22_X1 port map( A1 => n917, A2 => n1907, B1 => n884, B2 => n1908,
                           ZN => n2102);
   U1094 : NOR4_X1 port map( A1 => n2106, A2 => n2107, A3 => n2108, A4 => n2109
                           , ZN => n2090);
   U1095 : OAI22_X1 port map( A1 => n985, A2 => n1913, B1 => n951, B2 => n1914,
                           ZN => n2109);
   U1096 : OAI22_X1 port map( A1 => n1052, A2 => n1915, B1 => n1018, B2 => 
                           n1916, ZN => n2108);
   U1097 : OAI22_X1 port map( A1 => n93, A2 => n1917, B1 => n1085, B2 => n43, 
                           ZN => n2107);
   U1098 : OAI22_X1 port map( A1 => n167, A2 => n1919, B1 => n132, B2 => n45, 
                           ZN => n2106);
   U1099 : OAI22_X1 port map( A1 => n2110, A2 => n1867, B1 => n1868, B2 => 
                           n1348, ZN => N4532);
   U1100 : NOR4_X1 port map( A1 => n2115, A2 => n2116, A3 => n2117, A4 => n2118
                           , ZN => n2114);
   U1101 : OAI22_X1 port map( A1 => n189, A2 => n1877, B1 => n879, B2 => n1878,
                           ZN => n2118);
   U1102 : OAI22_X1 port map( A1 => n253, A2 => n1879, B1 => n221, B2 => n1880,
                           ZN => n2117);
   U1103 : OAI22_X1 port map( A1 => n317, A2 => n1881, B1 => n285, B2 => n1882,
                           ZN => n2116);
   U1104 : OAI22_X1 port map( A1 => n381, A2 => n1883, B1 => n349, B2 => n1884,
                           ZN => n2115);
   U1105 : NOR4_X1 port map( A1 => n2119, A2 => n2120, A3 => n2121, A4 => n2122
                           , ZN => n2113);
   U1106 : OAI22_X1 port map( A1 => n446, A2 => n1889, B1 => n413, B2 => n1890,
                           ZN => n2122);
   U1107 : OAI22_X1 port map( A1 => n513, A2 => n1891, B1 => n479, B2 => n1892,
                           ZN => n2121);
   U1108 : OAI22_X1 port map( A1 => n580, A2 => n1893, B1 => n547, B2 => n1894,
                           ZN => n2120);
   U1109 : OAI22_X1 port map( A1 => n647, A2 => n1895, B1 => n614, B2 => n1896,
                           ZN => n2119);
   U1110 : NOR4_X1 port map( A1 => n2123, A2 => n2124, A3 => n2125, A4 => n2126
                           , ZN => n2112);
   U1111 : OAI22_X1 port map( A1 => n715, A2 => n1901, B1 => n681, B2 => n1902,
                           ZN => n2126);
   U1112 : OAI22_X1 port map( A1 => n782, A2 => n1903, B1 => n748, B2 => n1904,
                           ZN => n2125);
   U1113 : OAI22_X1 port map( A1 => n849, A2 => n1905, B1 => n815, B2 => n1906,
                           ZN => n2124);
   U1114 : OAI22_X1 port map( A1 => n916, A2 => n1907, B1 => n883, B2 => n1908,
                           ZN => n2123);
   U1115 : NOR4_X1 port map( A1 => n2127, A2 => n2128, A3 => n2129, A4 => n2130
                           , ZN => n2111);
   U1116 : OAI22_X1 port map( A1 => n983, A2 => n1913, B1 => n950, B2 => n1914,
                           ZN => n2130);
   U1117 : OAI22_X1 port map( A1 => n1051, A2 => n1915, B1 => n1017, B2 => 
                           n1916, ZN => n2129);
   U1118 : OAI22_X1 port map( A1 => n91, A2 => n1917, B1 => n1084, B2 => n43, 
                           ZN => n2128);
   U1119 : OAI22_X1 port map( A1 => n166, A2 => n1919, B1 => n130, B2 => n45, 
                           ZN => n2127);
   U1120 : OAI22_X1 port map( A1 => n2131, A2 => n1867, B1 => n1868, B2 => 
                           n1370, ZN => N4530);
   U1121 : NOR4_X1 port map( A1 => n2136, A2 => n2137, A3 => n2138, A4 => n2139
                           , ZN => n2135);
   U1122 : OAI22_X1 port map( A1 => n188, A2 => n1877, B1 => n858, B2 => n1878,
                           ZN => n2139);
   U1123 : OAI22_X1 port map( A1 => n252, A2 => n1879, B1 => n220, B2 => n1880,
                           ZN => n2138);
   U1124 : OAI22_X1 port map( A1 => n316, A2 => n1881, B1 => n284, B2 => n1882,
                           ZN => n2137);
   U1125 : OAI22_X1 port map( A1 => n380, A2 => n1883, B1 => n348, B2 => n1884,
                           ZN => n2136);
   U1126 : NOR4_X1 port map( A1 => n2140, A2 => n2141, A3 => n2142, A4 => n2143
                           , ZN => n2134);
   U1127 : OAI22_X1 port map( A1 => n445, A2 => n1889, B1 => n412, B2 => n1890,
                           ZN => n2143);
   U1128 : OAI22_X1 port map( A1 => n512, A2 => n1891, B1 => n478, B2 => n1892,
                           ZN => n2142);
   U1129 : OAI22_X1 port map( A1 => n579, A2 => n1893, B1 => n546, B2 => n1894,
                           ZN => n2141);
   U1130 : OAI22_X1 port map( A1 => n646, A2 => n1895, B1 => n613, B2 => n1896,
                           ZN => n2140);
   U1131 : NOR4_X1 port map( A1 => n2144, A2 => n2145, A3 => n2146, A4 => n2147
                           , ZN => n2133);
   U1132 : OAI22_X1 port map( A1 => n714, A2 => n1901, B1 => n680, B2 => n1902,
                           ZN => n2147);
   U1133 : OAI22_X1 port map( A1 => n781, A2 => n1903, B1 => n747, B2 => n1904,
                           ZN => n2146);
   U1134 : OAI22_X1 port map( A1 => n848, A2 => n1905, B1 => n814, B2 => n1906,
                           ZN => n2145);
   U1135 : OAI22_X1 port map( A1 => n915, A2 => n1907, B1 => n882, B2 => n1908,
                           ZN => n2144);
   U1136 : NOR4_X1 port map( A1 => n2148, A2 => n2149, A3 => n2150, A4 => n2151
                           , ZN => n2132);
   U1137 : OAI22_X1 port map( A1 => n982, A2 => n1913, B1 => n949, B2 => n1914,
                           ZN => n2151);
   U1138 : OAI22_X1 port map( A1 => n1050, A2 => n1915, B1 => n1016, B2 => 
                           n1916, ZN => n2150);
   U1139 : OAI22_X1 port map( A1 => n89, A2 => n1917, B1 => n1083, B2 => n43, 
                           ZN => n2149);
   U1140 : OAI22_X1 port map( A1 => n165, A2 => n1919, B1 => n129, B2 => n1920,
                           ZN => n2148);
   U1141 : OAI22_X1 port map( A1 => n2152, A2 => n1867, B1 => n1868, B2 => 
                           n1392, ZN => N4528);
   U1142 : NOR4_X1 port map( A1 => n2157, A2 => n2158, A3 => n2159, A4 => n2160
                           , ZN => n2156);
   U1143 : OAI22_X1 port map( A1 => n187, A2 => n1877, B1 => n837, B2 => n1878,
                           ZN => n2160);
   U1144 : OAI22_X1 port map( A1 => n251, A2 => n1879, B1 => n219, B2 => n1880,
                           ZN => n2159);
   U1145 : OAI22_X1 port map( A1 => n315, A2 => n1881, B1 => n283, B2 => n1882,
                           ZN => n2158);
   U1146 : OAI22_X1 port map( A1 => n379, A2 => n1883, B1 => n347, B2 => n1884,
                           ZN => n2157);
   U1147 : NOR4_X1 port map( A1 => n2161, A2 => n2162, A3 => n2163, A4 => n2164
                           , ZN => n2155);
   U1148 : OAI22_X1 port map( A1 => n444, A2 => n1889, B1 => n411, B2 => n1890,
                           ZN => n2164);
   U1149 : OAI22_X1 port map( A1 => n511, A2 => n1891, B1 => n477, B2 => n1892,
                           ZN => n2163);
   U1150 : OAI22_X1 port map( A1 => n578, A2 => n1893, B1 => n545, B2 => n1894,
                           ZN => n2162);
   U1151 : OAI22_X1 port map( A1 => n645, A2 => n1895, B1 => n612, B2 => n1896,
                           ZN => n2161);
   U1152 : NOR4_X1 port map( A1 => n2165, A2 => n2166, A3 => n2167, A4 => n2168
                           , ZN => n2154);
   U1153 : OAI22_X1 port map( A1 => n713, A2 => n1901, B1 => n679, B2 => n1902,
                           ZN => n2168);
   U1154 : OAI22_X1 port map( A1 => n780, A2 => n1903, B1 => n746, B2 => n1904,
                           ZN => n2167);
   U1155 : OAI22_X1 port map( A1 => n847, A2 => n1905, B1 => n813, B2 => n1906,
                           ZN => n2166);
   U1156 : OAI22_X1 port map( A1 => n914, A2 => n1907, B1 => n881, B2 => n1908,
                           ZN => n2165);
   U1157 : NOR4_X1 port map( A1 => n2169, A2 => n2170, A3 => n2171, A4 => n2172
                           , ZN => n2153);
   U1158 : OAI22_X1 port map( A1 => n981, A2 => n1913, B1 => n948, B2 => n1914,
                           ZN => n2172);
   U1159 : OAI22_X1 port map( A1 => n1049, A2 => n1915, B1 => n1015, B2 => 
                           n1916, ZN => n2171);
   U1160 : OAI22_X1 port map( A1 => n87, A2 => n41, B1 => n1082, B2 => n43, ZN 
                           => n2170);
   U1161 : OAI22_X1 port map( A1 => n163, A2 => n1919, B1 => n128, B2 => n1920,
                           ZN => n2169);
   U1162 : OAI22_X1 port map( A1 => n2173, A2 => n1867, B1 => n1868, B2 => 
                           n1414, ZN => N4526);
   U1163 : NOR4_X1 port map( A1 => n2178, A2 => n2179, A3 => n2180, A4 => n2181
                           , ZN => n2177);
   U1164 : OAI22_X1 port map( A1 => n186, A2 => n1877, B1 => n816, B2 => n1878,
                           ZN => n2181);
   U1165 : OAI22_X1 port map( A1 => n250, A2 => n1879, B1 => n218, B2 => n1880,
                           ZN => n2180);
   U1166 : OAI22_X1 port map( A1 => n314, A2 => n1881, B1 => n282, B2 => n1882,
                           ZN => n2179);
   U1167 : OAI22_X1 port map( A1 => n378, A2 => n1883, B1 => n346, B2 => n1884,
                           ZN => n2178);
   U1168 : NOR4_X1 port map( A1 => n2182, A2 => n2183, A3 => n2184, A4 => n2185
                           , ZN => n2176);
   U1169 : OAI22_X1 port map( A1 => n443, A2 => n1889, B1 => n410, B2 => n1890,
                           ZN => n2185);
   U1170 : OAI22_X1 port map( A1 => n510, A2 => n1891, B1 => n476, B2 => n1892,
                           ZN => n2184);
   U1171 : OAI22_X1 port map( A1 => n577, A2 => n1893, B1 => n544, B2 => n1894,
                           ZN => n2183);
   U1172 : OAI22_X1 port map( A1 => n644, A2 => n1895, B1 => n611, B2 => n1896,
                           ZN => n2182);
   U1173 : NOR4_X1 port map( A1 => n2186, A2 => n2187, A3 => n2188, A4 => n2189
                           , ZN => n2175);
   U1174 : OAI22_X1 port map( A1 => n712, A2 => n1901, B1 => n678, B2 => n1902,
                           ZN => n2189);
   U1175 : OAI22_X1 port map( A1 => n779, A2 => n1903, B1 => n745, B2 => n1904,
                           ZN => n2188);
   U1176 : OAI22_X1 port map( A1 => n846, A2 => n1905, B1 => n812, B2 => n1906,
                           ZN => n2187);
   U1177 : OAI22_X1 port map( A1 => n913, A2 => n1907, B1 => n880, B2 => n1908,
                           ZN => n2186);
   U1178 : NOR4_X1 port map( A1 => n2190, A2 => n2191, A3 => n2192, A4 => n2193
                           , ZN => n2174);
   U1179 : OAI22_X1 port map( A1 => n980, A2 => n1913, B1 => n947, B2 => n1914,
                           ZN => n2193);
   U1180 : OAI22_X1 port map( A1 => n1048, A2 => n1915, B1 => n1014, B2 => 
                           n1916, ZN => n2192);
   U1181 : OAI22_X1 port map( A1 => n85, A2 => n41, B1 => n1081, B2 => n43, ZN 
                           => n2191);
   U1182 : OAI22_X1 port map( A1 => n162, A2 => n1919, B1 => n127, B2 => n1920,
                           ZN => n2190);
   U1183 : OAI22_X1 port map( A1 => n2194, A2 => n1867, B1 => n1868, B2 => 
                           n1436, ZN => N4524);
   U1184 : NOR4_X1 port map( A1 => n2199, A2 => n2200, A3 => n2201, A4 => n2202
                           , ZN => n2198);
   U1185 : OAI22_X1 port map( A1 => n185, A2 => n1877, B1 => n795, B2 => n1878,
                           ZN => n2202);
   U1186 : OAI22_X1 port map( A1 => n249, A2 => n1879, B1 => n217, B2 => n1880,
                           ZN => n2201);
   U1187 : OAI22_X1 port map( A1 => n313, A2 => n1881, B1 => n281, B2 => n1882,
                           ZN => n2200);
   U1188 : OAI22_X1 port map( A1 => n377, A2 => n1883, B1 => n345, B2 => n1884,
                           ZN => n2199);
   U1189 : NOR4_X1 port map( A1 => n2203, A2 => n2204, A3 => n2205, A4 => n2206
                           , ZN => n2197);
   U1190 : OAI22_X1 port map( A1 => n442, A2 => n1889, B1 => n409, B2 => n1890,
                           ZN => n2206);
   U1191 : OAI22_X1 port map( A1 => n509, A2 => n1891, B1 => n475, B2 => n1892,
                           ZN => n2205);
   U1192 : OAI22_X1 port map( A1 => n576, A2 => n1893, B1 => n542, B2 => n1894,
                           ZN => n2204);
   U1193 : OAI22_X1 port map( A1 => n643, A2 => n1895, B1 => n610, B2 => n1896,
                           ZN => n2203);
   U1194 : NOR4_X1 port map( A1 => n2207, A2 => n2208, A3 => n2209, A4 => n2210
                           , ZN => n2196);
   U1195 : OAI22_X1 port map( A1 => n710, A2 => n1901, B1 => n677, B2 => n1902,
                           ZN => n2210);
   U1196 : OAI22_X1 port map( A1 => n778, A2 => n1903, B1 => n744, B2 => n1904,
                           ZN => n2209);
   U1197 : OAI22_X1 port map( A1 => n845, A2 => n1905, B1 => n811, B2 => n1906,
                           ZN => n2208);
   U1198 : OAI22_X1 port map( A1 => n912, A2 => n1907, B1 => n878, B2 => n1908,
                           ZN => n2207);
   U1199 : NOR4_X1 port map( A1 => n2211, A2 => n2212, A3 => n2213, A4 => n2214
                           , ZN => n2195);
   U1200 : OAI22_X1 port map( A1 => n979, A2 => n1913, B1 => n946, B2 => n1914,
                           ZN => n2214);
   U1201 : OAI22_X1 port map( A1 => n1046, A2 => n1915, B1 => n1013, B2 => 
                           n1916, ZN => n2213);
   U1202 : OAI22_X1 port map( A1 => n83, A2 => n41, B1 => n1080, B2 => n43, ZN 
                           => n2212);
   U1203 : OAI22_X1 port map( A1 => n161, A2 => n1919, B1 => n126, B2 => n1920,
                           ZN => n2211);
   U1204 : OAI22_X1 port map( A1 => n2215, A2 => n1867, B1 => n1868, B2 => 
                           n1458, ZN => N4522);
   U1205 : NOR4_X1 port map( A1 => n2220, A2 => n2221, A3 => n2222, A4 => n2223
                           , ZN => n2219);
   U1206 : OAI22_X1 port map( A1 => n184, A2 => n1877, B1 => n774, B2 => n1878,
                           ZN => n2223);
   U1207 : OAI22_X1 port map( A1 => n248, A2 => n1879, B1 => n216, B2 => n1880,
                           ZN => n2222);
   U1208 : OAI22_X1 port map( A1 => n312, A2 => n1881, B1 => n280, B2 => n1882,
                           ZN => n2221);
   U1209 : OAI22_X1 port map( A1 => n376, A2 => n1883, B1 => n344, B2 => n1884,
                           ZN => n2220);
   U1210 : NOR4_X1 port map( A1 => n2224, A2 => n2225, A3 => n2226, A4 => n2227
                           , ZN => n2218);
   U1211 : OAI22_X1 port map( A1 => n441, A2 => n1889, B1 => n408, B2 => n1890,
                           ZN => n2227);
   U1212 : OAI22_X1 port map( A1 => n508, A2 => n1891, B1 => n474, B2 => n1892,
                           ZN => n2226);
   U1213 : OAI22_X1 port map( A1 => n575, A2 => n1893, B1 => n541, B2 => n1894,
                           ZN => n2225);
   U1214 : OAI22_X1 port map( A1 => n642, A2 => n1895, B1 => n609, B2 => n1896,
                           ZN => n2224);
   U1215 : NOR4_X1 port map( A1 => n2228, A2 => n2229, A3 => n2230, A4 => n2231
                           , ZN => n2217);
   U1216 : OAI22_X1 port map( A1 => n709, A2 => n1901, B1 => n676, B2 => n1902,
                           ZN => n2231);
   U1217 : OAI22_X1 port map( A1 => n777, A2 => n1903, B1 => n743, B2 => n1904,
                           ZN => n2230);
   U1218 : OAI22_X1 port map( A1 => n844, A2 => n1905, B1 => n810, B2 => n1906,
                           ZN => n2229);
   U1219 : OAI22_X1 port map( A1 => n911, A2 => n1907, B1 => n877, B2 => n1908,
                           ZN => n2228);
   U1220 : NOR4_X1 port map( A1 => n2232, A2 => n2233, A3 => n2234, A4 => n2235
                           , ZN => n2216);
   U1221 : OAI22_X1 port map( A1 => n978, A2 => n1913, B1 => n945, B2 => n1914,
                           ZN => n2235);
   U1222 : OAI22_X1 port map( A1 => n1045, A2 => n1915, B1 => n1012, B2 => 
                           n1916, ZN => n2234);
   U1223 : OAI22_X1 port map( A1 => n81, A2 => n41, B1 => n1079, B2 => n43, ZN 
                           => n2233);
   U1224 : OAI22_X1 port map( A1 => n160, A2 => n1919, B1 => n125, B2 => n1920,
                           ZN => n2232);
   U1225 : OAI22_X1 port map( A1 => n2236, A2 => n1867, B1 => n1868, B2 => 
                           n1480, ZN => N4520);
   U1226 : NOR4_X1 port map( A1 => n2241, A2 => n2242, A3 => n2243, A4 => n2244
                           , ZN => n2240);
   U1227 : OAI22_X1 port map( A1 => n183, A2 => n1877, B1 => n753, B2 => n1878,
                           ZN => n2244);
   U1228 : OAI22_X1 port map( A1 => n247, A2 => n1879, B1 => n215, B2 => n1880,
                           ZN => n2243);
   U1229 : OAI22_X1 port map( A1 => n311, A2 => n1881, B1 => n279, B2 => n1882,
                           ZN => n2242);
   U1230 : OAI22_X1 port map( A1 => n375, A2 => n1883, B1 => n343, B2 => n1884,
                           ZN => n2241);
   U1231 : NOR4_X1 port map( A1 => n2245, A2 => n2246, A3 => n2247, A4 => n2248
                           , ZN => n2239);
   U1232 : OAI22_X1 port map( A1 => n440, A2 => n1889, B1 => n407, B2 => n1890,
                           ZN => n2248);
   U1233 : OAI22_X1 port map( A1 => n507, A2 => n1891, B1 => n473, B2 => n1892,
                           ZN => n2247);
   U1234 : OAI22_X1 port map( A1 => n574, A2 => n1893, B1 => n540, B2 => n1894,
                           ZN => n2246);
   U1235 : OAI22_X1 port map( A1 => n641, A2 => n1895, B1 => n608, B2 => n1896,
                           ZN => n2245);
   U1236 : NOR4_X1 port map( A1 => n2249, A2 => n2250, A3 => n2251, A4 => n2252
                           , ZN => n2238);
   U1237 : OAI22_X1 port map( A1 => n708, A2 => n1901, B1 => n675, B2 => n1902,
                           ZN => n2252);
   U1238 : OAI22_X1 port map( A1 => n776, A2 => n1903, B1 => n742, B2 => n1904,
                           ZN => n2251);
   U1239 : OAI22_X1 port map( A1 => n843, A2 => n1905, B1 => n809, B2 => n1906,
                           ZN => n2250);
   U1240 : OAI22_X1 port map( A1 => n910, A2 => n1907, B1 => n876, B2 => n1908,
                           ZN => n2249);
   U1241 : NOR4_X1 port map( A1 => n2253, A2 => n2254, A3 => n2255, A4 => n2256
                           , ZN => n2237);
   U1242 : OAI22_X1 port map( A1 => n977, A2 => n1913, B1 => n944, B2 => n1914,
                           ZN => n2256);
   U1243 : OAI22_X1 port map( A1 => n1044, A2 => n1915, B1 => n1011, B2 => 
                           n1916, ZN => n2255);
   U1244 : OAI22_X1 port map( A1 => n79, A2 => n41, B1 => n1078, B2 => n43, ZN 
                           => n2254);
   U1245 : OAI22_X1 port map( A1 => n159, A2 => n1919, B1 => n124, B2 => n1920,
                           ZN => n2253);
   U1246 : OAI22_X1 port map( A1 => n2257, A2 => n1867, B1 => n1868, B2 => 
                           n1502, ZN => N4518);
   U1247 : NOR4_X1 port map( A1 => n2262, A2 => n2263, A3 => n2264, A4 => n2265
                           , ZN => n2261);
   U1248 : OAI22_X1 port map( A1 => n182, A2 => n1877, B1 => n732, B2 => n1878,
                           ZN => n2265);
   U1249 : OAI22_X1 port map( A1 => n246, A2 => n1879, B1 => n214, B2 => n1880,
                           ZN => n2264);
   U1250 : OAI22_X1 port map( A1 => n310, A2 => n1881, B1 => n278, B2 => n1882,
                           ZN => n2263);
   U1251 : OAI22_X1 port map( A1 => n374, A2 => n1883, B1 => n342, B2 => n1884,
                           ZN => n2262);
   U1252 : NOR4_X1 port map( A1 => n2266, A2 => n2267, A3 => n2268, A4 => n2269
                           , ZN => n2260);
   U1253 : OAI22_X1 port map( A1 => n439, A2 => n1889, B1 => n406, B2 => n1890,
                           ZN => n2269);
   U1254 : OAI22_X1 port map( A1 => n506, A2 => n1891, B1 => n472, B2 => n1892,
                           ZN => n2268);
   U1255 : OAI22_X1 port map( A1 => n573, A2 => n1893, B1 => n539, B2 => n1894,
                           ZN => n2267);
   U1256 : OAI22_X1 port map( A1 => n640, A2 => n1895, B1 => n607, B2 => n1896,
                           ZN => n2266);
   U1257 : NOR4_X1 port map( A1 => n2270, A2 => n2271, A3 => n2272, A4 => n2273
                           , ZN => n2259);
   U1258 : OAI22_X1 port map( A1 => n707, A2 => n1901, B1 => n674, B2 => n1902,
                           ZN => n2273);
   U1259 : OAI22_X1 port map( A1 => n775, A2 => n1903, B1 => n741, B2 => n1904,
                           ZN => n2272);
   U1260 : OAI22_X1 port map( A1 => n842, A2 => n1905, B1 => n808, B2 => n1906,
                           ZN => n2271);
   U1261 : OAI22_X1 port map( A1 => n909, A2 => n1907, B1 => n875, B2 => n1908,
                           ZN => n2270);
   U1262 : NOR4_X1 port map( A1 => n2274, A2 => n2275, A3 => n2276, A4 => n2277
                           , ZN => n2258);
   U1263 : OAI22_X1 port map( A1 => n976, A2 => n1913, B1 => n943, B2 => n1914,
                           ZN => n2277);
   U1264 : OAI22_X1 port map( A1 => n1043, A2 => n1915, B1 => n1010, B2 => 
                           n1916, ZN => n2276);
   U1265 : OAI22_X1 port map( A1 => n77, A2 => n41, B1 => n1077, B2 => n43, ZN 
                           => n2275);
   U1266 : OAI22_X1 port map( A1 => n158, A2 => n1919, B1 => n123, B2 => n1920,
                           ZN => n2274);
   U1267 : OAI22_X1 port map( A1 => n2278, A2 => n1867, B1 => n1868, B2 => 
                           n1524, ZN => N4516);
   U1268 : NOR4_X1 port map( A1 => n2283, A2 => n2284, A3 => n2285, A4 => n2286
                           , ZN => n2282);
   U1269 : OAI22_X1 port map( A1 => n181, A2 => n1877, B1 => n711, B2 => n1878,
                           ZN => n2286);
   U1270 : OAI22_X1 port map( A1 => n245, A2 => n1879, B1 => n213, B2 => n1880,
                           ZN => n2285);
   U1271 : OAI22_X1 port map( A1 => n309, A2 => n1881, B1 => n277, B2 => n1882,
                           ZN => n2284);
   U1272 : OAI22_X1 port map( A1 => n373, A2 => n1883, B1 => n341, B2 => n1884,
                           ZN => n2283);
   U1273 : NOR4_X1 port map( A1 => n2287, A2 => n2288, A3 => n2289, A4 => n2290
                           , ZN => n2281);
   U1274 : OAI22_X1 port map( A1 => n437, A2 => n1889, B1 => n405, B2 => n1890,
                           ZN => n2290);
   U1275 : OAI22_X1 port map( A1 => n505, A2 => n1891, B1 => n471, B2 => n1892,
                           ZN => n2289);
   U1276 : OAI22_X1 port map( A1 => n572, A2 => n1893, B1 => n538, B2 => n1894,
                           ZN => n2288);
   U1277 : OAI22_X1 port map( A1 => n639, A2 => n1895, B1 => n605, B2 => n1896,
                           ZN => n2287);
   U1278 : NOR4_X1 port map( A1 => n2291, A2 => n2292, A3 => n2293, A4 => n2294
                           , ZN => n2280);
   U1279 : OAI22_X1 port map( A1 => n706, A2 => n1901, B1 => n673, B2 => n1902,
                           ZN => n2294);
   U1280 : OAI22_X1 port map( A1 => n773, A2 => n1903, B1 => n740, B2 => n1904,
                           ZN => n2293);
   U1281 : OAI22_X1 port map( A1 => n841, A2 => n1905, B1 => n807, B2 => n1906,
                           ZN => n2292);
   U1282 : OAI22_X1 port map( A1 => n908, A2 => n1907, B1 => n874, B2 => n1908,
                           ZN => n2291);
   U1283 : NOR4_X1 port map( A1 => n2295, A2 => n2296, A3 => n2297, A4 => n2298
                           , ZN => n2279);
   U1284 : OAI22_X1 port map( A1 => n975, A2 => n1913, B1 => n941, B2 => n1914,
                           ZN => n2298);
   U1285 : OAI22_X1 port map( A1 => n1042, A2 => n1915, B1 => n1009, B2 => 
                           n1916, ZN => n2297);
   U1286 : OAI22_X1 port map( A1 => n73, A2 => n41, B1 => n1076, B2 => n43, ZN 
                           => n2296);
   U1287 : OAI22_X1 port map( A1 => n157, A2 => n1919, B1 => n122, B2 => n1920,
                           ZN => n2295);
   U1288 : OAI22_X1 port map( A1 => n2299, A2 => n1867, B1 => n1868, B2 => 
                           n1546, ZN => N4514);
   U1289 : NOR4_X1 port map( A1 => n2304, A2 => n2305, A3 => n2306, A4 => n2307
                           , ZN => n2303);
   U1290 : OAI22_X1 port map( A1 => n180, A2 => n1877, B1 => n690, B2 => n1878,
                           ZN => n2307);
   U1291 : OAI22_X1 port map( A1 => n244, A2 => n1879, B1 => n212, B2 => n1880,
                           ZN => n2306);
   U1292 : OAI22_X1 port map( A1 => n308, A2 => n1881, B1 => n276, B2 => n1882,
                           ZN => n2305);
   U1293 : OAI22_X1 port map( A1 => n372, A2 => n1883, B1 => n340, B2 => n1884,
                           ZN => n2304);
   U1294 : NOR4_X1 port map( A1 => n2308, A2 => n2309, A3 => n2310, A4 => n2311
                           , ZN => n2302);
   U1295 : OAI22_X1 port map( A1 => n436, A2 => n1889, B1 => n404, B2 => n1890,
                           ZN => n2311);
   U1296 : OAI22_X1 port map( A1 => n504, A2 => n1891, B1 => n470, B2 => n1892,
                           ZN => n2310);
   U1297 : OAI22_X1 port map( A1 => n571, A2 => n1893, B1 => n537, B2 => n1894,
                           ZN => n2309);
   U1298 : OAI22_X1 port map( A1 => n638, A2 => n1895, B1 => n604, B2 => n1896,
                           ZN => n2308);
   U1299 : NOR4_X1 port map( A1 => n2312, A2 => n2313, A3 => n2314, A4 => n2315
                           , ZN => n2301);
   U1300 : OAI22_X1 port map( A1 => n705, A2 => n1901, B1 => n672, B2 => n1902,
                           ZN => n2315);
   U1301 : OAI22_X1 port map( A1 => n772, A2 => n1903, B1 => n739, B2 => n1904,
                           ZN => n2314);
   U1302 : OAI22_X1 port map( A1 => n840, A2 => n1905, B1 => n806, B2 => n1906,
                           ZN => n2313);
   U1303 : OAI22_X1 port map( A1 => n907, A2 => n1907, B1 => n873, B2 => n1908,
                           ZN => n2312);
   U1304 : NOR4_X1 port map( A1 => n2316, A2 => n2317, A3 => n2318, A4 => n2319
                           , ZN => n2300);
   U1305 : OAI22_X1 port map( A1 => n974, A2 => n1913, B1 => n940, B2 => n1914,
                           ZN => n2319);
   U1306 : OAI22_X1 port map( A1 => n1041, A2 => n1915, B1 => n1008, B2 => 
                           n1916, ZN => n2318);
   U1307 : OAI22_X1 port map( A1 => n71, A2 => n41, B1 => n1075, B2 => n43, ZN 
                           => n2317);
   U1308 : OAI22_X1 port map( A1 => n156, A2 => n1919, B1 => n121, B2 => n1920,
                           ZN => n2316);
   U1309 : OAI22_X1 port map( A1 => n2320, A2 => n1867, B1 => n1868, B2 => 
                           n1568, ZN => N4512);
   U1310 : NOR4_X1 port map( A1 => n2325, A2 => n2326, A3 => n2327, A4 => n2328
                           , ZN => n2324);
   U1311 : OAI22_X1 port map( A1 => n179, A2 => n1877, B1 => n669, B2 => n1878,
                           ZN => n2328);
   U1312 : OAI22_X1 port map( A1 => n243, A2 => n1879, B1 => n211, B2 => n1880,
                           ZN => n2327);
   U1313 : OAI22_X1 port map( A1 => n307, A2 => n1881, B1 => n275, B2 => n1882,
                           ZN => n2326);
   U1314 : OAI22_X1 port map( A1 => n371, A2 => n1883, B1 => n339, B2 => n1884,
                           ZN => n2325);
   U1315 : NOR4_X1 port map( A1 => n2329, A2 => n2330, A3 => n2331, A4 => n2332
                           , ZN => n2323);
   U1316 : OAI22_X1 port map( A1 => n435, A2 => n1889, B1 => n403, B2 => n1890,
                           ZN => n2332);
   U1317 : OAI22_X1 port map( A1 => n503, A2 => n1891, B1 => n469, B2 => n1892,
                           ZN => n2331);
   U1318 : OAI22_X1 port map( A1 => n570, A2 => n1893, B1 => n536, B2 => n1894,
                           ZN => n2330);
   U1319 : OAI22_X1 port map( A1 => n637, A2 => n1895, B1 => n603, B2 => n1896,
                           ZN => n2329);
   U1320 : NOR4_X1 port map( A1 => n2333, A2 => n2334, A3 => n2335, A4 => n2336
                           , ZN => n2322);
   U1321 : OAI22_X1 port map( A1 => n704, A2 => n1901, B1 => n671, B2 => n1902,
                           ZN => n2336);
   U1322 : OAI22_X1 port map( A1 => n771, A2 => n1903, B1 => n738, B2 => n1904,
                           ZN => n2335);
   U1323 : OAI22_X1 port map( A1 => n839, A2 => n1905, B1 => n805, B2 => n1906,
                           ZN => n2334);
   U1324 : OAI22_X1 port map( A1 => n906, A2 => n39, B1 => n872, B2 => n1908, 
                           ZN => n2333);
   U1325 : NOR4_X1 port map( A1 => n2337, A2 => n2338, A3 => n2339, A4 => n2340
                           , ZN => n2321);
   U1326 : OAI22_X1 port map( A1 => n973, A2 => n1913, B1 => n939, B2 => n1914,
                           ZN => n2340);
   U1327 : OAI22_X1 port map( A1 => n1040, A2 => n1915, B1 => n1007, B2 => 
                           n1916, ZN => n2339);
   U1328 : OAI22_X1 port map( A1 => n69, A2 => n41, B1 => n1074, B2 => n1918, 
                           ZN => n2338);
   U1329 : OAI22_X1 port map( A1 => n155, A2 => n1919, B1 => n119, B2 => n1920,
                           ZN => n2337);
   U1330 : OAI22_X1 port map( A1 => n2341, A2 => n1867, B1 => n1868, B2 => 
                           n1590, ZN => N4510);
   U1331 : NOR4_X1 port map( A1 => n2346, A2 => n2347, A3 => n2348, A4 => n2349
                           , ZN => n2345);
   U1332 : OAI22_X1 port map( A1 => n178, A2 => n1877, B1 => n648, B2 => n1878,
                           ZN => n2349);
   U1333 : OAI22_X1 port map( A1 => n242, A2 => n1879, B1 => n210, B2 => n1880,
                           ZN => n2348);
   U1334 : OAI22_X1 port map( A1 => n306, A2 => n1881, B1 => n274, B2 => n1882,
                           ZN => n2347);
   U1335 : OAI22_X1 port map( A1 => n370, A2 => n1883, B1 => n338, B2 => n1884,
                           ZN => n2346);
   U1336 : NOR4_X1 port map( A1 => n2350, A2 => n2351, A3 => n2352, A4 => n2353
                           , ZN => n2344);
   U1337 : OAI22_X1 port map( A1 => n434, A2 => n1889, B1 => n402, B2 => n1890,
                           ZN => n2353);
   U1338 : OAI22_X1 port map( A1 => n502, A2 => n1891, B1 => n468, B2 => n1892,
                           ZN => n2352);
   U1339 : OAI22_X1 port map( A1 => n569, A2 => n1893, B1 => n535, B2 => n1894,
                           ZN => n2351);
   U1340 : OAI22_X1 port map( A1 => n636, A2 => n1895, B1 => n602, B2 => n1896,
                           ZN => n2350);
   U1341 : NOR4_X1 port map( A1 => n2354, A2 => n2355, A3 => n2356, A4 => n2357
                           , ZN => n2343);
   U1342 : OAI22_X1 port map( A1 => n703, A2 => n1901, B1 => n670, B2 => n1902,
                           ZN => n2357);
   U1343 : OAI22_X1 port map( A1 => n770, A2 => n1903, B1 => n737, B2 => n1904,
                           ZN => n2356);
   U1344 : OAI22_X1 port map( A1 => n838, A2 => n1905, B1 => n804, B2 => n1906,
                           ZN => n2355);
   U1345 : OAI22_X1 port map( A1 => n905, A2 => n39, B1 => n871, B2 => n1908, 
                           ZN => n2354);
   U1346 : NOR4_X1 port map( A1 => n2358, A2 => n2359, A3 => n2360, A4 => n2361
                           , ZN => n2342);
   U1347 : OAI22_X1 port map( A1 => n972, A2 => n1913, B1 => n938, B2 => n1914,
                           ZN => n2361);
   U1348 : OAI22_X1 port map( A1 => n1039, A2 => n1915, B1 => n1006, B2 => 
                           n1916, ZN => n2360);
   U1349 : OAI22_X1 port map( A1 => n67, A2 => n41, B1 => n1073, B2 => n1918, 
                           ZN => n2359);
   U1350 : OAI22_X1 port map( A1 => n154, A2 => n1919, B1 => n118, B2 => n1920,
                           ZN => n2358);
   U1351 : OAI22_X1 port map( A1 => n2362, A2 => n1867, B1 => n1868, B2 => 
                           n1612, ZN => N4508);
   U1352 : NOR4_X1 port map( A1 => n2367, A2 => n2368, A3 => n2369, A4 => n2370
                           , ZN => n2366);
   U1353 : OAI22_X1 port map( A1 => n175, A2 => n1877, B1 => n627, B2 => n1878,
                           ZN => n2370);
   U1354 : OAI22_X1 port map( A1 => n241, A2 => n1879, B1 => n209, B2 => n1880,
                           ZN => n2369);
   U1355 : OAI22_X1 port map( A1 => n305, A2 => n1881, B1 => n273, B2 => n1882,
                           ZN => n2368);
   U1356 : OAI22_X1 port map( A1 => n369, A2 => n1883, B1 => n337, B2 => n1884,
                           ZN => n2367);
   U1357 : NOR4_X1 port map( A1 => n2371, A2 => n2372, A3 => n2373, A4 => n2374
                           , ZN => n2365);
   U1358 : OAI22_X1 port map( A1 => n433, A2 => n1889, B1 => n401, B2 => n1890,
                           ZN => n2374);
   U1359 : OAI22_X1 port map( A1 => n500, A2 => n1891, B1 => n467, B2 => n1892,
                           ZN => n2373);
   U1360 : OAI22_X1 port map( A1 => n568, A2 => n1893, B1 => n534, B2 => n1894,
                           ZN => n2372);
   U1361 : OAI22_X1 port map( A1 => n635, A2 => n1895, B1 => n601, B2 => n1896,
                           ZN => n2371);
   U1362 : NOR4_X1 port map( A1 => n2375, A2 => n2376, A3 => n2377, A4 => n2378
                           , ZN => n2364);
   U1363 : OAI22_X1 port map( A1 => n702, A2 => n1901, B1 => n668, B2 => n1902,
                           ZN => n2378);
   U1364 : OAI22_X1 port map( A1 => n769, A2 => n1903, B1 => n736, B2 => n1904,
                           ZN => n2377);
   U1365 : OAI22_X1 port map( A1 => n836, A2 => n1905, B1 => n803, B2 => n1906,
                           ZN => n2376);
   U1366 : OAI22_X1 port map( A1 => n904, A2 => n39, B1 => n870, B2 => n1908, 
                           ZN => n2375);
   U1367 : NOR4_X1 port map( A1 => n2379, A2 => n2380, A3 => n2381, A4 => n2382
                           , ZN => n2363);
   U1368 : OAI22_X1 port map( A1 => n971, A2 => n1913, B1 => n937, B2 => n1914,
                           ZN => n2382);
   U1369 : OAI22_X1 port map( A1 => n1038, A2 => n1915, B1 => n1004, B2 => 
                           n1916, ZN => n2381);
   U1370 : OAI22_X1 port map( A1 => n65, A2 => n41, B1 => n1072, B2 => n1918, 
                           ZN => n2380);
   U1371 : OAI22_X1 port map( A1 => n152, A2 => n1919, B1 => n117, B2 => n1920,
                           ZN => n2379);
   U1372 : OAI22_X1 port map( A1 => n2383, A2 => n1867, B1 => n1868, B2 => 
                           n1634, ZN => N4506);
   U1373 : NOR4_X1 port map( A1 => n2388, A2 => n2389, A3 => n2390, A4 => n2391
                           , ZN => n2387);
   U1374 : OAI22_X1 port map( A1 => n164, A2 => n1877, B1 => n606, B2 => n1878,
                           ZN => n2391);
   U1375 : OAI22_X1 port map( A1 => n240, A2 => n1879, B1 => n208, B2 => n1880,
                           ZN => n2390);
   U1376 : OAI22_X1 port map( A1 => n304, A2 => n1881, B1 => n272, B2 => n1882,
                           ZN => n2389);
   U1377 : OAI22_X1 port map( A1 => n368, A2 => n1883, B1 => n336, B2 => n1884,
                           ZN => n2388);
   U1378 : NOR4_X1 port map( A1 => n2392, A2 => n2393, A3 => n2394, A4 => n2395
                           , ZN => n2386);
   U1379 : OAI22_X1 port map( A1 => n432, A2 => n1889, B1 => n400, B2 => n1890,
                           ZN => n2395);
   U1380 : OAI22_X1 port map( A1 => n499, A2 => n1891, B1 => n466, B2 => n1892,
                           ZN => n2394);
   U1381 : OAI22_X1 port map( A1 => n567, A2 => n1893, B1 => n533, B2 => n1894,
                           ZN => n2393);
   U1382 : OAI22_X1 port map( A1 => n634, A2 => n1895, B1 => n600, B2 => n1896,
                           ZN => n2392);
   U1383 : NOR4_X1 port map( A1 => n2396, A2 => n2397, A3 => n2398, A4 => n2399
                           , ZN => n2385);
   U1384 : OAI22_X1 port map( A1 => n701, A2 => n1901, B1 => n667, B2 => n1902,
                           ZN => n2399);
   U1385 : OAI22_X1 port map( A1 => n768, A2 => n1903, B1 => n735, B2 => n1904,
                           ZN => n2398);
   U1386 : OAI22_X1 port map( A1 => n835, A2 => n1905, B1 => n802, B2 => n1906,
                           ZN => n2397);
   U1387 : OAI22_X1 port map( A1 => n903, A2 => n39, B1 => n869, B2 => n1908, 
                           ZN => n2396);
   U1388 : NOR4_X1 port map( A1 => n2400, A2 => n2401, A3 => n2402, A4 => n2403
                           , ZN => n2384);
   U1389 : OAI22_X1 port map( A1 => n970, A2 => n1913, B1 => n936, B2 => n1914,
                           ZN => n2403);
   U1390 : OAI22_X1 port map( A1 => n1037, A2 => n1915, B1 => n1003, B2 => 
                           n1916, ZN => n2402);
   U1391 : OAI22_X1 port map( A1 => n63, A2 => n41, B1 => n1071, B2 => n1918, 
                           ZN => n2401);
   U1392 : OAI22_X1 port map( A1 => n151, A2 => n1919, B1 => n116, B2 => n45, 
                           ZN => n2400);
   U1393 : OAI22_X1 port map( A1 => n2404, A2 => n1867, B1 => n1868, B2 => 
                           n1656, ZN => N4504);
   U1394 : NOR4_X1 port map( A1 => n2409, A2 => n2410, A3 => n2411, A4 => n2412
                           , ZN => n2408);
   U1395 : OAI22_X1 port map( A1 => n153, A2 => n1877, B1 => n585, B2 => n1878,
                           ZN => n2412);
   U1396 : OAI22_X1 port map( A1 => n239, A2 => n1879, B1 => n207, B2 => n1880,
                           ZN => n2411);
   U1397 : OAI22_X1 port map( A1 => n303, A2 => n1881, B1 => n271, B2 => n1882,
                           ZN => n2410);
   U1398 : OAI22_X1 port map( A1 => n367, A2 => n1883, B1 => n335, B2 => n1884,
                           ZN => n2409);
   U1399 : NOR4_X1 port map( A1 => n2413, A2 => n2414, A3 => n2415, A4 => n2416
                           , ZN => n2407);
   U1400 : OAI22_X1 port map( A1 => n431, A2 => n1889, B1 => n399, B2 => n1890,
                           ZN => n2416);
   U1401 : OAI22_X1 port map( A1 => n498, A2 => n1891, B1 => n465, B2 => n1892,
                           ZN => n2415);
   U1402 : OAI22_X1 port map( A1 => n566, A2 => n1893, B1 => n532, B2 => n1894,
                           ZN => n2414);
   U1403 : OAI22_X1 port map( A1 => n633, A2 => n1895, B1 => n599, B2 => n1896,
                           ZN => n2413);
   U1404 : NOR4_X1 port map( A1 => n2417, A2 => n2418, A3 => n2419, A4 => n2420
                           , ZN => n2406);
   U1405 : OAI22_X1 port map( A1 => n700, A2 => n1901, B1 => n666, B2 => n1902,
                           ZN => n2420);
   U1406 : OAI22_X1 port map( A1 => n767, A2 => n1903, B1 => n734, B2 => n1904,
                           ZN => n2419);
   U1407 : OAI22_X1 port map( A1 => n834, A2 => n1905, B1 => n801, B2 => n1906,
                           ZN => n2418);
   U1408 : OAI22_X1 port map( A1 => n902, A2 => n39, B1 => n868, B2 => n1908, 
                           ZN => n2417);
   U1409 : NOR4_X1 port map( A1 => n2421, A2 => n2422, A3 => n2423, A4 => n2424
                           , ZN => n2405);
   U1410 : OAI22_X1 port map( A1 => n969, A2 => n1913, B1 => n935, B2 => n1914,
                           ZN => n2424);
   U1411 : OAI22_X1 port map( A1 => n1036, A2 => n1915, B1 => n1002, B2 => 
                           n1916, ZN => n2423);
   U1412 : OAI22_X1 port map( A1 => n61, A2 => n41, B1 => n1070, B2 => n1918, 
                           ZN => n2422);
   U1413 : OAI22_X1 port map( A1 => n150, A2 => n1919, B1 => n115, B2 => n1920,
                           ZN => n2421);
   U1414 : OAI22_X1 port map( A1 => n2425, A2 => n1867, B1 => n1868, B2 => 
                           n1678, ZN => N4502);
   U1415 : NOR4_X1 port map( A1 => n2430, A2 => n2431, A3 => n2432, A4 => n2433
                           , ZN => n2429);
   U1416 : OAI22_X1 port map( A1 => n142, A2 => n1877, B1 => n564, B2 => n1878,
                           ZN => n2433);
   U1417 : OAI22_X1 port map( A1 => n238, A2 => n1879, B1 => n206, B2 => n1880,
                           ZN => n2432);
   U1418 : OAI22_X1 port map( A1 => n302, A2 => n1881, B1 => n270, B2 => n1882,
                           ZN => n2431);
   U1419 : OAI22_X1 port map( A1 => n366, A2 => n1883, B1 => n334, B2 => n1884,
                           ZN => n2430);
   U1420 : NOR4_X1 port map( A1 => n2434, A2 => n2435, A3 => n2436, A4 => n2437
                           , ZN => n2428);
   U1421 : OAI22_X1 port map( A1 => n430, A2 => n1889, B1 => n398, B2 => n1890,
                           ZN => n2437);
   U1422 : OAI22_X1 port map( A1 => n497, A2 => n1891, B1 => n464, B2 => n1892,
                           ZN => n2436);
   U1423 : OAI22_X1 port map( A1 => n565, A2 => n1893, B1 => n531, B2 => n1894,
                           ZN => n2435);
   U1424 : OAI22_X1 port map( A1 => n632, A2 => n1895, B1 => n598, B2 => n1896,
                           ZN => n2434);
   U1425 : NOR4_X1 port map( A1 => n2438, A2 => n2439, A3 => n2440, A4 => n2441
                           , ZN => n2427);
   U1426 : OAI22_X1 port map( A1 => n699, A2 => n1901, B1 => n665, B2 => n1902,
                           ZN => n2441);
   U1427 : OAI22_X1 port map( A1 => n766, A2 => n1903, B1 => n733, B2 => n1904,
                           ZN => n2440);
   U1428 : OAI22_X1 port map( A1 => n833, A2 => n1905, B1 => n800, B2 => n1906,
                           ZN => n2439);
   U1429 : OAI22_X1 port map( A1 => n901, A2 => n39, B1 => n867, B2 => n1908, 
                           ZN => n2438);
   U1430 : NOR4_X1 port map( A1 => n2442, A2 => n2443, A3 => n2444, A4 => n2445
                           , ZN => n2426);
   U1431 : OAI22_X1 port map( A1 => n968, A2 => n1913, B1 => n934, B2 => n1914,
                           ZN => n2445);
   U1432 : OAI22_X1 port map( A1 => n1035, A2 => n1915, B1 => n1001, B2 => 
                           n1916, ZN => n2444);
   U1433 : OAI22_X1 port map( A1 => n59, A2 => n1917, B1 => n1069, B2 => n1918,
                           ZN => n2443);
   U1434 : OAI22_X1 port map( A1 => n149, A2 => n1919, B1 => n114, B2 => n45, 
                           ZN => n2442);
   U1435 : OAI22_X1 port map( A1 => n2446, A2 => n1867, B1 => n1868, B2 => 
                           n1700, ZN => N4500);
   U1436 : NOR4_X1 port map( A1 => n2451, A2 => n2452, A3 => n2453, A4 => n2454
                           , ZN => n2450);
   U1437 : OAI22_X1 port map( A1 => n131, A2 => n1877, B1 => n543, B2 => n1878,
                           ZN => n2454);
   U1438 : OAI22_X1 port map( A1 => n237, A2 => n1879, B1 => n205, B2 => n1880,
                           ZN => n2453);
   U1439 : OAI22_X1 port map( A1 => n301, A2 => n1881, B1 => n269, B2 => n1882,
                           ZN => n2452);
   U1440 : OAI22_X1 port map( A1 => n365, A2 => n1883, B1 => n333, B2 => n1884,
                           ZN => n2451);
   U1441 : NOR4_X1 port map( A1 => n2455, A2 => n2456, A3 => n2457, A4 => n2458
                           , ZN => n2449);
   U1442 : OAI22_X1 port map( A1 => n429, A2 => n1889, B1 => n397, B2 => n1890,
                           ZN => n2458);
   U1443 : OAI22_X1 port map( A1 => n496, A2 => n1891, B1 => n463, B2 => n1892,
                           ZN => n2457);
   U1444 : OAI22_X1 port map( A1 => n563, A2 => n1893, B1 => n530, B2 => n1894,
                           ZN => n2456);
   U1445 : OAI22_X1 port map( A1 => n631, A2 => n1895, B1 => n597, B2 => n1896,
                           ZN => n2455);
   U1446 : NOR4_X1 port map( A1 => n2459, A2 => n2460, A3 => n2461, A4 => n2462
                           , ZN => n2448);
   U1447 : OAI22_X1 port map( A1 => n698, A2 => n1901, B1 => n664, B2 => n1902,
                           ZN => n2462);
   U1448 : OAI22_X1 port map( A1 => n765, A2 => n1903, B1 => n731, B2 => n1904,
                           ZN => n2461);
   U1449 : OAI22_X1 port map( A1 => n832, A2 => n1905, B1 => n799, B2 => n1906,
                           ZN => n2460);
   U1450 : OAI22_X1 port map( A1 => n899, A2 => n39, B1 => n866, B2 => n1908, 
                           ZN => n2459);
   U1451 : NOR4_X1 port map( A1 => n2463, A2 => n2464, A3 => n2465, A4 => n2466
                           , ZN => n2447);
   U1452 : OAI22_X1 port map( A1 => n967, A2 => n1913, B1 => n933, B2 => n1914,
                           ZN => n2466);
   U1453 : OAI22_X1 port map( A1 => n1034, A2 => n1915, B1 => n1000, B2 => 
                           n1916, ZN => n2465);
   U1454 : OAI22_X1 port map( A1 => n57, A2 => n1917, B1 => n1067, B2 => n1918,
                           ZN => n2464);
   U1455 : OAI22_X1 port map( A1 => n148, A2 => n1919, B1 => n113, B2 => n1920,
                           ZN => n2463);
   U1456 : OAI22_X1 port map( A1 => n2467, A2 => n1867, B1 => n1868, B2 => 
                           n1722, ZN => N4498);
   U1457 : NOR4_X1 port map( A1 => n2472, A2 => n2473, A3 => n2474, A4 => n2475
                           , ZN => n2471);
   U1458 : OAI22_X1 port map( A1 => n120, A2 => n1877, B1 => n522, B2 => n1878,
                           ZN => n2475);
   U1459 : OAI22_X1 port map( A1 => n236, A2 => n1879, B1 => n204, B2 => n1880,
                           ZN => n2474);
   U1460 : OAI22_X1 port map( A1 => n300, A2 => n1881, B1 => n268, B2 => n1882,
                           ZN => n2473);
   U1461 : OAI22_X1 port map( A1 => n364, A2 => n1883, B1 => n332, B2 => n1884,
                           ZN => n2472);
   U1462 : NOR4_X1 port map( A1 => n2476, A2 => n2477, A3 => n2478, A4 => n2479
                           , ZN => n2470);
   U1463 : OAI22_X1 port map( A1 => n428, A2 => n1889, B1 => n396, B2 => n1890,
                           ZN => n2479);
   U1464 : OAI22_X1 port map( A1 => n495, A2 => n1891, B1 => n462, B2 => n1892,
                           ZN => n2478);
   U1465 : OAI22_X1 port map( A1 => n562, A2 => n1893, B1 => n529, B2 => n1894,
                           ZN => n2477);
   U1466 : OAI22_X1 port map( A1 => n630, A2 => n1895, B1 => n596, B2 => n1896,
                           ZN => n2476);
   U1467 : NOR4_X1 port map( A1 => n2480, A2 => n2481, A3 => n2482, A4 => n2483
                           , ZN => n2469);
   U1468 : OAI22_X1 port map( A1 => n697, A2 => n1901, B1 => n663, B2 => n1902,
                           ZN => n2483);
   U1469 : OAI22_X1 port map( A1 => n764, A2 => n1903, B1 => n730, B2 => n1904,
                           ZN => n2482);
   U1470 : OAI22_X1 port map( A1 => n831, A2 => n1905, B1 => n798, B2 => n1906,
                           ZN => n2481);
   U1471 : OAI22_X1 port map( A1 => n898, A2 => n39, B1 => n865, B2 => n1908, 
                           ZN => n2480);
   U1472 : NOR4_X1 port map( A1 => n2484, A2 => n2485, A3 => n2486, A4 => n2487
                           , ZN => n2468);
   U1473 : OAI22_X1 port map( A1 => n966, A2 => n1913, B1 => n932, B2 => n1914,
                           ZN => n2487);
   U1474 : OAI22_X1 port map( A1 => n1033, A2 => n1915, B1 => n999, B2 => n1916
                           , ZN => n2486);
   U1475 : OAI22_X1 port map( A1 => n55, A2 => n1917, B1 => n1066, B2 => n1918,
                           ZN => n2485);
   U1476 : OAI22_X1 port map( A1 => n147, A2 => n1919, B1 => n112, B2 => n1920,
                           ZN => n2484);
   U1477 : OAI22_X1 port map( A1 => n2488, A2 => n1867, B1 => n1868, B2 => 
                           n1744, ZN => N4496);
   U1478 : NOR4_X1 port map( A1 => n2489, A2 => n2490, A3 => n2491, A4 => n2492
                           , ZN => n2488);
   U1479 : OAI211_X1 port map( C1 => n1100, C2 => n1917, A => n2493, B => n2494
                           , ZN => n2492);
   U1480 : NOR4_X1 port map( A1 => n2495, A2 => n2496, A3 => n2497, A4 => n2498
                           , ZN => n2494);
   U1481 : OAI22_X1 port map( A1 => n109, A2 => n1877, B1 => n203, B2 => n1880,
                           ZN => n2498);
   U1482 : OAI22_X1 port map( A1 => n235, A2 => n1879, B1 => n267, B2 => n1882,
                           ZN => n2497);
   U1483 : OAI22_X1 port map( A1 => n299, A2 => n1881, B1 => n331, B2 => n1884,
                           ZN => n2496);
   U1484 : OAI22_X1 port map( A1 => n363, A2 => n1883, B1 => n395, B2 => n1890,
                           ZN => n2495);
   U1485 : NOR4_X1 port map( A1 => n2499, A2 => n2500, A3 => n2501, A4 => n2502
                           , ZN => n2493);
   U1486 : OAI22_X1 port map( A1 => n427, A2 => n1889, B1 => n461, B2 => n1892,
                           ZN => n2502);
   U1487 : OAI22_X1 port map( A1 => n494, A2 => n1891, B1 => n528, B2 => n1894,
                           ZN => n2501);
   U1488 : OAI22_X1 port map( A1 => n561, A2 => n1893, B1 => n595, B2 => n1896,
                           ZN => n2500);
   U1489 : OAI22_X1 port map( A1 => n629, A2 => n1895, B1 => n662, B2 => n1902,
                           ZN => n2499);
   U1490 : OAI211_X1 port map( C1 => n146, C2 => n1919, A => n2503_port, B => 
                           n2504, ZN => n2491);
   U1491 : NOR4_X1 port map( A1 => n2505, A2 => n2506, A3 => n2507, A4 => n2508
                           , ZN => n2504);
   U1492 : OAI22_X1 port map( A1 => n763, A2 => n1903, B1 => n797, B2 => n1906,
                           ZN => n2508);
   U1493 : OAI22_X1 port map( A1 => n696, A2 => n1901, B1 => n729, B2 => n1904,
                           ZN => n2507);
   U1494 : OAI22_X1 port map( A1 => n897, A2 => n39, B1 => n931, B2 => n1914, 
                           ZN => n2506);
   U1495 : OAI22_X1 port map( A1 => n830, A2 => n1905, B1 => n864, B2 => n1908,
                           ZN => n2505);
   U1496 : OAI22_X1 port map( A1 => n1878, A2 => n501, B1 => n45, B2 => n111, 
                           ZN => n2509);
   U1497 : OAI22_X1 port map( A1 => n1032, A2 => n1915, B1 => n1065, B2 => 
                           n1918, ZN => n2490);
   U1498 : OAI22_X1 port map( A1 => n965, A2 => n1913, B1 => n998, B2 => n1916,
                           ZN => n2489);
   U1499 : OAI22_X1 port map( A1 => n2510, A2 => n1867, B1 => n1868, B2 => 
                           n1766, ZN => N4494);
   U1500 : NOR4_X1 port map( A1 => n2515, A2 => n2516, A3 => n2517, A4 => n2518
                           , ZN => n2514);
   U1501 : OAI22_X1 port map( A1 => n97, A2 => n1877, B1 => n480, B2 => n1878, 
                           ZN => n2518);
   U1502 : OAI22_X1 port map( A1 => n234, A2 => n1879, B1 => n202, B2 => n1880,
                           ZN => n2517);
   U1503 : OAI22_X1 port map( A1 => n298, A2 => n1881, B1 => n266, B2 => n1882,
                           ZN => n2516);
   U1504 : OAI22_X1 port map( A1 => n362, A2 => n1883, B1 => n330, B2 => n1884,
                           ZN => n2515);
   U1505 : NOR4_X1 port map( A1 => n2519, A2 => n2520, A3 => n2521, A4 => n2522
                           , ZN => n2513);
   U1506 : OAI22_X1 port map( A1 => n426, A2 => n1889, B1 => n394, B2 => n1890,
                           ZN => n2522);
   U1507 : OAI22_X1 port map( A1 => n493, A2 => n1891, B1 => n460, B2 => n1892,
                           ZN => n2521);
   U1508 : OAI22_X1 port map( A1 => n560, A2 => n1893, B1 => n527, B2 => n1894,
                           ZN => n2520);
   U1509 : OAI22_X1 port map( A1 => n628, A2 => n1895, B1 => n594, B2 => n1896,
                           ZN => n2519);
   U1510 : NOR4_X1 port map( A1 => n2523, A2 => n2524, A3 => n2525, A4 => n2526
                           , ZN => n2512);
   U1511 : OAI22_X1 port map( A1 => n695, A2 => n1901, B1 => n661, B2 => n1902,
                           ZN => n2526);
   U1512 : OAI22_X1 port map( A1 => n762, A2 => n1903, B1 => n728, B2 => n1904,
                           ZN => n2525);
   U1513 : OAI22_X1 port map( A1 => n829, A2 => n1905, B1 => n796, B2 => n1906,
                           ZN => n2524);
   U1514 : OAI22_X1 port map( A1 => n896, A2 => n39, B1 => n863, B2 => n1908, 
                           ZN => n2523);
   U1515 : NOR4_X1 port map( A1 => n2527, A2 => n2528, A3 => n2529, A4 => n2530
                           , ZN => n2511);
   U1516 : OAI22_X1 port map( A1 => n964, A2 => n1913, B1 => n930, B2 => n1914,
                           ZN => n2530);
   U1517 : OAI22_X1 port map( A1 => n1031, A2 => n1915, B1 => n997, B2 => n1916
                           , ZN => n2529);
   U1518 : OAI22_X1 port map( A1 => n1099, A2 => n1917, B1 => n1064, B2 => 
                           n1918, ZN => n2528);
   U1519 : OAI22_X1 port map( A1 => n145, A2 => n1919, B1 => n110, B2 => n1920,
                           ZN => n2527);
   U1520 : OAI22_X1 port map( A1 => n2531, A2 => n1867, B1 => n1868, B2 => 
                           n1788, ZN => N4492);
   U1521 : NOR4_X1 port map( A1 => n2536, A2 => n2537, A3 => n2538, A4 => n2539
                           , ZN => n2535);
   U1522 : OAI22_X1 port map( A1 => n75, A2 => n1877, B1 => n459, B2 => n1878, 
                           ZN => n2539);
   U1523 : OAI22_X1 port map( A1 => n233, A2 => n1879, B1 => n201, B2 => n1880,
                           ZN => n2538);
   U1524 : OAI22_X1 port map( A1 => n297, A2 => n1881, B1 => n265, B2 => n1882,
                           ZN => n2537);
   U1525 : OAI22_X1 port map( A1 => n361, A2 => n1883, B1 => n329, B2 => n1884,
                           ZN => n2536);
   U1526 : NOR4_X1 port map( A1 => n2540, A2 => n2541, A3 => n2542, A4 => n2543
                           , ZN => n2534);
   U1527 : OAI22_X1 port map( A1 => n425, A2 => n1889, B1 => n393, B2 => n1890,
                           ZN => n2543);
   U1528 : OAI22_X1 port map( A1 => n492, A2 => n1891, B1 => n458, B2 => n1892,
                           ZN => n2542);
   U1529 : OAI22_X1 port map( A1 => n559, A2 => n1893, B1 => n526, B2 => n1894,
                           ZN => n2541);
   U1530 : OAI22_X1 port map( A1 => n626, A2 => n1895, B1 => n593, B2 => n1896,
                           ZN => n2540);
   U1531 : NOR4_X1 port map( A1 => n2544, A2 => n2545, A3 => n2546, A4 => n2547
                           , ZN => n2533);
   U1532 : OAI22_X1 port map( A1 => n694, A2 => n1901, B1 => n660, B2 => n1902,
                           ZN => n2547);
   U1533 : OAI22_X1 port map( A1 => n761, A2 => n1903, B1 => n727, B2 => n1904,
                           ZN => n2546);
   U1534 : OAI22_X1 port map( A1 => n828, A2 => n1905, B1 => n794, B2 => n1906,
                           ZN => n2545);
   U1535 : OAI22_X1 port map( A1 => n895, A2 => n39, B1 => n862, B2 => n1908, 
                           ZN => n2544);
   U1536 : NOR4_X1 port map( A1 => n2548, A2 => n2549, A3 => n2550, A4 => n2551
                           , ZN => n2532);
   U1537 : OAI22_X1 port map( A1 => n962, A2 => n1913, B1 => n929, B2 => n1914,
                           ZN => n2551);
   U1538 : OAI22_X1 port map( A1 => n1030, A2 => n1915, B1 => n996, B2 => n1916
                           , ZN => n2550);
   U1539 : OAI22_X1 port map( A1 => n1098, A2 => n1917, B1 => n1063, B2 => 
                           n1918, ZN => n2549);
   U1540 : OAI22_X1 port map( A1 => n144, A2 => n1919, B1 => n108, B2 => n1920,
                           ZN => n2548);
   U1541 : OAI22_X1 port map( A1 => n2552, A2 => n1867, B1 => n1868, B2 => 
                           n1810, ZN => N4490);
   U1542 : OAI221_X1 port map( B1 => n1825, B2 => ADD_RD1(2), C1 => n1826, C2 
                           => ADD_RD1(0), A => n2557, ZN => n2556);
   U1543 : AOI22_X1 port map( A1 => n1825, A2 => ADD_RD1(2), B1 => n1826, B2 =>
                           ADD_RD1(0), ZN => n2557);
   U1544 : AOI221_X1 port map( B1 => n2558, B2 => ADD_WR(4), C1 => n1829, C2 =>
                           ADD_RD1(3), A => n2559, ZN => n2553);
   U1545 : OAI22_X1 port map( A1 => ADD_WR(4), A2 => n2558, B1 => n1829, B2 => 
                           ADD_RD1(3), ZN => n2559);
   U1546 : NOR4_X1 port map( A1 => n2568, A2 => n2569, A3 => n2570, A4 => n2571
                           , ZN => n2567_port);
   U1547 : OAI22_X1 port map( A1 => n53, A2 => n1877, B1 => n438, B2 => n1878, 
                           ZN => n2571);
   U1548 : OAI22_X1 port map( A1 => n232, A2 => n1879, B1 => n200, B2 => n1880,
                           ZN => n2570);
   U1549 : OAI22_X1 port map( A1 => n296, A2 => n1881, B1 => n264, B2 => n1882,
                           ZN => n2569);
   U1550 : OAI22_X1 port map( A1 => n360, A2 => n1883, B1 => n328, B2 => n1884,
                           ZN => n2568);
   U1551 : NOR3_X1 port map( A1 => n2558, A2 => n2578, A3 => n2579, ZN => n2573
                           );
   U1552 : NAND2_X1 port map( A1 => ADD_RD1(4), A2 => ADD_RD1(3), ZN => n2580);
   U1553 : NOR4_X1 port map( A1 => n2581, A2 => n2582, A3 => n2583, A4 => n2584
                           , ZN => n2566);
   U1554 : OAI22_X1 port map( A1 => n424, A2 => n1889, B1 => n392, B2 => n1890,
                           ZN => n2584);
   U1555 : OAI22_X1 port map( A1 => n491, A2 => n1891, B1 => n457, B2 => n1892,
                           ZN => n2583);
   U1556 : OAI22_X1 port map( A1 => n558, A2 => n1893, B1 => n525, B2 => n1894,
                           ZN => n2582);
   U1557 : OAI22_X1 port map( A1 => n625, A2 => n1895, B1 => n592, B2 => n1896,
                           ZN => n2581);
   U1558 : NOR3_X1 port map( A1 => ADD_RD1(3), A2 => n2558, A3 => n2579, ZN => 
                           n2585);
   U1559 : NOR3_X1 port map( A1 => ADD_RD1(3), A2 => ADD_RD1(0), A3 => n2558, 
                           ZN => n2586);
   U1560 : NOR4_X1 port map( A1 => n2587, A2 => n2588, A3 => n2589, A4 => n2590
                           , ZN => n2565);
   U1561 : OAI22_X1 port map( A1 => n693, A2 => n1901, B1 => n659, B2 => n1902,
                           ZN => n2590);
   U1562 : OAI22_X1 port map( A1 => n760, A2 => n1903, B1 => n726, B2 => n1904,
                           ZN => n2589);
   U1563 : OAI22_X1 port map( A1 => n827, A2 => n1905, B1 => n793, B2 => n1906,
                           ZN => n2588);
   U1564 : OAI22_X1 port map( A1 => n894, A2 => n39, B1 => n861, B2 => n1908, 
                           ZN => n2587);
   U1565 : NOR3_X1 port map( A1 => ADD_RD1(4), A2 => n2578, A3 => n2579, ZN => 
                           n2591);
   U1566 : NAND2_X1 port map( A1 => n2577, A2 => n2592, ZN => n1907);
   U1567 : NOR3_X1 port map( A1 => ADD_RD1(4), A2 => ADD_RD1(0), A3 => n2578, 
                           ZN => n2592);
   U1568 : NOR4_X1 port map( A1 => n2593, A2 => n2594, A3 => n2595, A4 => n2596
                           , ZN => n2564);
   U1569 : OAI22_X1 port map( A1 => n961, A2 => n1913, B1 => n928, B2 => n1914,
                           ZN => n2596);
   U1570 : OAI22_X1 port map( A1 => n1029, A2 => n1915, B1 => n995, B2 => n1916
                           , ZN => n2595);
   U1571 : OAI22_X1 port map( A1 => n1097, A2 => n1917, B1 => n1062, B2 => 
                           n1918, ZN => n2594);
   U1572 : NAND2_X1 port map( A1 => n2576, A2 => n2597, ZN => n1918);
   U1573 : NAND2_X1 port map( A1 => n2598, A2 => n2576, ZN => n1917);
   U1574 : OAI22_X1 port map( A1 => n143, A2 => n1919, B1 => n107, B2 => n45, 
                           ZN => n2593);
   U1575 : NAND2_X1 port map( A1 => n2577, A2 => n2597, ZN => n1920);
   U1576 : NOR3_X1 port map( A1 => ADD_RD1(4), A2 => ADD_RD1(3), A3 => n2579, 
                           ZN => n2597);
   U1577 : NOR3_X1 port map( A1 => ADD_RD1(4), A2 => ADD_RD1(3), A3 => 
                           ADD_RD1(0), ZN => n2598);
   U1578 : OAI21_X1 port map( B1 => n2599, B2 => n2600, A => n47, ZN => N4423);
   U1579 : OAI21_X1 port map( B1 => n2600, B2 => n2601, A => n47, ZN => N4359);
   U1580 : OAI21_X1 port map( B1 => n2600, B2 => n2602, A => n47, ZN => N4295);
   U1581 : OAI21_X1 port map( B1 => n2600, B2 => n2603, A => n47, ZN => N4231);
   U1582 : OAI21_X1 port map( B1 => n2600, B2 => n2604, A => n47, ZN => N4167);
   U1583 : OAI21_X1 port map( B1 => n2600, B2 => n2605, A => n47, ZN => N4103);
   U1584 : OAI21_X1 port map( B1 => n2600, B2 => n2606, A => n47, ZN => N4039);
   U1585 : NAND2_X1 port map( A1 => n2561, A2 => WR, ZN => n2600);
   U1586 : OAI21_X1 port map( B1 => n2563, B2 => n2607, A => n49, ZN => N3975);
   U1587 : OAI21_X1 port map( B1 => n2599, B2 => n2607, A => n51, ZN => N3911);
   U1588 : OAI21_X1 port map( B1 => n2607, B2 => n2601, A => n49, ZN => N3847);
   U1589 : OAI21_X1 port map( B1 => n2607, B2 => n2602, A => n49, ZN => N3783);
   U1590 : OAI21_X1 port map( B1 => n2607, B2 => n2603, A => n49, ZN => N3719);
   U1591 : OAI21_X1 port map( B1 => n2607, B2 => n2604, A => n49, ZN => N3655);
   U1592 : OAI21_X1 port map( B1 => n2607, B2 => n2605, A => n49, ZN => N3591);
   U1593 : OAI21_X1 port map( B1 => n2607, B2 => n2606, A => n49, ZN => N3527);
   U1594 : INV_X1 port map( A => WR, ZN => n2562);
   U1595 : OAI21_X1 port map( B1 => n2563, B2 => n2608, A => n49, ZN => N3463);
   U1596 : OAI21_X1 port map( B1 => n2599, B2 => n2608, A => n47, ZN => N3399);
   U1597 : OAI21_X1 port map( B1 => n2608, B2 => n2601, A => n49, ZN => N3335);
   U1598 : OAI21_X1 port map( B1 => n2608, B2 => n2602, A => n49, ZN => N3271);
   U1599 : OAI21_X1 port map( B1 => n2608, B2 => n2603, A => n47, ZN => N3207);
   U1600 : OAI21_X1 port map( B1 => n2608, B2 => n2604, A => n47, ZN => N3143);
   U1601 : OAI21_X1 port map( B1 => n2608, B2 => n2605, A => n51, ZN => N3079);
   U1602 : OAI21_X1 port map( B1 => n2608, B2 => n2606, A => n49, ZN => N3015);
   U1603 : NAND3_X1 port map( A1 => ADD_WR(4), A2 => WR, A3 => n1829, ZN => 
                           n2608);
   U1604 : OAI21_X1 port map( B1 => n2563, B2 => n2609, A => n51, ZN => N2951);
   U1605 : OAI21_X1 port map( B1 => n2599, B2 => n2609, A => n49, ZN => N2887);
   U1606 : NAND3_X1 port map( A1 => ADD_WR(0), A2 => n1825, A3 => n1823, ZN => 
                           n2599);
   U1607 : OAI21_X1 port map( B1 => n2609, B2 => n2601, A => n47, ZN => N2823);
   U1608 : NAND3_X1 port map( A1 => ADD_WR(1), A2 => n1826, A3 => n1825, ZN => 
                           n2601);
   U1609 : OAI21_X1 port map( B1 => n2609, B2 => n2602, A => n47, ZN => N2759);
   U1610 : NAND3_X1 port map( A1 => ADD_WR(0), A2 => ADD_WR(1), A3 => n1825, ZN
                           => n2602);
   U1611 : OAI21_X1 port map( B1 => n2609, B2 => n2603, A => n51, ZN => N2695);
   U1612 : NAND3_X1 port map( A1 => ADD_WR(2), A2 => n1826, A3 => n1823, ZN => 
                           n2603);
   U1613 : OAI21_X1 port map( B1 => n2609, B2 => n2604, A => n49, ZN => N2631);
   U1614 : NAND3_X1 port map( A1 => ADD_WR(2), A2 => ADD_WR(0), A3 => n1823, ZN
                           => n2604);
   U1615 : OAI21_X1 port map( B1 => n2609, B2 => n2605, A => n49, ZN => N2567);
   U1616 : NAND3_X1 port map( A1 => ADD_WR(2), A2 => ADD_WR(1), A3 => n1826, ZN
                           => n2605);
   U1617 : OAI21_X1 port map( B1 => n2609, B2 => n2606, A => n51, ZN => N2503);
   U1618 : NAND3_X1 port map( A1 => ADD_WR(0), A2 => ADD_WR(2), A3 => ADD_WR(1)
                           , ZN => n2606);
   U1619 : NAND3_X1 port map( A1 => ADD_WR(4), A2 => ADD_WR(3), A3 => WR, ZN =>
                           n2609);

end SYN_A;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity 
   dlx_cu_MICROCODE_MEM_SIZE64_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE13 is

   port( Clk, Rst : in std_logic;  IR_IN : in std_logic_vector (31 downto 0);  
         stall_exe_i, mispredict_i : in std_logic;  D1_i, D2_i : in 
         std_logic_vector (4 downto 0);  S1_LATCH_EN, S2_LATCH_EN, S3_LATCH_EN 
         : out std_logic;  S_MUX_PC_BUS : out std_logic_vector (1 downto 0);  
         S_EXT, S_EXT_SIGN, S_EQ_NEQ : out std_logic;  S_MUX_DEST : out 
         std_logic_vector (1 downto 0);  S_MUX_LINK, S_MEM_W_R, S_MEM_EN, 
         S_RF_W_wb, S_RF_W_mem, S_RF_W_exe, S_MUX_ALUIN, stall_exe_o, 
         stall_dec_o, stall_fetch_o, stall_btb_o, was_branch_o, was_jmp_o : out
         std_logic;  ALU_WORD_o : out std_logic_vector (12 downto 0);  
         ALU_OPCODE : out std_logic_vector (0 to 4);  S_MUX_MEM_BAR : out 
         std_logic);

end dlx_cu_MICROCODE_MEM_SIZE64_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE13;

architecture SYN_dlx_cu_hw of 
   dlx_cu_MICROCODE_MEM_SIZE64_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE13 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X2
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFR_X2
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component 
      SNPS_CLOCK_GATE_HIGH_dlx_cu_MICROCODE_MEM_SIZE64_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE13_0
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component alu_ctrl
      port( OP : in std_logic_vector (0 to 4);  ALU_WORD : out std_logic_vector
            (12 downto 0));
   end component;
   
   component cw_mem_MICROCODE_MEM_SIZE64_OP_CODE_SIZE6_CW_SIZE13
      port( OPCODE_IN : in std_logic_vector (5 downto 0);  CW_OUT : out 
            std_logic_vector (12 downto 0));
   end component;
   
   component stall_logic_FUNC_SIZE11_OP_CODE_SIZE6
      port( OPCODE_i : in std_logic_vector (5 downto 0);  FUNC_i : in 
            std_logic_vector (10 downto 0);  rA_i, rB_i, D1_i, D2_i : in 
            std_logic_vector (4 downto 0);  S_mem_LOAD_i, S_exe_LOAD_i, 
            S_exe_WRITE_i : in std_logic;  S_MUX_PC_BUS_i : in std_logic_vector
            (1 downto 0);  mispredict_i : in std_logic;  bubble_dec_o, 
            bubble_exe_o, stall_exe_o, stall_dec_o, stall_btb_o, stall_fetch_o 
            : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFS_X1
      port( D, CK, SN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal S_MUX_PC_BUS_1_port, S_MUX_PC_BUS_0_port, S_MEM_W_R_port, n130, 
      S_MEM_LOAD, S_EXE_LOAD, next_bubble_dec, stall_dec_o_TEMP, 
      stall_btb_o_TEMP, stall_fetch_o_TEMP, cw_from_mem_12_port, 
      cw_from_mem_11_port, cw_from_mem_10_port, cw_from_mem_9_port, 
      cw_from_mem_8_port, cw_from_mem_7_port, cw_from_mem_6_port, 
      cw_from_mem_5_port, cw_from_mem_4_port, cw_from_mem_3_port, 
      cw_from_mem_2_port, cw_from_mem_1_port, cw_from_mem_0_port, 
      aluOpcode_d_4_port, aluOpcode_d_3_port, aluOpcode_d_2_port, 
      aluOpcode_d_1_port, aluOpcode_d_0_port, N20, N21, N22, N23, N24, N25, N26
      , N27, N29, N30, N31, N32, net3570, n2, n3, n4, n5, n15, n16, n17, n18, 
      n19, n20_port, n21_port, n22_port, n23_port, n24_port, n25_port, n26_port
      , n27_port, n28, n31_port, n33, n34, n37, n38, n39, n40, n41, n43, n44, 
      n45, n46, n47, n48, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60
      , n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n73, n74, n75, 
      n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n89, n90, n91
      , n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, 
      n105, n106, n111, n114, n115, n116, n117, n118, n120, n121, n123, n124, 
      n125, n1, n6, n7, n8, n9, n10, n11, n12, n13, n14, n29_port, n30_port, 
      n32_port, n35, n36, n42, n49, n72, n88, n107, n108, n109, n110, n112, 
      n113, n122, n126, n127, n128, n129, net47684, net47685, net47686, 
      net47687, net47688 : std_logic;

begin
   S_MUX_PC_BUS <= ( S_MUX_PC_BUS_1_port, S_MUX_PC_BUS_0_port );
   S_MEM_W_R <= S_MEM_W_R_port;
   stall_exe_o <= stall_exe_i;
   
   bubble_dec_reg : DFF_X1 port map( D => n123, CK => Clk, Q => n36, QN => n124
                           );
   cw_e_reg_0_inst : DFFR_X1 port map( D => N21, CK => net3570, RN => n49, Q =>
                           n130, QN => n2);
   cw_e_reg_5_inst : DFFR_X1 port map( D => N26, CK => net3570, RN => n49, Q =>
                           S_MUX_DEST(1), QN => n121);
   cw_e_reg_4_inst : DFFR_X1 port map( D => N25, CK => net3570, RN => n49, Q =>
                           S_MUX_DEST(0), QN => n120);
   cw_e_reg_3_inst : DFFR_X1 port map( D => N24, CK => net3570, RN => n49, Q =>
                           n3, QN => net47688);
   cw_m_reg_3_inst : DFFR_X1 port map( D => N32, CK => Clk, RN => n49, Q => 
                           S_MEM_EN, QN => n125);
   cw_m_reg_2_inst : DFFR_X1 port map( D => N31, CK => Clk, RN => n49, Q => 
                           S_MEM_W_R_port, QN => net47687);
   cw_m_reg_1_inst : DFFR_X1 port map( D => N30, CK => Clk, RN => n49, Q => 
                           net47686, QN => S_MUX_MEM_BAR);
   cw_m_reg_0_inst : DFFR_X1 port map( D => N29, CK => Clk, RN => n49, Q => 
                           S_RF_W_mem, QN => n118);
   cw_w_reg_0_inst : DFFS_X1 port map( D => n118, CK => Clk, SN => n49, Q => 
                           n117, QN => S_RF_W_wb);
   U3 : XOR2_X1 port map( A => S_MUX_PC_BUS_1_port, B => S_MUX_PC_BUS_0_port, Z
                           => was_jmp_o);
   U8 : MUX2_X1 port map( A => next_bubble_dec, B => n36, S => Rst, Z => n123);
   U59 : NAND3_X1 port map( A1 => IR_IN(3), A2 => n77, A3 => n78, ZN => n70);
   U67 : NAND3_X1 port map( A1 => IR_IN(4), A2 => IR_IN(5), A3 => IR_IN(0), ZN 
                           => n64);
   U71 : NAND3_X1 port map( A1 => IR_IN(4), A2 => n77, A3 => n91, ZN => n71);
   U82 : NAND3_X1 port map( A1 => n48, A2 => n101, A3 => n46, ZN => n76);
   U122 : NAND3_X1 port map( A1 => IR_IN(2), A2 => IR_IN(3), A3 => n63, ZN => 
                           n27_port);
   U128 : NAND3_X1 port map( A1 => n43, A2 => n114, A3 => n115, ZN => n93);
   STALL_L : stall_logic_FUNC_SIZE11_OP_CODE_SIZE6 port map( OPCODE_i(5) => 
                           IR_IN(31), OPCODE_i(4) => IR_IN(30), OPCODE_i(3) => 
                           IR_IN(29), OPCODE_i(2) => IR_IN(28), OPCODE_i(1) => 
                           IR_IN(27), OPCODE_i(0) => IR_IN(26), FUNC_i(10) => 
                           n72, FUNC_i(9) => n88, FUNC_i(8) => n107, FUNC_i(7) 
                           => n108, FUNC_i(6) => n109, FUNC_i(5) => n110, 
                           FUNC_i(4) => n112, FUNC_i(3) => n113, FUNC_i(2) => 
                           n122, FUNC_i(1) => n126, FUNC_i(0) => n127, rA_i(4) 
                           => IR_IN(25), rA_i(3) => IR_IN(24), rA_i(2) => 
                           IR_IN(23), rA_i(1) => IR_IN(22), rA_i(0) => 
                           IR_IN(21), rB_i(4) => IR_IN(20), rB_i(3) => 
                           IR_IN(19), rB_i(2) => IR_IN(18), rB_i(1) => 
                           IR_IN(17), rB_i(0) => IR_IN(16), D1_i(4) => D1_i(4),
                           D1_i(3) => D1_i(3), D1_i(2) => D1_i(2), D1_i(1) => 
                           D1_i(1), D1_i(0) => D1_i(0), D2_i(4) => D2_i(4), 
                           D2_i(3) => D2_i(3), D2_i(2) => D2_i(2), D2_i(1) => 
                           D2_i(1), D2_i(0) => D2_i(0), S_mem_LOAD_i => 
                           S_MEM_LOAD, S_exe_LOAD_i => S_EXE_LOAD, 
                           S_exe_WRITE_i => n130, S_MUX_PC_BUS_i(1) => n128, 
                           S_MUX_PC_BUS_i(0) => n129, mispredict_i => 
                           mispredict_i, bubble_dec_o => next_bubble_dec, 
                           bubble_exe_o => net47684, stall_exe_o => net47685, 
                           stall_dec_o => stall_dec_o_TEMP, stall_btb_o => 
                           stall_btb_o_TEMP, stall_fetch_o => 
                           stall_fetch_o_TEMP);
   CWM : cw_mem_MICROCODE_MEM_SIZE64_OP_CODE_SIZE6_CW_SIZE13 port map( 
                           OPCODE_IN(5) => IR_IN(31), OPCODE_IN(4) => IR_IN(30)
                           , OPCODE_IN(3) => IR_IN(29), OPCODE_IN(2) => 
                           IR_IN(28), OPCODE_IN(1) => IR_IN(27), OPCODE_IN(0) 
                           => IR_IN(26), CW_OUT(12) => cw_from_mem_12_port, 
                           CW_OUT(11) => cw_from_mem_11_port, CW_OUT(10) => 
                           cw_from_mem_10_port, CW_OUT(9) => cw_from_mem_9_port
                           , CW_OUT(8) => cw_from_mem_8_port, CW_OUT(7) => 
                           cw_from_mem_7_port, CW_OUT(6) => cw_from_mem_6_port,
                           CW_OUT(5) => cw_from_mem_5_port, CW_OUT(4) => 
                           cw_from_mem_4_port, CW_OUT(3) => cw_from_mem_3_port,
                           CW_OUT(2) => cw_from_mem_2_port, CW_OUT(1) => 
                           cw_from_mem_1_port, CW_OUT(0) => cw_from_mem_0_port)
                           ;
   ALU_C : alu_ctrl port map( OP(0) => aluOpcode_d_4_port, OP(1) => 
                           aluOpcode_d_3_port, OP(2) => aluOpcode_d_2_port, 
                           OP(3) => aluOpcode_d_1_port, OP(4) => 
                           aluOpcode_d_0_port, ALU_WORD(12) => ALU_WORD_o(12), 
                           ALU_WORD(11) => ALU_WORD_o(11), ALU_WORD(10) => 
                           ALU_WORD_o(10), ALU_WORD(9) => ALU_WORD_o(9), 
                           ALU_WORD(8) => ALU_WORD_o(8), ALU_WORD(7) => 
                           ALU_WORD_o(7), ALU_WORD(6) => ALU_WORD_o(6), 
                           ALU_WORD(5) => ALU_WORD_o(5), ALU_WORD(4) => 
                           ALU_WORD_o(4), ALU_WORD(3) => ALU_WORD_o(3), 
                           ALU_WORD(2) => ALU_WORD_o(2), ALU_WORD(1) => 
                           ALU_WORD_o(1), ALU_WORD(0) => ALU_WORD_o(0));
   clk_gate_cw_e_reg : 
                           SNPS_CLOCK_GATE_HIGH_dlx_cu_MICROCODE_MEM_SIZE64_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE13_0 
                           port map( CLK => Clk, EN => N20, ENCLK => net3570);
   U17 : AND2_X1 port map( A1 => n124, A2 => cw_from_mem_8_port, ZN => S_EQ_NEQ
                           );
   U12 : NOR2_X1 port map( A1 => n125, A2 => S_MEM_W_R_port, ZN => S_MEM_LOAD);
   U130 : NOR4_X1 port map( A1 => IR_IN(9), A2 => IR_IN(8), A3 => IR_IN(7), A4 
                           => IR_IN(6), ZN => n114);
   U129 : NOR2_X1 port map( A1 => IR_IN(31), A2 => IR_IN(10), ZN => n115);
   U91 : NAND2_X1 port map( A1 => n46, A2 => n91, ZN => n15);
   U126 : NAND2_X1 port map( A1 => IR_IN(4), A2 => IR_IN(5), ZN => n16);
   U105 : NAND2_X1 port map( A1 => IR_IN(30), A2 => IR_IN(29), ZN => n111);
   U103 : NAND2_X1 port map( A1 => IR_IN(31), A2 => n19, ZN => n24_port);
   U89 : NAND2_X1 port map( A1 => n105, A2 => IR_IN(2), ZN => n94);
   U72 : NOR3_X1 port map( A1 => IR_IN(29), A2 => IR_IN(0), A3 => n92, ZN => 
                           n77);
   U52 : OAI211_X1 port map( C1 => n24_port, C2 => n69, A => n70, B => n71, ZN 
                           => n20_port);
   U109 : INV_X1 port map( A => IR_IN(31), ZN => n22_port);
   U115 : NAND2_X1 port map( A1 => IR_IN(0), A2 => n48, ZN => n28);
   U23 : OAI211_X1 port map( C1 => n22_port, C2 => n23_port, A => n24_port, B 
                           => n25_port, ZN => n21_port);
   U22 : AOI211_X1 port map( C1 => IR_IN(26), C2 => n19, A => n20_port, B => 
                           n21_port, ZN => n17);
   U85 : NOR2_X1 port map( A1 => n91, A2 => IR_IN(2), ZN => n47);
   U84 : NAND2_X1 port map( A1 => IR_IN(1), A2 => n47, ZN => n38);
   U32 : AOI211_X1 port map( C1 => n27_port, C2 => n38, A => n26_port, B => n16
                           , ZN => n37);
   U21 : OAI211_X1 port map( C1 => n15, C2 => n16, A => n17, B => n18, ZN => 
                           aluOpcode_d_4_port);
   U48 : NOR2_X1 port map( A1 => n60, A2 => n15, ZN => n45);
   U118 : NAND2_X1 port map( A1 => n48, A2 => n104, ZN => n62);
   U53 : NOR2_X1 port map( A1 => n27_port, A2 => n62, ZN => n67);
   U51 : AOI211_X1 port map( C1 => n46, C2 => n67, A => n68, B => n20_port, ZN 
                           => n31_port);
   U46 : AOI221_X1 port map( B1 => n62, B2 => n63, C1 => n62, C2 => n64, A => 
                           IR_IN(3), ZN => n61);
   U41 : OAI21_X1 port map( B1 => IR_IN(26), B2 => n56, A => n23_port, ZN => 
                           n34);
   U108 : NAND2_X1 port map( A1 => IR_IN(29), A2 => n22_port, ZN => n44);
   U49 : AOI221_X1 port map( B1 => IR_IN(2), B2 => n64, C1 => n60, C2 => n28, A
                           => IR_IN(1), ZN => n65);
   U125 : NOR2_X1 port map( A1 => IR_IN(0), A2 => n16, ZN => n66);
   U47 : AOI22_X1 port map( A1 => n46, A2 => n65, B1 => n66, B2 => n45, ZN => 
                           n50);
   U114 : NOR2_X1 port map( A1 => IR_IN(2), A2 => n28, ZN => n58);
   U44 : AOI22_X1 port map( A1 => n58, A2 => n59, B1 => n33, B2 => n60, ZN => 
                           n51);
   U43 : NOR2_X1 port map( A1 => n57, A2 => n41, ZN => n53);
   U39 : AOI221_X1 port map( B1 => n53, B2 => IR_IN(31), C1 => n34, C2 => 
                           n22_port, A => n54, ZN => n52);
   U95 : NOR2_X1 port map( A1 => IR_IN(30), A2 => n44, ZN => n84);
   U93 : NOR4_X1 port map( A1 => IR_IN(31), A2 => IR_IN(29), A3 => n39, A4 => 
                           n40, ZN => n99);
   U92 : AOI22_X1 port map( A1 => n95, A2 => n84, B1 => n106, B2 => n99, ZN => 
                           n89);
   U88 : NOR2_X1 port map( A1 => IR_IN(4), A2 => n94, ZN => n87);
   U87 : OAI221_X1 port map( B1 => IR_IN(0), B2 => n63, C1 => n104, C2 => 
                           IR_IN(1), A => n87, ZN => n102);
   U86 : OAI211_X1 port map( C1 => IR_IN(1), C2 => n28, A => n102, B => n103, 
                           ZN => n96);
   U81 : NAND2_X1 port map( A1 => n101, A2 => n66, ZN => n100);
   U79 : OAI22_X1 port map( A1 => IR_IN(0), A2 => n76, B1 => n100, B2 => 
                           n26_port, ZN => n97);
   U76 : AOI22_X1 port map( A1 => IR_IN(26), A2 => n83, B1 => n23_port, B2 => 
                           n69, ZN => n98);
   U75 : AOI211_X1 port map( C1 => n59, C2 => n96, A => n97, B => n98, ZN => 
                           n90);
   U70 : NAND4_X1 port map( A1 => n73, A2 => n89, A3 => n90, A4 => n71, ZN => 
                           aluOpcode_d_0_port);
   U66 : NOR2_X1 port map( A1 => n38, A2 => n64, ZN => n79);
   U65 : NOR2_X1 port map( A1 => n86, A2 => n87, ZN => n85);
   U64 : AOI221_X1 port map( B1 => IR_IN(1), B2 => n85, C1 => n63, C2 => n64, A
                           => n15, ZN => n80);
   U62 : OAI221_X1 port map( B1 => IR_IN(26), B2 => n82, C1 => n69, C2 => 
                           n23_port, A => n83, ZN => n81);
   U61 : AOI211_X1 port map( C1 => n46, C2 => n79, A => n80, B => n81, ZN => 
                           n74);
   U57 : NAND2_X1 port map( A1 => IR_IN(0), A2 => n68, ZN => n75);
   U56 : NAND4_X1 port map( A1 => n73, A2 => n74, A3 => n70, A4 => n75, ZN => 
                           aluOpcode_d_1_port);
   U5 : OR2_X1 port map( A1 => stall_exe_i, A2 => stall_fetch_o_TEMP, ZN => 
                           stall_fetch_o);
   U133 : NOR2_X1 port map( A1 => n4, A2 => stall_exe_i, ZN => N31);
   U134 : NOR2_X1 port map( A1 => n5, A2 => stall_exe_i, ZN => N30);
   U135 : NOR2_X1 port map( A1 => n2, A2 => stall_exe_i, ZN => N29);
   U97 : INV_X1 port map( A => IR_IN(26), ZN => n69);
   U120 : NOR2_X1 port map( A1 => IR_IN(4), A2 => n105, ZN => n48);
   U38 : NAND4_X1 port map( A1 => n31_port, A2 => n50, A3 => n51, A4 => n52, ZN
                           => aluOpcode_d_2_port);
   U144 : NOR2_X1 port map( A1 => stall_dec_o_TEMP, A2 => n36, ZN => n116);
   U4 : AND2_X1 port map( A1 => S_MUX_PC_BUS_1_port, A2 => S_MUX_PC_BUS_0_port,
                           ZN => was_branch_o);
   U16 : AND2_X1 port map( A1 => n4, A2 => n3, ZN => S_EXE_LOAD);
   U6 : OR2_X1 port map( A1 => stall_exe_i, A2 => stall_dec_o_TEMP, ZN => 
                           stall_dec_o);
   U113 : INV_X1 port map( A => IR_IN(3), ZN => n91);
   U121 : INV_X1 port map( A => IR_IN(5), ZN => n105);
   U123 : INV_X1 port map( A => IR_IN(1), ZN => n63);
   U74 : INV_X1 port map( A => n95, ZN => n55);
   U73 : OR4_X1 port map( A1 => n93, A2 => n94, A3 => n63, A4 => n55, ZN => n92
                           );
   U60 : INV_X1 port map( A => IR_IN(4), ZN => n78);
   U80 : INV_X1 port map( A => n46, ZN => n26_port);
   U24 : OR3_X1 port map( A1 => n26_port, A2 => n27_port, A3 => n28, ZN => 
                           n25_port);
   U31 : INV_X1 port map( A => n37, ZN => n18);
   U50 : INV_X1 port map( A => IR_IN(2), ZN => n60);
   U119 : INV_X1 port map( A => IR_IN(0), ZN => n104);
   U83 : INV_X1 port map( A => n38, ZN => n101);
   U58 : INV_X1 port map( A => n76, ZN => n68);
   U45 : AND2_X1 port map( A1 => n61, A2 => n46, ZN => n33);
   U42 : INV_X1 port map( A => n19, ZN => n56);
   U110 : INV_X1 port map( A => IR_IN(30), ZN => n40);
   U90 : INV_X1 port map( A => n15, ZN => n59);
   U102 : INV_X1 port map( A => n43, ZN => n57);
   U124 : INV_X1 port map( A => n66, ZN => n103);
   U117 : INV_X1 port map( A => n62, ZN => n86);
   U139 : AND2_X1 port map( A1 => n116, A2 => cw_from_mem_4_port, ZN => N25);
   U138 : AND2_X1 port map( A1 => n116, A2 => cw_from_mem_5_port, ZN => N26);
   U141 : AND2_X1 port map( A1 => n116, A2 => cw_from_mem_2_port, ZN => N23);
   U142 : AND2_X1 port map( A1 => n116, A2 => cw_from_mem_1_port, ZN => N22);
   U143 : AND2_X1 port map( A1 => n116, A2 => cw_from_mem_0_port, ZN => N21);
   U137 : AND2_X1 port map( A1 => n116, A2 => cw_from_mem_6_port, ZN => N27);
   U140 : AND2_X1 port map( A1 => n116, A2 => cw_from_mem_3_port, ZN => N24);
   U132 : AND2_X1 port map( A1 => N20, A2 => n3, ZN => N32);
   cw_e_reg_6_inst : DFFR_X2 port map( D => N27, CK => net3570, RN => n49, Q =>
                           S_MUX_ALUIN, QN => n35);
   U10 : AND2_X1 port map( A1 => n124, A2 => cw_from_mem_11_port, ZN => 
                           S_MUX_PC_BUS_0_port);
   U7 : OR2_X1 port map( A1 => stall_exe_i, A2 => stall_btb_o_TEMP, ZN => 
                           stall_btb_o);
   cw_e_reg_2_inst : DFFR_X1 port map( D => N23, CK => net3570, RN => n49, Q =>
                           n32_port, QN => n4);
   cw_e_reg_1_inst : DFFR_X1 port map( D => N22, CK => net3570, RN => n49, Q =>
                           n30_port, QN => n5);
   U9 : OAI21_X1 port map( B1 => n44, B2 => n1, A => n18, ZN => n8);
   U11 : OR2_X1 port map( A1 => n43, A2 => n7, ZN => n1);
   U13 : OAI221_X1 port map( B1 => n45, B2 => n46, C1 => n45, C2 => n47, A => 
                           n48, ZN => n6);
   U14 : AOI21_X1 port map( B1 => n41, B2 => n40, A => n39, ZN => n7);
   U15 : AOI211_X1 port map( C1 => IR_IN(2), C2 => n33, A => n34, B => n8, ZN 
                           => n9);
   U18 : OAI211_X1 port map( C1 => IR_IN(1), C2 => n6, A => n31_port, B => n9, 
                           ZN => aluOpcode_d_3_port);
   U19 : NAND3_X1 port map( A1 => IR_IN(3), A2 => n63, A3 => n86, ZN => n10);
   U20 : OAI211_X1 port map( C1 => n66, C2 => n58, A => IR_IN(1), B => n91, ZN 
                           => n11);
   U25 : OAI211_X1 port map( C1 => n103, C2 => n27_port, A => n10, B => n11, ZN
                           => n12);
   U26 : NOR3_X1 port map( A1 => n44, A2 => n57, A3 => n41, ZN => n13);
   U27 : OR3_X1 port map( A1 => n42, A2 => n44, A3 => n40, ZN => n14);
   U28 : AOI21_X1 port map( B1 => n24_port, B2 => n14, A => IR_IN(26), ZN => 
                           n29_port);
   U29 : AOI211_X1 port map( C1 => n46, C2 => n12, A => n13, B => n29_port, ZN 
                           => n73);
   U30 : AND2_X1 port map( A1 => cw_from_mem_12_port, A2 => n124, ZN => 
                           S_MUX_PC_BUS_1_port);
   U33 : AND2_X2 port map( A1 => n124, A2 => cw_from_mem_7_port, ZN => 
                           S_MUX_LINK);
   U34 : AND2_X2 port map( A1 => cw_from_mem_10_port, A2 => n124, ZN => S_EXT);
   U35 : INV_X1 port map( A => Rst, ZN => n49);
   U36 : INV_X1 port map( A => stall_exe_i, ZN => N20);
   U37 : INV_X1 port map( A => IR_IN(28), ZN => n39);
   U40 : CLKBUF_X1 port map( A => IR_IN(27), Z => n42);
   U54 : AND2_X1 port map( A1 => cw_from_mem_9_port, A2 => n124, ZN => 
                           S_EXT_SIGN);
   U55 : NOR4_X2 port map( A1 => IR_IN(26), A2 => IR_IN(29), A3 => IR_IN(27), 
                           A4 => n93, ZN => n46);
   U63 : AOI211_X1 port map( C1 => IR_IN(30), C2 => n55, A => IR_IN(28), B => 
                           n44, ZN => n54);
   U68 : NOR2_X1 port map( A1 => IR_IN(30), A2 => IR_IN(28), ZN => n43);
   U69 : NOR2_X1 port map( A1 => IR_IN(26), A2 => n42, ZN => n106);
   U77 : NAND2_X1 port map( A1 => n42, A2 => n84, ZN => n82);
   U78 : NAND2_X1 port map( A1 => n42, A2 => n99, ZN => n83);
   U94 : NAND2_X1 port map( A1 => IR_IN(26), A2 => n42, ZN => n41);
   U96 : NAND4_X1 port map( A1 => IR_IN(30), A2 => IR_IN(29), A3 => n42, A4 => 
                           n39, ZN => n23_port);
   U98 : NOR3_X1 port map( A1 => n42, A2 => n39, A3 => n111, ZN => n19);
   U99 : NOR2_X1 port map( A1 => IR_IN(27), A2 => n69, ZN => n95);
   n72 <= '0';
   n88 <= '0';
   n107 <= '0';
   n108 <= '0';
   n109 <= '0';
   n110 <= '0';
   n112 <= '0';
   n113 <= '0';
   n122 <= '0';
   n126 <= '0';
   n127 <= '0';
   n128 <= '0';
   n129 <= '0';

end SYN_dlx_cu_hw;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity jump_logic is

   port( NPCF_i, IR_i, A_i : in std_logic_vector (31 downto 0);  A_o : out 
         std_logic_vector (31 downto 0);  rA_o, rB_o, rC_o : out 
         std_logic_vector (4 downto 0);  branch_target_o, sum_addr_o, 
         extended_imm : out std_logic_vector (31 downto 0);  taken_o : out 
         std_logic;  FW_X_i, FW_W_i : in std_logic_vector (31 downto 0);  
         S_FW_Adec_i : in std_logic_vector (1 downto 0);  S_EXT_i, S_EXT_SIGN_i
         , S_MUX_LINK_i, S_EQ_NEQ_i : in std_logic);

end jump_logic;

architecture SYN_struct of jump_logic is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component mux41_MUX_SIZE32_0
      port( IN0, IN1, IN2, IN3 : in std_logic_vector (31 downto 0);  CTRL : in 
            std_logic_vector (1 downto 0);  OUT1 : out std_logic_vector (31 
            downto 0));
   end component;
   
   component mux21_4
      port( IN0, IN1 : in std_logic_vector (31 downto 0);  CTRL : in std_logic;
            OUT1 : out std_logic_vector (31 downto 0));
   end component;
   
   component zerocheck
      port( IN0 : in std_logic_vector (31 downto 0);  CTRL : in std_logic;  
            OUT1 : out std_logic);
   end component;
   
   component mux21_0
      port( IN0, IN1 : in std_logic_vector (31 downto 0);  CTRL : in std_logic;
            OUT1 : out std_logic_vector (31 downto 0));
   end component;
   
   component p4add_N32_logN5_0
      port( A, B : in std_logic_vector (31 downto 0);  Cin, sign : in std_logic
            ;  S : out std_logic_vector (31 downto 0);  Cout : out std_logic);
   end component;
   
   component extender_32
      port( IN1 : in std_logic_vector (31 downto 0);  CTRL, SIGN : in std_logic
            ;  OUT1 : out std_logic_vector (31 downto 0));
   end component;
   
   signal X_Logic0_port, A_o_31_port, A_o_30_port, A_o_29_port, A_o_28_port, 
      A_o_27_port, A_o_26_port, A_o_25_port, A_o_24_port, A_o_23_port, 
      A_o_22_port, A_o_21_port, A_o_20_port, A_o_19_port, A_o_18_port, 
      A_o_17_port, A_o_16_port, A_o_15_port, A_o_14_port, A_o_13_port, 
      A_o_12_port, A_o_11_port, A_o_10_port, A_o_9_port, A_o_8_port, A_o_7_port
      , A_o_6_port, A_o_5_port, A_o_4_port, A_o_3_port, A_o_2_port, A_o_1_port,
      A_o_0_port, sum_addr_o_31_port, sum_addr_o_30_port, sum_addr_o_29_port, 
      sum_addr_o_28_port, sum_addr_o_27_port, sum_addr_o_26_port, 
      sum_addr_o_25_port, sum_addr_o_24_port, sum_addr_o_23_port, 
      sum_addr_o_22_port, sum_addr_o_21_port, sum_addr_o_20_port, 
      sum_addr_o_19_port, sum_addr_o_18_port, sum_addr_o_17_port, 
      sum_addr_o_16_port, sum_addr_o_15_port, sum_addr_o_14_port, 
      sum_addr_o_13_port, sum_addr_o_12_port, sum_addr_o_11_port, 
      sum_addr_o_10_port, sum_addr_o_9_port, sum_addr_o_8_port, 
      sum_addr_o_7_port, sum_addr_o_6_port, sum_addr_o_5_port, 
      sum_addr_o_4_port, sum_addr_o_3_port, sum_addr_o_2_port, 
      sum_addr_o_1_port, sum_addr_o_0_port, ext_imm_31_port, ext_imm_30_port, 
      ext_imm_29_port, ext_imm_28_port, ext_imm_27_port, ext_imm_26_port, 
      ext_imm_25_port, ext_imm_24_port, ext_imm_23_port, ext_imm_22_port, 
      ext_imm_21_port, ext_imm_20_port, ext_imm_19_port, ext_imm_18_port, 
      ext_imm_17_port, ext_imm_16_port, ext_imm_15_port, ext_imm_14_port, 
      ext_imm_13_port, ext_imm_12_port, ext_imm_11_port, ext_imm_10_port, 
      ext_imm_9_port, ext_imm_8_port, ext_imm_7_port, ext_imm_6_port, 
      ext_imm_5_port, ext_imm_4_port, ext_imm_3_port, ext_imm_2_port, 
      ext_imm_1_port, ext_imm_0_port, branch_sel, n1, n4, n5, n6, n7, n8, n9, 
      net47683 : std_logic;

begin
   A_o <= ( A_o_31_port, A_o_30_port, A_o_29_port, A_o_28_port, A_o_27_port, 
      A_o_26_port, A_o_25_port, A_o_24_port, A_o_23_port, A_o_22_port, 
      A_o_21_port, A_o_20_port, A_o_19_port, A_o_18_port, A_o_17_port, 
      A_o_16_port, A_o_15_port, A_o_14_port, A_o_13_port, A_o_12_port, 
      A_o_11_port, A_o_10_port, A_o_9_port, A_o_8_port, A_o_7_port, A_o_6_port,
      A_o_5_port, A_o_4_port, A_o_3_port, A_o_2_port, A_o_1_port, A_o_0_port );
   rA_o <= ( IR_i(25), IR_i(24), IR_i(23), IR_i(22), IR_i(21) );
   rB_o <= ( IR_i(20), IR_i(19), IR_i(18), IR_i(17), IR_i(16) );
   rC_o <= ( IR_i(15), IR_i(14), IR_i(13), IR_i(12), IR_i(11) );
   sum_addr_o <= ( sum_addr_o_31_port, sum_addr_o_30_port, sum_addr_o_29_port, 
      sum_addr_o_28_port, sum_addr_o_27_port, sum_addr_o_26_port, 
      sum_addr_o_25_port, sum_addr_o_24_port, sum_addr_o_23_port, 
      sum_addr_o_22_port, sum_addr_o_21_port, sum_addr_o_20_port, 
      sum_addr_o_19_port, sum_addr_o_18_port, sum_addr_o_17_port, 
      sum_addr_o_16_port, sum_addr_o_15_port, sum_addr_o_14_port, 
      sum_addr_o_13_port, sum_addr_o_12_port, sum_addr_o_11_port, 
      sum_addr_o_10_port, sum_addr_o_9_port, sum_addr_o_8_port, 
      sum_addr_o_7_port, sum_addr_o_6_port, sum_addr_o_5_port, 
      sum_addr_o_4_port, sum_addr_o_3_port, sum_addr_o_2_port, 
      sum_addr_o_1_port, sum_addr_o_0_port );
   
   X_Logic0_port <= '0';
   EXTENDER : extender_32 port map( IN1(31) => n4, IN1(30) => n5, IN1(29) => n6
                           , IN1(28) => n7, IN1(27) => n8, IN1(26) => n9, 
                           IN1(25) => IR_i(25), IN1(24) => IR_i(24), IN1(23) =>
                           IR_i(23), IN1(22) => IR_i(22), IN1(21) => IR_i(21), 
                           IN1(20) => IR_i(20), IN1(19) => IR_i(19), IN1(18) =>
                           IR_i(18), IN1(17) => IR_i(17), IN1(16) => IR_i(16), 
                           IN1(15) => IR_i(15), IN1(14) => IR_i(14), IN1(13) =>
                           IR_i(13), IN1(12) => IR_i(12), IN1(11) => IR_i(11), 
                           IN1(10) => IR_i(10), IN1(9) => IR_i(9), IN1(8) => 
                           IR_i(8), IN1(7) => IR_i(7), IN1(6) => IR_i(6), 
                           IN1(5) => IR_i(5), IN1(4) => IR_i(4), IN1(3) => 
                           IR_i(3), IN1(2) => IR_i(2), IN1(1) => IR_i(1), 
                           IN1(0) => IR_i(0), CTRL => S_EXT_i, SIGN => 
                           S_EXT_SIGN_i, OUT1(31) => ext_imm_31_port, OUT1(30) 
                           => ext_imm_30_port, OUT1(29) => ext_imm_29_port, 
                           OUT1(28) => ext_imm_28_port, OUT1(27) => 
                           ext_imm_27_port, OUT1(26) => ext_imm_26_port, 
                           OUT1(25) => ext_imm_25_port, OUT1(24) => 
                           ext_imm_24_port, OUT1(23) => ext_imm_23_port, 
                           OUT1(22) => ext_imm_22_port, OUT1(21) => 
                           ext_imm_21_port, OUT1(20) => ext_imm_20_port, 
                           OUT1(19) => ext_imm_19_port, OUT1(18) => 
                           ext_imm_18_port, OUT1(17) => ext_imm_17_port, 
                           OUT1(16) => ext_imm_16_port, OUT1(15) => 
                           ext_imm_15_port, OUT1(14) => ext_imm_14_port, 
                           OUT1(13) => ext_imm_13_port, OUT1(12) => 
                           ext_imm_12_port, OUT1(11) => ext_imm_11_port, 
                           OUT1(10) => ext_imm_10_port, OUT1(9) => 
                           ext_imm_9_port, OUT1(8) => ext_imm_8_port, OUT1(7) 
                           => ext_imm_7_port, OUT1(6) => ext_imm_6_port, 
                           OUT1(5) => ext_imm_5_port, OUT1(4) => ext_imm_4_port
                           , OUT1(3) => ext_imm_3_port, OUT1(2) => 
                           ext_imm_2_port, OUT1(1) => ext_imm_1_port, OUT1(0) 
                           => ext_imm_0_port);
   JUMPADDER : p4add_N32_logN5_0 port map( A(31) => NPCF_i(31), A(30) => 
                           NPCF_i(30), A(29) => NPCF_i(29), A(28) => NPCF_i(28)
                           , A(27) => NPCF_i(27), A(26) => NPCF_i(26), A(25) =>
                           NPCF_i(25), A(24) => NPCF_i(24), A(23) => NPCF_i(23)
                           , A(22) => NPCF_i(22), A(21) => NPCF_i(21), A(20) =>
                           NPCF_i(20), A(19) => NPCF_i(19), A(18) => NPCF_i(18)
                           , A(17) => NPCF_i(17), A(16) => NPCF_i(16), A(15) =>
                           NPCF_i(15), A(14) => NPCF_i(14), A(13) => NPCF_i(13)
                           , A(12) => NPCF_i(12), A(11) => NPCF_i(11), A(10) =>
                           NPCF_i(10), A(9) => NPCF_i(9), A(8) => NPCF_i(8), 
                           A(7) => NPCF_i(7), A(6) => NPCF_i(6), A(5) => 
                           NPCF_i(5), A(4) => NPCF_i(4), A(3) => NPCF_i(3), 
                           A(2) => NPCF_i(2), A(1) => NPCF_i(1), A(0) => 
                           NPCF_i(0), B(31) => ext_imm_31_port, B(30) => 
                           ext_imm_30_port, B(29) => ext_imm_29_port, B(28) => 
                           ext_imm_28_port, B(27) => ext_imm_27_port, B(26) => 
                           ext_imm_26_port, B(25) => ext_imm_25_port, B(24) => 
                           ext_imm_24_port, B(23) => ext_imm_23_port, B(22) => 
                           ext_imm_22_port, B(21) => ext_imm_21_port, B(20) => 
                           ext_imm_20_port, B(19) => ext_imm_19_port, B(18) => 
                           ext_imm_18_port, B(17) => ext_imm_17_port, B(16) => 
                           ext_imm_16_port, B(15) => ext_imm_15_port, B(14) => 
                           ext_imm_14_port, B(13) => ext_imm_13_port, B(12) => 
                           ext_imm_12_port, B(11) => ext_imm_11_port, B(10) => 
                           ext_imm_10_port, B(9) => ext_imm_9_port, B(8) => 
                           ext_imm_8_port, B(7) => ext_imm_7_port, B(6) => 
                           ext_imm_6_port, B(5) => ext_imm_5_port, B(4) => 
                           ext_imm_4_port, B(3) => ext_imm_3_port, B(2) => 
                           ext_imm_2_port, B(1) => ext_imm_1_port, B(0) => 
                           ext_imm_0_port, Cin => X_Logic0_port, sign => 
                           X_Logic0_port, S(31) => sum_addr_o_31_port, S(30) =>
                           sum_addr_o_30_port, S(29) => sum_addr_o_29_port, 
                           S(28) => sum_addr_o_28_port, S(27) => 
                           sum_addr_o_27_port, S(26) => sum_addr_o_26_port, 
                           S(25) => sum_addr_o_25_port, S(24) => 
                           sum_addr_o_24_port, S(23) => sum_addr_o_23_port, 
                           S(22) => sum_addr_o_22_port, S(21) => 
                           sum_addr_o_21_port, S(20) => sum_addr_o_20_port, 
                           S(19) => sum_addr_o_19_port, S(18) => 
                           sum_addr_o_18_port, S(17) => sum_addr_o_17_port, 
                           S(16) => sum_addr_o_16_port, S(15) => 
                           sum_addr_o_15_port, S(14) => sum_addr_o_14_port, 
                           S(13) => sum_addr_o_13_port, S(12) => 
                           sum_addr_o_12_port, S(11) => sum_addr_o_11_port, 
                           S(10) => sum_addr_o_10_port, S(9) => 
                           sum_addr_o_9_port, S(8) => sum_addr_o_8_port, S(7) 
                           => sum_addr_o_7_port, S(6) => sum_addr_o_6_port, 
                           S(5) => sum_addr_o_5_port, S(4) => sum_addr_o_4_port
                           , S(3) => sum_addr_o_3_port, S(2) => 
                           sum_addr_o_2_port, S(1) => sum_addr_o_1_port, S(0) 
                           => sum_addr_o_0_port, Cout => net47683);
   BRANCHMUX : mux21_0 port map( IN0(31) => sum_addr_o_31_port, IN0(30) => 
                           sum_addr_o_30_port, IN0(29) => sum_addr_o_29_port, 
                           IN0(28) => sum_addr_o_28_port, IN0(27) => 
                           sum_addr_o_27_port, IN0(26) => sum_addr_o_26_port, 
                           IN0(25) => sum_addr_o_25_port, IN0(24) => 
                           sum_addr_o_24_port, IN0(23) => sum_addr_o_23_port, 
                           IN0(22) => sum_addr_o_22_port, IN0(21) => 
                           sum_addr_o_21_port, IN0(20) => sum_addr_o_20_port, 
                           IN0(19) => sum_addr_o_19_port, IN0(18) => 
                           sum_addr_o_18_port, IN0(17) => sum_addr_o_17_port, 
                           IN0(16) => sum_addr_o_16_port, IN0(15) => 
                           sum_addr_o_15_port, IN0(14) => sum_addr_o_14_port, 
                           IN0(13) => sum_addr_o_13_port, IN0(12) => 
                           sum_addr_o_12_port, IN0(11) => sum_addr_o_11_port, 
                           IN0(10) => sum_addr_o_10_port, IN0(9) => 
                           sum_addr_o_9_port, IN0(8) => sum_addr_o_8_port, 
                           IN0(7) => sum_addr_o_7_port, IN0(6) => 
                           sum_addr_o_6_port, IN0(5) => sum_addr_o_5_port, 
                           IN0(4) => sum_addr_o_4_port, IN0(3) => 
                           sum_addr_o_3_port, IN0(2) => sum_addr_o_2_port, 
                           IN0(1) => sum_addr_o_1_port, IN0(0) => 
                           sum_addr_o_0_port, IN1(31) => NPCF_i(31), IN1(30) =>
                           NPCF_i(30), IN1(29) => NPCF_i(29), IN1(28) => 
                           NPCF_i(28), IN1(27) => NPCF_i(27), IN1(26) => 
                           NPCF_i(26), IN1(25) => NPCF_i(25), IN1(24) => 
                           NPCF_i(24), IN1(23) => NPCF_i(23), IN1(22) => 
                           NPCF_i(22), IN1(21) => NPCF_i(21), IN1(20) => 
                           NPCF_i(20), IN1(19) => NPCF_i(19), IN1(18) => 
                           NPCF_i(18), IN1(17) => NPCF_i(17), IN1(16) => 
                           NPCF_i(16), IN1(15) => NPCF_i(15), IN1(14) => 
                           NPCF_i(14), IN1(13) => NPCF_i(13), IN1(12) => 
                           NPCF_i(12), IN1(11) => NPCF_i(11), IN1(10) => 
                           NPCF_i(10), IN1(9) => NPCF_i(9), IN1(8) => NPCF_i(8)
                           , IN1(7) => NPCF_i(7), IN1(6) => NPCF_i(6), IN1(5) 
                           => NPCF_i(5), IN1(4) => NPCF_i(4), IN1(3) => 
                           NPCF_i(3), IN1(2) => NPCF_i(2), IN1(1) => NPCF_i(1),
                           IN1(0) => NPCF_i(0), CTRL => branch_sel, OUT1(31) =>
                           branch_target_o(31), OUT1(30) => branch_target_o(30)
                           , OUT1(29) => branch_target_o(29), OUT1(28) => 
                           branch_target_o(28), OUT1(27) => branch_target_o(27)
                           , OUT1(26) => branch_target_o(26), OUT1(25) => 
                           branch_target_o(25), OUT1(24) => branch_target_o(24)
                           , OUT1(23) => branch_target_o(23), OUT1(22) => 
                           branch_target_o(22), OUT1(21) => branch_target_o(21)
                           , OUT1(20) => branch_target_o(20), OUT1(19) => 
                           branch_target_o(19), OUT1(18) => branch_target_o(18)
                           , OUT1(17) => branch_target_o(17), OUT1(16) => 
                           branch_target_o(16), OUT1(15) => branch_target_o(15)
                           , OUT1(14) => branch_target_o(14), OUT1(13) => 
                           branch_target_o(13), OUT1(12) => branch_target_o(12)
                           , OUT1(11) => branch_target_o(11), OUT1(10) => 
                           branch_target_o(10), OUT1(9) => branch_target_o(9), 
                           OUT1(8) => branch_target_o(8), OUT1(7) => 
                           branch_target_o(7), OUT1(6) => branch_target_o(6), 
                           OUT1(5) => branch_target_o(5), OUT1(4) => 
                           branch_target_o(4), OUT1(3) => branch_target_o(3), 
                           OUT1(2) => branch_target_o(2), OUT1(1) => 
                           branch_target_o(1), OUT1(0) => branch_target_o(0));
   ZC : zerocheck port map( IN0(31) => A_o_31_port, IN0(30) => A_o_30_port, 
                           IN0(29) => A_o_29_port, IN0(28) => A_o_28_port, 
                           IN0(27) => A_o_27_port, IN0(26) => A_o_26_port, 
                           IN0(25) => A_o_25_port, IN0(24) => A_o_24_port, 
                           IN0(23) => A_o_23_port, IN0(22) => A_o_22_port, 
                           IN0(21) => A_o_21_port, IN0(20) => A_o_20_port, 
                           IN0(19) => A_o_19_port, IN0(18) => A_o_18_port, 
                           IN0(17) => A_o_17_port, IN0(16) => A_o_16_port, 
                           IN0(15) => A_o_15_port, IN0(14) => A_o_14_port, 
                           IN0(13) => A_o_13_port, IN0(12) => A_o_12_port, 
                           IN0(11) => A_o_11_port, IN0(10) => A_o_10_port, 
                           IN0(9) => A_o_9_port, IN0(8) => A_o_8_port, IN0(7) 
                           => A_o_7_port, IN0(6) => A_o_6_port, IN0(5) => 
                           A_o_5_port, IN0(4) => A_o_4_port, IN0(3) => 
                           A_o_3_port, IN0(2) => A_o_2_port, IN0(1) => 
                           A_o_1_port, IN0(0) => A_o_0_port, CTRL => S_EQ_NEQ_i
                           , OUT1 => branch_sel);
   MUXLINK : mux21_4 port map( IN0(31) => ext_imm_31_port, IN0(30) => 
                           ext_imm_30_port, IN0(29) => ext_imm_29_port, IN0(28)
                           => ext_imm_28_port, IN0(27) => ext_imm_27_port, 
                           IN0(26) => ext_imm_26_port, IN0(25) => 
                           ext_imm_25_port, IN0(24) => ext_imm_24_port, IN0(23)
                           => ext_imm_23_port, IN0(22) => ext_imm_22_port, 
                           IN0(21) => ext_imm_21_port, IN0(20) => 
                           ext_imm_20_port, IN0(19) => ext_imm_19_port, IN0(18)
                           => ext_imm_18_port, IN0(17) => ext_imm_17_port, 
                           IN0(16) => ext_imm_16_port, IN0(15) => 
                           ext_imm_15_port, IN0(14) => ext_imm_14_port, IN0(13)
                           => ext_imm_13_port, IN0(12) => ext_imm_12_port, 
                           IN0(11) => ext_imm_11_port, IN0(10) => 
                           ext_imm_10_port, IN0(9) => ext_imm_9_port, IN0(8) =>
                           ext_imm_8_port, IN0(7) => ext_imm_7_port, IN0(6) => 
                           ext_imm_6_port, IN0(5) => ext_imm_5_port, IN0(4) => 
                           ext_imm_4_port, IN0(3) => ext_imm_3_port, IN0(2) => 
                           ext_imm_2_port, IN0(1) => ext_imm_1_port, IN0(0) => 
                           ext_imm_0_port, IN1(31) => NPCF_i(31), IN1(30) => 
                           NPCF_i(30), IN1(29) => NPCF_i(29), IN1(28) => 
                           NPCF_i(28), IN1(27) => NPCF_i(27), IN1(26) => 
                           NPCF_i(26), IN1(25) => NPCF_i(25), IN1(24) => 
                           NPCF_i(24), IN1(23) => NPCF_i(23), IN1(22) => 
                           NPCF_i(22), IN1(21) => NPCF_i(21), IN1(20) => 
                           NPCF_i(20), IN1(19) => NPCF_i(19), IN1(18) => 
                           NPCF_i(18), IN1(17) => NPCF_i(17), IN1(16) => 
                           NPCF_i(16), IN1(15) => NPCF_i(15), IN1(14) => 
                           NPCF_i(14), IN1(13) => NPCF_i(13), IN1(12) => 
                           NPCF_i(12), IN1(11) => NPCF_i(11), IN1(10) => 
                           NPCF_i(10), IN1(9) => NPCF_i(9), IN1(8) => NPCF_i(8)
                           , IN1(7) => NPCF_i(7), IN1(6) => NPCF_i(6), IN1(5) 
                           => NPCF_i(5), IN1(4) => NPCF_i(4), IN1(3) => 
                           NPCF_i(3), IN1(2) => NPCF_i(2), IN1(1) => NPCF_i(1),
                           IN1(0) => NPCF_i(0), CTRL => S_MUX_LINK_i, OUT1(31) 
                           => extended_imm(31), OUT1(30) => extended_imm(30), 
                           OUT1(29) => extended_imm(29), OUT1(28) => 
                           extended_imm(28), OUT1(27) => extended_imm(27), 
                           OUT1(26) => extended_imm(26), OUT1(25) => 
                           extended_imm(25), OUT1(24) => extended_imm(24), 
                           OUT1(23) => extended_imm(23), OUT1(22) => 
                           extended_imm(22), OUT1(21) => extended_imm(21), 
                           OUT1(20) => extended_imm(20), OUT1(19) => 
                           extended_imm(19), OUT1(18) => extended_imm(18), 
                           OUT1(17) => extended_imm(17), OUT1(16) => 
                           extended_imm(16), OUT1(15) => extended_imm(15), 
                           OUT1(14) => extended_imm(14), OUT1(13) => 
                           extended_imm(13), OUT1(12) => extended_imm(12), 
                           OUT1(11) => extended_imm(11), OUT1(10) => 
                           extended_imm(10), OUT1(9) => extended_imm(9), 
                           OUT1(8) => extended_imm(8), OUT1(7) => 
                           extended_imm(7), OUT1(6) => extended_imm(6), OUT1(5)
                           => extended_imm(5), OUT1(4) => extended_imm(4), 
                           OUT1(3) => extended_imm(3), OUT1(2) => 
                           extended_imm(2), OUT1(1) => extended_imm(1), OUT1(0)
                           => extended_imm(0));
   MUX_FWA : mux41_MUX_SIZE32_0 port map( IN0(31) => A_i(31), IN0(30) => 
                           A_i(30), IN0(29) => A_i(29), IN0(28) => A_i(28), 
                           IN0(27) => A_i(27), IN0(26) => A_i(26), IN0(25) => 
                           A_i(25), IN0(24) => A_i(24), IN0(23) => A_i(23), 
                           IN0(22) => A_i(22), IN0(21) => A_i(21), IN0(20) => 
                           A_i(20), IN0(19) => A_i(19), IN0(18) => A_i(18), 
                           IN0(17) => A_i(17), IN0(16) => A_i(16), IN0(15) => 
                           A_i(15), IN0(14) => A_i(14), IN0(13) => A_i(13), 
                           IN0(12) => A_i(12), IN0(11) => A_i(11), IN0(10) => 
                           A_i(10), IN0(9) => A_i(9), IN0(8) => A_i(8), IN0(7) 
                           => A_i(7), IN0(6) => A_i(6), IN0(5) => A_i(5), 
                           IN0(4) => A_i(4), IN0(3) => A_i(3), IN0(2) => A_i(2)
                           , IN0(1) => A_i(1), IN0(0) => A_i(0), IN1(31) => 
                           FW_X_i(31), IN1(30) => FW_X_i(30), IN1(29) => 
                           FW_X_i(29), IN1(28) => FW_X_i(28), IN1(27) => 
                           FW_X_i(27), IN1(26) => FW_X_i(26), IN1(25) => 
                           FW_X_i(25), IN1(24) => FW_X_i(24), IN1(23) => 
                           FW_X_i(23), IN1(22) => FW_X_i(22), IN1(21) => 
                           FW_X_i(21), IN1(20) => FW_X_i(20), IN1(19) => 
                           FW_X_i(19), IN1(18) => FW_X_i(18), IN1(17) => 
                           FW_X_i(17), IN1(16) => FW_X_i(16), IN1(15) => 
                           FW_X_i(15), IN1(14) => FW_X_i(14), IN1(13) => 
                           FW_X_i(13), IN1(12) => FW_X_i(12), IN1(11) => 
                           FW_X_i(11), IN1(10) => FW_X_i(10), IN1(9) => 
                           FW_X_i(9), IN1(8) => FW_X_i(8), IN1(7) => FW_X_i(7),
                           IN1(6) => FW_X_i(6), IN1(5) => FW_X_i(5), IN1(4) => 
                           FW_X_i(4), IN1(3) => FW_X_i(3), IN1(2) => FW_X_i(2),
                           IN1(1) => FW_X_i(1), IN1(0) => FW_X_i(0), IN2(31) =>
                           FW_W_i(31), IN2(30) => FW_W_i(30), IN2(29) => 
                           FW_W_i(29), IN2(28) => FW_W_i(28), IN2(27) => 
                           FW_W_i(27), IN2(26) => FW_W_i(26), IN2(25) => 
                           FW_W_i(25), IN2(24) => FW_W_i(24), IN2(23) => 
                           FW_W_i(23), IN2(22) => FW_W_i(22), IN2(21) => 
                           FW_W_i(21), IN2(20) => FW_W_i(20), IN2(19) => 
                           FW_W_i(19), IN2(18) => FW_W_i(18), IN2(17) => 
                           FW_W_i(17), IN2(16) => FW_W_i(16), IN2(15) => 
                           FW_W_i(15), IN2(14) => FW_W_i(14), IN2(13) => 
                           FW_W_i(13), IN2(12) => FW_W_i(12), IN2(11) => 
                           FW_W_i(11), IN2(10) => FW_W_i(10), IN2(9) => 
                           FW_W_i(9), IN2(8) => FW_W_i(8), IN2(7) => FW_W_i(7),
                           IN2(6) => FW_W_i(6), IN2(5) => FW_W_i(5), IN2(4) => 
                           FW_W_i(4), IN2(3) => FW_W_i(3), IN2(2) => FW_W_i(2),
                           IN2(1) => FW_W_i(1), IN2(0) => FW_W_i(0), IN3(31) =>
                           X_Logic0_port, IN3(30) => X_Logic0_port, IN3(29) => 
                           X_Logic0_port, IN3(28) => X_Logic0_port, IN3(27) => 
                           X_Logic0_port, IN3(26) => X_Logic0_port, IN3(25) => 
                           X_Logic0_port, IN3(24) => X_Logic0_port, IN3(23) => 
                           X_Logic0_port, IN3(22) => X_Logic0_port, IN3(21) => 
                           X_Logic0_port, IN3(20) => X_Logic0_port, IN3(19) => 
                           X_Logic0_port, IN3(18) => X_Logic0_port, IN3(17) => 
                           X_Logic0_port, IN3(16) => X_Logic0_port, IN3(15) => 
                           X_Logic0_port, IN3(14) => X_Logic0_port, IN3(13) => 
                           X_Logic0_port, IN3(12) => X_Logic0_port, IN3(11) => 
                           X_Logic0_port, IN3(10) => X_Logic0_port, IN3(9) => 
                           X_Logic0_port, IN3(8) => X_Logic0_port, IN3(7) => 
                           X_Logic0_port, IN3(6) => X_Logic0_port, IN3(5) => 
                           X_Logic0_port, IN3(4) => X_Logic0_port, IN3(3) => 
                           X_Logic0_port, IN3(2) => X_Logic0_port, IN3(1) => 
                           X_Logic0_port, IN3(0) => X_Logic0_port, CTRL(1) => 
                           S_FW_Adec_i(1), CTRL(0) => S_FW_Adec_i(0), OUT1(31) 
                           => A_o_31_port, OUT1(30) => A_o_30_port, OUT1(29) =>
                           A_o_29_port, OUT1(28) => A_o_28_port, OUT1(27) => 
                           A_o_27_port, OUT1(26) => A_o_26_port, OUT1(25) => 
                           A_o_25_port, OUT1(24) => A_o_24_port, OUT1(23) => 
                           A_o_23_port, OUT1(22) => A_o_22_port, OUT1(21) => 
                           A_o_21_port, OUT1(20) => A_o_20_port, OUT1(19) => 
                           A_o_19_port, OUT1(18) => A_o_18_port, OUT1(17) => 
                           A_o_17_port, OUT1(16) => A_o_16_port, OUT1(15) => 
                           A_o_15_port, OUT1(14) => A_o_14_port, OUT1(13) => 
                           A_o_13_port, OUT1(12) => A_o_12_port, OUT1(11) => 
                           A_o_11_port, OUT1(10) => A_o_10_port, OUT1(9) => 
                           A_o_9_port, OUT1(8) => A_o_8_port, OUT1(7) => 
                           A_o_7_port, OUT1(6) => A_o_6_port, OUT1(5) => 
                           A_o_5_port, OUT1(4) => A_o_4_port, OUT1(3) => 
                           A_o_3_port, OUT1(2) => A_o_2_port, OUT1(1) => 
                           A_o_1_port, OUT1(0) => A_o_0_port);
   U2 : CLKBUF_X1 port map( A => branch_sel, Z => n1);
   U3 : INV_X1 port map( A => n1, ZN => taken_o);
   n4 <= '0';
   n5 <= '0';
   n6 <= '0';
   n7 <= '0';
   n8 <= '0';
   n9 <= '0';

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity fetch_regs is

   port( NPCF_i, IR_i : in std_logic_vector (31 downto 0);  NPCF_o, IR_o : out 
         std_logic_vector (31 downto 0);  stall_i, clk, rst : in std_logic);

end fetch_regs;

architecture SYN_struct of fetch_regs is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component ff32_en_IR
      port( D : in std_logic_vector (31 downto 0);  en, clk, rst : in std_logic
            ;  Q : out std_logic_vector (31 downto 0));
   end component;
   
   component ff32_en_1
      port( D : in std_logic_vector (31 downto 0);  en, clk, rst : in std_logic
            ;  Q : out std_logic_vector (31 downto 0));
   end component;
   
   signal enable : std_logic;

begin
   
   NPCF : ff32_en_1 port map( D(31) => NPCF_i(31), D(30) => NPCF_i(30), D(29) 
                           => NPCF_i(29), D(28) => NPCF_i(28), D(27) => 
                           NPCF_i(27), D(26) => NPCF_i(26), D(25) => NPCF_i(25)
                           , D(24) => NPCF_i(24), D(23) => NPCF_i(23), D(22) =>
                           NPCF_i(22), D(21) => NPCF_i(21), D(20) => NPCF_i(20)
                           , D(19) => NPCF_i(19), D(18) => NPCF_i(18), D(17) =>
                           NPCF_i(17), D(16) => NPCF_i(16), D(15) => NPCF_i(15)
                           , D(14) => NPCF_i(14), D(13) => NPCF_i(13), D(12) =>
                           NPCF_i(12), D(11) => NPCF_i(11), D(10) => NPCF_i(10)
                           , D(9) => NPCF_i(9), D(8) => NPCF_i(8), D(7) => 
                           NPCF_i(7), D(6) => NPCF_i(6), D(5) => NPCF_i(5), 
                           D(4) => NPCF_i(4), D(3) => NPCF_i(3), D(2) => 
                           NPCF_i(2), D(1) => NPCF_i(1), D(0) => NPCF_i(0), en 
                           => enable, clk => clk, rst => rst, Q(31) => 
                           NPCF_o(31), Q(30) => NPCF_o(30), Q(29) => NPCF_o(29)
                           , Q(28) => NPCF_o(28), Q(27) => NPCF_o(27), Q(26) =>
                           NPCF_o(26), Q(25) => NPCF_o(25), Q(24) => NPCF_o(24)
                           , Q(23) => NPCF_o(23), Q(22) => NPCF_o(22), Q(21) =>
                           NPCF_o(21), Q(20) => NPCF_o(20), Q(19) => NPCF_o(19)
                           , Q(18) => NPCF_o(18), Q(17) => NPCF_o(17), Q(16) =>
                           NPCF_o(16), Q(15) => NPCF_o(15), Q(14) => NPCF_o(14)
                           , Q(13) => NPCF_o(13), Q(12) => NPCF_o(12), Q(11) =>
                           NPCF_o(11), Q(10) => NPCF_o(10), Q(9) => NPCF_o(9), 
                           Q(8) => NPCF_o(8), Q(7) => NPCF_o(7), Q(6) => 
                           NPCF_o(6), Q(5) => NPCF_o(5), Q(4) => NPCF_o(4), 
                           Q(3) => NPCF_o(3), Q(2) => NPCF_o(2), Q(1) => 
                           NPCF_o(1), Q(0) => NPCF_o(0));
   IR : ff32_en_IR port map( D(31) => IR_i(31), D(30) => IR_i(30), D(29) => 
                           IR_i(29), D(28) => IR_i(28), D(27) => IR_i(27), 
                           D(26) => IR_i(26), D(25) => IR_i(25), D(24) => 
                           IR_i(24), D(23) => IR_i(23), D(22) => IR_i(22), 
                           D(21) => IR_i(21), D(20) => IR_i(20), D(19) => 
                           IR_i(19), D(18) => IR_i(18), D(17) => IR_i(17), 
                           D(16) => IR_i(16), D(15) => IR_i(15), D(14) => 
                           IR_i(14), D(13) => IR_i(13), D(12) => IR_i(12), 
                           D(11) => IR_i(11), D(10) => IR_i(10), D(9) => 
                           IR_i(9), D(8) => IR_i(8), D(7) => IR_i(7), D(6) => 
                           IR_i(6), D(5) => IR_i(5), D(4) => IR_i(4), D(3) => 
                           IR_i(3), D(2) => IR_i(2), D(1) => IR_i(1), D(0) => 
                           IR_i(0), en => enable, clk => clk, rst => rst, Q(31)
                           => IR_o(31), Q(30) => IR_o(30), Q(29) => IR_o(29), 
                           Q(28) => IR_o(28), Q(27) => IR_o(27), Q(26) => 
                           IR_o(26), Q(25) => IR_o(25), Q(24) => IR_o(24), 
                           Q(23) => IR_o(23), Q(22) => IR_o(22), Q(21) => 
                           IR_o(21), Q(20) => IR_o(20), Q(19) => IR_o(19), 
                           Q(18) => IR_o(18), Q(17) => IR_o(17), Q(16) => 
                           IR_o(16), Q(15) => IR_o(15), Q(14) => IR_o(14), 
                           Q(13) => IR_o(13), Q(12) => IR_o(12), Q(11) => 
                           IR_o(11), Q(10) => IR_o(10), Q(9) => IR_o(9), Q(8) 
                           => IR_o(8), Q(7) => IR_o(7), Q(6) => IR_o(6), Q(5) 
                           => IR_o(5), Q(4) => IR_o(4), Q(3) => IR_o(3), Q(2) 
                           => IR_o(2), Q(1) => IR_o(1), Q(0) => IR_o(0));
   U1 : INV_X1 port map( A => stall_i, ZN => enable);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity btb_N_LINES4_SIZE32 is

   port( clock, reset, stall_i : in std_logic;  TAG_i : in std_logic_vector (3 
         downto 0);  target_PC_i : in std_logic_vector (31 downto 0);  
         was_taken_i : in std_logic;  predicted_next_PC_o : out 
         std_logic_vector (31 downto 0);  taken_o, mispredict_o : out std_logic
         );

end btb_N_LINES4_SIZE32;

architecture SYN_bhe of btb_N_LINES4_SIZE32 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND4_X2
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X2
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_1
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_2
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_3
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_4
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_5
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_6
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_7
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_8
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_9
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_10
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_11
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_12
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_13
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_14
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_15
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_16
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_0
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component predictor_2_1
      port( clock, reset, enable, taken_i : in std_logic;  prediction_o : out 
            std_logic);
   end component;
   
   component predictor_2_2
      port( clock, reset, enable, taken_i : in std_logic;  prediction_o : out 
            std_logic);
   end component;
   
   component predictor_2_3
      port( clock, reset, enable, taken_i : in std_logic;  prediction_o : out 
            std_logic);
   end component;
   
   component predictor_2_4
      port( clock, reset, enable, taken_i : in std_logic;  prediction_o : out 
            std_logic);
   end component;
   
   component predictor_2_5
      port( clock, reset, enable, taken_i : in std_logic;  prediction_o : out 
            std_logic);
   end component;
   
   component predictor_2_6
      port( clock, reset, enable, taken_i : in std_logic;  prediction_o : out 
            std_logic);
   end component;
   
   component predictor_2_7
      port( clock, reset, enable, taken_i : in std_logic;  prediction_o : out 
            std_logic);
   end component;
   
   component predictor_2_8
      port( clock, reset, enable, taken_i : in std_logic;  prediction_o : out 
            std_logic);
   end component;
   
   component predictor_2_9
      port( clock, reset, enable, taken_i : in std_logic;  prediction_o : out 
            std_logic);
   end component;
   
   component predictor_2_10
      port( clock, reset, enable, taken_i : in std_logic;  prediction_o : out 
            std_logic);
   end component;
   
   component predictor_2_11
      port( clock, reset, enable, taken_i : in std_logic;  prediction_o : out 
            std_logic);
   end component;
   
   component predictor_2_12
      port( clock, reset, enable, taken_i : in std_logic;  prediction_o : out 
            std_logic);
   end component;
   
   component predictor_2_13
      port( clock, reset, enable, taken_i : in std_logic;  prediction_o : out 
            std_logic);
   end component;
   
   component predictor_2_14
      port( clock, reset, enable, taken_i : in std_logic;  prediction_o : out 
            std_logic);
   end component;
   
   component predictor_2_15
      port( clock, reset, enable, taken_i : in std_logic;  prediction_o : out 
            std_logic);
   end component;
   
   component predictor_2_0
      port( clock, reset, enable, taken_i : in std_logic;  prediction_o : out 
            std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFS_X1
      port( D, CK, SN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal predicted_next_PC_o_31_port, predicted_next_PC_o_30_port, 
      predicted_next_PC_o_29_port, predicted_next_PC_o_28_port, 
      predicted_next_PC_o_27_port, predicted_next_PC_o_26_port, 
      predicted_next_PC_o_25_port, predicted_next_PC_o_24_port, 
      predicted_next_PC_o_23_port, predicted_next_PC_o_22_port, 
      predicted_next_PC_o_21_port, predicted_next_PC_o_20_port, 
      predicted_next_PC_o_19_port, predicted_next_PC_o_18_port, 
      predicted_next_PC_o_17_port, predicted_next_PC_o_16_port, 
      predicted_next_PC_o_15_port, predicted_next_PC_o_14_port, 
      predicted_next_PC_o_13_port, predicted_next_PC_o_12_port, 
      predicted_next_PC_o_11_port, predicted_next_PC_o_10_port, 
      predicted_next_PC_o_9_port, predicted_next_PC_o_8_port, 
      predicted_next_PC_o_7_port, predicted_next_PC_o_6_port, 
      predicted_next_PC_o_5_port, predicted_next_PC_o_4_port, 
      predicted_next_PC_o_3_port, predicted_next_PC_o_2_port, 
      predicted_next_PC_o_1_port, predicted_next_PC_o_0_port, taken_o_port, 
      mispredict_o_port, taken_15_port, taken_14_port, taken_13_port, 
      taken_12_port, taken_11_port, taken_10_port, taken_9_port, taken_8_port, 
      taken_7_port, taken_6_port, taken_5_port, taken_4_port, taken_3_port, 
      taken_2_port, taken_1_port, taken_0_port, write_enable_15_port, 
      write_enable_14_port, write_enable_13_port, write_enable_12_port, 
      write_enable_11_port, write_enable_10_port, write_enable_9_port, 
      write_enable_8_port, write_enable_7_port, write_enable_6_port, 
      write_enable_5_port, write_enable_4_port, write_enable_3_port, 
      write_enable_2_port, write_enable_1_port, write_enable_0_port, 
      predict_PC_0_31_port, predict_PC_0_30_port, predict_PC_0_29_port, 
      predict_PC_0_28_port, predict_PC_0_27_port, predict_PC_0_26_port, 
      predict_PC_0_25_port, predict_PC_0_24_port, predict_PC_0_23_port, 
      predict_PC_0_22_port, predict_PC_0_21_port, predict_PC_0_20_port, 
      predict_PC_0_19_port, predict_PC_0_18_port, predict_PC_0_17_port, 
      predict_PC_0_16_port, predict_PC_0_15_port, predict_PC_0_14_port, 
      predict_PC_0_13_port, predict_PC_0_12_port, predict_PC_0_11_port, 
      predict_PC_0_10_port, predict_PC_0_9_port, predict_PC_0_8_port, 
      predict_PC_0_7_port, predict_PC_0_6_port, predict_PC_0_5_port, 
      predict_PC_0_4_port, predict_PC_0_3_port, predict_PC_0_2_port, 
      predict_PC_0_1_port, predict_PC_0_0_port, predict_PC_1_31_port, 
      predict_PC_1_30_port, predict_PC_1_29_port, predict_PC_1_28_port, 
      predict_PC_1_27_port, predict_PC_1_26_port, predict_PC_1_25_port, 
      predict_PC_1_24_port, predict_PC_1_23_port, predict_PC_1_22_port, 
      predict_PC_1_21_port, predict_PC_1_20_port, predict_PC_1_19_port, 
      predict_PC_1_18_port, predict_PC_1_17_port, predict_PC_1_16_port, 
      predict_PC_1_15_port, predict_PC_1_14_port, predict_PC_1_13_port, 
      predict_PC_1_12_port, predict_PC_1_11_port, predict_PC_1_10_port, 
      predict_PC_1_9_port, predict_PC_1_8_port, predict_PC_1_7_port, 
      predict_PC_1_6_port, predict_PC_1_5_port, predict_PC_1_4_port, 
      predict_PC_1_3_port, predict_PC_1_2_port, predict_PC_1_1_port, 
      predict_PC_1_0_port, predict_PC_2_31_port, predict_PC_2_30_port, 
      predict_PC_2_29_port, predict_PC_2_28_port, predict_PC_2_27_port, 
      predict_PC_2_26_port, predict_PC_2_25_port, predict_PC_2_24_port, 
      predict_PC_2_23_port, predict_PC_2_22_port, predict_PC_2_21_port, 
      predict_PC_2_20_port, predict_PC_2_19_port, predict_PC_2_18_port, 
      predict_PC_2_17_port, predict_PC_2_16_port, predict_PC_2_15_port, 
      predict_PC_2_14_port, predict_PC_2_13_port, predict_PC_2_12_port, 
      predict_PC_2_11_port, predict_PC_2_10_port, predict_PC_2_9_port, 
      predict_PC_2_8_port, predict_PC_2_7_port, predict_PC_2_6_port, 
      predict_PC_2_5_port, predict_PC_2_4_port, predict_PC_2_3_port, 
      predict_PC_2_2_port, predict_PC_2_1_port, predict_PC_2_0_port, 
      predict_PC_3_31_port, predict_PC_3_30_port, predict_PC_3_29_port, 
      predict_PC_3_28_port, predict_PC_3_27_port, predict_PC_3_26_port, 
      predict_PC_3_25_port, predict_PC_3_24_port, predict_PC_3_23_port, 
      predict_PC_3_22_port, predict_PC_3_21_port, predict_PC_3_20_port, 
      predict_PC_3_19_port, predict_PC_3_18_port, predict_PC_3_17_port, 
      predict_PC_3_16_port, predict_PC_3_15_port, predict_PC_3_14_port, 
      predict_PC_3_13_port, predict_PC_3_12_port, predict_PC_3_11_port, 
      predict_PC_3_10_port, predict_PC_3_9_port, predict_PC_3_8_port, 
      predict_PC_3_7_port, predict_PC_3_6_port, predict_PC_3_5_port, 
      predict_PC_3_4_port, predict_PC_3_3_port, predict_PC_3_2_port, 
      predict_PC_3_1_port, predict_PC_3_0_port, predict_PC_4_31_port, 
      predict_PC_4_30_port, predict_PC_4_29_port, predict_PC_4_28_port, 
      predict_PC_4_27_port, predict_PC_4_26_port, predict_PC_4_25_port, 
      predict_PC_4_24_port, predict_PC_4_23_port, predict_PC_4_22_port, 
      predict_PC_4_21_port, predict_PC_4_20_port, predict_PC_4_19_port, 
      predict_PC_4_18_port, predict_PC_4_17_port, predict_PC_4_16_port, 
      predict_PC_4_15_port, predict_PC_4_14_port, predict_PC_4_13_port, 
      predict_PC_4_12_port, predict_PC_4_11_port, predict_PC_4_10_port, 
      predict_PC_4_9_port, predict_PC_4_8_port, predict_PC_4_7_port, 
      predict_PC_4_6_port, predict_PC_4_5_port, predict_PC_4_4_port, 
      predict_PC_4_3_port, predict_PC_4_2_port, predict_PC_4_1_port, 
      predict_PC_4_0_port, predict_PC_5_31_port, predict_PC_5_30_port, 
      predict_PC_5_29_port, predict_PC_5_28_port, predict_PC_5_27_port, 
      predict_PC_5_26_port, predict_PC_5_25_port, predict_PC_5_24_port, 
      predict_PC_5_23_port, predict_PC_5_22_port, predict_PC_5_21_port, 
      predict_PC_5_20_port, predict_PC_5_19_port, predict_PC_5_18_port, 
      predict_PC_5_17_port, predict_PC_5_16_port, predict_PC_5_15_port, 
      predict_PC_5_14_port, predict_PC_5_13_port, predict_PC_5_12_port, 
      predict_PC_5_11_port, predict_PC_5_10_port, predict_PC_5_9_port, 
      predict_PC_5_8_port, predict_PC_5_7_port, predict_PC_5_6_port, 
      predict_PC_5_5_port, predict_PC_5_4_port, predict_PC_5_3_port, 
      predict_PC_5_2_port, predict_PC_5_1_port, predict_PC_5_0_port, 
      predict_PC_6_31_port, predict_PC_6_30_port, predict_PC_6_29_port, 
      predict_PC_6_28_port, predict_PC_6_27_port, predict_PC_6_26_port, 
      predict_PC_6_25_port, predict_PC_6_24_port, predict_PC_6_23_port, 
      predict_PC_6_22_port, predict_PC_6_21_port, predict_PC_6_20_port, 
      predict_PC_6_19_port, predict_PC_6_18_port, predict_PC_6_17_port, 
      predict_PC_6_16_port, predict_PC_6_15_port, predict_PC_6_14_port, 
      predict_PC_6_13_port, predict_PC_6_12_port, predict_PC_6_11_port, 
      predict_PC_6_10_port, predict_PC_6_9_port, predict_PC_6_8_port, 
      predict_PC_6_7_port, predict_PC_6_6_port, predict_PC_6_5_port, 
      predict_PC_6_4_port, predict_PC_6_3_port, predict_PC_6_2_port, 
      predict_PC_6_1_port, predict_PC_6_0_port, predict_PC_7_31_port, 
      predict_PC_7_30_port, predict_PC_7_29_port, predict_PC_7_28_port, 
      predict_PC_7_27_port, predict_PC_7_26_port, predict_PC_7_25_port, 
      predict_PC_7_24_port, predict_PC_7_23_port, predict_PC_7_22_port, 
      predict_PC_7_21_port, predict_PC_7_20_port, predict_PC_7_19_port, 
      predict_PC_7_18_port, predict_PC_7_17_port, predict_PC_7_16_port, 
      predict_PC_7_15_port, predict_PC_7_14_port, predict_PC_7_13_port, 
      predict_PC_7_12_port, predict_PC_7_11_port, predict_PC_7_10_port, 
      predict_PC_7_9_port, predict_PC_7_8_port, predict_PC_7_7_port, 
      predict_PC_7_6_port, predict_PC_7_5_port, predict_PC_7_4_port, 
      predict_PC_7_3_port, predict_PC_7_2_port, predict_PC_7_1_port, 
      predict_PC_7_0_port, predict_PC_8_31_port, predict_PC_8_30_port, 
      predict_PC_8_29_port, predict_PC_8_28_port, predict_PC_8_27_port, 
      predict_PC_8_26_port, predict_PC_8_25_port, predict_PC_8_24_port, 
      predict_PC_8_23_port, predict_PC_8_22_port, predict_PC_8_21_port, 
      predict_PC_8_20_port, predict_PC_8_19_port, predict_PC_8_18_port, 
      predict_PC_8_17_port, predict_PC_8_16_port, predict_PC_8_15_port, 
      predict_PC_8_14_port, predict_PC_8_13_port, predict_PC_8_12_port, 
      predict_PC_8_11_port, predict_PC_8_10_port, predict_PC_8_9_port, 
      predict_PC_8_8_port, predict_PC_8_7_port, predict_PC_8_6_port, 
      predict_PC_8_5_port, predict_PC_8_4_port, predict_PC_8_3_port, 
      predict_PC_8_2_port, predict_PC_8_1_port, predict_PC_8_0_port, 
      predict_PC_9_31_port, predict_PC_9_30_port, predict_PC_9_29_port, 
      predict_PC_9_28_port, predict_PC_9_27_port, predict_PC_9_26_port, 
      predict_PC_9_25_port, predict_PC_9_24_port, predict_PC_9_23_port, 
      predict_PC_9_22_port, predict_PC_9_21_port, predict_PC_9_20_port, 
      predict_PC_9_19_port, predict_PC_9_18_port, predict_PC_9_17_port, 
      predict_PC_9_16_port, predict_PC_9_15_port, predict_PC_9_14_port, 
      predict_PC_9_13_port, predict_PC_9_12_port, predict_PC_9_11_port, 
      predict_PC_9_10_port, predict_PC_9_9_port, predict_PC_9_8_port, 
      predict_PC_9_7_port, predict_PC_9_6_port, predict_PC_9_5_port, 
      predict_PC_9_4_port, predict_PC_9_3_port, predict_PC_9_2_port, 
      predict_PC_9_1_port, predict_PC_9_0_port, predict_PC_10_31_port, 
      predict_PC_10_30_port, predict_PC_10_29_port, predict_PC_10_28_port, 
      predict_PC_10_27_port, predict_PC_10_26_port, predict_PC_10_25_port, 
      predict_PC_10_24_port, predict_PC_10_23_port, predict_PC_10_22_port, 
      predict_PC_10_21_port, predict_PC_10_20_port, predict_PC_10_19_port, 
      predict_PC_10_18_port, predict_PC_10_17_port, predict_PC_10_16_port, 
      predict_PC_10_15_port, predict_PC_10_14_port, predict_PC_10_13_port, 
      predict_PC_10_12_port, predict_PC_10_11_port, predict_PC_10_10_port, 
      predict_PC_10_9_port, predict_PC_10_8_port, predict_PC_10_7_port, 
      predict_PC_10_6_port, predict_PC_10_5_port, predict_PC_10_4_port, 
      predict_PC_10_3_port, predict_PC_10_2_port, predict_PC_10_1_port, 
      predict_PC_10_0_port, predict_PC_11_31_port, predict_PC_11_30_port, 
      predict_PC_11_29_port, predict_PC_11_28_port, predict_PC_11_27_port, 
      predict_PC_11_26_port, predict_PC_11_25_port, predict_PC_11_24_port, 
      predict_PC_11_23_port, predict_PC_11_22_port, predict_PC_11_21_port, 
      predict_PC_11_20_port, predict_PC_11_19_port, predict_PC_11_18_port, 
      predict_PC_11_17_port, predict_PC_11_16_port, predict_PC_11_15_port, 
      predict_PC_11_14_port, predict_PC_11_13_port, predict_PC_11_12_port, 
      predict_PC_11_11_port, predict_PC_11_10_port, predict_PC_11_9_port, 
      predict_PC_11_8_port, predict_PC_11_7_port, predict_PC_11_6_port, 
      predict_PC_11_5_port, predict_PC_11_4_port, predict_PC_11_3_port, 
      predict_PC_11_2_port, predict_PC_11_1_port, predict_PC_11_0_port, 
      predict_PC_12_31_port, predict_PC_12_30_port, predict_PC_12_29_port, 
      predict_PC_12_28_port, predict_PC_12_27_port, predict_PC_12_26_port, 
      predict_PC_12_25_port, predict_PC_12_24_port, predict_PC_12_23_port, 
      predict_PC_12_22_port, predict_PC_12_21_port, predict_PC_12_20_port, 
      predict_PC_12_19_port, predict_PC_12_18_port, predict_PC_12_17_port, 
      predict_PC_12_16_port, predict_PC_12_15_port, predict_PC_12_14_port, 
      predict_PC_12_13_port, predict_PC_12_12_port, predict_PC_12_11_port, 
      predict_PC_12_10_port, predict_PC_12_9_port, predict_PC_12_8_port, 
      predict_PC_12_7_port, predict_PC_12_6_port, predict_PC_12_5_port, 
      predict_PC_12_4_port, predict_PC_12_3_port, predict_PC_12_2_port, 
      predict_PC_12_1_port, predict_PC_12_0_port, predict_PC_13_31_port, 
      predict_PC_13_30_port, predict_PC_13_29_port, predict_PC_13_28_port, 
      predict_PC_13_27_port, predict_PC_13_26_port, predict_PC_13_25_port, 
      predict_PC_13_24_port, predict_PC_13_23_port, predict_PC_13_22_port, 
      predict_PC_13_21_port, predict_PC_13_20_port, predict_PC_13_19_port, 
      predict_PC_13_18_port, predict_PC_13_17_port, predict_PC_13_16_port, 
      predict_PC_13_15_port, predict_PC_13_14_port, predict_PC_13_13_port, 
      predict_PC_13_12_port, predict_PC_13_11_port, predict_PC_13_10_port, 
      predict_PC_13_9_port, predict_PC_13_8_port, predict_PC_13_7_port, 
      predict_PC_13_6_port, predict_PC_13_5_port, predict_PC_13_4_port, 
      predict_PC_13_3_port, predict_PC_13_2_port, predict_PC_13_1_port, 
      predict_PC_13_0_port, predict_PC_14_31_port, predict_PC_14_30_port, 
      predict_PC_14_29_port, predict_PC_14_28_port, predict_PC_14_27_port, 
      predict_PC_14_26_port, predict_PC_14_25_port, predict_PC_14_24_port, 
      predict_PC_14_23_port, predict_PC_14_22_port, predict_PC_14_21_port, 
      predict_PC_14_20_port, predict_PC_14_19_port, predict_PC_14_18_port, 
      predict_PC_14_17_port, predict_PC_14_16_port, predict_PC_14_15_port, 
      predict_PC_14_14_port, predict_PC_14_13_port, predict_PC_14_12_port, 
      predict_PC_14_11_port, predict_PC_14_10_port, predict_PC_14_9_port, 
      predict_PC_14_8_port, predict_PC_14_7_port, predict_PC_14_6_port, 
      predict_PC_14_5_port, predict_PC_14_4_port, predict_PC_14_3_port, 
      predict_PC_14_2_port, predict_PC_14_1_port, predict_PC_14_0_port, 
      predict_PC_15_31_port, predict_PC_15_30_port, predict_PC_15_29_port, 
      predict_PC_15_28_port, predict_PC_15_27_port, predict_PC_15_26_port, 
      predict_PC_15_25_port, predict_PC_15_24_port, predict_PC_15_23_port, 
      predict_PC_15_22_port, predict_PC_15_21_port, predict_PC_15_20_port, 
      predict_PC_15_19_port, predict_PC_15_18_port, predict_PC_15_17_port, 
      predict_PC_15_16_port, predict_PC_15_15_port, predict_PC_15_14_port, 
      predict_PC_15_13_port, predict_PC_15_12_port, predict_PC_15_11_port, 
      predict_PC_15_10_port, predict_PC_15_9_port, predict_PC_15_8_port, 
      predict_PC_15_7_port, predict_PC_15_6_port, predict_PC_15_5_port, 
      predict_PC_15_4_port, predict_PC_15_3_port, predict_PC_15_2_port, 
      predict_PC_15_1_port, predict_PC_15_0_port, N38, N39, N40, N41, N42, N43,
      N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N86, N118, N150, N182, 
      N214, N246, N278, N310, N342, N374, N406, N438, N470, N502, N534, N566, 
      N567, net3621, net3626, net3631, net3636, net3641, net3646, net3651, 
      net3656, net3661, net3666, net3671, net3676, net3681, net3686, net3691, 
      net3696, net3701, n483, n485, n487, n489, n491, n493, n495, n497, n499, 
      n501, n503, n505, n507, n509, n511, n513, n515, n517, n519, n521, n523, 
      n525, n527, n529, n531, n533, n535, n537, n539, n541, n543, n545, n546, 
      n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, 
      n559, n560, n561, n562, n563, n564, n565, n566_port, n567_port, n568, 
      n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, 
      n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, 
      n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, 
      n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, 
      n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, 
      n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, 
      n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, 
      n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, 
      n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, 
      n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, 
      n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, 
      n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, 
      n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, 
      n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, 
      n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, 
      n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, 
      n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, 
      n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, 
      n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, 
      n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, 
      n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, 
      n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, 
      n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, 
      n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, 
      n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, 
      n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, 
      n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, 
      n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n943, 
      n944, n945, n946, n947, n948, n949, n951, n955, n956, n957, n958, n959, 
      n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, 
      n972, n973, n974, n975, n976, n977, n978, n979, n942, n941, n940, n939, 
      n938, n937, n936, n935, n934, n933, n932, n931, n930, n929, n928, n927, 
      n926, n925, n924, n923, n922, n921, n920, n919, n918, n917, n916, n915, 
      n914, n913, n912, n911, n906, n905, n1, n2, n3, n4, n5, n6, n7, n8, n9, 
      n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24
      , n25, n26, n27, n28, n29, n30, n31, n32, n33, n35, n36, n37, n38_port, 
      n39_port, n40_port, n41_port, n42_port, n43_port, n44_port, n45_port, 
      n46_port, n47_port, n48_port, n49_port, n50_port, n51_port, n52_port, 
      n53_port, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66
      , n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, 
      n81, n82, n83, n84, n85, n86_port, n87, n88, n89, n90, n91, n92, n93, n94
      , n95, n96, n97, n98, n99, n100, net47171, net47172, net47173, net47174, 
      net47175, net47176, net47177, net47178, net47179, net47180, net47181, 
      net47182, net47183, net47184, net47185, net47186, net47187, net47188, 
      net47189, net47190, net47191, net47192, net47193, net47194, net47195, 
      net47196, net47197, net47198, net47199, net47200, net47201, net47202, 
      net47203, net47204, net47205, net47206, net47207, net47208, net47209, 
      net47210, net47211, net47212, net47213, net47214, net47215, net47216, 
      net47217, net47218, net47219, net47220, net47221, net47222, net47223, 
      net47224, net47225, net47226, net47227, net47228, net47229, net47230, 
      net47231, net47232, net47233, net47234, net47235, net47236, net47237, 
      net47238, net47239, net47240, net47241, net47242, net47243, net47244, 
      net47245, net47246, net47247, net47248, net47249, net47250, net47251, 
      net47252, net47253, net47254, net47255, net47256, net47257, net47258, 
      net47259, net47260, net47261, net47262, net47263, net47264, net47265, 
      net47266, net47267, net47268, net47269, net47270, net47271, net47272, 
      net47273, net47274, net47275, net47276, net47277, net47278, net47279, 
      net47280, net47281, net47282, net47283, net47284, net47285, net47286, 
      net47287, net47288, net47289, net47290, net47291, net47292, net47293, 
      net47294, net47295, net47296, net47297, net47298, net47299, net47300, 
      net47301, net47302, net47303, net47304, net47305, net47306, net47307, 
      net47308, net47309, net47310, net47311, net47312, net47313, net47314, 
      net47315, net47316, net47317, net47318, net47319, net47320, net47321, 
      net47322, net47323, net47324, net47325, net47326, net47327, net47328, 
      net47329, net47330, net47331, net47332, net47333, net47334, net47335, 
      net47336, net47337, net47338, net47339, net47340, net47341, net47342, 
      net47343, net47344, net47345, net47346, net47347, net47348, net47349, 
      net47350, net47351, net47352, net47353, net47354, net47355, net47356, 
      net47357, net47358, net47359, net47360, net47361, net47362, net47363, 
      net47364, net47365, net47366, net47367, net47368, net47369, net47370, 
      net47371, net47372, net47373, net47374, net47375, net47376, net47377, 
      net47378, net47379, net47380, net47381, net47382, net47383, net47384, 
      net47385, net47386, net47387, net47388, net47389, net47390, net47391, 
      net47392, net47393, net47394, net47395, net47396, net47397, net47398, 
      net47399, net47400, net47401, net47402, net47403, net47404, net47405, 
      net47406, net47407, net47408, net47409, net47410, net47411, net47412, 
      net47413, net47414, net47415, net47416, net47417, net47418, net47419, 
      net47420, net47421, net47422, net47423, net47424, net47425, net47426, 
      net47427, net47428, net47429, net47430, net47431, net47432, net47433, 
      net47434, net47435, net47436, net47437, net47438, net47439, net47440, 
      net47441, net47442, net47443, net47444, net47445, net47446, net47447, 
      net47448, net47449, net47450, net47451, net47452, net47453, net47454, 
      net47455, net47456, net47457, net47458, net47459, net47460, net47461, 
      net47462, net47463, net47464, net47465, net47466, net47467, net47468, 
      net47469, net47470, net47471, net47472, net47473, net47474, net47475, 
      net47476, net47477, net47478, net47479, net47480, net47481, net47482, 
      net47483, net47484, net47485, net47486, net47487, net47488, net47489, 
      net47490, net47491, net47492, net47493, net47494, net47495, net47496, 
      net47497, net47498, net47499, net47500, net47501, net47502, net47503, 
      net47504, net47505, net47506, net47507, net47508, net47509, net47510, 
      net47511, net47512, net47513, net47514, net47515, net47516, net47517, 
      net47518, net47519, net47520, net47521, net47522, net47523, net47524, 
      net47525, net47526, net47527, net47528, net47529, net47530, net47531, 
      net47532, net47533, net47534, net47535, net47536, net47537, net47538, 
      net47539, net47540, net47541, net47542, net47543, net47544, net47545, 
      net47546, net47547, net47548, net47549, net47550, net47551, net47552, 
      net47553, net47554, net47555, net47556, net47557, net47558, net47559, 
      net47560, net47561, net47562, net47563, net47564, net47565, net47566, 
      net47567, net47568, net47569, net47570, net47571, net47572, net47573, 
      net47574, net47575, net47576, net47577, net47578, net47579, net47580, 
      net47581, net47582, net47583, net47584, net47585, net47586, net47587, 
      net47588, net47589, net47590, net47591, net47592, net47593, net47594, 
      net47595, net47596, net47597, net47598, net47599, net47600, net47601, 
      net47602, net47603, net47604, net47605, net47606, net47607, net47608, 
      net47609, net47610, net47611, net47612, net47613, net47614, net47615, 
      net47616, net47617, net47618, net47619, net47620, net47621, net47622, 
      net47623, net47624, net47625, net47626, net47627, net47628, net47629, 
      net47630, net47631, net47632, net47633, net47634, net47635, net47636, 
      net47637, net47638, net47639, net47640, net47641, net47642, net47643, 
      net47644, net47645, net47646, net47647, net47648, net47649, net47650, 
      net47651, net47652, net47653, net47654, net47655, net47656, net47657, 
      net47658, net47659, net47660, net47661, net47662, net47663, net47664, 
      net47665, net47666, net47667, net47668, net47669, net47670, net47671, 
      net47672, net47673, net47674, net47675, net47676, net47677, net47678, 
      net47679, net47680, net47681, net47682 : std_logic;

begin
   predicted_next_PC_o <= ( predicted_next_PC_o_31_port, 
      predicted_next_PC_o_30_port, predicted_next_PC_o_29_port, 
      predicted_next_PC_o_28_port, predicted_next_PC_o_27_port, 
      predicted_next_PC_o_26_port, predicted_next_PC_o_25_port, 
      predicted_next_PC_o_24_port, predicted_next_PC_o_23_port, 
      predicted_next_PC_o_22_port, predicted_next_PC_o_21_port, 
      predicted_next_PC_o_20_port, predicted_next_PC_o_19_port, 
      predicted_next_PC_o_18_port, predicted_next_PC_o_17_port, 
      predicted_next_PC_o_16_port, predicted_next_PC_o_15_port, 
      predicted_next_PC_o_14_port, predicted_next_PC_o_13_port, 
      predicted_next_PC_o_12_port, predicted_next_PC_o_11_port, 
      predicted_next_PC_o_10_port, predicted_next_PC_o_9_port, 
      predicted_next_PC_o_8_port, predicted_next_PC_o_7_port, 
      predicted_next_PC_o_6_port, predicted_next_PC_o_5_port, 
      predicted_next_PC_o_4_port, predicted_next_PC_o_3_port, 
      predicted_next_PC_o_2_port, predicted_next_PC_o_1_port, 
      predicted_next_PC_o_0_port );
   taken_o <= taken_o_port;
   mispredict_o <= mispredict_o_port;
   
   last_TAG_reg_3_inst : DFFS_X1 port map( D => n972, CK => net3621, SN => 
                           n86_port, Q => n977, QN => n53_port);
   last_TAG_reg_2_inst : DFFS_X1 port map( D => n973, CK => net3621, SN => n77,
                           Q => n976, QN => n51_port);
   last_TAG_reg_1_inst : DFFS_X1 port map( D => n974, CK => net3621, SN => n79,
                           Q => n979, QN => n52_port);
   last_TAG_reg_0_inst : DFFR_X1 port map( D => TAG_i(0), CK => net3621, RN => 
                           n87, Q => n50_port, QN => n978);
   write_enable_reg_15_inst : DFFR_X1 port map( D => N53, CK => net3621, RN => 
                           n81, Q => write_enable_15_port, QN => n971);
   write_enable_reg_14_inst : DFFR_X1 port map( D => N52, CK => net3621, RN => 
                           n79, Q => write_enable_14_port, QN => n970);
   write_enable_reg_13_inst : DFFR_X1 port map( D => N51, CK => net3621, RN => 
                           n82, Q => write_enable_13_port, QN => n969);
   write_enable_reg_12_inst : DFFR_X1 port map( D => N50, CK => net3621, RN => 
                           n83, Q => write_enable_12_port, QN => n968);
   write_enable_reg_11_inst : DFFR_X1 port map( D => N49, CK => net3621, RN => 
                           n85, Q => write_enable_11_port, QN => n967);
   write_enable_reg_10_inst : DFFR_X1 port map( D => N48, CK => net3621, RN => 
                           n86_port, Q => write_enable_10_port, QN => n966);
   write_enable_reg_9_inst : DFFR_X1 port map( D => N47, CK => net3621, RN => 
                           n85, Q => write_enable_9_port, QN => n965);
   write_enable_reg_8_inst : DFFR_X1 port map( D => N46, CK => net3621, RN => 
                           n84, Q => write_enable_8_port, QN => n964);
   write_enable_reg_7_inst : DFFR_X1 port map( D => N45, CK => net3621, RN => 
                           n87, Q => write_enable_7_port, QN => n963);
   write_enable_reg_6_inst : DFFR_X1 port map( D => N44, CK => net3621, RN => 
                           n84, Q => write_enable_6_port, QN => n962);
   write_enable_reg_5_inst : DFFR_X1 port map( D => N43, CK => net3621, RN => 
                           n86_port, Q => write_enable_5_port, QN => n961);
   write_enable_reg_4_inst : DFFR_X1 port map( D => N42, CK => net3621, RN => 
                           n85, Q => write_enable_4_port, QN => n960);
   write_enable_reg_3_inst : DFFR_X1 port map( D => N41, CK => net3621, RN => 
                           n84, Q => write_enable_3_port, QN => n959);
   write_enable_reg_2_inst : DFFR_X1 port map( D => N40, CK => net3621, RN => 
                           n87, Q => write_enable_2_port, QN => n958);
   write_enable_reg_1_inst : DFFR_X1 port map( D => N39, CK => net3621, RN => 
                           n87, Q => write_enable_1_port, QN => n957);
   write_enable_reg_0_inst : DFFR_X1 port map( D => N38, CK => net3621, RN => 
                           n86_port, Q => write_enable_0_port, QN => n956);
   last_taken_reg : DFF_X1 port map( D => n955, CK => clock, Q => n54, QN => 
                           n975);
   predict_PC_reg_0_31_inst : DFFR_X1 port map( D => n59, CK => net3626, RN => 
                           n87, Q => predict_PC_0_31_port, QN => net47682);
   predict_PC_reg_0_30_inst : DFFR_X1 port map( D => n38_port, CK => net3626, 
                           RN => n84, Q => predict_PC_0_30_port, QN => net47681
                           );
   predict_PC_reg_0_29_inst : DFFR_X1 port map( D => n58, CK => net3626, RN => 
                           n85, Q => predict_PC_0_29_port, QN => net47680);
   predict_PC_reg_0_28_inst : DFFR_X1 port map( D => n39_port, CK => net3626, 
                           RN => n86_port, Q => predict_PC_0_28_port, QN => 
                           net47679);
   predict_PC_reg_0_27_inst : DFFR_X1 port map( D => n60, CK => net3626, RN => 
                           n87, Q => predict_PC_0_27_port, QN => net47678);
   predict_PC_reg_0_26_inst : DFFR_X1 port map( D => n37, CK => net3626, RN => 
                           n84, Q => predict_PC_0_26_port, QN => net47677);
   predict_PC_reg_0_25_inst : DFFR_X1 port map( D => n35, CK => net3626, RN => 
                           n85, Q => predict_PC_0_25_port, QN => net47676);
   predict_PC_reg_0_24_inst : DFFR_X1 port map( D => n36, CK => net3626, RN => 
                           n86_port, Q => predict_PC_0_24_port, QN => net47675)
                           ;
   predict_PC_reg_0_23_inst : DFFR_X1 port map( D => target_PC_i(23), CK => 
                           net3626, RN => n87, Q => predict_PC_0_23_port, QN =>
                           net47674);
   predict_PC_reg_0_22_inst : DFFR_X1 port map( D => target_PC_i(22), CK => 
                           net3626, RN => n84, Q => predict_PC_0_22_port, QN =>
                           net47673);
   predict_PC_reg_0_21_inst : DFFR_X1 port map( D => target_PC_i(21), CK => 
                           net3626, RN => n85, Q => predict_PC_0_21_port, QN =>
                           net47672);
   predict_PC_reg_0_20_inst : DFFR_X1 port map( D => target_PC_i(20), CK => 
                           net3626, RN => n86_port, Q => predict_PC_0_20_port, 
                           QN => net47671);
   predict_PC_reg_0_19_inst : DFFR_X1 port map( D => target_PC_i(19), CK => 
                           net3626, RN => n84, Q => predict_PC_0_19_port, QN =>
                           net47670);
   predict_PC_reg_0_18_inst : DFFR_X1 port map( D => target_PC_i(18), CK => 
                           net3626, RN => n84, Q => predict_PC_0_18_port, QN =>
                           net47669);
   predict_PC_reg_0_17_inst : DFFR_X1 port map( D => target_PC_i(17), CK => 
                           net3626, RN => n84, Q => predict_PC_0_17_port, QN =>
                           net47668);
   predict_PC_reg_0_16_inst : DFFR_X1 port map( D => target_PC_i(16), CK => 
                           net3626, RN => n84, Q => predict_PC_0_16_port, QN =>
                           net47667);
   predict_PC_reg_0_15_inst : DFFR_X1 port map( D => target_PC_i(15), CK => 
                           net3626, RN => n84, Q => predict_PC_0_15_port, QN =>
                           net47666);
   predict_PC_reg_0_14_inst : DFFR_X1 port map( D => target_PC_i(14), CK => 
                           net3626, RN => n84, Q => predict_PC_0_14_port, QN =>
                           net47665);
   predict_PC_reg_0_13_inst : DFFR_X1 port map( D => target_PC_i(13), CK => 
                           net3626, RN => n84, Q => predict_PC_0_13_port, QN =>
                           net47664);
   predict_PC_reg_0_12_inst : DFFR_X1 port map( D => target_PC_i(12), CK => 
                           net3626, RN => n84, Q => predict_PC_0_12_port, QN =>
                           net47663);
   predict_PC_reg_0_11_inst : DFFR_X1 port map( D => target_PC_i(11), CK => 
                           net3626, RN => n84, Q => predict_PC_0_11_port, QN =>
                           net47662);
   predict_PC_reg_0_10_inst : DFFR_X1 port map( D => target_PC_i(10), CK => 
                           net3626, RN => n84, Q => predict_PC_0_10_port, QN =>
                           net47661);
   predict_PC_reg_0_9_inst : DFFR_X1 port map( D => target_PC_i(9), CK => 
                           net3626, RN => n84, Q => predict_PC_0_9_port, QN => 
                           net47660);
   predict_PC_reg_0_8_inst : DFFR_X1 port map( D => target_PC_i(8), CK => 
                           net3626, RN => n84, Q => predict_PC_0_8_port, QN => 
                           net47659);
   predict_PC_reg_0_7_inst : DFFR_X1 port map( D => target_PC_i(7), CK => 
                           net3626, RN => n85, Q => predict_PC_0_7_port, QN => 
                           net47658);
   predict_PC_reg_0_6_inst : DFFR_X1 port map( D => target_PC_i(6), CK => 
                           net3626, RN => n85, Q => predict_PC_0_6_port, QN => 
                           net47657);
   predict_PC_reg_0_5_inst : DFFR_X1 port map( D => target_PC_i(5), CK => 
                           net3626, RN => n85, Q => predict_PC_0_5_port, QN => 
                           net47656);
   predict_PC_reg_0_4_inst : DFFR_X1 port map( D => target_PC_i(4), CK => 
                           net3626, RN => n85, Q => predict_PC_0_4_port, QN => 
                           net47655);
   predict_PC_reg_0_3_inst : DFFR_X1 port map( D => target_PC_i(3), CK => 
                           net3626, RN => n85, Q => predict_PC_0_3_port, QN => 
                           net47654);
   predict_PC_reg_0_2_inst : DFFR_X1 port map( D => target_PC_i(2), CK => 
                           net3626, RN => n85, Q => predict_PC_0_2_port, QN => 
                           net47653);
   predict_PC_reg_0_1_inst : DFFR_X1 port map( D => target_PC_i(1), CK => 
                           net3626, RN => n85, Q => predict_PC_0_1_port, QN => 
                           net47652);
   predict_PC_reg_0_0_inst : DFFR_X1 port map( D => target_PC_i(0), CK => 
                           net3626, RN => n85, Q => predict_PC_0_0_port, QN => 
                           net47651);
   predict_PC_reg_1_31_inst : DFFR_X1 port map( D => n59, CK => net3631, RN => 
                           n85, Q => predict_PC_1_31_port, QN => net47650);
   predict_PC_reg_1_30_inst : DFFR_X1 port map( D => n38_port, CK => net3631, 
                           RN => n85, Q => predict_PC_1_30_port, QN => net47649
                           );
   predict_PC_reg_1_29_inst : DFFR_X1 port map( D => n58, CK => net3631, RN => 
                           n85, Q => predict_PC_1_29_port, QN => net47648);
   predict_PC_reg_1_28_inst : DFFR_X1 port map( D => n39_port, CK => net3631, 
                           RN => n85, Q => predict_PC_1_28_port, QN => net47647
                           );
   predict_PC_reg_1_27_inst : DFFR_X1 port map( D => n60, CK => net3631, RN => 
                           n86_port, Q => predict_PC_1_27_port, QN => net47646)
                           ;
   predict_PC_reg_1_26_inst : DFFR_X1 port map( D => n37, CK => net3631, RN => 
                           n86_port, Q => predict_PC_1_26_port, QN => net47645)
                           ;
   predict_PC_reg_1_25_inst : DFFR_X1 port map( D => n35, CK => net3631, RN => 
                           n86_port, Q => predict_PC_1_25_port, QN => net47644)
                           ;
   predict_PC_reg_1_24_inst : DFFR_X1 port map( D => n36, CK => net3631, RN => 
                           n86_port, Q => predict_PC_1_24_port, QN => net47643)
                           ;
   predict_PC_reg_1_23_inst : DFFR_X1 port map( D => target_PC_i(23), CK => 
                           net3631, RN => n86_port, Q => predict_PC_1_23_port, 
                           QN => net47642);
   predict_PC_reg_1_22_inst : DFFR_X1 port map( D => target_PC_i(22), CK => 
                           net3631, RN => n86_port, Q => predict_PC_1_22_port, 
                           QN => net47641);
   predict_PC_reg_1_21_inst : DFFR_X1 port map( D => target_PC_i(21), CK => 
                           net3631, RN => n86_port, Q => predict_PC_1_21_port, 
                           QN => net47640);
   predict_PC_reg_1_20_inst : DFFR_X1 port map( D => target_PC_i(20), CK => 
                           net3631, RN => n86_port, Q => predict_PC_1_20_port, 
                           QN => net47639);
   predict_PC_reg_1_19_inst : DFFR_X1 port map( D => target_PC_i(19), CK => 
                           net3631, RN => n86_port, Q => predict_PC_1_19_port, 
                           QN => net47638);
   predict_PC_reg_1_18_inst : DFFR_X1 port map( D => target_PC_i(18), CK => 
                           net3631, RN => n86_port, Q => predict_PC_1_18_port, 
                           QN => net47637);
   predict_PC_reg_1_17_inst : DFFR_X1 port map( D => target_PC_i(17), CK => 
                           net3631, RN => n86_port, Q => predict_PC_1_17_port, 
                           QN => net47636);
   predict_PC_reg_1_16_inst : DFFR_X1 port map( D => target_PC_i(16), CK => 
                           net3631, RN => n86_port, Q => predict_PC_1_16_port, 
                           QN => net47635);
   predict_PC_reg_1_15_inst : DFFR_X1 port map( D => target_PC_i(15), CK => 
                           net3631, RN => n87, Q => predict_PC_1_15_port, QN =>
                           net47634);
   predict_PC_reg_1_14_inst : DFFR_X1 port map( D => target_PC_i(14), CK => 
                           net3631, RN => n87, Q => predict_PC_1_14_port, QN =>
                           net47633);
   predict_PC_reg_1_13_inst : DFFR_X1 port map( D => target_PC_i(13), CK => 
                           net3631, RN => n87, Q => predict_PC_1_13_port, QN =>
                           net47632);
   predict_PC_reg_1_12_inst : DFFR_X1 port map( D => target_PC_i(12), CK => 
                           net3631, RN => n87, Q => predict_PC_1_12_port, QN =>
                           net47631);
   predict_PC_reg_1_11_inst : DFFR_X1 port map( D => target_PC_i(11), CK => 
                           net3631, RN => n87, Q => predict_PC_1_11_port, QN =>
                           net47630);
   predict_PC_reg_1_10_inst : DFFR_X1 port map( D => target_PC_i(10), CK => 
                           net3631, RN => n87, Q => predict_PC_1_10_port, QN =>
                           net47629);
   predict_PC_reg_1_9_inst : DFFR_X1 port map( D => target_PC_i(9), CK => 
                           net3631, RN => n87, Q => predict_PC_1_9_port, QN => 
                           net47628);
   predict_PC_reg_1_8_inst : DFFR_X1 port map( D => target_PC_i(8), CK => 
                           net3631, RN => n87, Q => predict_PC_1_8_port, QN => 
                           net47627);
   predict_PC_reg_1_7_inst : DFFR_X1 port map( D => target_PC_i(7), CK => 
                           net3631, RN => n87, Q => predict_PC_1_7_port, QN => 
                           net47626);
   predict_PC_reg_1_6_inst : DFFR_X1 port map( D => target_PC_i(6), CK => 
                           net3631, RN => n87, Q => predict_PC_1_6_port, QN => 
                           net47625);
   predict_PC_reg_1_5_inst : DFFR_X1 port map( D => target_PC_i(5), CK => 
                           net3631, RN => n87, Q => predict_PC_1_5_port, QN => 
                           net47624);
   predict_PC_reg_1_4_inst : DFFR_X1 port map( D => target_PC_i(4), CK => 
                           net3631, RN => n88, Q => predict_PC_1_4_port, QN => 
                           net47623);
   predict_PC_reg_1_3_inst : DFFR_X1 port map( D => target_PC_i(3), CK => 
                           net3631, RN => n88, Q => predict_PC_1_3_port, QN => 
                           net47622);
   predict_PC_reg_1_2_inst : DFFR_X1 port map( D => target_PC_i(2), CK => 
                           net3631, RN => n88, Q => predict_PC_1_2_port, QN => 
                           net47621);
   predict_PC_reg_1_1_inst : DFFR_X1 port map( D => target_PC_i(1), CK => 
                           net3631, RN => n88, Q => predict_PC_1_1_port, QN => 
                           net47620);
   predict_PC_reg_1_0_inst : DFFR_X1 port map( D => target_PC_i(0), CK => 
                           net3631, RN => n88, Q => predict_PC_1_0_port, QN => 
                           net47619);
   predict_PC_reg_2_31_inst : DFFR_X1 port map( D => n59, CK => net3636, RN => 
                           n88, Q => predict_PC_2_31_port, QN => net47618);
   predict_PC_reg_2_30_inst : DFFR_X1 port map( D => n38_port, CK => net3636, 
                           RN => n88, Q => predict_PC_2_30_port, QN => net47617
                           );
   predict_PC_reg_2_29_inst : DFFR_X1 port map( D => n58, CK => net3636, RN => 
                           n88, Q => predict_PC_2_29_port, QN => net47616);
   predict_PC_reg_2_28_inst : DFFR_X1 port map( D => n39_port, CK => net3636, 
                           RN => n88, Q => predict_PC_2_28_port, QN => net47615
                           );
   predict_PC_reg_2_27_inst : DFFR_X1 port map( D => n60, CK => net3636, RN => 
                           n88, Q => predict_PC_2_27_port, QN => net47614);
   predict_PC_reg_2_26_inst : DFFR_X1 port map( D => n37, CK => net3636, RN => 
                           n88, Q => predict_PC_2_26_port, QN => net47613);
   predict_PC_reg_2_25_inst : DFFR_X1 port map( D => n35, CK => net3636, RN => 
                           n88, Q => predict_PC_2_25_port, QN => net47612);
   predict_PC_reg_2_24_inst : DFFR_X1 port map( D => n36, CK => net3636, RN => 
                           n89, Q => predict_PC_2_24_port, QN => net47611);
   predict_PC_reg_2_23_inst : DFFR_X1 port map( D => target_PC_i(23), CK => 
                           net3636, RN => n89, Q => predict_PC_2_23_port, QN =>
                           net47610);
   predict_PC_reg_2_22_inst : DFFR_X1 port map( D => target_PC_i(22), CK => 
                           net3636, RN => n89, Q => predict_PC_2_22_port, QN =>
                           net47609);
   predict_PC_reg_2_21_inst : DFFR_X1 port map( D => target_PC_i(21), CK => 
                           net3636, RN => n89, Q => predict_PC_2_21_port, QN =>
                           net47608);
   predict_PC_reg_2_20_inst : DFFR_X1 port map( D => target_PC_i(20), CK => 
                           net3636, RN => n89, Q => predict_PC_2_20_port, QN =>
                           net47607);
   predict_PC_reg_2_19_inst : DFFR_X1 port map( D => target_PC_i(19), CK => 
                           net3636, RN => n89, Q => predict_PC_2_19_port, QN =>
                           net47606);
   predict_PC_reg_2_18_inst : DFFR_X1 port map( D => target_PC_i(18), CK => 
                           net3636, RN => n89, Q => predict_PC_2_18_port, QN =>
                           net47605);
   predict_PC_reg_2_17_inst : DFFR_X1 port map( D => target_PC_i(17), CK => 
                           net3636, RN => n89, Q => predict_PC_2_17_port, QN =>
                           net47604);
   predict_PC_reg_2_16_inst : DFFR_X1 port map( D => target_PC_i(16), CK => 
                           net3636, RN => n89, Q => predict_PC_2_16_port, QN =>
                           net47603);
   predict_PC_reg_2_15_inst : DFFR_X1 port map( D => target_PC_i(15), CK => 
                           net3636, RN => n89, Q => predict_PC_2_15_port, QN =>
                           net47602);
   predict_PC_reg_2_14_inst : DFFR_X1 port map( D => target_PC_i(14), CK => 
                           net3636, RN => n89, Q => predict_PC_2_14_port, QN =>
                           net47601);
   predict_PC_reg_2_13_inst : DFFR_X1 port map( D => target_PC_i(13), CK => 
                           net3636, RN => n89, Q => predict_PC_2_13_port, QN =>
                           net47600);
   predict_PC_reg_2_12_inst : DFFR_X1 port map( D => target_PC_i(12), CK => 
                           net3636, RN => n90, Q => predict_PC_2_12_port, QN =>
                           net47599);
   predict_PC_reg_2_11_inst : DFFR_X1 port map( D => target_PC_i(11), CK => 
                           net3636, RN => n90, Q => predict_PC_2_11_port, QN =>
                           net47598);
   predict_PC_reg_2_10_inst : DFFR_X1 port map( D => target_PC_i(10), CK => 
                           net3636, RN => n90, Q => predict_PC_2_10_port, QN =>
                           net47597);
   predict_PC_reg_2_9_inst : DFFR_X1 port map( D => target_PC_i(9), CK => 
                           net3636, RN => n90, Q => predict_PC_2_9_port, QN => 
                           net47596);
   predict_PC_reg_2_8_inst : DFFR_X1 port map( D => target_PC_i(8), CK => 
                           net3636, RN => n90, Q => predict_PC_2_8_port, QN => 
                           net47595);
   predict_PC_reg_2_7_inst : DFFR_X1 port map( D => target_PC_i(7), CK => 
                           net3636, RN => n90, Q => predict_PC_2_7_port, QN => 
                           net47594);
   predict_PC_reg_2_6_inst : DFFR_X1 port map( D => target_PC_i(6), CK => 
                           net3636, RN => n90, Q => predict_PC_2_6_port, QN => 
                           net47593);
   predict_PC_reg_2_5_inst : DFFR_X1 port map( D => target_PC_i(5), CK => 
                           net3636, RN => n90, Q => predict_PC_2_5_port, QN => 
                           net47592);
   predict_PC_reg_2_4_inst : DFFR_X1 port map( D => target_PC_i(4), CK => 
                           net3636, RN => n90, Q => predict_PC_2_4_port, QN => 
                           net47591);
   predict_PC_reg_2_3_inst : DFFR_X1 port map( D => target_PC_i(3), CK => 
                           net3636, RN => n90, Q => predict_PC_2_3_port, QN => 
                           net47590);
   predict_PC_reg_2_2_inst : DFFR_X1 port map( D => target_PC_i(2), CK => 
                           net3636, RN => n90, Q => predict_PC_2_2_port, QN => 
                           net47589);
   predict_PC_reg_2_1_inst : DFFR_X1 port map( D => target_PC_i(1), CK => 
                           net3636, RN => n90, Q => predict_PC_2_1_port, QN => 
                           net47588);
   predict_PC_reg_2_0_inst : DFFR_X1 port map( D => target_PC_i(0), CK => 
                           net3636, RN => n91, Q => predict_PC_2_0_port, QN => 
                           net47587);
   predict_PC_reg_3_31_inst : DFFR_X1 port map( D => n59, CK => net3641, RN => 
                           n91, Q => predict_PC_3_31_port, QN => net47586);
   predict_PC_reg_3_30_inst : DFFR_X1 port map( D => target_PC_i(30), CK => 
                           net3641, RN => n91, Q => predict_PC_3_30_port, QN =>
                           net47585);
   predict_PC_reg_3_29_inst : DFFR_X1 port map( D => n58, CK => net3641, RN => 
                           n91, Q => predict_PC_3_29_port, QN => net47584);
   predict_PC_reg_3_28_inst : DFFR_X1 port map( D => n39_port, CK => net3641, 
                           RN => n91, Q => predict_PC_3_28_port, QN => net47583
                           );
   predict_PC_reg_3_27_inst : DFFR_X1 port map( D => target_PC_i(27), CK => 
                           net3641, RN => n91, Q => predict_PC_3_27_port, QN =>
                           net47582);
   predict_PC_reg_3_26_inst : DFFR_X1 port map( D => n37, CK => net3641, RN => 
                           n91, Q => predict_PC_3_26_port, QN => net47581);
   predict_PC_reg_3_25_inst : DFFR_X1 port map( D => n35, CK => net3641, RN => 
                           n91, Q => predict_PC_3_25_port, QN => net47580);
   predict_PC_reg_3_24_inst : DFFR_X1 port map( D => n36, CK => net3641, RN => 
                           n91, Q => predict_PC_3_24_port, QN => net47579);
   predict_PC_reg_3_23_inst : DFFR_X1 port map( D => target_PC_i(23), CK => 
                           net3641, RN => n91, Q => predict_PC_3_23_port, QN =>
                           net47578);
   predict_PC_reg_3_22_inst : DFFR_X1 port map( D => target_PC_i(22), CK => 
                           net3641, RN => n91, Q => predict_PC_3_22_port, QN =>
                           net47577);
   predict_PC_reg_3_21_inst : DFFR_X1 port map( D => target_PC_i(21), CK => 
                           net3641, RN => n91, Q => predict_PC_3_21_port, QN =>
                           net47576);
   predict_PC_reg_3_20_inst : DFFR_X1 port map( D => target_PC_i(20), CK => 
                           net3641, RN => n92, Q => predict_PC_3_20_port, QN =>
                           net47575);
   predict_PC_reg_3_19_inst : DFFR_X1 port map( D => target_PC_i(19), CK => 
                           net3641, RN => n92, Q => predict_PC_3_19_port, QN =>
                           net47574);
   predict_PC_reg_3_18_inst : DFFR_X1 port map( D => target_PC_i(18), CK => 
                           net3641, RN => n92, Q => predict_PC_3_18_port, QN =>
                           net47573);
   predict_PC_reg_3_17_inst : DFFR_X1 port map( D => target_PC_i(17), CK => 
                           net3641, RN => n92, Q => predict_PC_3_17_port, QN =>
                           net47572);
   predict_PC_reg_3_16_inst : DFFR_X1 port map( D => target_PC_i(16), CK => 
                           net3641, RN => n92, Q => predict_PC_3_16_port, QN =>
                           net47571);
   predict_PC_reg_3_15_inst : DFFR_X1 port map( D => target_PC_i(15), CK => 
                           net3641, RN => n92, Q => predict_PC_3_15_port, QN =>
                           net47570);
   predict_PC_reg_3_14_inst : DFFR_X1 port map( D => target_PC_i(14), CK => 
                           net3641, RN => n92, Q => predict_PC_3_14_port, QN =>
                           net47569);
   predict_PC_reg_3_13_inst : DFFR_X1 port map( D => target_PC_i(13), CK => 
                           net3641, RN => n92, Q => predict_PC_3_13_port, QN =>
                           net47568);
   predict_PC_reg_3_12_inst : DFFR_X1 port map( D => target_PC_i(12), CK => 
                           net3641, RN => n92, Q => predict_PC_3_12_port, QN =>
                           net47567);
   predict_PC_reg_3_11_inst : DFFR_X1 port map( D => target_PC_i(11), CK => 
                           net3641, RN => n92, Q => predict_PC_3_11_port, QN =>
                           net47566);
   predict_PC_reg_3_10_inst : DFFR_X1 port map( D => target_PC_i(10), CK => 
                           net3641, RN => n92, Q => predict_PC_3_10_port, QN =>
                           net47565);
   predict_PC_reg_3_9_inst : DFFR_X1 port map( D => target_PC_i(9), CK => 
                           net3641, RN => n92, Q => predict_PC_3_9_port, QN => 
                           net47564);
   predict_PC_reg_3_8_inst : DFFR_X1 port map( D => target_PC_i(8), CK => 
                           net3641, RN => n93, Q => predict_PC_3_8_port, QN => 
                           net47563);
   predict_PC_reg_3_7_inst : DFFR_X1 port map( D => target_PC_i(7), CK => 
                           net3641, RN => n93, Q => predict_PC_3_7_port, QN => 
                           net47562);
   predict_PC_reg_3_6_inst : DFFR_X1 port map( D => target_PC_i(6), CK => 
                           net3641, RN => n93, Q => predict_PC_3_6_port, QN => 
                           net47561);
   predict_PC_reg_3_5_inst : DFFR_X1 port map( D => target_PC_i(5), CK => 
                           net3641, RN => n93, Q => predict_PC_3_5_port, QN => 
                           net47560);
   predict_PC_reg_3_4_inst : DFFR_X1 port map( D => target_PC_i(4), CK => 
                           net3641, RN => n93, Q => predict_PC_3_4_port, QN => 
                           net47559);
   predict_PC_reg_3_3_inst : DFFR_X1 port map( D => target_PC_i(3), CK => 
                           net3641, RN => n93, Q => predict_PC_3_3_port, QN => 
                           net47558);
   predict_PC_reg_3_2_inst : DFFR_X1 port map( D => target_PC_i(2), CK => 
                           net3641, RN => n80, Q => predict_PC_3_2_port, QN => 
                           net47557);
   predict_PC_reg_3_1_inst : DFFR_X1 port map( D => target_PC_i(1), CK => 
                           net3641, RN => n77, Q => predict_PC_3_1_port, QN => 
                           net47556);
   predict_PC_reg_3_0_inst : DFFR_X1 port map( D => target_PC_i(0), CK => 
                           net3641, RN => n78, Q => predict_PC_3_0_port, QN => 
                           net47555);
   predict_PC_reg_4_31_inst : DFFR_X1 port map( D => n59, CK => net3646, RN => 
                           n78, Q => predict_PC_4_31_port, QN => net47554);
   predict_PC_reg_4_30_inst : DFFR_X1 port map( D => n38_port, CK => net3646, 
                           RN => n79, Q => predict_PC_4_30_port, QN => net47553
                           );
   predict_PC_reg_4_29_inst : DFFR_X1 port map( D => n58, CK => net3646, RN => 
                           n77, Q => predict_PC_4_29_port, QN => net47552);
   predict_PC_reg_4_28_inst : DFFR_X1 port map( D => n39_port, CK => net3646, 
                           RN => n79, Q => predict_PC_4_28_port, QN => net47551
                           );
   predict_PC_reg_4_27_inst : DFFR_X1 port map( D => n60, CK => net3646, RN => 
                           n78, Q => predict_PC_4_27_port, QN => net47550);
   predict_PC_reg_4_26_inst : DFFR_X1 port map( D => target_PC_i(26), CK => 
                           net3646, RN => n79, Q => predict_PC_4_26_port, QN =>
                           net47549);
   predict_PC_reg_4_25_inst : DFFR_X1 port map( D => n35, CK => net3646, RN => 
                           n77, Q => predict_PC_4_25_port, QN => net47548);
   predict_PC_reg_4_24_inst : DFFR_X1 port map( D => target_PC_i(24), CK => 
                           net3646, RN => n77, Q => predict_PC_4_24_port, QN =>
                           net47547);
   predict_PC_reg_4_23_inst : DFFR_X1 port map( D => target_PC_i(23), CK => 
                           net3646, RN => n78, Q => predict_PC_4_23_port, QN =>
                           net47546);
   predict_PC_reg_4_22_inst : DFFR_X1 port map( D => target_PC_i(22), CK => 
                           net3646, RN => n78, Q => predict_PC_4_22_port, QN =>
                           net47545);
   predict_PC_reg_4_21_inst : DFFR_X1 port map( D => target_PC_i(21), CK => 
                           net3646, RN => n77, Q => predict_PC_4_21_port, QN =>
                           net47544);
   predict_PC_reg_4_20_inst : DFFR_X1 port map( D => target_PC_i(20), CK => 
                           net3646, RN => n78, Q => predict_PC_4_20_port, QN =>
                           net47543);
   predict_PC_reg_4_19_inst : DFFR_X1 port map( D => target_PC_i(19), CK => 
                           net3646, RN => n79, Q => predict_PC_4_19_port, QN =>
                           net47542);
   predict_PC_reg_4_18_inst : DFFR_X1 port map( D => target_PC_i(18), CK => 
                           net3646, RN => n77, Q => predict_PC_4_18_port, QN =>
                           net47541);
   predict_PC_reg_4_17_inst : DFFR_X1 port map( D => target_PC_i(17), CK => 
                           net3646, RN => n78, Q => predict_PC_4_17_port, QN =>
                           net47540);
   predict_PC_reg_4_16_inst : DFFR_X1 port map( D => target_PC_i(16), CK => 
                           net3646, RN => n79, Q => predict_PC_4_16_port, QN =>
                           net47539);
   predict_PC_reg_4_15_inst : DFFR_X1 port map( D => target_PC_i(15), CK => 
                           net3646, RN => n77, Q => predict_PC_4_15_port, QN =>
                           net47538);
   predict_PC_reg_4_14_inst : DFFR_X1 port map( D => target_PC_i(14), CK => 
                           net3646, RN => n78, Q => predict_PC_4_14_port, QN =>
                           net47537);
   predict_PC_reg_4_13_inst : DFFR_X1 port map( D => target_PC_i(13), CK => 
                           net3646, RN => n79, Q => predict_PC_4_13_port, QN =>
                           net47536);
   predict_PC_reg_4_12_inst : DFFR_X1 port map( D => target_PC_i(12), CK => 
                           net3646, RN => n77, Q => predict_PC_4_12_port, QN =>
                           net47535);
   predict_PC_reg_4_11_inst : DFFR_X1 port map( D => target_PC_i(11), CK => 
                           net3646, RN => n78, Q => predict_PC_4_11_port, QN =>
                           net47534);
   predict_PC_reg_4_10_inst : DFFR_X1 port map( D => target_PC_i(10), CK => 
                           net3646, RN => n77, Q => predict_PC_4_10_port, QN =>
                           net47533);
   predict_PC_reg_4_9_inst : DFFR_X1 port map( D => target_PC_i(9), CK => 
                           net3646, RN => n77, Q => predict_PC_4_9_port, QN => 
                           net47532);
   predict_PC_reg_4_8_inst : DFFR_X1 port map( D => target_PC_i(8), CK => 
                           net3646, RN => n77, Q => predict_PC_4_8_port, QN => 
                           net47531);
   predict_PC_reg_4_7_inst : DFFR_X1 port map( D => target_PC_i(7), CK => 
                           net3646, RN => n77, Q => predict_PC_4_7_port, QN => 
                           net47530);
   predict_PC_reg_4_6_inst : DFFR_X1 port map( D => target_PC_i(6), CK => 
                           net3646, RN => n77, Q => predict_PC_4_6_port, QN => 
                           net47529);
   predict_PC_reg_4_5_inst : DFFR_X1 port map( D => target_PC_i(5), CK => 
                           net3646, RN => n77, Q => predict_PC_4_5_port, QN => 
                           net47528);
   predict_PC_reg_4_4_inst : DFFR_X1 port map( D => target_PC_i(4), CK => 
                           net3646, RN => n77, Q => predict_PC_4_4_port, QN => 
                           net47527);
   predict_PC_reg_4_3_inst : DFFR_X1 port map( D => target_PC_i(3), CK => 
                           net3646, RN => n77, Q => predict_PC_4_3_port, QN => 
                           net47526);
   predict_PC_reg_4_2_inst : DFFR_X1 port map( D => target_PC_i(2), CK => 
                           net3646, RN => n77, Q => predict_PC_4_2_port, QN => 
                           net47525);
   predict_PC_reg_4_1_inst : DFFR_X1 port map( D => target_PC_i(1), CK => 
                           net3646, RN => n77, Q => predict_PC_4_1_port, QN => 
                           net47524);
   predict_PC_reg_4_0_inst : DFFR_X1 port map( D => target_PC_i(0), CK => 
                           net3646, RN => n77, Q => predict_PC_4_0_port, QN => 
                           net47523);
   predict_PC_reg_5_31_inst : DFFR_X1 port map( D => n59, CK => net3651, RN => 
                           n77, Q => predict_PC_5_31_port, QN => net47522);
   predict_PC_reg_5_30_inst : DFFR_X1 port map( D => n38_port, CK => net3651, 
                           RN => n78, Q => predict_PC_5_30_port, QN => net47521
                           );
   predict_PC_reg_5_29_inst : DFFR_X1 port map( D => n58, CK => net3651, RN => 
                           n78, Q => predict_PC_5_29_port, QN => net47520);
   predict_PC_reg_5_28_inst : DFFR_X1 port map( D => n39_port, CK => net3651, 
                           RN => n78, Q => predict_PC_5_28_port, QN => net47519
                           );
   predict_PC_reg_5_27_inst : DFFR_X1 port map( D => n60, CK => net3651, RN => 
                           n78, Q => predict_PC_5_27_port, QN => net47518);
   predict_PC_reg_5_26_inst : DFFR_X1 port map( D => n37, CK => net3651, RN => 
                           n78, Q => predict_PC_5_26_port, QN => net47517);
   predict_PC_reg_5_25_inst : DFFR_X1 port map( D => n35, CK => net3651, RN => 
                           n78, Q => predict_PC_5_25_port, QN => net47516);
   predict_PC_reg_5_24_inst : DFFR_X1 port map( D => n36, CK => net3651, RN => 
                           n78, Q => predict_PC_5_24_port, QN => net47515);
   predict_PC_reg_5_23_inst : DFFR_X1 port map( D => target_PC_i(23), CK => 
                           net3651, RN => n78, Q => predict_PC_5_23_port, QN =>
                           net47514);
   predict_PC_reg_5_22_inst : DFFR_X1 port map( D => target_PC_i(22), CK => 
                           net3651, RN => n78, Q => predict_PC_5_22_port, QN =>
                           net47513);
   predict_PC_reg_5_21_inst : DFFR_X1 port map( D => target_PC_i(21), CK => 
                           net3651, RN => n78, Q => predict_PC_5_21_port, QN =>
                           net47512);
   predict_PC_reg_5_20_inst : DFFR_X1 port map( D => target_PC_i(20), CK => 
                           net3651, RN => n78, Q => predict_PC_5_20_port, QN =>
                           net47511);
   predict_PC_reg_5_19_inst : DFFR_X1 port map( D => target_PC_i(19), CK => 
                           net3651, RN => n78, Q => predict_PC_5_19_port, QN =>
                           net47510);
   predict_PC_reg_5_18_inst : DFFR_X1 port map( D => target_PC_i(18), CK => 
                           net3651, RN => n79, Q => predict_PC_5_18_port, QN =>
                           net47509);
   predict_PC_reg_5_17_inst : DFFR_X1 port map( D => target_PC_i(17), CK => 
                           net3651, RN => n79, Q => predict_PC_5_17_port, QN =>
                           net47508);
   predict_PC_reg_5_16_inst : DFFR_X1 port map( D => target_PC_i(16), CK => 
                           net3651, RN => n79, Q => predict_PC_5_16_port, QN =>
                           net47507);
   predict_PC_reg_5_15_inst : DFFR_X1 port map( D => target_PC_i(15), CK => 
                           net3651, RN => n79, Q => predict_PC_5_15_port, QN =>
                           net47506);
   predict_PC_reg_5_14_inst : DFFR_X1 port map( D => target_PC_i(14), CK => 
                           net3651, RN => n79, Q => predict_PC_5_14_port, QN =>
                           net47505);
   predict_PC_reg_5_13_inst : DFFR_X1 port map( D => target_PC_i(13), CK => 
                           net3651, RN => n79, Q => predict_PC_5_13_port, QN =>
                           net47504);
   predict_PC_reg_5_12_inst : DFFR_X1 port map( D => target_PC_i(12), CK => 
                           net3651, RN => n79, Q => predict_PC_5_12_port, QN =>
                           net47503);
   predict_PC_reg_5_11_inst : DFFR_X1 port map( D => target_PC_i(11), CK => 
                           net3651, RN => n79, Q => predict_PC_5_11_port, QN =>
                           net47502);
   predict_PC_reg_5_10_inst : DFFR_X1 port map( D => target_PC_i(10), CK => 
                           net3651, RN => n79, Q => predict_PC_5_10_port, QN =>
                           net47501);
   predict_PC_reg_5_9_inst : DFFR_X1 port map( D => target_PC_i(9), CK => 
                           net3651, RN => n79, Q => predict_PC_5_9_port, QN => 
                           net47500);
   predict_PC_reg_5_8_inst : DFFR_X1 port map( D => target_PC_i(8), CK => 
                           net3651, RN => n79, Q => predict_PC_5_8_port, QN => 
                           net47499);
   predict_PC_reg_5_7_inst : DFFR_X1 port map( D => target_PC_i(7), CK => 
                           net3651, RN => n79, Q => predict_PC_5_7_port, QN => 
                           net47498);
   predict_PC_reg_5_6_inst : DFFR_X1 port map( D => target_PC_i(6), CK => 
                           net3651, RN => n80, Q => predict_PC_5_6_port, QN => 
                           net47497);
   predict_PC_reg_5_5_inst : DFFR_X1 port map( D => target_PC_i(5), CK => 
                           net3651, RN => n81, Q => predict_PC_5_5_port, QN => 
                           net47496);
   predict_PC_reg_5_4_inst : DFFR_X1 port map( D => target_PC_i(4), CK => 
                           net3651, RN => n82, Q => predict_PC_5_4_port, QN => 
                           net47495);
   predict_PC_reg_5_3_inst : DFFR_X1 port map( D => target_PC_i(3), CK => 
                           net3651, RN => n83, Q => predict_PC_5_3_port, QN => 
                           net47494);
   predict_PC_reg_5_2_inst : DFFR_X1 port map( D => target_PC_i(2), CK => 
                           net3651, RN => n83, Q => predict_PC_5_2_port, QN => 
                           net47493);
   predict_PC_reg_5_1_inst : DFFR_X1 port map( D => target_PC_i(1), CK => 
                           net3651, RN => n80, Q => predict_PC_5_1_port, QN => 
                           net47492);
   predict_PC_reg_5_0_inst : DFFR_X1 port map( D => target_PC_i(0), CK => 
                           net3651, RN => n81, Q => predict_PC_5_0_port, QN => 
                           net47491);
   predict_PC_reg_6_31_inst : DFFR_X1 port map( D => n59, CK => net3656, RN => 
                           n82, Q => predict_PC_6_31_port, QN => net47490);
   predict_PC_reg_6_30_inst : DFFR_X1 port map( D => n38_port, CK => net3656, 
                           RN => n83, Q => predict_PC_6_30_port, QN => net47489
                           );
   predict_PC_reg_6_29_inst : DFFR_X1 port map( D => n58, CK => net3656, RN => 
                           n83, Q => predict_PC_6_29_port, QN => net47488);
   predict_PC_reg_6_28_inst : DFFR_X1 port map( D => n39_port, CK => net3656, 
                           RN => n81, Q => predict_PC_6_28_port, QN => net47487
                           );
   predict_PC_reg_6_27_inst : DFFR_X1 port map( D => n60, CK => net3656, RN => 
                           n81, Q => predict_PC_6_27_port, QN => net47486);
   predict_PC_reg_6_26_inst : DFFR_X1 port map( D => n37, CK => net3656, RN => 
                           n82, Q => predict_PC_6_26_port, QN => net47485);
   predict_PC_reg_6_25_inst : DFFR_X1 port map( D => n35, CK => net3656, RN => 
                           n83, Q => predict_PC_6_25_port, QN => net47484);
   predict_PC_reg_6_24_inst : DFFR_X1 port map( D => n36, CK => net3656, RN => 
                           n80, Q => predict_PC_6_24_port, QN => net47483);
   predict_PC_reg_6_23_inst : DFFR_X1 port map( D => target_PC_i(23), CK => 
                           net3656, RN => n81, Q => predict_PC_6_23_port, QN =>
                           net47482);
   predict_PC_reg_6_22_inst : DFFR_X1 port map( D => target_PC_i(22), CK => 
                           net3656, RN => n82, Q => predict_PC_6_22_port, QN =>
                           net47481);
   predict_PC_reg_6_21_inst : DFFR_X1 port map( D => target_PC_i(21), CK => 
                           net3656, RN => n83, Q => predict_PC_6_21_port, QN =>
                           net47480);
   predict_PC_reg_6_20_inst : DFFR_X1 port map( D => target_PC_i(20), CK => 
                           net3656, RN => n80, Q => predict_PC_6_20_port, QN =>
                           net47479);
   predict_PC_reg_6_19_inst : DFFR_X1 port map( D => target_PC_i(19), CK => 
                           net3656, RN => n81, Q => predict_PC_6_19_port, QN =>
                           net47478);
   predict_PC_reg_6_18_inst : DFFR_X1 port map( D => target_PC_i(18), CK => 
                           net3656, RN => n82, Q => predict_PC_6_18_port, QN =>
                           net47477);
   predict_PC_reg_6_17_inst : DFFR_X1 port map( D => target_PC_i(17), CK => 
                           net3656, RN => n83, Q => predict_PC_6_17_port, QN =>
                           net47476);
   predict_PC_reg_6_16_inst : DFFR_X1 port map( D => target_PC_i(16), CK => 
                           net3656, RN => n80, Q => predict_PC_6_16_port, QN =>
                           net47475);
   predict_PC_reg_6_15_inst : DFFR_X1 port map( D => target_PC_i(15), CK => 
                           net3656, RN => n80, Q => predict_PC_6_15_port, QN =>
                           net47474);
   predict_PC_reg_6_14_inst : DFFR_X1 port map( D => target_PC_i(14), CK => 
                           net3656, RN => n80, Q => predict_PC_6_14_port, QN =>
                           net47473);
   predict_PC_reg_6_13_inst : DFFR_X1 port map( D => target_PC_i(13), CK => 
                           net3656, RN => n80, Q => predict_PC_6_13_port, QN =>
                           net47472);
   predict_PC_reg_6_12_inst : DFFR_X1 port map( D => target_PC_i(12), CK => 
                           net3656, RN => n80, Q => predict_PC_6_12_port, QN =>
                           net47471);
   predict_PC_reg_6_11_inst : DFFR_X1 port map( D => target_PC_i(11), CK => 
                           net3656, RN => n80, Q => predict_PC_6_11_port, QN =>
                           net47470);
   predict_PC_reg_6_10_inst : DFFR_X1 port map( D => target_PC_i(10), CK => 
                           net3656, RN => n80, Q => predict_PC_6_10_port, QN =>
                           net47469);
   predict_PC_reg_6_9_inst : DFFR_X1 port map( D => target_PC_i(9), CK => 
                           net3656, RN => n80, Q => predict_PC_6_9_port, QN => 
                           net47468);
   predict_PC_reg_6_8_inst : DFFR_X1 port map( D => target_PC_i(8), CK => 
                           net3656, RN => n80, Q => predict_PC_6_8_port, QN => 
                           net47467);
   predict_PC_reg_6_7_inst : DFFR_X1 port map( D => target_PC_i(7), CK => 
                           net3656, RN => n80, Q => predict_PC_6_7_port, QN => 
                           net47466);
   predict_PC_reg_6_6_inst : DFFR_X1 port map( D => target_PC_i(6), CK => 
                           net3656, RN => n80, Q => predict_PC_6_6_port, QN => 
                           net47465);
   predict_PC_reg_6_5_inst : DFFR_X1 port map( D => target_PC_i(5), CK => 
                           net3656, RN => n80, Q => predict_PC_6_5_port, QN => 
                           net47464);
   predict_PC_reg_6_4_inst : DFFR_X1 port map( D => target_PC_i(4), CK => 
                           net3656, RN => n80, Q => predict_PC_6_4_port, QN => 
                           net47463);
   predict_PC_reg_6_3_inst : DFFR_X1 port map( D => target_PC_i(3), CK => 
                           net3656, RN => n81, Q => predict_PC_6_3_port, QN => 
                           net47462);
   predict_PC_reg_6_2_inst : DFFR_X1 port map( D => target_PC_i(2), CK => 
                           net3656, RN => n81, Q => predict_PC_6_2_port, QN => 
                           net47461);
   predict_PC_reg_6_1_inst : DFFR_X1 port map( D => target_PC_i(1), CK => 
                           net3656, RN => n81, Q => predict_PC_6_1_port, QN => 
                           net47460);
   predict_PC_reg_6_0_inst : DFFR_X1 port map( D => target_PC_i(0), CK => 
                           net3656, RN => n81, Q => predict_PC_6_0_port, QN => 
                           net47459);
   predict_PC_reg_7_31_inst : DFFR_X1 port map( D => n59, CK => net3661, RN => 
                           n81, Q => predict_PC_7_31_port, QN => net47458);
   predict_PC_reg_7_30_inst : DFFR_X1 port map( D => n38_port, CK => net3661, 
                           RN => n81, Q => predict_PC_7_30_port, QN => net47457
                           );
   predict_PC_reg_7_29_inst : DFFR_X1 port map( D => n58, CK => net3661, RN => 
                           n81, Q => predict_PC_7_29_port, QN => net47456);
   predict_PC_reg_7_28_inst : DFFR_X1 port map( D => n39_port, CK => net3661, 
                           RN => n81, Q => predict_PC_7_28_port, QN => net47455
                           );
   predict_PC_reg_7_27_inst : DFFR_X1 port map( D => n60, CK => net3661, RN => 
                           n81, Q => predict_PC_7_27_port, QN => net47454);
   predict_PC_reg_7_26_inst : DFFR_X1 port map( D => n37, CK => net3661, RN => 
                           n81, Q => predict_PC_7_26_port, QN => net47453);
   predict_PC_reg_7_25_inst : DFFR_X1 port map( D => n35, CK => net3661, RN => 
                           n81, Q => predict_PC_7_25_port, QN => net47452);
   predict_PC_reg_7_24_inst : DFFR_X1 port map( D => n36, CK => net3661, RN => 
                           n81, Q => predict_PC_7_24_port, QN => net47451);
   predict_PC_reg_7_23_inst : DFFR_X1 port map( D => target_PC_i(23), CK => 
                           net3661, RN => n82, Q => predict_PC_7_23_port, QN =>
                           net47450);
   predict_PC_reg_7_22_inst : DFFR_X1 port map( D => target_PC_i(22), CK => 
                           net3661, RN => n82, Q => predict_PC_7_22_port, QN =>
                           net47449);
   predict_PC_reg_7_21_inst : DFFR_X1 port map( D => target_PC_i(21), CK => 
                           net3661, RN => n82, Q => predict_PC_7_21_port, QN =>
                           net47448);
   predict_PC_reg_7_20_inst : DFFR_X1 port map( D => target_PC_i(20), CK => 
                           net3661, RN => n82, Q => predict_PC_7_20_port, QN =>
                           net47447);
   predict_PC_reg_7_19_inst : DFFR_X1 port map( D => target_PC_i(19), CK => 
                           net3661, RN => n82, Q => predict_PC_7_19_port, QN =>
                           net47446);
   predict_PC_reg_7_18_inst : DFFR_X1 port map( D => target_PC_i(18), CK => 
                           net3661, RN => n82, Q => predict_PC_7_18_port, QN =>
                           net47445);
   predict_PC_reg_7_17_inst : DFFR_X1 port map( D => target_PC_i(17), CK => 
                           net3661, RN => n82, Q => predict_PC_7_17_port, QN =>
                           net47444);
   predict_PC_reg_7_16_inst : DFFR_X1 port map( D => target_PC_i(16), CK => 
                           net3661, RN => n82, Q => predict_PC_7_16_port, QN =>
                           net47443);
   predict_PC_reg_7_15_inst : DFFR_X1 port map( D => target_PC_i(15), CK => 
                           net3661, RN => n82, Q => predict_PC_7_15_port, QN =>
                           net47442);
   predict_PC_reg_7_14_inst : DFFR_X1 port map( D => target_PC_i(14), CK => 
                           net3661, RN => n82, Q => predict_PC_7_14_port, QN =>
                           net47441);
   predict_PC_reg_7_13_inst : DFFR_X1 port map( D => target_PC_i(13), CK => 
                           net3661, RN => n82, Q => predict_PC_7_13_port, QN =>
                           net47440);
   predict_PC_reg_7_12_inst : DFFR_X1 port map( D => target_PC_i(12), CK => 
                           net3661, RN => n82, Q => predict_PC_7_12_port, QN =>
                           net47439);
   predict_PC_reg_7_11_inst : DFFR_X1 port map( D => target_PC_i(11), CK => 
                           net3661, RN => n83, Q => predict_PC_7_11_port, QN =>
                           net47438);
   predict_PC_reg_7_10_inst : DFFR_X1 port map( D => target_PC_i(10), CK => 
                           net3661, RN => n83, Q => predict_PC_7_10_port, QN =>
                           net47437);
   predict_PC_reg_7_9_inst : DFFR_X1 port map( D => target_PC_i(9), CK => 
                           net3661, RN => n83, Q => predict_PC_7_9_port, QN => 
                           net47436);
   predict_PC_reg_7_8_inst : DFFR_X1 port map( D => target_PC_i(8), CK => 
                           net3661, RN => n83, Q => predict_PC_7_8_port, QN => 
                           net47435);
   predict_PC_reg_7_7_inst : DFFR_X1 port map( D => target_PC_i(7), CK => 
                           net3661, RN => n83, Q => predict_PC_7_7_port, QN => 
                           net47434);
   predict_PC_reg_7_6_inst : DFFR_X1 port map( D => target_PC_i(6), CK => 
                           net3661, RN => n83, Q => predict_PC_7_6_port, QN => 
                           net47433);
   predict_PC_reg_7_5_inst : DFFR_X1 port map( D => target_PC_i(5), CK => 
                           net3661, RN => n83, Q => predict_PC_7_5_port, QN => 
                           net47432);
   predict_PC_reg_7_4_inst : DFFR_X1 port map( D => target_PC_i(4), CK => 
                           net3661, RN => n83, Q => predict_PC_7_4_port, QN => 
                           net47431);
   predict_PC_reg_7_3_inst : DFFR_X1 port map( D => target_PC_i(3), CK => 
                           net3661, RN => n83, Q => predict_PC_7_3_port, QN => 
                           net47430);
   predict_PC_reg_7_2_inst : DFFR_X1 port map( D => target_PC_i(2), CK => 
                           net3661, RN => n83, Q => predict_PC_7_2_port, QN => 
                           net47429);
   predict_PC_reg_7_1_inst : DFFR_X1 port map( D => target_PC_i(1), CK => 
                           net3661, RN => n83, Q => predict_PC_7_1_port, QN => 
                           net47428);
   predict_PC_reg_7_0_inst : DFFR_X1 port map( D => target_PC_i(0), CK => 
                           net3661, RN => n83, Q => predict_PC_7_0_port, QN => 
                           net47427);
   predict_PC_reg_8_31_inst : DFFR_X1 port map( D => n59, CK => net3666, RN => 
                           n82, Q => predict_PC_8_31_port, QN => net47426);
   predict_PC_reg_8_30_inst : DFFR_X1 port map( D => target_PC_i(30), CK => 
                           net3666, RN => n81, Q => predict_PC_8_30_port, QN =>
                           net47425);
   predict_PC_reg_8_29_inst : DFFR_X1 port map( D => n58, CK => net3666, RN => 
                           n80, Q => predict_PC_8_29_port, QN => net47424);
   predict_PC_reg_8_28_inst : DFFR_X1 port map( D => n39_port, CK => net3666, 
                           RN => n81, Q => predict_PC_8_28_port, QN => net47423
                           );
   predict_PC_reg_8_27_inst : DFFR_X1 port map( D => target_PC_i(27), CK => 
                           net3666, RN => n82, Q => predict_PC_8_27_port, QN =>
                           net47422);
   predict_PC_reg_8_26_inst : DFFR_X1 port map( D => n37, CK => net3666, RN => 
                           n83, Q => predict_PC_8_26_port, QN => net47421);
   predict_PC_reg_8_25_inst : DFFR_X1 port map( D => n35, CK => net3666, RN => 
                           n80, Q => predict_PC_8_25_port, QN => net47420);
   predict_PC_reg_8_24_inst : DFFR_X1 port map( D => n36, CK => net3666, RN => 
                           n82, Q => predict_PC_8_24_port, QN => net47419);
   predict_PC_reg_8_23_inst : DFFR_X1 port map( D => target_PC_i(23), CK => 
                           net3666, RN => n80, Q => predict_PC_8_23_port, QN =>
                           net47418);
   predict_PC_reg_8_22_inst : DFFR_X1 port map( D => target_PC_i(22), CK => 
                           net3666, RN => n97, Q => predict_PC_8_22_port, QN =>
                           net47417);
   predict_PC_reg_8_21_inst : DFFR_X1 port map( D => target_PC_i(21), CK => 
                           net3666, RN => n97, Q => predict_PC_8_21_port, QN =>
                           net47416);
   predict_PC_reg_8_20_inst : DFFR_X1 port map( D => target_PC_i(20), CK => 
                           net3666, RN => n85, Q => predict_PC_8_20_port, QN =>
                           net47415);
   predict_PC_reg_8_19_inst : DFFR_X1 port map( D => target_PC_i(19), CK => 
                           net3666, RN => n91, Q => predict_PC_8_19_port, QN =>
                           net47414);
   predict_PC_reg_8_18_inst : DFFR_X1 port map( D => target_PC_i(18), CK => 
                           net3666, RN => n90, Q => predict_PC_8_18_port, QN =>
                           net47413);
   predict_PC_reg_8_17_inst : DFFR_X1 port map( D => target_PC_i(17), CK => 
                           net3666, RN => n89, Q => predict_PC_8_17_port, QN =>
                           net47412);
   predict_PC_reg_8_16_inst : DFFR_X1 port map( D => target_PC_i(16), CK => 
                           net3666, RN => n88, Q => predict_PC_8_16_port, QN =>
                           net47411);
   predict_PC_reg_8_15_inst : DFFR_X1 port map( D => target_PC_i(15), CK => 
                           net3666, RN => n93, Q => predict_PC_8_15_port, QN =>
                           net47410);
   predict_PC_reg_8_14_inst : DFFR_X1 port map( D => target_PC_i(14), CK => 
                           net3666, RN => n92, Q => predict_PC_8_14_port, QN =>
                           net47409);
   predict_PC_reg_8_13_inst : DFFR_X1 port map( D => target_PC_i(13), CK => 
                           net3666, RN => n94, Q => predict_PC_8_13_port, QN =>
                           net47408);
   predict_PC_reg_8_12_inst : DFFR_X1 port map( D => target_PC_i(12), CK => 
                           net3666, RN => n87, Q => predict_PC_8_12_port, QN =>
                           net47407);
   predict_PC_reg_8_11_inst : DFFR_X1 port map( D => target_PC_i(11), CK => 
                           net3666, RN => n99, Q => predict_PC_8_11_port, QN =>
                           net47406);
   predict_PC_reg_8_10_inst : DFFR_X1 port map( D => target_PC_i(10), CK => 
                           net3666, RN => n91, Q => predict_PC_8_10_port, QN =>
                           net47405);
   predict_PC_reg_8_9_inst : DFFR_X1 port map( D => target_PC_i(9), CK => 
                           net3666, RN => n92, Q => predict_PC_8_9_port, QN => 
                           net47404);
   predict_PC_reg_8_8_inst : DFFR_X1 port map( D => target_PC_i(8), CK => 
                           net3666, RN => n92, Q => predict_PC_8_8_port, QN => 
                           net47403);
   predict_PC_reg_8_7_inst : DFFR_X1 port map( D => target_PC_i(7), CK => 
                           net3666, RN => n82, Q => predict_PC_8_7_port, QN => 
                           net47402);
   predict_PC_reg_8_6_inst : DFFR_X1 port map( D => target_PC_i(6), CK => 
                           net3666, RN => n90, Q => predict_PC_8_6_port, QN => 
                           net47401);
   predict_PC_reg_8_5_inst : DFFR_X1 port map( D => target_PC_i(5), CK => 
                           net3666, RN => n98, Q => predict_PC_8_5_port, QN => 
                           net47400);
   predict_PC_reg_8_4_inst : DFFR_X1 port map( D => target_PC_i(4), CK => 
                           net3666, RN => n96, Q => predict_PC_8_4_port, QN => 
                           net47399);
   predict_PC_reg_8_3_inst : DFFR_X1 port map( D => target_PC_i(3), CK => 
                           net3666, RN => n92, Q => predict_PC_8_3_port, QN => 
                           net47398);
   predict_PC_reg_8_2_inst : DFFR_X1 port map( D => target_PC_i(2), CK => 
                           net3666, RN => n84, Q => predict_PC_8_2_port, QN => 
                           net47397);
   predict_PC_reg_8_1_inst : DFFR_X1 port map( D => target_PC_i(1), CK => 
                           net3666, RN => n93, Q => predict_PC_8_1_port, QN => 
                           net47396);
   predict_PC_reg_8_0_inst : DFFR_X1 port map( D => target_PC_i(0), CK => 
                           net3666, RN => n83, Q => predict_PC_8_0_port, QN => 
                           net47395);
   predict_PC_reg_9_31_inst : DFFR_X1 port map( D => n59, CK => net3671, RN => 
                           n97, Q => predict_PC_9_31_port, QN => net47394);
   predict_PC_reg_9_30_inst : DFFR_X1 port map( D => n38_port, CK => net3671, 
                           RN => n97, Q => predict_PC_9_30_port, QN => net47393
                           );
   predict_PC_reg_9_29_inst : DFFR_X1 port map( D => n58, CK => net3671, RN => 
                           n97, Q => predict_PC_9_29_port, QN => net47392);
   predict_PC_reg_9_28_inst : DFFR_X1 port map( D => n39_port, CK => net3671, 
                           RN => n97, Q => predict_PC_9_28_port, QN => net47391
                           );
   predict_PC_reg_9_27_inst : DFFR_X1 port map( D => n60, CK => net3671, RN => 
                           n97, Q => predict_PC_9_27_port, QN => net47390);
   predict_PC_reg_9_26_inst : DFFR_X1 port map( D => n37, CK => net3671, RN => 
                           n97, Q => predict_PC_9_26_port, QN => net47389);
   predict_PC_reg_9_25_inst : DFFR_X1 port map( D => n35, CK => net3671, RN => 
                           n97, Q => predict_PC_9_25_port, QN => net47388);
   predict_PC_reg_9_24_inst : DFFR_X1 port map( D => n36, CK => net3671, RN => 
                           n97, Q => predict_PC_9_24_port, QN => net47387);
   predict_PC_reg_9_23_inst : DFFR_X1 port map( D => target_PC_i(23), CK => 
                           net3671, RN => n97, Q => predict_PC_9_23_port, QN =>
                           net47386);
   predict_PC_reg_9_22_inst : DFFR_X1 port map( D => target_PC_i(22), CK => 
                           net3671, RN => n97, Q => predict_PC_9_22_port, QN =>
                           net47385);
   predict_PC_reg_9_21_inst : DFFR_X1 port map( D => target_PC_i(21), CK => 
                           net3671, RN => n97, Q => predict_PC_9_21_port, QN =>
                           net47384);
   predict_PC_reg_9_20_inst : DFFR_X1 port map( D => target_PC_i(20), CK => 
                           net3671, RN => n97, Q => predict_PC_9_20_port, QN =>
                           net47383);
   predict_PC_reg_9_19_inst : DFFR_X1 port map( D => target_PC_i(19), CK => 
                           net3671, RN => n98, Q => predict_PC_9_19_port, QN =>
                           net47382);
   predict_PC_reg_9_18_inst : DFFR_X1 port map( D => target_PC_i(18), CK => 
                           net3671, RN => n98, Q => predict_PC_9_18_port, QN =>
                           net47381);
   predict_PC_reg_9_17_inst : DFFR_X1 port map( D => target_PC_i(17), CK => 
                           net3671, RN => n98, Q => predict_PC_9_17_port, QN =>
                           net47380);
   predict_PC_reg_9_16_inst : DFFR_X1 port map( D => target_PC_i(16), CK => 
                           net3671, RN => n98, Q => predict_PC_9_16_port, QN =>
                           net47379);
   predict_PC_reg_9_15_inst : DFFR_X1 port map( D => target_PC_i(15), CK => 
                           net3671, RN => n98, Q => predict_PC_9_15_port, QN =>
                           net47378);
   predict_PC_reg_9_14_inst : DFFR_X1 port map( D => target_PC_i(14), CK => 
                           net3671, RN => n98, Q => predict_PC_9_14_port, QN =>
                           net47377);
   predict_PC_reg_9_13_inst : DFFR_X1 port map( D => target_PC_i(13), CK => 
                           net3671, RN => n98, Q => predict_PC_9_13_port, QN =>
                           net47376);
   predict_PC_reg_9_12_inst : DFFR_X1 port map( D => target_PC_i(12), CK => 
                           net3671, RN => n98, Q => predict_PC_9_12_port, QN =>
                           net47375);
   predict_PC_reg_9_11_inst : DFFR_X1 port map( D => target_PC_i(11), CK => 
                           net3671, RN => n98, Q => predict_PC_9_11_port, QN =>
                           net47374);
   predict_PC_reg_9_10_inst : DFFR_X1 port map( D => target_PC_i(10), CK => 
                           net3671, RN => n98, Q => predict_PC_9_10_port, QN =>
                           net47373);
   predict_PC_reg_9_9_inst : DFFR_X1 port map( D => target_PC_i(9), CK => 
                           net3671, RN => n98, Q => predict_PC_9_9_port, QN => 
                           net47372);
   predict_PC_reg_9_8_inst : DFFR_X1 port map( D => target_PC_i(8), CK => 
                           net3671, RN => n98, Q => predict_PC_9_8_port, QN => 
                           net47371);
   predict_PC_reg_9_7_inst : DFFR_X1 port map( D => target_PC_i(7), CK => 
                           net3671, RN => n83, Q => predict_PC_9_7_port, QN => 
                           net47370);
   predict_PC_reg_9_6_inst : DFFR_X1 port map( D => target_PC_i(6), CK => 
                           net3671, RN => n91, Q => predict_PC_9_6_port, QN => 
                           net47369);
   predict_PC_reg_9_5_inst : DFFR_X1 port map( D => target_PC_i(5), CK => 
                           net3671, RN => n90, Q => predict_PC_9_5_port, QN => 
                           net47368);
   predict_PC_reg_9_4_inst : DFFR_X1 port map( D => target_PC_i(4), CK => 
                           net3671, RN => n89, Q => predict_PC_9_4_port, QN => 
                           net47367);
   predict_PC_reg_9_3_inst : DFFR_X1 port map( D => target_PC_i(3), CK => 
                           net3671, RN => n88, Q => predict_PC_9_3_port, QN => 
                           net47366);
   predict_PC_reg_9_2_inst : DFFR_X1 port map( D => target_PC_i(2), CK => 
                           net3671, RN => n93, Q => predict_PC_9_2_port, QN => 
                           net47365);
   predict_PC_reg_9_1_inst : DFFR_X1 port map( D => target_PC_i(1), CK => 
                           net3671, RN => n92, Q => predict_PC_9_1_port, QN => 
                           net47364);
   predict_PC_reg_9_0_inst : DFFR_X1 port map( D => target_PC_i(0), CK => 
                           net3671, RN => n94, Q => predict_PC_9_0_port, QN => 
                           net47363);
   predict_PC_reg_10_31_inst : DFFR_X1 port map( D => n59, CK => net3676, RN =>
                           n88, Q => predict_PC_10_31_port, QN => net47362);
   predict_PC_reg_10_30_inst : DFFR_X1 port map( D => n38_port, CK => net3676, 
                           RN => n90, Q => predict_PC_10_30_port, QN => 
                           net47361);
   predict_PC_reg_10_29_inst : DFFR_X1 port map( D => n58, CK => net3676, RN =>
                           n100, Q => predict_PC_10_29_port, QN => net47360);
   predict_PC_reg_10_28_inst : DFFR_X1 port map( D => n39_port, CK => net3676, 
                           RN => n99, Q => predict_PC_10_28_port, QN => 
                           net47359);
   predict_PC_reg_10_27_inst : DFFR_X1 port map( D => target_PC_i(27), CK => 
                           net3676, RN => n96, Q => predict_PC_10_27_port, QN 
                           => net47358);
   predict_PC_reg_10_26_inst : DFFR_X1 port map( D => n37, CK => net3676, RN =>
                           n95, Q => predict_PC_10_26_port, QN => net47357);
   predict_PC_reg_10_25_inst : DFFR_X1 port map( D => n35, CK => net3676, RN =>
                           n81, Q => predict_PC_10_25_port, QN => net47356);
   predict_PC_reg_10_24_inst : DFFR_X1 port map( D => n36, CK => net3676, RN =>
                           n98, Q => predict_PC_10_24_port, QN => net47355);
   predict_PC_reg_10_23_inst : DFFR_X1 port map( D => target_PC_i(23), CK => 
                           net3676, RN => n97, Q => predict_PC_10_23_port, QN 
                           => net47354);
   predict_PC_reg_10_22_inst : DFFR_X1 port map( D => target_PC_i(22), CK => 
                           net3676, RN => n91, Q => predict_PC_10_22_port, QN 
                           => net47353);
   predict_PC_reg_10_21_inst : DFFR_X1 port map( D => target_PC_i(21), CK => 
                           net3676, RN => n90, Q => predict_PC_10_21_port, QN 
                           => net47352);
   predict_PC_reg_10_20_inst : DFFR_X1 port map( D => target_PC_i(20), CK => 
                           net3676, RN => n89, Q => predict_PC_10_20_port, QN 
                           => net47351);
   predict_PC_reg_10_19_inst : DFFR_X1 port map( D => target_PC_i(19), CK => 
                           net3676, RN => n88, Q => predict_PC_10_19_port, QN 
                           => net47350);
   predict_PC_reg_10_18_inst : DFFR_X1 port map( D => target_PC_i(18), CK => 
                           net3676, RN => n93, Q => predict_PC_10_18_port, QN 
                           => net47349);
   predict_PC_reg_10_17_inst : DFFR_X1 port map( D => target_PC_i(17), CK => 
                           net3676, RN => n92, Q => predict_PC_10_17_port, QN 
                           => net47348);
   predict_PC_reg_10_16_inst : DFFR_X1 port map( D => target_PC_i(16), CK => 
                           net3676, RN => n94, Q => predict_PC_10_16_port, QN 
                           => net47347);
   predict_PC_reg_10_15_inst : DFFR_X1 port map( D => target_PC_i(15), CK => 
                           net3676, RN => n85, Q => predict_PC_10_15_port, QN 
                           => net47346);
   predict_PC_reg_10_14_inst : DFFR_X1 port map( D => target_PC_i(14), CK => 
                           net3676, RN => n89, Q => predict_PC_10_14_port, QN 
                           => net47345);
   predict_PC_reg_10_13_inst : DFFR_X1 port map( D => target_PC_i(13), CK => 
                           net3676, RN => n89, Q => predict_PC_10_13_port, QN 
                           => net47344);
   predict_PC_reg_10_12_inst : DFFR_X1 port map( D => target_PC_i(12), CK => 
                           net3676, RN => n94, Q => predict_PC_10_12_port, QN 
                           => net47343);
   predict_PC_reg_10_11_inst : DFFR_X1 port map( D => target_PC_i(11), CK => 
                           net3676, RN => n99, Q => predict_PC_10_11_port, QN 
                           => net47342);
   predict_PC_reg_10_10_inst : DFFR_X1 port map( D => target_PC_i(10), CK => 
                           net3676, RN => n96, Q => predict_PC_10_10_port, QN 
                           => net47341);
   predict_PC_reg_10_9_inst : DFFR_X1 port map( D => target_PC_i(9), CK => 
                           net3676, RN => n88, Q => predict_PC_10_9_port, QN =>
                           net47340);
   predict_PC_reg_10_8_inst : DFFR_X1 port map( D => target_PC_i(8), CK => 
                           net3676, RN => n93, Q => predict_PC_10_8_port, QN =>
                           net47339);
   predict_PC_reg_10_7_inst : DFFR_X1 port map( D => target_PC_i(7), CK => 
                           net3676, RN => n98, Q => predict_PC_10_7_port, QN =>
                           net47338);
   predict_PC_reg_10_6_inst : DFFR_X1 port map( D => target_PC_i(6), CK => 
                           net3676, RN => n95, Q => predict_PC_10_6_port, QN =>
                           net47337);
   predict_PC_reg_10_5_inst : DFFR_X1 port map( D => target_PC_i(5), CK => 
                           net3676, RN => n100, Q => predict_PC_10_5_port, QN 
                           => net47336);
   predict_PC_reg_10_4_inst : DFFR_X1 port map( D => target_PC_i(4), CK => 
                           net3676, RN => n82, Q => predict_PC_10_4_port, QN =>
                           net47335);
   predict_PC_reg_10_3_inst : DFFR_X1 port map( D => target_PC_i(3), CK => 
                           net3676, RN => n82, Q => predict_PC_10_3_port, QN =>
                           net47334);
   predict_PC_reg_10_2_inst : DFFR_X1 port map( D => target_PC_i(2), CK => 
                           net3676, RN => n95, Q => predict_PC_10_2_port, QN =>
                           net47333);
   predict_PC_reg_10_1_inst : DFFR_X1 port map( D => target_PC_i(1), CK => 
                           net3676, RN => n84, Q => predict_PC_10_1_port, QN =>
                           net47332);
   predict_PC_reg_10_0_inst : DFFR_X1 port map( D => target_PC_i(0), CK => 
                           net3676, RN => n98, Q => predict_PC_10_0_port, QN =>
                           net47331);
   predict_PC_reg_11_31_inst : DFFR_X1 port map( D => n59, CK => net3681, RN =>
                           n97, Q => predict_PC_11_31_port, QN => net47330);
   predict_PC_reg_11_30_inst : DFFR_X1 port map( D => n38_port, CK => net3681, 
                           RN => n85, Q => predict_PC_11_30_port, QN => 
                           net47329);
   predict_PC_reg_11_29_inst : DFFR_X1 port map( D => n58, CK => net3681, RN =>
                           n87, Q => predict_PC_11_29_port, QN => net47328);
   predict_PC_reg_11_28_inst : DFFR_X1 port map( D => target_PC_i(28), CK => 
                           net3681, RN => n84, Q => predict_PC_11_28_port, QN 
                           => net47327);
   predict_PC_reg_11_27_inst : DFFR_X1 port map( D => target_PC_i(27), CK => 
                           net3681, RN => n91, Q => predict_PC_11_27_port, QN 
                           => net47326);
   predict_PC_reg_11_26_inst : DFFR_X1 port map( D => n37, CK => net3681, RN =>
                           n90, Q => predict_PC_11_26_port, QN => net47325);
   predict_PC_reg_11_25_inst : DFFR_X1 port map( D => target_PC_i(25), CK => 
                           net3681, RN => n92, Q => predict_PC_11_25_port, QN 
                           => net47324);
   predict_PC_reg_11_24_inst : DFFR_X1 port map( D => n36, CK => net3681, RN =>
                           n99, Q => predict_PC_11_24_port, QN => net47323);
   predict_PC_reg_11_23_inst : DFFR_X1 port map( D => target_PC_i(23), CK => 
                           net3681, RN => n96, Q => predict_PC_11_23_port, QN 
                           => net47322);
   predict_PC_reg_11_22_inst : DFFR_X1 port map( D => target_PC_i(22), CK => 
                           net3681, RN => n81, Q => predict_PC_11_22_port, QN 
                           => net47321);
   predict_PC_reg_11_21_inst : DFFR_X1 port map( D => target_PC_i(21), CK => 
                           net3681, RN => n81, Q => predict_PC_11_21_port, QN 
                           => net47320);
   predict_PC_reg_11_20_inst : DFFR_X1 port map( D => target_PC_i(20), CK => 
                           net3681, RN => n95, Q => predict_PC_11_20_port, QN 
                           => net47319);
   predict_PC_reg_11_19_inst : DFFR_X1 port map( D => target_PC_i(19), CK => 
                           net3681, RN => n80, Q => predict_PC_11_19_port, QN 
                           => net47318);
   predict_PC_reg_11_18_inst : DFFR_X1 port map( D => target_PC_i(18), CK => 
                           net3681, RN => n98, Q => predict_PC_11_18_port, QN 
                           => net47317);
   predict_PC_reg_11_17_inst : DFFR_X1 port map( D => target_PC_i(17), CK => 
                           net3681, RN => n97, Q => predict_PC_11_17_port, QN 
                           => net47316);
   predict_PC_reg_11_16_inst : DFFR_X1 port map( D => target_PC_i(16), CK => 
                           net3681, RN => n86_port, Q => predict_PC_11_16_port,
                           QN => net47315);
   predict_PC_reg_11_15_inst : DFFR_X1 port map( D => target_PC_i(15), CK => 
                           net3681, RN => n85, Q => predict_PC_11_15_port, QN 
                           => net47314);
   predict_PC_reg_11_14_inst : DFFR_X1 port map( D => target_PC_i(14), CK => 
                           net3681, RN => n87, Q => predict_PC_11_14_port, QN 
                           => net47313);
   predict_PC_reg_11_13_inst : DFFR_X1 port map( D => target_PC_i(13), CK => 
                           net3681, RN => n99, Q => predict_PC_11_13_port, QN 
                           => net47312);
   predict_PC_reg_11_12_inst : DFFR_X1 port map( D => target_PC_i(12), CK => 
                           net3681, RN => n99, Q => predict_PC_11_12_port, QN 
                           => net47311);
   predict_PC_reg_11_11_inst : DFFR_X1 port map( D => target_PC_i(11), CK => 
                           net3681, RN => n99, Q => predict_PC_11_11_port, QN 
                           => net47310);
   predict_PC_reg_11_10_inst : DFFR_X1 port map( D => target_PC_i(10), CK => 
                           net3681, RN => n99, Q => predict_PC_11_10_port, QN 
                           => net47309);
   predict_PC_reg_11_9_inst : DFFR_X1 port map( D => target_PC_i(9), CK => 
                           net3681, RN => n99, Q => predict_PC_11_9_port, QN =>
                           net47308);
   predict_PC_reg_11_8_inst : DFFR_X1 port map( D => target_PC_i(8), CK => 
                           net3681, RN => n99, Q => predict_PC_11_8_port, QN =>
                           net47307);
   predict_PC_reg_11_7_inst : DFFR_X1 port map( D => target_PC_i(7), CK => 
                           net3681, RN => n99, Q => predict_PC_11_7_port, QN =>
                           net47306);
   predict_PC_reg_11_6_inst : DFFR_X1 port map( D => target_PC_i(6), CK => 
                           net3681, RN => n99, Q => predict_PC_11_6_port, QN =>
                           net47305);
   predict_PC_reg_11_5_inst : DFFR_X1 port map( D => target_PC_i(5), CK => 
                           net3681, RN => n84, Q => predict_PC_11_5_port, QN =>
                           net47304);
   predict_PC_reg_11_4_inst : DFFR_X1 port map( D => target_PC_i(4), CK => 
                           net3681, RN => n99, Q => predict_PC_11_4_port, QN =>
                           net47303);
   predict_PC_reg_11_3_inst : DFFR_X1 port map( D => target_PC_i(3), CK => 
                           net3681, RN => n99, Q => predict_PC_11_3_port, QN =>
                           net47302);
   predict_PC_reg_11_2_inst : DFFR_X1 port map( D => target_PC_i(2), CK => 
                           net3681, RN => n99, Q => predict_PC_11_2_port, QN =>
                           net47301);
   predict_PC_reg_11_1_inst : DFFR_X1 port map( D => target_PC_i(1), CK => 
                           net3681, RN => n100, Q => predict_PC_11_1_port, QN 
                           => net47300);
   predict_PC_reg_11_0_inst : DFFR_X1 port map( D => target_PC_i(0), CK => 
                           net3681, RN => n100, Q => predict_PC_11_0_port, QN 
                           => net47299);
   predict_PC_reg_12_31_inst : DFFR_X1 port map( D => n59, CK => net3686, RN =>
                           n100, Q => predict_PC_12_31_port, QN => net47298);
   predict_PC_reg_12_30_inst : DFFR_X1 port map( D => n38_port, CK => net3686, 
                           RN => n100, Q => predict_PC_12_30_port, QN => 
                           net47297);
   predict_PC_reg_12_29_inst : DFFR_X1 port map( D => n58, CK => net3686, RN =>
                           n100, Q => predict_PC_12_29_port, QN => net47296);
   predict_PC_reg_12_28_inst : DFFR_X1 port map( D => n39_port, CK => net3686, 
                           RN => n100, Q => predict_PC_12_28_port, QN => 
                           net47295);
   predict_PC_reg_12_27_inst : DFFR_X1 port map( D => target_PC_i(27), CK => 
                           net3686, RN => n100, Q => predict_PC_12_27_port, QN 
                           => net47294);
   predict_PC_reg_12_26_inst : DFFR_X1 port map( D => n37, CK => net3686, RN =>
                           n100, Q => predict_PC_12_26_port, QN => net47293);
   predict_PC_reg_12_25_inst : DFFR_X1 port map( D => n35, CK => net3686, RN =>
                           n100, Q => predict_PC_12_25_port, QN => net47292);
   predict_PC_reg_12_24_inst : DFFR_X1 port map( D => n36, CK => net3686, RN =>
                           n100, Q => predict_PC_12_24_port, QN => net47291);
   predict_PC_reg_12_23_inst : DFFR_X1 port map( D => target_PC_i(23), CK => 
                           net3686, RN => n99, Q => predict_PC_12_23_port, QN 
                           => net47290);
   predict_PC_reg_12_22_inst : DFFR_X1 port map( D => target_PC_i(22), CK => 
                           net3686, RN => n100, Q => predict_PC_12_22_port, QN 
                           => net47289);
   predict_PC_reg_12_21_inst : DFFR_X1 port map( D => target_PC_i(21), CK => 
                           net3686, RN => n79, Q => predict_PC_12_21_port, QN 
                           => net47288);
   predict_PC_reg_12_20_inst : DFFR_X1 port map( D => target_PC_i(20), CK => 
                           net3686, RN => n79, Q => predict_PC_12_20_port, QN 
                           => net47287);
   predict_PC_reg_12_19_inst : DFFR_X1 port map( D => target_PC_i(19), CK => 
                           net3686, RN => n78, Q => predict_PC_12_19_port, QN 
                           => net47286);
   predict_PC_reg_12_18_inst : DFFR_X1 port map( D => target_PC_i(18), CK => 
                           net3686, RN => n78, Q => predict_PC_12_18_port, QN 
                           => net47285);
   predict_PC_reg_12_17_inst : DFFR_X1 port map( D => target_PC_i(17), CK => 
                           net3686, RN => n79, Q => predict_PC_12_17_port, QN 
                           => net47284);
   predict_PC_reg_12_16_inst : DFFR_X1 port map( D => target_PC_i(16), CK => 
                           net3686, RN => n77, Q => predict_PC_12_16_port, QN 
                           => net47283);
   predict_PC_reg_12_15_inst : DFFR_X1 port map( D => target_PC_i(15), CK => 
                           net3686, RN => n77, Q => predict_PC_12_15_port, QN 
                           => net47282);
   predict_PC_reg_12_14_inst : DFFR_X1 port map( D => target_PC_i(14), CK => 
                           net3686, RN => n77, Q => predict_PC_12_14_port, QN 
                           => net47281);
   predict_PC_reg_12_13_inst : DFFR_X1 port map( D => target_PC_i(13), CK => 
                           net3686, RN => n78, Q => predict_PC_12_13_port, QN 
                           => net47280);
   predict_PC_reg_12_12_inst : DFFR_X1 port map( D => target_PC_i(12), CK => 
                           net3686, RN => n79, Q => predict_PC_12_12_port, QN 
                           => net47279);
   predict_PC_reg_12_11_inst : DFFR_X1 port map( D => target_PC_i(11), CK => 
                           net3686, RN => n100, Q => predict_PC_12_11_port, QN 
                           => net47278);
   predict_PC_reg_12_10_inst : DFFR_X1 port map( D => target_PC_i(10), CK => 
                           net3686, RN => n99, Q => predict_PC_12_10_port, QN 
                           => net47277);
   predict_PC_reg_12_9_inst : DFFR_X1 port map( D => target_PC_i(9), CK => 
                           net3686, RN => n93, Q => predict_PC_12_9_port, QN =>
                           net47276);
   predict_PC_reg_12_8_inst : DFFR_X1 port map( D => target_PC_i(8), CK => 
                           net3686, RN => n93, Q => predict_PC_12_8_port, QN =>
                           net47275);
   predict_PC_reg_12_7_inst : DFFR_X1 port map( D => target_PC_i(7), CK => 
                           net3686, RN => n93, Q => predict_PC_12_7_port, QN =>
                           net47274);
   predict_PC_reg_12_6_inst : DFFR_X1 port map( D => target_PC_i(6), CK => 
                           net3686, RN => n93, Q => predict_PC_12_6_port, QN =>
                           net47273);
   predict_PC_reg_12_5_inst : DFFR_X1 port map( D => target_PC_i(5), CK => 
                           net3686, RN => n93, Q => predict_PC_12_5_port, QN =>
                           net47272);
   predict_PC_reg_12_4_inst : DFFR_X1 port map( D => target_PC_i(4), CK => 
                           net3686, RN => n93, Q => predict_PC_12_4_port, QN =>
                           net47271);
   predict_PC_reg_12_3_inst : DFFR_X1 port map( D => target_PC_i(3), CK => 
                           net3686, RN => n94, Q => predict_PC_12_3_port, QN =>
                           net47270);
   predict_PC_reg_12_2_inst : DFFR_X1 port map( D => target_PC_i(2), CK => 
                           net3686, RN => n94, Q => predict_PC_12_2_port, QN =>
                           net47269);
   predict_PC_reg_12_1_inst : DFFR_X1 port map( D => target_PC_i(1), CK => 
                           net3686, RN => n94, Q => predict_PC_12_1_port, QN =>
                           net47268);
   predict_PC_reg_12_0_inst : DFFR_X1 port map( D => target_PC_i(0), CK => 
                           net3686, RN => n94, Q => predict_PC_12_0_port, QN =>
                           net47267);
   predict_PC_reg_13_31_inst : DFFR_X1 port map( D => n59, CK => net3691, RN =>
                           n94, Q => predict_PC_13_31_port, QN => net47266);
   predict_PC_reg_13_30_inst : DFFR_X1 port map( D => n38_port, CK => net3691, 
                           RN => n94, Q => predict_PC_13_30_port, QN => 
                           net47265);
   predict_PC_reg_13_29_inst : DFFR_X1 port map( D => n58, CK => net3691, RN =>
                           n94, Q => predict_PC_13_29_port, QN => net47264);
   predict_PC_reg_13_28_inst : DFFR_X1 port map( D => n39_port, CK => net3691, 
                           RN => n94, Q => predict_PC_13_28_port, QN => 
                           net47263);
   predict_PC_reg_13_27_inst : DFFR_X1 port map( D => n60, CK => net3691, RN =>
                           n94, Q => predict_PC_13_27_port, QN => net47262);
   predict_PC_reg_13_26_inst : DFFR_X1 port map( D => n37, CK => net3691, RN =>
                           n94, Q => predict_PC_13_26_port, QN => net47261);
   predict_PC_reg_13_25_inst : DFFR_X1 port map( D => n35, CK => net3691, RN =>
                           n94, Q => predict_PC_13_25_port, QN => net47260);
   predict_PC_reg_13_24_inst : DFFR_X1 port map( D => n36, CK => net3691, RN =>
                           n94, Q => predict_PC_13_24_port, QN => net47259);
   predict_PC_reg_13_23_inst : DFFR_X1 port map( D => target_PC_i(23), CK => 
                           net3691, RN => n90, Q => predict_PC_13_23_port, QN 
                           => net47258);
   predict_PC_reg_13_22_inst : DFFR_X1 port map( D => target_PC_i(22), CK => 
                           net3691, RN => n92, Q => predict_PC_13_22_port, QN 
                           => net47257);
   predict_PC_reg_13_21_inst : DFFR_X1 port map( D => target_PC_i(21), CK => 
                           net3691, RN => n94, Q => predict_PC_13_21_port, QN 
                           => net47256);
   predict_PC_reg_13_20_inst : DFFR_X1 port map( D => target_PC_i(20), CK => 
                           net3691, RN => n100, Q => predict_PC_13_20_port, QN 
                           => net47255);
   predict_PC_reg_13_19_inst : DFFR_X1 port map( D => target_PC_i(19), CK => 
                           net3691, RN => n99, Q => predict_PC_13_19_port, QN 
                           => net47254);
   predict_PC_reg_13_18_inst : DFFR_X1 port map( D => target_PC_i(18), CK => 
                           net3691, RN => n96, Q => predict_PC_13_18_port, QN 
                           => net47253);
   predict_PC_reg_13_17_inst : DFFR_X1 port map( D => target_PC_i(17), CK => 
                           net3691, RN => n84, Q => predict_PC_13_17_port, QN 
                           => net47252);
   predict_PC_reg_13_16_inst : DFFR_X1 port map( D => target_PC_i(16), CK => 
                           net3691, RN => n84, Q => predict_PC_13_16_port, QN 
                           => net47251);
   predict_PC_reg_13_15_inst : DFFR_X1 port map( D => target_PC_i(15), CK => 
                           net3691, RN => n95, Q => predict_PC_13_15_port, QN 
                           => net47250);
   predict_PC_reg_13_14_inst : DFFR_X1 port map( D => target_PC_i(14), CK => 
                           net3691, RN => n98, Q => predict_PC_13_14_port, QN 
                           => net47249);
   predict_PC_reg_13_13_inst : DFFR_X1 port map( D => target_PC_i(13), CK => 
                           net3691, RN => n97, Q => predict_PC_13_13_port, QN 
                           => net47248);
   predict_PC_reg_13_12_inst : DFFR_X1 port map( D => target_PC_i(12), CK => 
                           net3691, RN => n86_port, Q => predict_PC_13_12_port,
                           QN => net47247);
   predict_PC_reg_13_11_inst : DFFR_X1 port map( D => target_PC_i(11), CK => 
                           net3691, RN => n95, Q => predict_PC_13_11_port, QN 
                           => net47246);
   predict_PC_reg_13_10_inst : DFFR_X1 port map( D => target_PC_i(10), CK => 
                           net3691, RN => n95, Q => predict_PC_13_10_port, QN 
                           => net47245);
   predict_PC_reg_13_9_inst : DFFR_X1 port map( D => target_PC_i(9), CK => 
                           net3691, RN => n95, Q => predict_PC_13_9_port, QN =>
                           net47244);
   predict_PC_reg_13_8_inst : DFFR_X1 port map( D => target_PC_i(8), CK => 
                           net3691, RN => n95, Q => predict_PC_13_8_port, QN =>
                           net47243);
   predict_PC_reg_13_7_inst : DFFR_X1 port map( D => target_PC_i(7), CK => 
                           net3691, RN => n95, Q => predict_PC_13_7_port, QN =>
                           net47242);
   predict_PC_reg_13_6_inst : DFFR_X1 port map( D => target_PC_i(6), CK => 
                           net3691, RN => n95, Q => predict_PC_13_6_port, QN =>
                           net47241);
   predict_PC_reg_13_5_inst : DFFR_X1 port map( D => target_PC_i(5), CK => 
                           net3691, RN => n95, Q => predict_PC_13_5_port, QN =>
                           net47240);
   predict_PC_reg_13_4_inst : DFFR_X1 port map( D => target_PC_i(4), CK => 
                           net3691, RN => n95, Q => predict_PC_13_4_port, QN =>
                           net47239);
   predict_PC_reg_13_3_inst : DFFR_X1 port map( D => target_PC_i(3), CK => 
                           net3691, RN => n95, Q => predict_PC_13_3_port, QN =>
                           net47238);
   predict_PC_reg_13_2_inst : DFFR_X1 port map( D => target_PC_i(2), CK => 
                           net3691, RN => n95, Q => predict_PC_13_2_port, QN =>
                           net47237);
   predict_PC_reg_13_1_inst : DFFR_X1 port map( D => target_PC_i(1), CK => 
                           net3691, RN => n95, Q => predict_PC_13_1_port, QN =>
                           net47236);
   predict_PC_reg_13_0_inst : DFFR_X1 port map( D => target_PC_i(0), CK => 
                           net3691, RN => n95, Q => predict_PC_13_0_port, QN =>
                           net47235);
   predict_PC_reg_14_31_inst : DFFR_X1 port map( D => n59, CK => net3696, RN =>
                           n95, Q => predict_PC_14_31_port, QN => net47234);
   predict_PC_reg_14_30_inst : DFFR_X1 port map( D => n38_port, CK => net3696, 
                           RN => n98, Q => predict_PC_14_30_port, QN => 
                           net47233);
   predict_PC_reg_14_29_inst : DFFR_X1 port map( D => n58, CK => net3696, RN =>
                           n91, Q => predict_PC_14_29_port, QN => net47232);
   predict_PC_reg_14_28_inst : DFFR_X1 port map( D => n39_port, CK => net3696, 
                           RN => n89, Q => predict_PC_14_28_port, QN => 
                           net47231);
   predict_PC_reg_14_27_inst : DFFR_X1 port map( D => n60, CK => net3696, RN =>
                           n88, Q => predict_PC_14_27_port, QN => net47230);
   predict_PC_reg_14_26_inst : DFFR_X1 port map( D => n37, CK => net3696, RN =>
                           n93, Q => predict_PC_14_26_port, QN => net47229);
   predict_PC_reg_14_25_inst : DFFR_X1 port map( D => n35, CK => net3696, RN =>
                           n92, Q => predict_PC_14_25_port, QN => net47228);
   predict_PC_reg_14_24_inst : DFFR_X1 port map( D => n36, CK => net3696, RN =>
                           n94, Q => predict_PC_14_24_port, QN => net47227);
   predict_PC_reg_14_23_inst : DFFR_X1 port map( D => target_PC_i(23), CK => 
                           net3696, RN => n100, Q => predict_PC_14_23_port, QN 
                           => net47226);
   predict_PC_reg_14_22_inst : DFFR_X1 port map( D => target_PC_i(22), CK => 
                           net3696, RN => n99, Q => predict_PC_14_22_port, QN 
                           => net47225);
   predict_PC_reg_14_21_inst : DFFR_X1 port map( D => target_PC_i(21), CK => 
                           net3696, RN => n96, Q => predict_PC_14_21_port, QN 
                           => net47224);
   predict_PC_reg_14_20_inst : DFFR_X1 port map( D => target_PC_i(20), CK => 
                           net3696, RN => n91, Q => predict_PC_14_20_port, QN 
                           => net47223);
   predict_PC_reg_14_19_inst : DFFR_X1 port map( D => target_PC_i(19), CK => 
                           net3696, RN => n90, Q => predict_PC_14_19_port, QN 
                           => net47222);
   predict_PC_reg_14_18_inst : DFFR_X1 port map( D => target_PC_i(18), CK => 
                           net3696, RN => n90, Q => predict_PC_14_18_port, QN 
                           => net47221);
   predict_PC_reg_14_17_inst : DFFR_X1 port map( D => target_PC_i(17), CK => 
                           net3696, RN => n89, Q => predict_PC_14_17_port, QN 
                           => net47220);
   predict_PC_reg_14_16_inst : DFFR_X1 port map( D => target_PC_i(16), CK => 
                           net3696, RN => n88, Q => predict_PC_14_16_port, QN 
                           => net47219);
   predict_PC_reg_14_15_inst : DFFR_X1 port map( D => target_PC_i(15), CK => 
                           net3696, RN => n93, Q => predict_PC_14_15_port, QN 
                           => net47218);
   predict_PC_reg_14_14_inst : DFFR_X1 port map( D => target_PC_i(14), CK => 
                           net3696, RN => n92, Q => predict_PC_14_14_port, QN 
                           => net47217);
   predict_PC_reg_14_13_inst : DFFR_X1 port map( D => target_PC_i(13), CK => 
                           net3696, RN => n94, Q => predict_PC_14_13_port, QN 
                           => net47216);
   predict_PC_reg_14_12_inst : DFFR_X1 port map( D => target_PC_i(12), CK => 
                           net3696, RN => n100, Q => predict_PC_14_12_port, QN 
                           => net47215);
   predict_PC_reg_14_11_inst : DFFR_X1 port map( D => target_PC_i(11), CK => 
                           net3696, RN => n99, Q => predict_PC_14_11_port, QN 
                           => net47214);
   predict_PC_reg_14_10_inst : DFFR_X1 port map( D => target_PC_i(10), CK => 
                           net3696, RN => n96, Q => predict_PC_14_10_port, QN 
                           => net47213);
   predict_PC_reg_14_9_inst : DFFR_X1 port map( D => target_PC_i(9), CK => 
                           net3696, RN => n95, Q => predict_PC_14_9_port, QN =>
                           net47212);
   predict_PC_reg_14_8_inst : DFFR_X1 port map( D => target_PC_i(8), CK => 
                           net3696, RN => n98, Q => predict_PC_14_8_port, QN =>
                           net47211);
   predict_PC_reg_14_7_inst : DFFR_X1 port map( D => target_PC_i(7), CK => 
                           net3696, RN => n93, Q => predict_PC_14_7_port, QN =>
                           net47210);
   predict_PC_reg_14_6_inst : DFFR_X1 port map( D => target_PC_i(6), CK => 
                           net3696, RN => n94, Q => predict_PC_14_6_port, QN =>
                           net47209);
   predict_PC_reg_14_5_inst : DFFR_X1 port map( D => target_PC_i(5), CK => 
                           net3696, RN => n100, Q => predict_PC_14_5_port, QN 
                           => net47208);
   predict_PC_reg_14_4_inst : DFFR_X1 port map( D => target_PC_i(4), CK => 
                           net3696, RN => n96, Q => predict_PC_14_4_port, QN =>
                           net47207);
   predict_PC_reg_14_3_inst : DFFR_X1 port map( D => target_PC_i(3), CK => 
                           net3696, RN => n91, Q => predict_PC_14_3_port, QN =>
                           net47206);
   predict_PC_reg_14_2_inst : DFFR_X1 port map( D => target_PC_i(2), CK => 
                           net3696, RN => n80, Q => predict_PC_14_2_port, QN =>
                           net47205);
   predict_PC_reg_14_1_inst : DFFR_X1 port map( D => target_PC_i(1), CK => 
                           net3696, RN => n80, Q => predict_PC_14_1_port, QN =>
                           net47204);
   predict_PC_reg_14_0_inst : DFFR_X1 port map( D => target_PC_i(0), CK => 
                           net3696, RN => n95, Q => predict_PC_14_0_port, QN =>
                           net47203);
   predict_PC_reg_15_31_inst : DFFR_X1 port map( D => n59, CK => net3701, RN =>
                           n91, Q => predict_PC_15_31_port, QN => net47202);
   predict_PC_reg_15_30_inst : DFFR_X1 port map( D => n38_port, CK => net3701, 
                           RN => n98, Q => predict_PC_15_30_port, QN => 
                           net47201);
   predict_PC_reg_15_29_inst : DFFR_X1 port map( D => n58, CK => net3701, RN =>
                           n97, Q => predict_PC_15_29_port, QN => net47200);
   predict_PC_reg_15_28_inst : DFFR_X1 port map( D => n39_port, CK => net3701, 
                           RN => n94, Q => predict_PC_15_28_port, QN => 
                           net47199);
   predict_PC_reg_15_27_inst : DFFR_X1 port map( D => n60, CK => net3701, RN =>
                           n91, Q => predict_PC_15_27_port, QN => net47198);
   predict_PC_reg_15_26_inst : DFFR_X1 port map( D => n37, CK => net3701, RN =>
                           n100, Q => predict_PC_15_26_port, QN => net47197);
   predict_PC_reg_15_25_inst : DFFR_X1 port map( D => n35, CK => net3701, RN =>
                           n99, Q => predict_PC_15_25_port, QN => net47196);
   predict_PC_reg_15_24_inst : DFFR_X1 port map( D => n36, CK => net3701, RN =>
                           n89, Q => predict_PC_15_24_port, QN => net47195);
   predict_PC_reg_15_23_inst : DFFR_X1 port map( D => target_PC_i(23), CK => 
                           net3701, RN => n97, Q => predict_PC_15_23_port, QN 
                           => net47194);
   predict_PC_reg_15_22_inst : DFFR_X1 port map( D => target_PC_i(22), CK => 
                           net3701, RN => n88, Q => predict_PC_15_22_port, QN 
                           => net47193);
   predict_PC_reg_15_21_inst : DFFR_X1 port map( D => target_PC_i(21), CK => 
                           net3701, RN => n100, Q => predict_PC_15_21_port, QN 
                           => net47192);
   predict_PC_reg_15_20_inst : DFFR_X1 port map( D => target_PC_i(20), CK => 
                           net3701, RN => n88, Q => predict_PC_15_20_port, QN 
                           => net47191);
   predict_PC_reg_15_19_inst : DFFR_X1 port map( D => target_PC_i(19), CK => 
                           net3701, RN => n96, Q => predict_PC_15_19_port, QN 
                           => net47190);
   predict_PC_reg_15_18_inst : DFFR_X1 port map( D => target_PC_i(18), CK => 
                           net3701, RN => n93, Q => predict_PC_15_18_port, QN 
                           => net47189);
   predict_PC_reg_15_17_inst : DFFR_X1 port map( D => target_PC_i(17), CK => 
                           net3701, RN => n96, Q => predict_PC_15_17_port, QN 
                           => net47188);
   predict_PC_reg_15_16_inst : DFFR_X1 port map( D => target_PC_i(16), CK => 
                           net3701, RN => n91, Q => predict_PC_15_16_port, QN 
                           => net47187);
   predict_PC_reg_15_15_inst : DFFR_X1 port map( D => target_PC_i(15), CK => 
                           net3701, RN => n90, Q => predict_PC_15_15_port, QN 
                           => net47186);
   predict_PC_reg_15_14_inst : DFFR_X1 port map( D => target_PC_i(14), CK => 
                           net3701, RN => n89, Q => predict_PC_15_14_port, QN 
                           => net47185);
   predict_PC_reg_15_13_inst : DFFR_X1 port map( D => target_PC_i(13), CK => 
                           net3701, RN => n88, Q => predict_PC_15_13_port, QN 
                           => net47184);
   predict_PC_reg_15_12_inst : DFFR_X1 port map( D => target_PC_i(12), CK => 
                           net3701, RN => n93, Q => predict_PC_15_12_port, QN 
                           => net47183);
   predict_PC_reg_15_11_inst : DFFR_X1 port map( D => target_PC_i(11), CK => 
                           net3701, RN => n92, Q => predict_PC_15_11_port, QN 
                           => net47182);
   predict_PC_reg_15_10_inst : DFFR_X1 port map( D => target_PC_i(10), CK => 
                           net3701, RN => n96, Q => predict_PC_15_10_port, QN 
                           => net47181);
   predict_PC_reg_15_9_inst : DFFR_X1 port map( D => target_PC_i(9), CK => 
                           net3701, RN => n98, Q => predict_PC_15_9_port, QN =>
                           net47180);
   predict_PC_reg_15_8_inst : DFFR_X1 port map( D => target_PC_i(8), CK => 
                           net3701, RN => n85, Q => predict_PC_15_8_port, QN =>
                           net47179);
   predict_PC_reg_15_7_inst : DFFR_X1 port map( D => target_PC_i(7), CK => 
                           net3701, RN => n85, Q => predict_PC_15_7_port, QN =>
                           net47178);
   predict_PC_reg_15_6_inst : DFFR_X1 port map( D => target_PC_i(6), CK => 
                           net3701, RN => n95, Q => predict_PC_15_6_port, QN =>
                           net47177);
   predict_PC_reg_15_5_inst : DFFR_X1 port map( D => target_PC_i(5), CK => 
                           net3701, RN => n96, Q => predict_PC_15_5_port, QN =>
                           net47176);
   predict_PC_reg_15_4_inst : DFFR_X1 port map( D => target_PC_i(4), CK => 
                           net3701, RN => n96, Q => predict_PC_15_4_port, QN =>
                           net47175);
   predict_PC_reg_15_3_inst : DFFR_X1 port map( D => target_PC_i(3), CK => 
                           net3701, RN => n96, Q => predict_PC_15_3_port, QN =>
                           net47174);
   predict_PC_reg_15_2_inst : DFFR_X1 port map( D => target_PC_i(2), CK => 
                           net3701, RN => n96, Q => predict_PC_15_2_port, QN =>
                           net47173);
   predict_PC_reg_15_1_inst : DFFR_X1 port map( D => target_PC_i(1), CK => 
                           net3701, RN => n96, Q => predict_PC_15_1_port, QN =>
                           net47172);
   predict_PC_reg_15_0_inst : DFFR_X1 port map( D => target_PC_i(0), CK => 
                           net3701, RN => n96, Q => predict_PC_15_0_port, QN =>
                           net47171);
   pred_x_0 : predictor_2_0 port map( clock => clock, reset => reset, enable =>
                           write_enable_0_port, taken_i => was_taken_i, 
                           prediction_o => taken_0_port);
   pred_x_1 : predictor_2_15 port map( clock => clock, reset => reset, enable 
                           => write_enable_1_port, taken_i => was_taken_i, 
                           prediction_o => taken_1_port);
   pred_x_2 : predictor_2_14 port map( clock => clock, reset => reset, enable 
                           => write_enable_2_port, taken_i => was_taken_i, 
                           prediction_o => taken_2_port);
   pred_x_3 : predictor_2_13 port map( clock => clock, reset => reset, enable 
                           => write_enable_3_port, taken_i => was_taken_i, 
                           prediction_o => taken_3_port);
   pred_x_4 : predictor_2_12 port map( clock => clock, reset => reset, enable 
                           => write_enable_4_port, taken_i => was_taken_i, 
                           prediction_o => taken_4_port);
   pred_x_5 : predictor_2_11 port map( clock => clock, reset => reset, enable 
                           => write_enable_5_port, taken_i => was_taken_i, 
                           prediction_o => taken_5_port);
   pred_x_6 : predictor_2_10 port map( clock => clock, reset => reset, enable 
                           => write_enable_6_port, taken_i => was_taken_i, 
                           prediction_o => taken_6_port);
   pred_x_7 : predictor_2_9 port map( clock => clock, reset => reset, enable =>
                           write_enable_7_port, taken_i => was_taken_i, 
                           prediction_o => taken_7_port);
   pred_x_8 : predictor_2_8 port map( clock => clock, reset => reset, enable =>
                           write_enable_8_port, taken_i => was_taken_i, 
                           prediction_o => taken_8_port);
   pred_x_9 : predictor_2_7 port map( clock => clock, reset => reset, enable =>
                           write_enable_9_port, taken_i => was_taken_i, 
                           prediction_o => taken_9_port);
   pred_x_10 : predictor_2_6 port map( clock => clock, reset => reset, enable 
                           => write_enable_10_port, taken_i => was_taken_i, 
                           prediction_o => taken_10_port);
   pred_x_11 : predictor_2_5 port map( clock => clock, reset => reset, enable 
                           => write_enable_11_port, taken_i => was_taken_i, 
                           prediction_o => taken_11_port);
   pred_x_12 : predictor_2_4 port map( clock => clock, reset => reset, enable 
                           => write_enable_12_port, taken_i => was_taken_i, 
                           prediction_o => taken_12_port);
   pred_x_13 : predictor_2_3 port map( clock => clock, reset => reset, enable 
                           => write_enable_13_port, taken_i => was_taken_i, 
                           prediction_o => taken_13_port);
   pred_x_14 : predictor_2_2 port map( clock => clock, reset => reset, enable 
                           => write_enable_14_port, taken_i => was_taken_i, 
                           prediction_o => taken_14_port);
   pred_x_15 : predictor_2_1 port map( clock => clock, reset => reset, enable 
                           => write_enable_15_port, taken_i => was_taken_i, 
                           prediction_o => taken_15_port);
   clk_gate_last_TAG_reg : SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_0 port map(
                           CLK => clock, EN => N567, ENCLK => net3621);
   clk_gate_predict_PC_reg_0_inst : SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_16
                           port map( CLK => clock, EN => N566, ENCLK => net3626
                           );
   clk_gate_predict_PC_reg_1_inst : SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_15
                           port map( CLK => clock, EN => N534, ENCLK => net3631
                           );
   clk_gate_predict_PC_reg_2_inst : SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_14
                           port map( CLK => clock, EN => N502, ENCLK => net3636
                           );
   clk_gate_predict_PC_reg_3_inst : SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_13
                           port map( CLK => clock, EN => N470, ENCLK => net3641
                           );
   clk_gate_predict_PC_reg_4_inst : SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_12
                           port map( CLK => clock, EN => N438, ENCLK => net3646
                           );
   clk_gate_predict_PC_reg_5_inst : SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_11
                           port map( CLK => clock, EN => N406, ENCLK => net3651
                           );
   clk_gate_predict_PC_reg_6_inst : SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_10
                           port map( CLK => clock, EN => N374, ENCLK => net3656
                           );
   clk_gate_predict_PC_reg_7_inst : SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_9 
                           port map( CLK => clock, EN => N342, ENCLK => net3661
                           );
   clk_gate_predict_PC_reg_8_inst : SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_8 
                           port map( CLK => clock, EN => N310, ENCLK => net3666
                           );
   clk_gate_predict_PC_reg_9_inst : SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_7 
                           port map( CLK => clock, EN => N278, ENCLK => net3671
                           );
   clk_gate_predict_PC_reg_10_inst : SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_6
                           port map( CLK => clock, EN => N246, ENCLK => net3676
                           );
   clk_gate_predict_PC_reg_11_inst : SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_5
                           port map( CLK => clock, EN => N214, ENCLK => net3681
                           );
   clk_gate_predict_PC_reg_12_inst : SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_4
                           port map( CLK => clock, EN => N182, ENCLK => net3686
                           );
   clk_gate_predict_PC_reg_13_inst : SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_3
                           port map( CLK => clock, EN => N150, ENCLK => net3691
                           );
   clk_gate_predict_PC_reg_14_inst : SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_2
                           port map( CLK => clock, EN => N118, ENCLK => net3696
                           );
   clk_gate_predict_PC_reg_15_inst : SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_1
                           port map( CLK => clock, EN => N86, ENCLK => net3701)
                           ;
   U391 : NAND2_X1 port map( A1 => TAG_i(1), A2 => n903, ZN => n895);
   U390 : NAND2_X1 port map( A1 => TAG_i(3), A2 => n973, ZN => n902);
   U386 : AOI22_X1 port map( A1 => n557, A2 => taken_10_port, B1 => n558, B2 =>
                           taken_11_port, ZN => n897);
   U381 : AOI22_X1 port map( A1 => n559, A2 => taken_8_port, B1 => n69, B2 => 
                           taken_9_port, ZN => n898);
   U380 : NAND2_X1 port map( A1 => TAG_i(2), A2 => TAG_i(3), ZN => n901);
   U377 : AOI22_X1 port map( A1 => n553, A2 => taken_14_port, B1 => n554, B2 =>
                           taken_15_port, ZN => n899);
   U374 : AOI22_X1 port map( A1 => n555, A2 => taken_12_port, B1 => n556, B2 =>
                           taken_13_port, ZN => n900);
   U369 : AOI22_X1 port map( A1 => n64, A2 => taken_2_port, B1 => n63, B2 => 
                           taken_3_port, ZN => n887);
   U366 : AOI22_X1 port map( A1 => n62, A2 => taken_0_port, B1 => n61, B2 => 
                           taken_1_port, ZN => n888);
   U365 : NAND2_X1 port map( A1 => TAG_i(2), A2 => n972, ZN => n892);
   U362 : AOI22_X1 port map( A1 => n68, A2 => taken_6_port, B1 => n67, B2 => 
                           taken_7_port, ZN => n889);
   U359 : AOI22_X1 port map( A1 => n66, A2 => taken_4_port, B1 => n65, B2 => 
                           taken_5_port, ZN => n890);
   U430 : OAI22_X1 port map( A1 => target_PC_i(17), A2 => n511, B1 => 
                           target_PC_i(16), B2 => n513, ZN => n940);
   U429 : AOI221_X1 port map( B1 => target_PC_i(17), B2 => n511, C1 => n513, C2
                           => target_PC_i(16), A => n940, ZN => n937);
   U428 : OAI22_X1 port map( A1 => target_PC_i(11), A2 => n523, B1 => 
                           target_PC_i(10), B2 => n525, ZN => n939);
   U188 : AOI22_X1 port map( A1 => n62, A2 => predict_PC_0_23_port, B1 => n61, 
                           B2 => predict_PC_1_23_port, ZN => n729);
   U187 : AOI22_X1 port map( A1 => n64, A2 => predict_PC_2_23_port, B1 => n63, 
                           B2 => predict_PC_3_23_port, ZN => n730);
   U186 : AOI22_X1 port map( A1 => n66, A2 => predict_PC_4_23_port, B1 => n65, 
                           B2 => predict_PC_5_23_port, ZN => n731);
   U185 : AOI22_X1 port map( A1 => n68, A2 => predict_PC_6_23_port, B1 => n67, 
                           B2 => predict_PC_7_23_port, ZN => n732);
   U184 : NAND4_X1 port map( A1 => n729, A2 => n730, A3 => n731, A4 => n732, ZN
                           => n723);
   U183 : AOI22_X1 port map( A1 => n70, A2 => predict_PC_8_23_port, B1 => n69, 
                           B2 => predict_PC_9_23_port, ZN => n725);
   U182 : AOI22_X1 port map( A1 => n72, A2 => predict_PC_10_23_port, B1 => n71,
                           B2 => predict_PC_11_23_port, ZN => n726);
   U181 : AOI22_X1 port map( A1 => n74, A2 => predict_PC_12_23_port, B1 => n73,
                           B2 => predict_PC_13_23_port, ZN => n727);
   U180 : AOI22_X1 port map( A1 => n76, A2 => predict_PC_14_23_port, B1 => n75,
                           B2 => predict_PC_15_23_port, ZN => n728);
   U179 : NAND4_X1 port map( A1 => n725, A2 => n726, A3 => n727, A4 => n728, ZN
                           => n724);
   U133 : AOI22_X1 port map( A1 => n62, A2 => predict_PC_0_28_port, B1 => n61, 
                           B2 => predict_PC_1_28_port, ZN => n679);
   U132 : AOI22_X1 port map( A1 => n64, A2 => predict_PC_2_28_port, B1 => n63, 
                           B2 => predict_PC_3_28_port, ZN => n680);
   U131 : AOI22_X1 port map( A1 => n66, A2 => predict_PC_4_28_port, B1 => n65, 
                           B2 => predict_PC_5_28_port, ZN => n681);
   U130 : AOI22_X1 port map( A1 => n68, A2 => predict_PC_6_28_port, B1 => n67, 
                           B2 => predict_PC_7_28_port, ZN => n682);
   U129 : NAND4_X1 port map( A1 => n679, A2 => n680, A3 => n681, A4 => n682, ZN
                           => n673);
   U128 : AOI22_X1 port map( A1 => n70, A2 => predict_PC_8_28_port, B1 => n69, 
                           B2 => predict_PC_9_28_port, ZN => n675);
   U127 : AOI22_X1 port map( A1 => n72, A2 => predict_PC_10_28_port, B1 => n71,
                           B2 => predict_PC_11_28_port, ZN => n676);
   U126 : AOI22_X1 port map( A1 => n74, A2 => predict_PC_12_28_port, B1 => n73,
                           B2 => predict_PC_13_28_port, ZN => n677);
   U125 : AOI22_X1 port map( A1 => n76, A2 => predict_PC_14_28_port, B1 => n75,
                           B2 => predict_PC_15_28_port, ZN => n678);
   U124 : NAND4_X1 port map( A1 => n675, A2 => n676, A3 => n677, A4 => n678, ZN
                           => n674);
   U111 : AOI22_X1 port map( A1 => n62, A2 => predict_PC_0_2_port, B1 => n61, 
                           B2 => predict_PC_1_2_port, ZN => n659);
   U110 : AOI22_X1 port map( A1 => n64, A2 => predict_PC_2_2_port, B1 => n63, 
                           B2 => predict_PC_3_2_port, ZN => n660);
   U109 : AOI22_X1 port map( A1 => n66, A2 => predict_PC_4_2_port, B1 => n65, 
                           B2 => predict_PC_5_2_port, ZN => n661);
   U108 : AOI22_X1 port map( A1 => n68, A2 => predict_PC_6_2_port, B1 => n67, 
                           B2 => predict_PC_7_2_port, ZN => n662);
   U107 : NAND4_X1 port map( A1 => n659, A2 => n660, A3 => n661, A4 => n662, ZN
                           => n653);
   U106 : AOI22_X1 port map( A1 => n70, A2 => predict_PC_8_2_port, B1 => n69, 
                           B2 => predict_PC_9_2_port, ZN => n655);
   U105 : AOI22_X1 port map( A1 => n72, A2 => predict_PC_10_2_port, B1 => n71, 
                           B2 => predict_PC_11_2_port, ZN => n656);
   U104 : AOI22_X1 port map( A1 => n74, A2 => predict_PC_12_2_port, B1 => n73, 
                           B2 => predict_PC_13_2_port, ZN => n657);
   U103 : AOI22_X1 port map( A1 => n76, A2 => predict_PC_14_2_port, B1 => n75, 
                           B2 => predict_PC_15_2_port, ZN => n658);
   U102 : NAND4_X1 port map( A1 => n655, A2 => n656, A3 => n657, A4 => n658, ZN
                           => n654);
   U45 : AOI22_X1 port map( A1 => n62, A2 => predict_PC_0_6_port, B1 => n61, B2
                           => predict_PC_1_6_port, ZN => n599);
   U44 : AOI22_X1 port map( A1 => n64, A2 => predict_PC_2_6_port, B1 => n63, B2
                           => predict_PC_3_6_port, ZN => n600);
   U43 : AOI22_X1 port map( A1 => n66, A2 => predict_PC_4_6_port, B1 => n65, B2
                           => predict_PC_5_6_port, ZN => n601);
   U42 : AOI22_X1 port map( A1 => n68, A2 => predict_PC_6_6_port, B1 => n67, B2
                           => predict_PC_7_6_port, ZN => n602);
   U41 : NAND4_X1 port map( A1 => n599, A2 => n600, A3 => n601, A4 => n602, ZN 
                           => n593);
   U40 : AOI22_X1 port map( A1 => n70, A2 => predict_PC_8_6_port, B1 => n69, B2
                           => predict_PC_9_6_port, ZN => n595);
   U39 : AOI22_X1 port map( A1 => n72, A2 => predict_PC_10_6_port, B1 => n71, 
                           B2 => predict_PC_11_6_port, ZN => n596);
   U38 : AOI22_X1 port map( A1 => n74, A2 => predict_PC_12_6_port, B1 => n73, 
                           B2 => predict_PC_13_6_port, ZN => n597);
   U37 : AOI22_X1 port map( A1 => n76, A2 => predict_PC_14_6_port, B1 => n75, 
                           B2 => predict_PC_15_6_port, ZN => n598);
   U36 : NAND4_X1 port map( A1 => n595, A2 => n596, A3 => n597, A4 => n598, ZN 
                           => n594);
   U67 : AOI22_X1 port map( A1 => n62, A2 => predict_PC_0_4_port, B1 => n61, B2
                           => predict_PC_1_4_port, ZN => n619);
   U66 : AOI22_X1 port map( A1 => n64, A2 => predict_PC_2_4_port, B1 => n63, B2
                           => predict_PC_3_4_port, ZN => n620);
   U65 : AOI22_X1 port map( A1 => n66, A2 => predict_PC_4_4_port, B1 => n65, B2
                           => predict_PC_5_4_port, ZN => n621);
   U64 : AOI22_X1 port map( A1 => n68, A2 => predict_PC_6_4_port, B1 => n67, B2
                           => predict_PC_7_4_port, ZN => n622);
   U63 : NAND4_X1 port map( A1 => n619, A2 => n620, A3 => n621, A4 => n622, ZN 
                           => n613);
   U62 : AOI22_X1 port map( A1 => n70, A2 => predict_PC_8_4_port, B1 => n69, B2
                           => predict_PC_9_4_port, ZN => n615);
   U61 : AOI22_X1 port map( A1 => n72, A2 => predict_PC_10_4_port, B1 => n71, 
                           B2 => predict_PC_11_4_port, ZN => n616);
   U60 : AOI22_X1 port map( A1 => n74, A2 => predict_PC_12_4_port, B1 => n73, 
                           B2 => predict_PC_13_4_port, ZN => n617);
   U59 : AOI22_X1 port map( A1 => n76, A2 => predict_PC_14_4_port, B1 => n75, 
                           B2 => predict_PC_15_4_port, ZN => n618);
   U58 : NAND4_X1 port map( A1 => n615, A2 => n616, A3 => n617, A4 => n618, ZN 
                           => n614);
   U56 : AOI22_X1 port map( A1 => n62, A2 => predict_PC_0_5_port, B1 => n61, B2
                           => predict_PC_1_5_port, ZN => n609);
   U55 : AOI22_X1 port map( A1 => n64, A2 => predict_PC_2_5_port, B1 => n63, B2
                           => predict_PC_3_5_port, ZN => n610);
   U54 : AOI22_X1 port map( A1 => n66, A2 => predict_PC_4_5_port, B1 => n65, B2
                           => predict_PC_5_5_port, ZN => n611);
   U53 : AOI22_X1 port map( A1 => n68, A2 => predict_PC_6_5_port, B1 => n67, B2
                           => predict_PC_7_5_port, ZN => n612);
   U52 : NAND4_X1 port map( A1 => n609, A2 => n610, A3 => n611, A4 => n612, ZN 
                           => n603);
   U51 : AOI22_X1 port map( A1 => n70, A2 => predict_PC_8_5_port, B1 => n69, B2
                           => predict_PC_9_5_port, ZN => n605);
   U50 : AOI22_X1 port map( A1 => n72, A2 => predict_PC_10_5_port, B1 => n71, 
                           B2 => predict_PC_11_5_port, ZN => n606);
   U49 : AOI22_X1 port map( A1 => n74, A2 => predict_PC_12_5_port, B1 => n73, 
                           B2 => predict_PC_13_5_port, ZN => n607);
   U48 : AOI22_X1 port map( A1 => n76, A2 => predict_PC_14_5_port, B1 => n75, 
                           B2 => predict_PC_15_5_port, ZN => n608);
   U47 : NAND4_X1 port map( A1 => n605, A2 => n606, A3 => n607, A4 => n608, ZN 
                           => n604);
   U12 : AOI22_X1 port map( A1 => n62, A2 => predict_PC_0_9_port, B1 => n572, 
                           B2 => predict_PC_1_9_port, ZN => n561);
   U11 : AOI22_X1 port map( A1 => n64, A2 => predict_PC_2_9_port, B1 => n570, 
                           B2 => predict_PC_3_9_port, ZN => n562);
   U10 : AOI22_X1 port map( A1 => n66, A2 => predict_PC_4_9_port, B1 => n568, 
                           B2 => predict_PC_5_9_port, ZN => n563);
   U9 : AOI22_X1 port map( A1 => n68, A2 => predict_PC_6_9_port, B1 => 
                           n566_port, B2 => predict_PC_7_9_port, ZN => n564);
   U8 : NAND4_X1 port map( A1 => n561, A2 => n562, A3 => n563, A4 => n564, ZN 
                           => n547);
   U7 : AOI22_X1 port map( A1 => n70, A2 => predict_PC_8_9_port, B1 => n560, B2
                           => predict_PC_9_9_port, ZN => n549);
   U6 : AOI22_X1 port map( A1 => n72, A2 => predict_PC_10_9_port, B1 => n71, B2
                           => predict_PC_11_9_port, ZN => n550);
   U5 : AOI22_X1 port map( A1 => n74, A2 => predict_PC_12_9_port, B1 => n73, B2
                           => predict_PC_13_9_port, ZN => n551);
   U4 : AOI22_X1 port map( A1 => n76, A2 => predict_PC_14_9_port, B1 => n75, B2
                           => predict_PC_15_9_port, ZN => n552);
   U3 : NAND4_X1 port map( A1 => n549, A2 => n550, A3 => n551, A4 => n552, ZN 
                           => n548);
   U34 : AOI22_X1 port map( A1 => n62, A2 => predict_PC_0_7_port, B1 => n61, B2
                           => predict_PC_1_7_port, ZN => n589);
   U33 : AOI22_X1 port map( A1 => n64, A2 => predict_PC_2_7_port, B1 => n63, B2
                           => predict_PC_3_7_port, ZN => n590);
   U32 : AOI22_X1 port map( A1 => n66, A2 => predict_PC_4_7_port, B1 => n65, B2
                           => predict_PC_5_7_port, ZN => n591);
   U31 : AOI22_X1 port map( A1 => n68, A2 => predict_PC_6_7_port, B1 => n67, B2
                           => predict_PC_7_7_port, ZN => n592);
   U30 : NAND4_X1 port map( A1 => n589, A2 => n590, A3 => n591, A4 => n592, ZN 
                           => n583);
   U29 : AOI22_X1 port map( A1 => n70, A2 => predict_PC_8_7_port, B1 => n69, B2
                           => predict_PC_9_7_port, ZN => n585);
   U28 : AOI22_X1 port map( A1 => n72, A2 => predict_PC_10_7_port, B1 => n71, 
                           B2 => predict_PC_11_7_port, ZN => n586);
   U27 : AOI22_X1 port map( A1 => n74, A2 => predict_PC_12_7_port, B1 => n73, 
                           B2 => predict_PC_13_7_port, ZN => n587);
   U26 : AOI22_X1 port map( A1 => n76, A2 => predict_PC_14_7_port, B1 => n75, 
                           B2 => predict_PC_15_7_port, ZN => n588);
   U25 : NAND4_X1 port map( A1 => n585, A2 => n586, A3 => n587, A4 => n588, ZN 
                           => n584);
   U23 : AOI22_X1 port map( A1 => n62, A2 => predict_PC_0_8_port, B1 => n61, B2
                           => predict_PC_1_8_port, ZN => n579);
   U22 : AOI22_X1 port map( A1 => n64, A2 => predict_PC_2_8_port, B1 => n63, B2
                           => predict_PC_3_8_port, ZN => n580);
   U21 : AOI22_X1 port map( A1 => n66, A2 => predict_PC_4_8_port, B1 => n65, B2
                           => predict_PC_5_8_port, ZN => n581);
   U20 : AOI22_X1 port map( A1 => n68, A2 => predict_PC_6_8_port, B1 => n67, B2
                           => predict_PC_7_8_port, ZN => n582);
   U19 : NAND4_X1 port map( A1 => n579, A2 => n580, A3 => n581, A4 => n582, ZN 
                           => n573);
   U18 : AOI22_X1 port map( A1 => n70, A2 => predict_PC_8_8_port, B1 => n69, B2
                           => predict_PC_9_8_port, ZN => n575);
   U17 : AOI22_X1 port map( A1 => n72, A2 => predict_PC_10_8_port, B1 => n71, 
                           B2 => predict_PC_11_8_port, ZN => n576);
   U16 : AOI22_X1 port map( A1 => n74, A2 => predict_PC_12_8_port, B1 => n73, 
                           B2 => predict_PC_13_8_port, ZN => n577);
   U15 : AOI22_X1 port map( A1 => n76, A2 => predict_PC_14_8_port, B1 => n75, 
                           B2 => predict_PC_15_8_port, ZN => n578);
   U14 : NAND4_X1 port map( A1 => n575, A2 => n576, A3 => n577, A4 => n578, ZN 
                           => n574);
   U78 : AOI22_X1 port map( A1 => n62, A2 => predict_PC_0_3_port, B1 => n61, B2
                           => predict_PC_1_3_port, ZN => n629);
   U77 : AOI22_X1 port map( A1 => n64, A2 => predict_PC_2_3_port, B1 => n63, B2
                           => predict_PC_3_3_port, ZN => n630);
   U76 : AOI22_X1 port map( A1 => n66, A2 => predict_PC_4_3_port, B1 => n65, B2
                           => predict_PC_5_3_port, ZN => n631);
   U75 : AOI22_X1 port map( A1 => n68, A2 => predict_PC_6_3_port, B1 => n67, B2
                           => predict_PC_7_3_port, ZN => n632);
   U74 : NAND4_X1 port map( A1 => n629, A2 => n630, A3 => n631, A4 => n632, ZN 
                           => n623);
   U73 : AOI22_X1 port map( A1 => n70, A2 => predict_PC_8_3_port, B1 => n69, B2
                           => predict_PC_9_3_port, ZN => n625);
   U72 : AOI22_X1 port map( A1 => n72, A2 => predict_PC_10_3_port, B1 => n71, 
                           B2 => predict_PC_11_3_port, ZN => n626);
   U71 : AOI22_X1 port map( A1 => n74, A2 => predict_PC_12_3_port, B1 => n73, 
                           B2 => predict_PC_13_3_port, ZN => n627);
   U70 : AOI22_X1 port map( A1 => n76, A2 => predict_PC_14_3_port, B1 => n75, 
                           B2 => predict_PC_15_3_port, ZN => n628);
   U69 : NAND4_X1 port map( A1 => n625, A2 => n626, A3 => n627, A4 => n628, ZN 
                           => n624);
   U122 : AOI22_X1 port map( A1 => n62, A2 => predict_PC_0_29_port, B1 => n61, 
                           B2 => predict_PC_1_29_port, ZN => n669);
   U121 : AOI22_X1 port map( A1 => n64, A2 => predict_PC_2_29_port, B1 => n63, 
                           B2 => predict_PC_3_29_port, ZN => n670);
   U120 : AOI22_X1 port map( A1 => n66, A2 => predict_PC_4_29_port, B1 => n65, 
                           B2 => predict_PC_5_29_port, ZN => n671);
   U119 : AOI22_X1 port map( A1 => n68, A2 => predict_PC_6_29_port, B1 => n67, 
                           B2 => predict_PC_7_29_port, ZN => n672);
   U118 : NAND4_X1 port map( A1 => n669, A2 => n670, A3 => n671, A4 => n672, ZN
                           => n663);
   U117 : AOI22_X1 port map( A1 => n70, A2 => predict_PC_8_29_port, B1 => n69, 
                           B2 => predict_PC_9_29_port, ZN => n665);
   U116 : AOI22_X1 port map( A1 => n72, A2 => predict_PC_10_29_port, B1 => n71,
                           B2 => predict_PC_11_29_port, ZN => n666);
   U115 : AOI22_X1 port map( A1 => n74, A2 => predict_PC_12_29_port, B1 => n73,
                           B2 => predict_PC_13_29_port, ZN => n667);
   U114 : AOI22_X1 port map( A1 => n76, A2 => predict_PC_14_29_port, B1 => n75,
                           B2 => predict_PC_15_29_port, ZN => n668);
   U113 : NAND4_X1 port map( A1 => n665, A2 => n666, A3 => n667, A4 => n668, ZN
                           => n664);
   U100 : AOI22_X1 port map( A1 => n62, A2 => predict_PC_0_30_port, B1 => n61, 
                           B2 => predict_PC_1_30_port, ZN => n649);
   U99 : AOI22_X1 port map( A1 => n64, A2 => predict_PC_2_30_port, B1 => n63, 
                           B2 => predict_PC_3_30_port, ZN => n650);
   U98 : AOI22_X1 port map( A1 => n66, A2 => predict_PC_4_30_port, B1 => n65, 
                           B2 => predict_PC_5_30_port, ZN => n651);
   U97 : AOI22_X1 port map( A1 => n68, A2 => predict_PC_6_30_port, B1 => n67, 
                           B2 => predict_PC_7_30_port, ZN => n652);
   U96 : NAND4_X1 port map( A1 => n649, A2 => n650, A3 => n651, A4 => n652, ZN 
                           => n643);
   U95 : AOI22_X1 port map( A1 => n70, A2 => predict_PC_8_30_port, B1 => n69, 
                           B2 => predict_PC_9_30_port, ZN => n645);
   U94 : AOI22_X1 port map( A1 => n72, A2 => predict_PC_10_30_port, B1 => n71, 
                           B2 => predict_PC_11_30_port, ZN => n646);
   U93 : AOI22_X1 port map( A1 => n74, A2 => predict_PC_12_30_port, B1 => n73, 
                           B2 => predict_PC_13_30_port, ZN => n647);
   U92 : AOI22_X1 port map( A1 => n76, A2 => predict_PC_14_30_port, B1 => n75, 
                           B2 => predict_PC_15_30_port, ZN => n648);
   U91 : NAND4_X1 port map( A1 => n645, A2 => n646, A3 => n647, A4 => n648, ZN 
                           => n644);
   U89 : AOI22_X1 port map( A1 => n62, A2 => predict_PC_0_31_port, B1 => n61, 
                           B2 => predict_PC_1_31_port, ZN => n639);
   U88 : AOI22_X1 port map( A1 => n64, A2 => predict_PC_2_31_port, B1 => n63, 
                           B2 => predict_PC_3_31_port, ZN => n640);
   U87 : AOI22_X1 port map( A1 => n66, A2 => predict_PC_4_31_port, B1 => n65, 
                           B2 => predict_PC_5_31_port, ZN => n641);
   U86 : AOI22_X1 port map( A1 => n68, A2 => predict_PC_6_31_port, B1 => n67, 
                           B2 => predict_PC_7_31_port, ZN => n642);
   U85 : NAND4_X1 port map( A1 => n639, A2 => n640, A3 => n641, A4 => n642, ZN 
                           => n633);
   U84 : AOI22_X1 port map( A1 => n70, A2 => predict_PC_8_31_port, B1 => n69, 
                           B2 => predict_PC_9_31_port, ZN => n635);
   U83 : AOI22_X1 port map( A1 => n72, A2 => predict_PC_10_31_port, B1 => n71, 
                           B2 => predict_PC_11_31_port, ZN => n636);
   U82 : AOI22_X1 port map( A1 => n74, A2 => predict_PC_12_31_port, B1 => n73, 
                           B2 => predict_PC_13_31_port, ZN => n637);
   U81 : AOI22_X1 port map( A1 => n76, A2 => predict_PC_14_31_port, B1 => n75, 
                           B2 => predict_PC_15_31_port, ZN => n638);
   U80 : NAND4_X1 port map( A1 => n635, A2 => n636, A3 => n637, A4 => n638, ZN 
                           => n634);
   U265 : AOI22_X1 port map( A1 => n62, A2 => predict_PC_0_17_port, B1 => n61, 
                           B2 => predict_PC_1_17_port, ZN => n799);
   U264 : AOI22_X1 port map( A1 => n64, A2 => predict_PC_2_17_port, B1 => n63, 
                           B2 => predict_PC_3_17_port, ZN => n800);
   U263 : AOI22_X1 port map( A1 => n66, A2 => predict_PC_4_17_port, B1 => n65, 
                           B2 => predict_PC_5_17_port, ZN => n801);
   U262 : AOI22_X1 port map( A1 => n68, A2 => predict_PC_6_17_port, B1 => n67, 
                           B2 => predict_PC_7_17_port, ZN => n802);
   U261 : NAND4_X1 port map( A1 => n799, A2 => n800, A3 => n801, A4 => n802, ZN
                           => n793);
   U260 : AOI22_X1 port map( A1 => n70, A2 => predict_PC_8_17_port, B1 => n69, 
                           B2 => predict_PC_9_17_port, ZN => n795);
   U259 : AOI22_X1 port map( A1 => n72, A2 => predict_PC_10_17_port, B1 => n71,
                           B2 => predict_PC_11_17_port, ZN => n796);
   U258 : AOI22_X1 port map( A1 => n74, A2 => predict_PC_12_17_port, B1 => n73,
                           B2 => predict_PC_13_17_port, ZN => n797);
   U257 : AOI22_X1 port map( A1 => n76, A2 => predict_PC_14_17_port, B1 => n75,
                           B2 => predict_PC_15_17_port, ZN => n798);
   U256 : NAND4_X1 port map( A1 => n795, A2 => n796, A3 => n797, A4 => n798, ZN
                           => n794);
   U232 : AOI22_X1 port map( A1 => n571, A2 => predict_PC_0_1_port, B1 => n572,
                           B2 => predict_PC_1_1_port, ZN => n769);
   U231 : AOI22_X1 port map( A1 => n569, A2 => predict_PC_2_1_port, B1 => n570,
                           B2 => predict_PC_3_1_port, ZN => n770);
   U230 : AOI22_X1 port map( A1 => n567_port, A2 => predict_PC_4_1_port, B1 => 
                           n568, B2 => predict_PC_5_1_port, ZN => n771);
   U229 : AOI22_X1 port map( A1 => n565, A2 => predict_PC_6_1_port, B1 => 
                           n566_port, B2 => predict_PC_7_1_port, ZN => n772);
   U228 : NAND4_X1 port map( A1 => n769, A2 => n770, A3 => n771, A4 => n772, ZN
                           => n763);
   U227 : AOI22_X1 port map( A1 => n70, A2 => predict_PC_8_1_port, B1 => n560, 
                           B2 => predict_PC_9_1_port, ZN => n765);
   U226 : AOI22_X1 port map( A1 => n72, A2 => predict_PC_10_1_port, B1 => n71, 
                           B2 => predict_PC_11_1_port, ZN => n766);
   U225 : AOI22_X1 port map( A1 => n74, A2 => predict_PC_12_1_port, B1 => n73, 
                           B2 => predict_PC_13_1_port, ZN => n767);
   U224 : AOI22_X1 port map( A1 => n76, A2 => predict_PC_14_1_port, B1 => n75, 
                           B2 => predict_PC_15_1_port, ZN => n768);
   U223 : NAND4_X1 port map( A1 => n765, A2 => n766, A3 => n767, A4 => n768, ZN
                           => n764);
   U177 : AOI22_X1 port map( A1 => n571, A2 => predict_PC_0_24_port, B1 => n572
                           , B2 => predict_PC_1_24_port, ZN => n719);
   U176 : AOI22_X1 port map( A1 => n569, A2 => predict_PC_2_24_port, B1 => n570
                           , B2 => predict_PC_3_24_port, ZN => n720);
   U175 : AOI22_X1 port map( A1 => n567_port, A2 => predict_PC_4_24_port, B1 =>
                           n568, B2 => predict_PC_5_24_port, ZN => n721);
   U174 : AOI22_X1 port map( A1 => n565, A2 => predict_PC_6_24_port, B1 => 
                           n566_port, B2 => predict_PC_7_24_port, ZN => n722);
   U173 : NAND4_X1 port map( A1 => n719, A2 => n720, A3 => n721, A4 => n722, ZN
                           => n713);
   U172 : AOI22_X1 port map( A1 => n70, A2 => predict_PC_8_24_port, B1 => n560,
                           B2 => predict_PC_9_24_port, ZN => n715);
   U171 : AOI22_X1 port map( A1 => n72, A2 => predict_PC_10_24_port, B1 => n71,
                           B2 => predict_PC_11_24_port, ZN => n716);
   U170 : AOI22_X1 port map( A1 => n74, A2 => predict_PC_12_24_port, B1 => n73,
                           B2 => predict_PC_13_24_port, ZN => n717);
   U169 : AOI22_X1 port map( A1 => n76, A2 => predict_PC_14_24_port, B1 => n75,
                           B2 => predict_PC_15_24_port, ZN => n718);
   U168 : NAND4_X1 port map( A1 => n715, A2 => n716, A3 => n717, A4 => n718, ZN
                           => n714);
   U221 : AOI22_X1 port map( A1 => n62, A2 => predict_PC_0_20_port, B1 => n61, 
                           B2 => predict_PC_1_20_port, ZN => n759);
   U220 : AOI22_X1 port map( A1 => n64, A2 => predict_PC_2_20_port, B1 => n63, 
                           B2 => predict_PC_3_20_port, ZN => n760);
   U219 : AOI22_X1 port map( A1 => n66, A2 => predict_PC_4_20_port, B1 => n65, 
                           B2 => predict_PC_5_20_port, ZN => n761);
   U218 : AOI22_X1 port map( A1 => n68, A2 => predict_PC_6_20_port, B1 => n67, 
                           B2 => predict_PC_7_20_port, ZN => n762);
   U217 : NAND4_X1 port map( A1 => n759, A2 => n760, A3 => n761, A4 => n762, ZN
                           => n753);
   U216 : AOI22_X1 port map( A1 => n70, A2 => predict_PC_8_20_port, B1 => n69, 
                           B2 => predict_PC_9_20_port, ZN => n755);
   U215 : AOI22_X1 port map( A1 => n72, A2 => predict_PC_10_20_port, B1 => n71,
                           B2 => predict_PC_11_20_port, ZN => n756);
   U214 : AOI22_X1 port map( A1 => n74, A2 => predict_PC_12_20_port, B1 => n73,
                           B2 => predict_PC_13_20_port, ZN => n757);
   U213 : AOI22_X1 port map( A1 => n76, A2 => predict_PC_14_20_port, B1 => n75,
                           B2 => predict_PC_15_20_port, ZN => n758);
   U212 : NAND4_X1 port map( A1 => n755, A2 => n756, A3 => n757, A4 => n758, ZN
                           => n754);
   U155 : AOI22_X1 port map( A1 => n571, A2 => predict_PC_0_26_port, B1 => n572
                           , B2 => predict_PC_1_26_port, ZN => n699);
   U154 : AOI22_X1 port map( A1 => n569, A2 => predict_PC_2_26_port, B1 => n570
                           , B2 => predict_PC_3_26_port, ZN => n700);
   U153 : AOI22_X1 port map( A1 => n567_port, A2 => predict_PC_4_26_port, B1 =>
                           n568, B2 => predict_PC_5_26_port, ZN => n701);
   U152 : AOI22_X1 port map( A1 => n565, A2 => predict_PC_6_26_port, B1 => 
                           n566_port, B2 => predict_PC_7_26_port, ZN => n702);
   U151 : NAND4_X1 port map( A1 => n699, A2 => n700, A3 => n701, A4 => n702, ZN
                           => n693);
   U150 : AOI22_X1 port map( A1 => n70, A2 => predict_PC_8_26_port, B1 => n560,
                           B2 => predict_PC_9_26_port, ZN => n695);
   U149 : AOI22_X1 port map( A1 => n72, A2 => predict_PC_10_26_port, B1 => n71,
                           B2 => predict_PC_11_26_port, ZN => n696);
   U148 : AOI22_X1 port map( A1 => n74, A2 => predict_PC_12_26_port, B1 => n73,
                           B2 => predict_PC_13_26_port, ZN => n697);
   U147 : AOI22_X1 port map( A1 => n76, A2 => predict_PC_14_26_port, B1 => n75,
                           B2 => predict_PC_15_26_port, ZN => n698);
   U146 : NAND4_X1 port map( A1 => n695, A2 => n696, A3 => n697, A4 => n698, ZN
                           => n694);
   U254 : AOI22_X1 port map( A1 => n571, A2 => predict_PC_0_18_port, B1 => n572
                           , B2 => predict_PC_1_18_port, ZN => n789);
   U253 : AOI22_X1 port map( A1 => n569, A2 => predict_PC_2_18_port, B1 => n570
                           , B2 => predict_PC_3_18_port, ZN => n790);
   U252 : AOI22_X1 port map( A1 => n567_port, A2 => predict_PC_4_18_port, B1 =>
                           n568, B2 => predict_PC_5_18_port, ZN => n791);
   U251 : AOI22_X1 port map( A1 => n565, A2 => predict_PC_6_18_port, B1 => 
                           n566_port, B2 => predict_PC_7_18_port, ZN => n792);
   U250 : NAND4_X1 port map( A1 => n789, A2 => n790, A3 => n791, A4 => n792, ZN
                           => n783);
   U249 : AOI22_X1 port map( A1 => n70, A2 => predict_PC_8_18_port, B1 => n69, 
                           B2 => predict_PC_9_18_port, ZN => n785);
   U248 : AOI22_X1 port map( A1 => n72, A2 => predict_PC_10_18_port, B1 => n71,
                           B2 => predict_PC_11_18_port, ZN => n786);
   U247 : AOI22_X1 port map( A1 => n74, A2 => predict_PC_12_18_port, B1 => n73,
                           B2 => predict_PC_13_18_port, ZN => n787);
   U246 : AOI22_X1 port map( A1 => n76, A2 => predict_PC_14_18_port, B1 => n75,
                           B2 => predict_PC_15_18_port, ZN => n788);
   U245 : NAND4_X1 port map( A1 => n785, A2 => n786, A3 => n787, A4 => n788, ZN
                           => n784);
   U199 : AOI22_X1 port map( A1 => n571, A2 => predict_PC_0_22_port, B1 => n61,
                           B2 => predict_PC_1_22_port, ZN => n739);
   U198 : AOI22_X1 port map( A1 => n569, A2 => predict_PC_2_22_port, B1 => n63,
                           B2 => predict_PC_3_22_port, ZN => n740);
   U197 : AOI22_X1 port map( A1 => n567_port, A2 => predict_PC_4_22_port, B1 =>
                           n65, B2 => predict_PC_5_22_port, ZN => n741);
   U196 : AOI22_X1 port map( A1 => n565, A2 => predict_PC_6_22_port, B1 => n67,
                           B2 => predict_PC_7_22_port, ZN => n742);
   U195 : NAND4_X1 port map( A1 => n739, A2 => n740, A3 => n741, A4 => n742, ZN
                           => n733);
   U194 : AOI22_X1 port map( A1 => n70, A2 => predict_PC_8_22_port, B1 => n69, 
                           B2 => predict_PC_9_22_port, ZN => n735);
   U193 : AOI22_X1 port map( A1 => n72, A2 => predict_PC_10_22_port, B1 => n71,
                           B2 => predict_PC_11_22_port, ZN => n736);
   U192 : AOI22_X1 port map( A1 => n74, A2 => predict_PC_12_22_port, B1 => n73,
                           B2 => predict_PC_13_22_port, ZN => n737);
   U191 : AOI22_X1 port map( A1 => n76, A2 => predict_PC_14_22_port, B1 => n75,
                           B2 => predict_PC_15_22_port, ZN => n738);
   U190 : NAND4_X1 port map( A1 => n735, A2 => n736, A3 => n737, A4 => n738, ZN
                           => n734);
   U210 : AOI22_X1 port map( A1 => n571, A2 => predict_PC_0_21_port, B1 => n572
                           , B2 => predict_PC_1_21_port, ZN => n749);
   U209 : AOI22_X1 port map( A1 => n569, A2 => predict_PC_2_21_port, B1 => n570
                           , B2 => predict_PC_3_21_port, ZN => n750);
   U208 : AOI22_X1 port map( A1 => n567_port, A2 => predict_PC_4_21_port, B1 =>
                           n568, B2 => predict_PC_5_21_port, ZN => n751);
   U207 : AOI22_X1 port map( A1 => n565, A2 => predict_PC_6_21_port, B1 => 
                           n566_port, B2 => predict_PC_7_21_port, ZN => n752);
   U206 : NAND4_X1 port map( A1 => n749, A2 => n750, A3 => n751, A4 => n752, ZN
                           => n743);
   U205 : AOI22_X1 port map( A1 => n70, A2 => predict_PC_8_21_port, B1 => n560,
                           B2 => predict_PC_9_21_port, ZN => n745);
   U204 : AOI22_X1 port map( A1 => n72, A2 => predict_PC_10_21_port, B1 => n71,
                           B2 => predict_PC_11_21_port, ZN => n746);
   U203 : AOI22_X1 port map( A1 => n74, A2 => predict_PC_12_21_port, B1 => n73,
                           B2 => predict_PC_13_21_port, ZN => n747);
   U202 : AOI22_X1 port map( A1 => n76, A2 => predict_PC_14_21_port, B1 => n75,
                           B2 => predict_PC_15_21_port, ZN => n748);
   U201 : NAND4_X1 port map( A1 => n745, A2 => n746, A3 => n747, A4 => n748, ZN
                           => n744);
   U243 : AOI22_X1 port map( A1 => n62, A2 => predict_PC_0_19_port, B1 => n61, 
                           B2 => predict_PC_1_19_port, ZN => n779);
   U242 : AOI22_X1 port map( A1 => n64, A2 => predict_PC_2_19_port, B1 => n63, 
                           B2 => predict_PC_3_19_port, ZN => n780);
   U241 : AOI22_X1 port map( A1 => n66, A2 => predict_PC_4_19_port, B1 => n65, 
                           B2 => predict_PC_5_19_port, ZN => n781);
   U240 : AOI22_X1 port map( A1 => n68, A2 => predict_PC_6_19_port, B1 => n67, 
                           B2 => predict_PC_7_19_port, ZN => n782);
   U239 : NAND4_X1 port map( A1 => n779, A2 => n780, A3 => n781, A4 => n782, ZN
                           => n773);
   U238 : AOI22_X1 port map( A1 => n70, A2 => predict_PC_8_19_port, B1 => n69, 
                           B2 => predict_PC_9_19_port, ZN => n775);
   U237 : AOI22_X1 port map( A1 => n72, A2 => predict_PC_10_19_port, B1 => n71,
                           B2 => predict_PC_11_19_port, ZN => n776);
   U236 : AOI22_X1 port map( A1 => n74, A2 => predict_PC_12_19_port, B1 => n73,
                           B2 => predict_PC_13_19_port, ZN => n777);
   U235 : AOI22_X1 port map( A1 => n76, A2 => predict_PC_14_19_port, B1 => n75,
                           B2 => predict_PC_15_19_port, ZN => n778);
   U234 : NAND4_X1 port map( A1 => n775, A2 => n776, A3 => n777, A4 => n778, ZN
                           => n774);
   U166 : AOI22_X1 port map( A1 => n62, A2 => predict_PC_0_25_port, B1 => n572,
                           B2 => predict_PC_1_25_port, ZN => n709);
   U165 : AOI22_X1 port map( A1 => n64, A2 => predict_PC_2_25_port, B1 => n570,
                           B2 => predict_PC_3_25_port, ZN => n710);
   U164 : AOI22_X1 port map( A1 => n66, A2 => predict_PC_4_25_port, B1 => n568,
                           B2 => predict_PC_5_25_port, ZN => n711);
   U163 : AOI22_X1 port map( A1 => n68, A2 => predict_PC_6_25_port, B1 => 
                           n566_port, B2 => predict_PC_7_25_port, ZN => n712);
   U162 : NAND4_X1 port map( A1 => n709, A2 => n710, A3 => n711, A4 => n712, ZN
                           => n703);
   U161 : AOI22_X1 port map( A1 => n70, A2 => predict_PC_8_25_port, B1 => n560,
                           B2 => predict_PC_9_25_port, ZN => n705);
   U160 : AOI22_X1 port map( A1 => n72, A2 => predict_PC_10_25_port, B1 => n71,
                           B2 => predict_PC_11_25_port, ZN => n706);
   U159 : AOI22_X1 port map( A1 => n74, A2 => predict_PC_12_25_port, B1 => n73,
                           B2 => predict_PC_13_25_port, ZN => n707);
   U158 : AOI22_X1 port map( A1 => n76, A2 => predict_PC_14_25_port, B1 => n75,
                           B2 => predict_PC_15_25_port, ZN => n708);
   U157 : NAND4_X1 port map( A1 => n705, A2 => n706, A3 => n707, A4 => n708, ZN
                           => n704);
   U144 : AOI22_X1 port map( A1 => n62, A2 => predict_PC_0_27_port, B1 => n61, 
                           B2 => predict_PC_1_27_port, ZN => n689);
   U143 : AOI22_X1 port map( A1 => n64, A2 => predict_PC_2_27_port, B1 => n63, 
                           B2 => predict_PC_3_27_port, ZN => n690);
   U142 : AOI22_X1 port map( A1 => n66, A2 => predict_PC_4_27_port, B1 => n65, 
                           B2 => predict_PC_5_27_port, ZN => n691);
   U141 : AOI22_X1 port map( A1 => n68, A2 => predict_PC_6_27_port, B1 => n67, 
                           B2 => predict_PC_7_27_port, ZN => n692);
   U140 : NAND4_X1 port map( A1 => n689, A2 => n690, A3 => n691, A4 => n692, ZN
                           => n683);
   U139 : AOI22_X1 port map( A1 => n70, A2 => predict_PC_8_27_port, B1 => n560,
                           B2 => predict_PC_9_27_port, ZN => n685);
   U138 : AOI22_X1 port map( A1 => n72, A2 => predict_PC_10_27_port, B1 => n71,
                           B2 => predict_PC_11_27_port, ZN => n686);
   U137 : AOI22_X1 port map( A1 => n74, A2 => predict_PC_12_27_port, B1 => n73,
                           B2 => predict_PC_13_27_port, ZN => n687);
   U136 : AOI22_X1 port map( A1 => n76, A2 => predict_PC_14_27_port, B1 => n75,
                           B2 => predict_PC_15_27_port, ZN => n688);
   U135 : NAND4_X1 port map( A1 => n685, A2 => n686, A3 => n687, A4 => n688, ZN
                           => n684);
   U353 : AOI22_X1 port map( A1 => n62, A2 => predict_PC_0_0_port, B1 => n61, 
                           B2 => predict_PC_1_0_port, ZN => n879);
   U352 : AOI22_X1 port map( A1 => n64, A2 => predict_PC_2_0_port, B1 => n63, 
                           B2 => predict_PC_3_0_port, ZN => n880);
   U351 : AOI22_X1 port map( A1 => n66, A2 => predict_PC_4_0_port, B1 => n65, 
                           B2 => predict_PC_5_0_port, ZN => n881);
   U350 : AOI22_X1 port map( A1 => n68, A2 => predict_PC_6_0_port, B1 => n67, 
                           B2 => predict_PC_7_0_port, ZN => n882);
   U349 : NAND4_X1 port map( A1 => n879, A2 => n880, A3 => n881, A4 => n882, ZN
                           => n873);
   U348 : AOI22_X1 port map( A1 => n70, A2 => predict_PC_8_0_port, B1 => n69, 
                           B2 => predict_PC_9_0_port, ZN => n875);
   U347 : AOI22_X1 port map( A1 => n557, A2 => predict_PC_10_0_port, B1 => n558
                           , B2 => predict_PC_11_0_port, ZN => n876);
   U346 : AOI22_X1 port map( A1 => n74, A2 => predict_PC_12_0_port, B1 => n73, 
                           B2 => predict_PC_13_0_port, ZN => n877);
   U345 : AOI22_X1 port map( A1 => n553, A2 => predict_PC_14_0_port, B1 => n554
                           , B2 => predict_PC_15_0_port, ZN => n878);
   U344 : NAND4_X1 port map( A1 => n875, A2 => n876, A3 => n877, A4 => n878, ZN
                           => n874);
   U331 : AOI22_X1 port map( A1 => n62, A2 => predict_PC_0_11_port, B1 => n61, 
                           B2 => predict_PC_1_11_port, ZN => n859);
   U330 : AOI22_X1 port map( A1 => n64, A2 => predict_PC_2_11_port, B1 => n63, 
                           B2 => predict_PC_3_11_port, ZN => n860);
   U329 : AOI22_X1 port map( A1 => n66, A2 => predict_PC_4_11_port, B1 => n65, 
                           B2 => predict_PC_5_11_port, ZN => n861);
   U328 : AOI22_X1 port map( A1 => n68, A2 => predict_PC_6_11_port, B1 => n67, 
                           B2 => predict_PC_7_11_port, ZN => n862);
   U327 : NAND4_X1 port map( A1 => n859, A2 => n860, A3 => n861, A4 => n862, ZN
                           => n853);
   U326 : AOI22_X1 port map( A1 => n70, A2 => predict_PC_8_11_port, B1 => n69, 
                           B2 => predict_PC_9_11_port, ZN => n855);
   U325 : AOI22_X1 port map( A1 => n557, A2 => predict_PC_10_11_port, B1 => 
                           n558, B2 => predict_PC_11_11_port, ZN => n856);
   U324 : AOI22_X1 port map( A1 => n74, A2 => predict_PC_12_11_port, B1 => n73,
                           B2 => predict_PC_13_11_port, ZN => n857);
   U323 : AOI22_X1 port map( A1 => n553, A2 => predict_PC_14_11_port, B1 => 
                           n554, B2 => predict_PC_15_11_port, ZN => n858);
   U322 : NAND4_X1 port map( A1 => n855, A2 => n856, A3 => n857, A4 => n858, ZN
                           => n854);
   U320 : AOI22_X1 port map( A1 => n62, A2 => predict_PC_0_12_port, B1 => n61, 
                           B2 => predict_PC_1_12_port, ZN => n849);
   U319 : AOI22_X1 port map( A1 => n64, A2 => predict_PC_2_12_port, B1 => n63, 
                           B2 => predict_PC_3_12_port, ZN => n850);
   U318 : AOI22_X1 port map( A1 => n66, A2 => predict_PC_4_12_port, B1 => n65, 
                           B2 => predict_PC_5_12_port, ZN => n851);
   U317 : AOI22_X1 port map( A1 => n68, A2 => predict_PC_6_12_port, B1 => n67, 
                           B2 => predict_PC_7_12_port, ZN => n852);
   U316 : NAND4_X1 port map( A1 => n849, A2 => n850, A3 => n851, A4 => n852, ZN
                           => n843);
   U315 : AOI22_X1 port map( A1 => n70, A2 => predict_PC_8_12_port, B1 => n69, 
                           B2 => predict_PC_9_12_port, ZN => n845);
   U314 : AOI22_X1 port map( A1 => n557, A2 => predict_PC_10_12_port, B1 => 
                           n558, B2 => predict_PC_11_12_port, ZN => n846);
   U313 : AOI22_X1 port map( A1 => n74, A2 => predict_PC_12_12_port, B1 => n73,
                           B2 => predict_PC_13_12_port, ZN => n847);
   U312 : AOI22_X1 port map( A1 => n553, A2 => predict_PC_14_12_port, B1 => 
                           n554, B2 => predict_PC_15_12_port, ZN => n848);
   U311 : NAND4_X1 port map( A1 => n845, A2 => n846, A3 => n847, A4 => n848, ZN
                           => n844);
   U342 : AOI22_X1 port map( A1 => n62, A2 => predict_PC_0_10_port, B1 => n61, 
                           B2 => predict_PC_1_10_port, ZN => n869);
   U341 : AOI22_X1 port map( A1 => n64, A2 => predict_PC_2_10_port, B1 => n63, 
                           B2 => predict_PC_3_10_port, ZN => n870);
   U340 : AOI22_X1 port map( A1 => n66, A2 => predict_PC_4_10_port, B1 => n65, 
                           B2 => predict_PC_5_10_port, ZN => n871);
   U339 : AOI22_X1 port map( A1 => n68, A2 => predict_PC_6_10_port, B1 => n67, 
                           B2 => predict_PC_7_10_port, ZN => n872);
   U338 : NAND4_X1 port map( A1 => n869, A2 => n870, A3 => n871, A4 => n872, ZN
                           => n863);
   U337 : AOI22_X1 port map( A1 => n70, A2 => predict_PC_8_10_port, B1 => n69, 
                           B2 => predict_PC_9_10_port, ZN => n865);
   U336 : AOI22_X1 port map( A1 => n557, A2 => predict_PC_10_10_port, B1 => 
                           n558, B2 => predict_PC_11_10_port, ZN => n866);
   U335 : AOI22_X1 port map( A1 => n74, A2 => predict_PC_12_10_port, B1 => n73,
                           B2 => predict_PC_13_10_port, ZN => n867);
   U334 : AOI22_X1 port map( A1 => n553, A2 => predict_PC_14_10_port, B1 => 
                           n554, B2 => predict_PC_15_10_port, ZN => n868);
   U333 : NAND4_X1 port map( A1 => n865, A2 => n866, A3 => n867, A4 => n868, ZN
                           => n864);
   U276 : AOI22_X1 port map( A1 => n62, A2 => predict_PC_0_16_port, B1 => n61, 
                           B2 => predict_PC_1_16_port, ZN => n809);
   U275 : AOI22_X1 port map( A1 => n64, A2 => predict_PC_2_16_port, B1 => n63, 
                           B2 => predict_PC_3_16_port, ZN => n810);
   U274 : AOI22_X1 port map( A1 => n66, A2 => predict_PC_4_16_port, B1 => n65, 
                           B2 => predict_PC_5_16_port, ZN => n811);
   U273 : AOI22_X1 port map( A1 => n68, A2 => predict_PC_6_16_port, B1 => n67, 
                           B2 => predict_PC_7_16_port, ZN => n812);
   U272 : NAND4_X1 port map( A1 => n809, A2 => n810, A3 => n811, A4 => n812, ZN
                           => n803);
   U271 : AOI22_X1 port map( A1 => n70, A2 => predict_PC_8_16_port, B1 => n69, 
                           B2 => predict_PC_9_16_port, ZN => n805);
   U270 : AOI22_X1 port map( A1 => n557, A2 => predict_PC_10_16_port, B1 => 
                           n558, B2 => predict_PC_11_16_port, ZN => n806);
   U269 : AOI22_X1 port map( A1 => n74, A2 => predict_PC_12_16_port, B1 => n73,
                           B2 => predict_PC_13_16_port, ZN => n807);
   U268 : AOI22_X1 port map( A1 => n553, A2 => predict_PC_14_16_port, B1 => 
                           n554, B2 => predict_PC_15_16_port, ZN => n808);
   U267 : NAND4_X1 port map( A1 => n805, A2 => n806, A3 => n807, A4 => n808, ZN
                           => n804);
   U287 : AOI22_X1 port map( A1 => n62, A2 => predict_PC_0_15_port, B1 => n61, 
                           B2 => predict_PC_1_15_port, ZN => n819);
   U286 : AOI22_X1 port map( A1 => n64, A2 => predict_PC_2_15_port, B1 => n63, 
                           B2 => predict_PC_3_15_port, ZN => n820);
   U285 : AOI22_X1 port map( A1 => n66, A2 => predict_PC_4_15_port, B1 => n65, 
                           B2 => predict_PC_5_15_port, ZN => n821);
   U284 : AOI22_X1 port map( A1 => n68, A2 => predict_PC_6_15_port, B1 => n67, 
                           B2 => predict_PC_7_15_port, ZN => n822);
   U283 : NAND4_X1 port map( A1 => n819, A2 => n820, A3 => n821, A4 => n822, ZN
                           => n813);
   U282 : AOI22_X1 port map( A1 => n70, A2 => predict_PC_8_15_port, B1 => n69, 
                           B2 => predict_PC_9_15_port, ZN => n815);
   U281 : AOI22_X1 port map( A1 => n557, A2 => predict_PC_10_15_port, B1 => 
                           n558, B2 => predict_PC_11_15_port, ZN => n816);
   U280 : AOI22_X1 port map( A1 => n74, A2 => predict_PC_12_15_port, B1 => n73,
                           B2 => predict_PC_13_15_port, ZN => n817);
   U279 : AOI22_X1 port map( A1 => n553, A2 => predict_PC_14_15_port, B1 => 
                           n554, B2 => predict_PC_15_15_port, ZN => n818);
   U278 : NAND4_X1 port map( A1 => n815, A2 => n816, A3 => n817, A4 => n818, ZN
                           => n814);
   U298 : AOI22_X1 port map( A1 => n62, A2 => predict_PC_0_14_port, B1 => n61, 
                           B2 => predict_PC_1_14_port, ZN => n829);
   U297 : AOI22_X1 port map( A1 => n64, A2 => predict_PC_2_14_port, B1 => n63, 
                           B2 => predict_PC_3_14_port, ZN => n830);
   U296 : AOI22_X1 port map( A1 => n66, A2 => predict_PC_4_14_port, B1 => n65, 
                           B2 => predict_PC_5_14_port, ZN => n831);
   U295 : AOI22_X1 port map( A1 => n68, A2 => predict_PC_6_14_port, B1 => n67, 
                           B2 => predict_PC_7_14_port, ZN => n832);
   U294 : NAND4_X1 port map( A1 => n829, A2 => n830, A3 => n831, A4 => n832, ZN
                           => n823);
   U293 : AOI22_X1 port map( A1 => n70, A2 => predict_PC_8_14_port, B1 => n69, 
                           B2 => predict_PC_9_14_port, ZN => n825);
   U292 : AOI22_X1 port map( A1 => n557, A2 => predict_PC_10_14_port, B1 => 
                           n558, B2 => predict_PC_11_14_port, ZN => n826);
   U291 : AOI22_X1 port map( A1 => n74, A2 => predict_PC_12_14_port, B1 => n73,
                           B2 => predict_PC_13_14_port, ZN => n827);
   U290 : AOI22_X1 port map( A1 => n553, A2 => predict_PC_14_14_port, B1 => 
                           n554, B2 => predict_PC_15_14_port, ZN => n828);
   U289 : NAND4_X1 port map( A1 => n825, A2 => n826, A3 => n827, A4 => n828, ZN
                           => n824);
   U309 : AOI22_X1 port map( A1 => n62, A2 => predict_PC_0_13_port, B1 => n61, 
                           B2 => predict_PC_1_13_port, ZN => n839);
   U308 : AOI22_X1 port map( A1 => n64, A2 => predict_PC_2_13_port, B1 => n63, 
                           B2 => predict_PC_3_13_port, ZN => n840);
   U307 : AOI22_X1 port map( A1 => n66, A2 => predict_PC_4_13_port, B1 => n65, 
                           B2 => predict_PC_5_13_port, ZN => n841);
   U306 : AOI22_X1 port map( A1 => n68, A2 => predict_PC_6_13_port, B1 => n67, 
                           B2 => predict_PC_7_13_port, ZN => n842);
   U305 : NAND4_X1 port map( A1 => n839, A2 => n840, A3 => n841, A4 => n842, ZN
                           => n833);
   U304 : AOI22_X1 port map( A1 => n70, A2 => predict_PC_8_13_port, B1 => n69, 
                           B2 => predict_PC_9_13_port, ZN => n835);
   U303 : AOI22_X1 port map( A1 => n557, A2 => predict_PC_10_13_port, B1 => 
                           n558, B2 => predict_PC_11_13_port, ZN => n836);
   U302 : AOI22_X1 port map( A1 => n74, A2 => predict_PC_12_13_port, B1 => n73,
                           B2 => predict_PC_13_13_port, ZN => n837);
   U301 : AOI22_X1 port map( A1 => n553, A2 => predict_PC_14_13_port, B1 => 
                           n554, B2 => predict_PC_15_13_port, ZN => n838);
   U300 : NAND4_X1 port map( A1 => n835, A2 => n836, A3 => n837, A4 => n838, ZN
                           => n834);
   U477 : NAND2_X1 port map( A1 => n978, A2 => n52_port, ZN => n949);
   U465 : NAND2_X1 port map( A1 => n976, A2 => n53_port, ZN => n951);
   U462 : NOR2_X1 port map( A1 => n949, A2 => n951, ZN => N48);
   U469 : NAND2_X1 port map( A1 => n979, A2 => n978, ZN => n945);
   U458 : NOR2_X1 port map( A1 => n945, A2 => n951, ZN => N46);
   U479 : NAND2_X1 port map( A1 => n53_port, A2 => n51_port, ZN => n943);
   U476 : NOR2_X1 port map( A1 => n943, A2 => n949, ZN => N52);
   U456 : NAND2_X1 port map( A1 => n977, A2 => n51_port, ZN => n946);
   U444 : NOR2_X1 port map( A1 => n945, A2 => n946, ZN => N42);
   U448 : NOR2_X1 port map( A1 => n949, A2 => n947, ZN => N40);
   U466 : NAND2_X1 port map( A1 => n52_port, A2 => n50_port, ZN => n944);
   U455 : NOR2_X1 port map( A1 => n944, A2 => n946, ZN => N45);
   U453 : NOR2_X1 port map( A1 => n949, A2 => n946, ZN => N44);
   U464 : NOR2_X1 port map( A1 => n944, A2 => n951, ZN => N49);
   U449 : NOR2_X1 port map( A1 => n948, A2 => n947, ZN => N39);
   U460 : NOR2_X1 port map( A1 => n948, A2 => n951, ZN => N47);
   U447 : NOR2_X1 port map( A1 => n948, A2 => n946, ZN => N43);
   U471 : NOR2_X1 port map( A1 => n943, A2 => n948, ZN => N51);
   U440 : NOR2_X1 port map( A1 => n943, A2 => n944, ZN => N53);
   U450 : NOR2_X1 port map( A1 => n945, A2 => n947, ZN => N38);
   U468 : NOR2_X1 port map( A1 => n943, A2 => n945, ZN => N50);
   U445 : NOR2_X1 port map( A1 => n944, A2 => n947, ZN => N41);
   U355 : NOR2_X1 port map( A1 => stall_i, A2 => reset, ZN => n884);
   U354 : OAI22_X1 port map( A1 => stall_i, A2 => n883, B1 => n884, B2 => n975,
                           ZN => n955);
   U451 : NAND2_X1 port map( A1 => n977, A2 => n976, ZN => n947);
   U472 : NAND2_X1 port map( A1 => n979, A2 => n50_port, ZN => n948);
   U393 : INV_X1 port map( A => TAG_i(1), ZN => n974);
   U394 : INV_X1 port map( A => TAG_i(2), ZN => n973);
   U385 : NAND2_X1 port map( A1 => n903, A2 => n974, ZN => n893);
   U395 : INV_X1 port map( A => TAG_i(3), ZN => n972);
   U372 : NAND2_X1 port map( A1 => n973, A2 => n972, ZN => n896);
   U371 : NOR2_X1 port map( A1 => n895, A2 => n896, ZN => n569);
   U370 : NOR2_X1 port map( A1 => n894, A2 => n896, ZN => n570);
   U368 : NOR2_X1 port map( A1 => n893, A2 => n896, ZN => n571);
   U367 : NOR2_X1 port map( A1 => n891, A2 => n896, ZN => n572);
   U364 : NOR2_X1 port map( A1 => n895, A2 => n892, ZN => n565);
   U363 : NOR2_X1 port map( A1 => n894, A2 => n892, ZN => n566_port);
   U361 : NOR2_X1 port map( A1 => n893, A2 => n892, ZN => n567_port);
   U360 : NOR2_X1 port map( A1 => n891, A2 => n892, ZN => n568);
   U382 : NOR2_X1 port map( A1 => n902, A2 => n891, ZN => n560);
   U397 : OAI21_X1 port map( B1 => was_taken_i, B2 => n54, A => n546, ZN => 
                           n906);
   U373 : AND4_X1 port map( A1 => n897, A2 => n898, A3 => n899, A4 => n900, ZN 
                           => n885);
   U358 : AND4_X1 port map( A1 => n887, A2 => n888, A3 => n889, A4 => n890, ZN 
                           => n886);
   U178 : OR2_X1 port map( A1 => n723, A2 => n724, ZN => 
                           predicted_next_PC_o_23_port);
   U123 : OR2_X1 port map( A1 => n673, A2 => n674, ZN => 
                           predicted_next_PC_o_28_port);
   U101 : OR2_X1 port map( A1 => n653, A2 => n654, ZN => 
                           predicted_next_PC_o_2_port);
   U35 : OR2_X1 port map( A1 => n593, A2 => n594, ZN => 
                           predicted_next_PC_o_6_port);
   U57 : OR2_X1 port map( A1 => n613, A2 => n614, ZN => 
                           predicted_next_PC_o_4_port);
   U46 : OR2_X1 port map( A1 => n603, A2 => n604, ZN => 
                           predicted_next_PC_o_5_port);
   U2 : OR2_X1 port map( A1 => n547, A2 => n548, ZN => 
                           predicted_next_PC_o_9_port);
   U24 : OR2_X1 port map( A1 => n583, A2 => n584, ZN => 
                           predicted_next_PC_o_7_port);
   U13 : OR2_X1 port map( A1 => n573, A2 => n574, ZN => 
                           predicted_next_PC_o_8_port);
   U68 : OR2_X1 port map( A1 => n623, A2 => n624, ZN => 
                           predicted_next_PC_o_3_port);
   U112 : OR2_X1 port map( A1 => n663, A2 => n664, ZN => 
                           predicted_next_PC_o_29_port);
   U90 : OR2_X1 port map( A1 => n643, A2 => n644, ZN => 
                           predicted_next_PC_o_30_port);
   U79 : OR2_X1 port map( A1 => n633, A2 => n634, ZN => 
                           predicted_next_PC_o_31_port);
   U255 : OR2_X1 port map( A1 => n793, A2 => n794, ZN => 
                           predicted_next_PC_o_17_port);
   U222 : OR2_X1 port map( A1 => n763, A2 => n764, ZN => 
                           predicted_next_PC_o_1_port);
   U167 : OR2_X1 port map( A1 => n713, A2 => n714, ZN => 
                           predicted_next_PC_o_24_port);
   U211 : OR2_X1 port map( A1 => n753, A2 => n754, ZN => 
                           predicted_next_PC_o_20_port);
   U145 : OR2_X1 port map( A1 => n693, A2 => n694, ZN => 
                           predicted_next_PC_o_26_port);
   U244 : OR2_X1 port map( A1 => n783, A2 => n784, ZN => 
                           predicted_next_PC_o_18_port);
   U189 : OR2_X1 port map( A1 => n733, A2 => n734, ZN => 
                           predicted_next_PC_o_22_port);
   U200 : OR2_X1 port map( A1 => n743, A2 => n744, ZN => 
                           predicted_next_PC_o_21_port);
   U233 : OR2_X1 port map( A1 => n773, A2 => n774, ZN => 
                           predicted_next_PC_o_19_port);
   U156 : OR2_X1 port map( A1 => n703, A2 => n704, ZN => 
                           predicted_next_PC_o_25_port);
   U134 : OR2_X1 port map( A1 => n683, A2 => n684, ZN => 
                           predicted_next_PC_o_27_port);
   U343 : OR2_X1 port map( A1 => n873, A2 => n874, ZN => 
                           predicted_next_PC_o_0_port);
   U321 : OR2_X1 port map( A1 => n853, A2 => n854, ZN => 
                           predicted_next_PC_o_11_port);
   U310 : OR2_X1 port map( A1 => n843, A2 => n844, ZN => 
                           predicted_next_PC_o_12_port);
   U332 : OR2_X1 port map( A1 => n863, A2 => n864, ZN => 
                           predicted_next_PC_o_10_port);
   U266 : OR2_X1 port map( A1 => n803, A2 => n804, ZN => 
                           predicted_next_PC_o_16_port);
   U277 : OR2_X1 port map( A1 => n813, A2 => n814, ZN => 
                           predicted_next_PC_o_15_port);
   U288 : OR2_X1 port map( A1 => n823, A2 => n824, ZN => 
                           predicted_next_PC_o_14_port);
   U299 : OR2_X1 port map( A1 => n833, A2 => n834, ZN => 
                           predicted_next_PC_o_13_port);
   U475 : INV_X1 port map( A => stall_i, ZN => N567);
   U461 : AND2_X1 port map( A1 => N48, A2 => N567, ZN => N246);
   U457 : AND2_X1 port map( A1 => N46, A2 => N567, ZN => N310);
   U474 : AND2_X1 port map( A1 => N52, A2 => N567, ZN => N118);
   U443 : AND2_X1 port map( A1 => N42, A2 => N567, ZN => N438);
   U441 : AND2_X1 port map( A1 => N40, A2 => N567, ZN => N502);
   U454 : AND2_X1 port map( A1 => N45, A2 => N567, ZN => N342);
   U452 : AND2_X1 port map( A1 => N44, A2 => N567, ZN => N374);
   U463 : AND2_X1 port map( A1 => N49, A2 => N567, ZN => N214);
   U439 : AND2_X1 port map( A1 => N39, A2 => N567, ZN => N534);
   U459 : AND2_X1 port map( A1 => N47, A2 => N567, ZN => N278);
   U446 : AND2_X1 port map( A1 => N43, A2 => N567, ZN => N406);
   U470 : AND2_X1 port map( A1 => N51, A2 => N567, ZN => N150);
   U436 : AND2_X1 port map( A1 => N53, A2 => N567, ZN => N86);
   U438 : AND2_X1 port map( A1 => N38, A2 => N567, ZN => N566);
   U467 : AND2_X1 port map( A1 => N50, A2 => N567, ZN => N182);
   U442 : AND2_X1 port map( A1 => N41, A2 => N567, ZN => N470);
   U356 : INV_X1 port map( A => taken_o_port, ZN => n883);
   last_PC_reg_16_inst : DFFR_X1 port map( D => predicted_next_PC_o_16_port, CK
                           => net3621, RN => n99, Q => n33, QN => n513);
   last_PC_reg_15_inst : DFFR_X1 port map( D => predicted_next_PC_o_15_port, CK
                           => net3621, RN => n94, Q => n32, QN => n515);
   last_PC_reg_14_inst : DFFR_X1 port map( D => predicted_next_PC_o_14_port, CK
                           => net3621, RN => n96, Q => n31, QN => n517);
   last_PC_reg_13_inst : DFFR_X1 port map( D => predicted_next_PC_o_13_port, CK
                           => net3621, RN => n99, Q => n30, QN => n519);
   last_PC_reg_12_inst : DFFR_X1 port map( D => predicted_next_PC_o_12_port, CK
                           => net3621, RN => n96, Q => n29, QN => n521);
   last_PC_reg_11_inst : DFFR_X1 port map( D => predicted_next_PC_o_11_port, CK
                           => net3621, RN => n96, Q => n28, QN => n523);
   last_PC_reg_10_inst : DFFR_X1 port map( D => predicted_next_PC_o_10_port, CK
                           => net3621, RN => n86_port, Q => n27, QN => n525);
   last_PC_reg_0_inst : DFFR_X1 port map( D => predicted_next_PC_o_0_port, CK 
                           => net3621, RN => n97, Q => n26, QN => n545);
   last_PC_reg_28_inst : DFFR_X1 port map( D => predicted_next_PC_o_28_port, CK
                           => net3621, RN => n90, Q => n25, QN => n489);
   last_PC_reg_23_inst : DFFR_X1 port map( D => predicted_next_PC_o_23_port, CK
                           => net3621, RN => n86_port, Q => n24, QN => n499);
   last_PC_reg_31_inst : DFFR_X1 port map( D => predicted_next_PC_o_31_port, CK
                           => net3621, RN => n83, Q => n23, QN => n483);
   last_PC_reg_30_inst : DFFR_X1 port map( D => predicted_next_PC_o_30_port, CK
                           => net3621, RN => n96, Q => n22, QN => n485);
   last_PC_reg_29_inst : DFFR_X1 port map( D => predicted_next_PC_o_29_port, CK
                           => net3621, RN => n91, Q => n21, QN => n487);
   last_PC_reg_27_inst : DFFR_X1 port map( D => predicted_next_PC_o_27_port, CK
                           => net3621, RN => n100, Q => n20, QN => n491);
   last_PC_reg_26_inst : DFFR_X1 port map( D => predicted_next_PC_o_26_port, CK
                           => net3621, RN => n86_port, Q => n19, QN => n493);
   last_PC_reg_25_inst : DFFR_X1 port map( D => predicted_next_PC_o_25_port, CK
                           => net3621, RN => n100, Q => n18, QN => n495);
   last_PC_reg_24_inst : DFFR_X1 port map( D => predicted_next_PC_o_24_port, CK
                           => net3621, RN => n97, Q => n17, QN => n497);
   last_PC_reg_22_inst : DFFR_X1 port map( D => predicted_next_PC_o_22_port, CK
                           => net3621, RN => n96, Q => n16, QN => n501);
   last_PC_reg_21_inst : DFFR_X1 port map( D => predicted_next_PC_o_21_port, CK
                           => net3621, RN => n90, Q => n15, QN => n503);
   last_PC_reg_20_inst : DFFR_X1 port map( D => predicted_next_PC_o_20_port, CK
                           => net3621, RN => n93, Q => n14, QN => n505);
   last_PC_reg_19_inst : DFFR_X1 port map( D => predicted_next_PC_o_19_port, CK
                           => net3621, RN => n95, Q => n13, QN => n507);
   last_PC_reg_18_inst : DFFR_X1 port map( D => predicted_next_PC_o_18_port, CK
                           => net3621, RN => n87, Q => n12, QN => n509);
   last_PC_reg_17_inst : DFFR_X1 port map( D => predicted_next_PC_o_17_port, CK
                           => net3621, RN => n89, Q => n11, QN => n511);
   last_PC_reg_9_inst : DFFR_X1 port map( D => predicted_next_PC_o_9_port, CK 
                           => net3621, RN => n100, Q => n10, QN => n527);
   last_PC_reg_8_inst : DFFR_X1 port map( D => predicted_next_PC_o_8_port, CK 
                           => net3621, RN => n96, Q => n9, QN => n529);
   last_PC_reg_7_inst : DFFR_X1 port map( D => predicted_next_PC_o_7_port, CK 
                           => net3621, RN => n89, Q => n8, QN => n531);
   last_PC_reg_6_inst : DFFR_X1 port map( D => predicted_next_PC_o_6_port, CK 
                           => net3621, RN => n94, Q => n7, QN => n533);
   last_PC_reg_5_inst : DFFR_X1 port map( D => predicted_next_PC_o_5_port, CK 
                           => net3621, RN => n87, Q => n6, QN => n535);
   last_PC_reg_4_inst : DFFR_X1 port map( D => predicted_next_PC_o_4_port, CK 
                           => net3621, RN => n88, Q => n5, QN => n537);
   last_PC_reg_3_inst : DFFR_X1 port map( D => predicted_next_PC_o_3_port, CK 
                           => net3621, RN => n87, Q => n4, QN => n539);
   last_PC_reg_2_inst : DFFR_X1 port map( D => predicted_next_PC_o_2_port, CK 
                           => net3621, RN => n97, Q => n3, QN => n541);
   last_PC_reg_1_inst : DFFR_X1 port map( D => predicted_next_PC_o_1_port, CK 
                           => net3621, RN => n98, Q => n2, QN => n543);
   last_mispredict_reg : DFFR_X1 port map( D => mispredict_o_port, CK => 
                           net3621, RN => n95, Q => n1, QN => n546);
   U357 : AOI21_X2 port map( B1 => n905, B2 => n54, A => n906, ZN => 
                           mispredict_o_port);
   U375 : AND4_X2 port map( A1 => n46_port, A2 => n47_port, A3 => n48_port, A4 
                           => n49_port, ZN => n905);
   U376 : NOR2_X1 port map( A1 => n895, A2 => n901, ZN => n553);
   U378 : BUF_X1 port map( A => target_PC_i(29), Z => n58);
   U379 : BUF_X1 port map( A => target_PC_i(28), Z => n39_port);
   U383 : BUF_X1 port map( A => target_PC_i(27), Z => n60);
   U384 : BUF_X1 port map( A => n560, Z => n69);
   U387 : BUF_X2 port map( A => n569, Z => n64);
   U388 : BUF_X2 port map( A => n559, Z => n70);
   U389 : BUF_X1 port map( A => n557, Z => n72);
   U392 : BUF_X1 port map( A => n558, Z => n71);
   U396 : BUF_X2 port map( A => n555, Z => n74);
   U398 : BUF_X2 port map( A => n556, Z => n73);
   U399 : BUF_X1 port map( A => n553, Z => n76);
   U400 : BUF_X1 port map( A => n568, Z => n65);
   U401 : BUF_X2 port map( A => n567_port, Z => n66);
   U402 : BUF_X1 port map( A => n566_port, Z => n67);
   U403 : BUF_X2 port map( A => n565, Z => n68);
   U404 : BUF_X1 port map( A => n572, Z => n61);
   U405 : BUF_X2 port map( A => n571, Z => n62);
   U406 : BUF_X1 port map( A => n570, Z => n63);
   U407 : BUF_X1 port map( A => n554, Z => n75);
   U408 : BUF_X1 port map( A => target_PC_i(25), Z => n35);
   U409 : BUF_X1 port map( A => target_PC_i(24), Z => n36);
   U410 : BUF_X1 port map( A => target_PC_i(26), Z => n37);
   U411 : CLKBUF_X1 port map( A => target_PC_i(30), Z => n38_port);
   U412 : AND2_X1 port map( A1 => target_PC_i(15), A2 => n515, ZN => n40_port);
   U413 : AND2_X1 port map( A1 => n517, A2 => target_PC_i(14), ZN => n41_port);
   U414 : NOR3_X1 port map( A1 => n40_port, A2 => n41_port, A3 => n933, ZN => 
                           n928);
   U415 : AND2_X1 port map( A1 => target_PC_i(13), A2 => n519, ZN => n42_port);
   U416 : AND2_X1 port map( A1 => n521, A2 => target_PC_i(12), ZN => n43_port);
   U417 : NOR3_X1 port map( A1 => n42_port, A2 => n43_port, A3 => n932, ZN => 
                           n929);
   U418 : AND2_X1 port map( A1 => target_PC_i(11), A2 => n523, ZN => n44_port);
   U419 : AND2_X1 port map( A1 => target_PC_i(10), A2 => n525, ZN => n45_port);
   U420 : NOR3_X1 port map( A1 => n44_port, A2 => n45_port, A3 => n939, ZN => 
                           n938);
   U421 : AND4_X1 port map( A1 => n935, A2 => n936, A3 => n937, A4 => n938, ZN 
                           => n46_port);
   U422 : AND4_X1 port map( A1 => n913, A2 => n912, A3 => n914, A4 => n911, ZN 
                           => n47_port);
   U423 : AND4_X1 port map( A1 => n919, A2 => n922, A3 => n921, A4 => n920, ZN 
                           => n48_port);
   U424 : AND4_X1 port map( A1 => n927, A2 => n928, A3 => n929, A4 => n930, ZN 
                           => n49_port);
   U425 : INV_X1 port map( A => reset, ZN => n97);
   U426 : INV_X1 port map( A => reset, ZN => n98);
   U427 : INV_X1 port map( A => reset, ZN => n95);
   U431 : INV_X1 port map( A => reset, ZN => n96);
   U432 : INV_X1 port map( A => reset, ZN => n99);
   U433 : INV_X1 port map( A => reset, ZN => n100);
   U434 : INV_X1 port map( A => reset, ZN => n94);
   U435 : INV_X1 port map( A => reset, ZN => n92);
   U437 : INV_X1 port map( A => reset, ZN => n93);
   U473 : INV_X1 port map( A => reset, ZN => n88);
   U478 : INV_X1 port map( A => reset, ZN => n89);
   U480 : INV_X1 port map( A => reset, ZN => n90);
   U481 : INV_X1 port map( A => reset, ZN => n91);
   U482 : INV_X1 port map( A => reset, ZN => n84);
   U483 : INV_X1 port map( A => reset, ZN => n80);
   U484 : INV_X1 port map( A => reset, ZN => n81);
   U485 : INV_X1 port map( A => reset, ZN => n82);
   U486 : INV_X1 port map( A => reset, ZN => n83);
   U487 : INV_X1 port map( A => reset, ZN => n77);
   U488 : INV_X1 port map( A => reset, ZN => n78);
   U489 : INV_X1 port map( A => reset, ZN => n79);
   U490 : INV_X1 port map( A => reset, ZN => n87);
   U491 : INV_X1 port map( A => reset, ZN => n85);
   U492 : INV_X1 port map( A => reset, ZN => n86_port);
   U493 : CLKBUF_X1 port map( A => target_PC_i(31), Z => n59);
   U494 : AND3_X1 port map( A1 => n55, A2 => n56, A3 => n57, ZN => n911);
   U495 : INV_X1 port map( A => n918, ZN => n57);
   U496 : AOI21_X1 port map( B1 => n885, B2 => n886, A => reset, ZN => 
                           taken_o_port);
   U497 : INV_X1 port map( A => TAG_i(0), ZN => n903);
   U498 : NOR2_X1 port map( A1 => n902, A2 => n893, ZN => n559);
   U499 : NOR2_X1 port map( A1 => n895, A2 => n902, ZN => n557);
   U500 : NOR2_X1 port map( A1 => n893, A2 => n901, ZN => n555);
   U501 : NOR2_X1 port map( A1 => n902, A2 => n894, ZN => n558);
   U502 : NOR2_X1 port map( A1 => n894, A2 => n901, ZN => n554);
   U503 : NOR2_X1 port map( A1 => n891, A2 => n901, ZN => n556);
   U504 : OAI22_X1 port map( A1 => target_PC_i(29), A2 => n487, B1 => 
                           target_PC_i(28), B2 => n489, ZN => n942);
   U505 : OAI22_X1 port map( A1 => target_PC_i(31), A2 => n483, B1 => 
                           target_PC_i(30), B2 => n485, ZN => n918);
   U506 : OAI22_X1 port map( A1 => target_PC_i(3), A2 => n539, B1 => 
                           target_PC_i(2), B2 => n541, ZN => n931);
   U507 : OAI22_X1 port map( A1 => target_PC_i(13), A2 => n519, B1 => 
                           target_PC_i(12), B2 => n521, ZN => n932);
   U508 : OAI22_X1 port map( A1 => target_PC_i(15), A2 => n515, B1 => 
                           target_PC_i(14), B2 => n517, ZN => n933);
   U509 : OAI22_X1 port map( A1 => target_PC_i(9), A2 => n527, B1 => 
                           target_PC_i(8), B2 => n529, ZN => n934);
   U510 : OAI22_X1 port map( A1 => target_PC_i(23), A2 => n499, B1 => 
                           target_PC_i(22), B2 => n501, ZN => n923);
   U511 : OAI22_X1 port map( A1 => target_PC_i(5), A2 => n535, B1 => 
                           target_PC_i(4), B2 => n537, ZN => n924);
   U512 : OAI22_X1 port map( A1 => target_PC_i(7), A2 => n531, B1 => 
                           target_PC_i(6), B2 => n533, ZN => n925);
   U513 : OAI22_X1 port map( A1 => target_PC_i(1), A2 => n543, B1 => 
                           target_PC_i(0), B2 => n545, ZN => n926);
   U514 : OAI22_X1 port map( A1 => target_PC_i(21), A2 => n503, B1 => 
                           target_PC_i(20), B2 => n505, ZN => n915);
   U515 : OAI22_X1 port map( A1 => target_PC_i(25), A2 => n495, B1 => 
                           target_PC_i(24), B2 => n497, ZN => n916);
   U516 : OAI22_X1 port map( A1 => target_PC_i(27), A2 => n491, B1 => 
                           target_PC_i(26), B2 => n493, ZN => n917);
   U517 : NAND2_X1 port map( A1 => n485, A2 => target_PC_i(30), ZN => n56);
   U518 : NAND2_X1 port map( A1 => target_PC_i(31), A2 => n483, ZN => n55);
   U519 : OAI22_X1 port map( A1 => target_PC_i(19), A2 => n507, B1 => 
                           target_PC_i(18), B2 => n509, ZN => n941);
   U520 : AOI221_X1 port map( B1 => target_PC_i(3), B2 => n539, C1 => n541, C2 
                           => target_PC_i(2), A => n931, ZN => n930);
   U521 : AOI221_X1 port map( B1 => target_PC_i(9), B2 => n527, C1 => 
                           target_PC_i(8), C2 => n529, A => n934, ZN => n927);
   U522 : AOI221_X1 port map( B1 => target_PC_i(23), B2 => n499, C1 => n501, C2
                           => target_PC_i(22), A => n923, ZN => n922);
   U523 : AOI221_X1 port map( B1 => target_PC_i(5), B2 => n535, C1 => n537, C2 
                           => target_PC_i(4), A => n924, ZN => n921);
   U524 : AOI221_X1 port map( B1 => target_PC_i(7), B2 => n531, C1 => n533, C2 
                           => target_PC_i(6), A => n925, ZN => n920);
   U525 : AOI221_X1 port map( B1 => target_PC_i(1), B2 => n543, C1 => n545, C2 
                           => target_PC_i(0), A => n926, ZN => n919);
   U526 : AOI221_X1 port map( B1 => target_PC_i(21), B2 => n503, C1 => n505, C2
                           => target_PC_i(20), A => n915, ZN => n914);
   U527 : AOI221_X1 port map( B1 => target_PC_i(25), B2 => n495, C1 => n497, C2
                           => target_PC_i(24), A => n916, ZN => n913);
   U528 : AOI221_X1 port map( B1 => target_PC_i(27), B2 => n491, C1 => n493, C2
                           => target_PC_i(26), A => n917, ZN => n912);
   U529 : AOI221_X1 port map( B1 => target_PC_i(19), B2 => n507, C1 => n509, C2
                           => target_PC_i(18), A => n941, ZN => n936);
   U530 : AOI221_X1 port map( B1 => target_PC_i(29), B2 => n487, C1 => n489, C2
                           => target_PC_i(28), A => n942, ZN => n935);
   U531 : NAND2_X1 port map( A1 => TAG_i(0), A2 => TAG_i(1), ZN => n894);
   U532 : NAND2_X1 port map( A1 => TAG_i(0), A2 => n974, ZN => n891);

end SYN_bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity fetch_block is

   port( branch_target_i, sum_addr_i, A_i, NPC4_i : in std_logic_vector (31 
         downto 0);  S_MUX_PC_BUS_i : in std_logic_vector (1 downto 0);  PC_o, 
         PC4_o, PC_BUS_pre_BTB : out std_logic_vector (31 downto 0);  stall_i, 
         take_prediction_i, mispredict_i : in std_logic;  predicted_PC : in 
         std_logic_vector (31 downto 0);  clk, rst : in std_logic);

end fetch_block;

architecture SYN_Struct of fetch_block is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component mux41_1
      port( IN0, IN1, IN2, IN3 : in std_logic_vector (31 downto 0);  CTRL : in 
            std_logic_vector (1 downto 0);  OUT1 : out std_logic_vector (31 
            downto 0));
   end component;
   
   component mux41_0
      port( IN0, IN1, IN2, IN3 : in std_logic_vector (31 downto 0);  CTRL : in 
            std_logic_vector (1 downto 0);  OUT1 : out std_logic_vector (31 
            downto 0));
   end component;
   
   component add4
      port( IN1 : in std_logic_vector (31 downto 0);  OUT1 : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component ff32_en_0
      port( D : in std_logic_vector (31 downto 0);  en, clk, rst : in std_logic
            ;  Q : out std_logic_vector (31 downto 0));
   end component;
   
   signal PC_o_31_port, PC_o_30_port, PC_o_29_port, PC_o_28_port, PC_o_27_port,
      PC_o_26_port, PC_o_25_port, PC_o_24_port, PC_o_23_port, PC_o_22_port, 
      PC_o_21_port, PC_o_20_port, PC_o_19_port, PC_o_18_port, PC_o_17_port, 
      PC_o_16_port, PC_o_15_port, PC_o_14_port, PC_o_13_port, PC_o_12_port, 
      PC_o_11_port, PC_o_10_port, PC_o_9_port, PC_o_8_port, PC_o_7_port, 
      PC_o_6_port, PC_o_5_port, PC_o_4_port, PC_o_3_port, PC_o_2_port, 
      PC_o_1_port, PC_o_0_port, PC4_o_31_port, PC4_o_30_port, PC4_o_29_port, 
      PC4_o_28_port, PC4_o_27_port, PC4_o_26_port, PC4_o_25_port, PC4_o_24_port
      , PC4_o_23_port, PC4_o_22_port, PC4_o_21_port, PC4_o_20_port, 
      PC4_o_19_port, PC4_o_18_port, PC4_o_17_port, PC4_o_16_port, PC4_o_15_port
      , PC4_o_14_port, PC4_o_13_port, PC4_o_12_port, PC4_o_11_port, 
      PC4_o_10_port, PC4_o_9_port, PC4_o_8_port, PC4_o_7_port, PC4_o_6_port, 
      PC4_o_5_port, PC4_o_4_port, PC4_o_3_port, PC4_o_2_port, PC4_o_1_port, 
      PC4_o_0_port, PC_BUS_pre_BTB_31_port, PC_BUS_pre_BTB_30_port, 
      PC_BUS_pre_BTB_28_port, PC_BUS_pre_BTB_27_port, PC_BUS_pre_BTB_26_port, 
      PC_BUS_pre_BTB_25_port, PC_BUS_pre_BTB_24_port, PC_BUS_pre_BTB_23_port, 
      PC_BUS_pre_BTB_22_port, PC_BUS_pre_BTB_21_port, PC_BUS_pre_BTB_20_port, 
      PC_BUS_pre_BTB_19_port, PC_BUS_pre_BTB_18_port, PC_BUS_pre_BTB_17_port, 
      PC_BUS_pre_BTB_16_port, PC_BUS_pre_BTB_15_port, PC_BUS_pre_BTB_14_port, 
      PC_BUS_pre_BTB_13_port, PC_BUS_pre_BTB_12_port, PC_BUS_pre_BTB_11_port, 
      PC_BUS_pre_BTB_10_port, PC_BUS_pre_BTB_9_port, PC_BUS_pre_BTB_8_port, 
      PC_BUS_pre_BTB_7_port, PC_BUS_pre_BTB_6_port, PC_BUS_pre_BTB_5_port, 
      PC_BUS_pre_BTB_4_port, PC_BUS_pre_BTB_3_port, PC_BUS_pre_BTB_2_port, 
      PC_BUS_pre_BTB_1_port, PC_BUS_pre_BTB_0_port, en_IR, PC_BUS_31_port, 
      PC_BUS_30_port, PC_BUS_29_port, PC_BUS_28_port, PC_BUS_27_port, 
      PC_BUS_26_port, PC_BUS_25_port, PC_BUS_24_port, PC_BUS_23_port, 
      PC_BUS_22_port, PC_BUS_21_port, PC_BUS_20_port, PC_BUS_19_port, 
      PC_BUS_18_port, PC_BUS_17_port, PC_BUS_16_port, PC_BUS_15_port, 
      PC_BUS_14_port, PC_BUS_13_port, PC_BUS_12_port, PC_BUS_11_port, 
      PC_BUS_10_port, PC_BUS_9_port, PC_BUS_8_port, PC_BUS_7_port, 
      PC_BUS_6_port, PC_BUS_5_port, PC_BUS_4_port, PC_BUS_3_port, PC_BUS_2_port
      , PC_BUS_1_port, PC_BUS_0_port, n1, PC_BUS_pre_BTB_29_port : std_logic;

begin
   PC_o <= ( PC_o_31_port, PC_o_30_port, PC_o_29_port, PC_o_28_port, 
      PC_o_27_port, PC_o_26_port, PC_o_25_port, PC_o_24_port, PC_o_23_port, 
      PC_o_22_port, PC_o_21_port, PC_o_20_port, PC_o_19_port, PC_o_18_port, 
      PC_o_17_port, PC_o_16_port, PC_o_15_port, PC_o_14_port, PC_o_13_port, 
      PC_o_12_port, PC_o_11_port, PC_o_10_port, PC_o_9_port, PC_o_8_port, 
      PC_o_7_port, PC_o_6_port, PC_o_5_port, PC_o_4_port, PC_o_3_port, 
      PC_o_2_port, PC_o_1_port, PC_o_0_port );
   PC4_o <= ( PC4_o_31_port, PC4_o_30_port, PC4_o_29_port, PC4_o_28_port, 
      PC4_o_27_port, PC4_o_26_port, PC4_o_25_port, PC4_o_24_port, PC4_o_23_port
      , PC4_o_22_port, PC4_o_21_port, PC4_o_20_port, PC4_o_19_port, 
      PC4_o_18_port, PC4_o_17_port, PC4_o_16_port, PC4_o_15_port, PC4_o_14_port
      , PC4_o_13_port, PC4_o_12_port, PC4_o_11_port, PC4_o_10_port, 
      PC4_o_9_port, PC4_o_8_port, PC4_o_7_port, PC4_o_6_port, PC4_o_5_port, 
      PC4_o_4_port, PC4_o_3_port, PC4_o_2_port, PC4_o_1_port, PC4_o_0_port );
   PC_BUS_pre_BTB <= ( PC_BUS_pre_BTB_31_port, PC_BUS_pre_BTB_30_port, 
      PC_BUS_pre_BTB_29_port, PC_BUS_pre_BTB_28_port, PC_BUS_pre_BTB_27_port, 
      PC_BUS_pre_BTB_26_port, PC_BUS_pre_BTB_25_port, PC_BUS_pre_BTB_24_port, 
      PC_BUS_pre_BTB_23_port, PC_BUS_pre_BTB_22_port, PC_BUS_pre_BTB_21_port, 
      PC_BUS_pre_BTB_20_port, PC_BUS_pre_BTB_19_port, PC_BUS_pre_BTB_18_port, 
      PC_BUS_pre_BTB_17_port, PC_BUS_pre_BTB_16_port, PC_BUS_pre_BTB_15_port, 
      PC_BUS_pre_BTB_14_port, PC_BUS_pre_BTB_13_port, PC_BUS_pre_BTB_12_port, 
      PC_BUS_pre_BTB_11_port, PC_BUS_pre_BTB_10_port, PC_BUS_pre_BTB_9_port, 
      PC_BUS_pre_BTB_8_port, PC_BUS_pre_BTB_7_port, PC_BUS_pre_BTB_6_port, 
      PC_BUS_pre_BTB_5_port, PC_BUS_pre_BTB_4_port, PC_BUS_pre_BTB_3_port, 
      PC_BUS_pre_BTB_2_port, PC_BUS_pre_BTB_1_port, PC_BUS_pre_BTB_0_port );
   
   PC : ff32_en_0 port map( D(31) => PC_BUS_31_port, D(30) => PC_BUS_30_port, 
                           D(29) => PC_BUS_29_port, D(28) => PC_BUS_28_port, 
                           D(27) => PC_BUS_27_port, D(26) => PC_BUS_26_port, 
                           D(25) => PC_BUS_25_port, D(24) => PC_BUS_24_port, 
                           D(23) => PC_BUS_23_port, D(22) => PC_BUS_22_port, 
                           D(21) => PC_BUS_21_port, D(20) => PC_BUS_20_port, 
                           D(19) => PC_BUS_19_port, D(18) => PC_BUS_18_port, 
                           D(17) => PC_BUS_17_port, D(16) => PC_BUS_16_port, 
                           D(15) => PC_BUS_15_port, D(14) => PC_BUS_14_port, 
                           D(13) => PC_BUS_13_port, D(12) => PC_BUS_12_port, 
                           D(11) => PC_BUS_11_port, D(10) => PC_BUS_10_port, 
                           D(9) => PC_BUS_9_port, D(8) => PC_BUS_8_port, D(7) 
                           => PC_BUS_7_port, D(6) => PC_BUS_6_port, D(5) => 
                           PC_BUS_5_port, D(4) => PC_BUS_4_port, D(3) => 
                           PC_BUS_3_port, D(2) => PC_BUS_2_port, D(1) => 
                           PC_BUS_1_port, D(0) => PC_BUS_0_port, en => en_IR, 
                           clk => clk, rst => rst, Q(31) => PC_o_31_port, Q(30)
                           => PC_o_30_port, Q(29) => PC_o_29_port, Q(28) => 
                           PC_o_28_port, Q(27) => PC_o_27_port, Q(26) => 
                           PC_o_26_port, Q(25) => PC_o_25_port, Q(24) => 
                           PC_o_24_port, Q(23) => PC_o_23_port, Q(22) => 
                           PC_o_22_port, Q(21) => PC_o_21_port, Q(20) => 
                           PC_o_20_port, Q(19) => PC_o_19_port, Q(18) => 
                           PC_o_18_port, Q(17) => PC_o_17_port, Q(16) => 
                           PC_o_16_port, Q(15) => PC_o_15_port, Q(14) => 
                           PC_o_14_port, Q(13) => PC_o_13_port, Q(12) => 
                           PC_o_12_port, Q(11) => PC_o_11_port, Q(10) => 
                           PC_o_10_port, Q(9) => PC_o_9_port, Q(8) => 
                           PC_o_8_port, Q(7) => PC_o_7_port, Q(6) => 
                           PC_o_6_port, Q(5) => PC_o_5_port, Q(4) => 
                           PC_o_4_port, Q(3) => PC_o_3_port, Q(2) => 
                           PC_o_2_port, Q(1) => PC_o_1_port, Q(0) => 
                           PC_o_0_port);
   PCADD : add4 port map( IN1(31) => PC_o_31_port, IN1(30) => PC_o_30_port, 
                           IN1(29) => PC_o_29_port, IN1(28) => PC_o_28_port, 
                           IN1(27) => PC_o_27_port, IN1(26) => PC_o_26_port, 
                           IN1(25) => PC_o_25_port, IN1(24) => PC_o_24_port, 
                           IN1(23) => PC_o_23_port, IN1(22) => PC_o_22_port, 
                           IN1(21) => PC_o_21_port, IN1(20) => PC_o_20_port, 
                           IN1(19) => PC_o_19_port, IN1(18) => PC_o_18_port, 
                           IN1(17) => PC_o_17_port, IN1(16) => PC_o_16_port, 
                           IN1(15) => PC_o_15_port, IN1(14) => PC_o_14_port, 
                           IN1(13) => PC_o_13_port, IN1(12) => PC_o_12_port, 
                           IN1(11) => PC_o_11_port, IN1(10) => PC_o_10_port, 
                           IN1(9) => PC_o_9_port, IN1(8) => PC_o_8_port, IN1(7)
                           => PC_o_7_port, IN1(6) => PC_o_6_port, IN1(5) => 
                           PC_o_5_port, IN1(4) => PC_o_4_port, IN1(3) => 
                           PC_o_3_port, IN1(2) => PC_o_2_port, IN1(1) => 
                           PC_o_1_port, IN1(0) => PC_o_0_port, OUT1(31) => 
                           PC4_o_31_port, OUT1(30) => PC4_o_30_port, OUT1(29) 
                           => PC4_o_29_port, OUT1(28) => PC4_o_28_port, 
                           OUT1(27) => PC4_o_27_port, OUT1(26) => PC4_o_26_port
                           , OUT1(25) => PC4_o_25_port, OUT1(24) => 
                           PC4_o_24_port, OUT1(23) => PC4_o_23_port, OUT1(22) 
                           => PC4_o_22_port, OUT1(21) => PC4_o_21_port, 
                           OUT1(20) => PC4_o_20_port, OUT1(19) => PC4_o_19_port
                           , OUT1(18) => PC4_o_18_port, OUT1(17) => 
                           PC4_o_17_port, OUT1(16) => PC4_o_16_port, OUT1(15) 
                           => PC4_o_15_port, OUT1(14) => PC4_o_14_port, 
                           OUT1(13) => PC4_o_13_port, OUT1(12) => PC4_o_12_port
                           , OUT1(11) => PC4_o_11_port, OUT1(10) => 
                           PC4_o_10_port, OUT1(9) => PC4_o_9_port, OUT1(8) => 
                           PC4_o_8_port, OUT1(7) => PC4_o_7_port, OUT1(6) => 
                           PC4_o_6_port, OUT1(5) => PC4_o_5_port, OUT1(4) => 
                           PC4_o_4_port, OUT1(3) => PC4_o_3_port, OUT1(2) => 
                           PC4_o_2_port, OUT1(1) => PC4_o_1_port, OUT1(0) => 
                           PC4_o_0_port);
   MUXTARGET : mux41_0 port map( IN0(31) => NPC4_i(31), IN0(30) => NPC4_i(30), 
                           IN0(29) => NPC4_i(29), IN0(28) => NPC4_i(28), 
                           IN0(27) => NPC4_i(27), IN0(26) => NPC4_i(26), 
                           IN0(25) => NPC4_i(25), IN0(24) => NPC4_i(24), 
                           IN0(23) => NPC4_i(23), IN0(22) => NPC4_i(22), 
                           IN0(21) => NPC4_i(21), IN0(20) => NPC4_i(20), 
                           IN0(19) => NPC4_i(19), IN0(18) => NPC4_i(18), 
                           IN0(17) => NPC4_i(17), IN0(16) => NPC4_i(16), 
                           IN0(15) => NPC4_i(15), IN0(14) => NPC4_i(14), 
                           IN0(13) => NPC4_i(13), IN0(12) => NPC4_i(12), 
                           IN0(11) => NPC4_i(11), IN0(10) => NPC4_i(10), IN0(9)
                           => NPC4_i(9), IN0(8) => NPC4_i(8), IN0(7) => 
                           NPC4_i(7), IN0(6) => NPC4_i(6), IN0(5) => NPC4_i(5),
                           IN0(4) => NPC4_i(4), IN0(3) => NPC4_i(3), IN0(2) => 
                           NPC4_i(2), IN0(1) => NPC4_i(1), IN0(0) => NPC4_i(0),
                           IN1(31) => A_i(31), IN1(30) => A_i(30), IN1(29) => 
                           A_i(29), IN1(28) => A_i(28), IN1(27) => A_i(27), 
                           IN1(26) => A_i(26), IN1(25) => A_i(25), IN1(24) => 
                           A_i(24), IN1(23) => A_i(23), IN1(22) => A_i(22), 
                           IN1(21) => A_i(21), IN1(20) => A_i(20), IN1(19) => 
                           A_i(19), IN1(18) => A_i(18), IN1(17) => A_i(17), 
                           IN1(16) => A_i(16), IN1(15) => A_i(15), IN1(14) => 
                           A_i(14), IN1(13) => A_i(13), IN1(12) => A_i(12), 
                           IN1(11) => A_i(11), IN1(10) => A_i(10), IN1(9) => 
                           A_i(9), IN1(8) => A_i(8), IN1(7) => A_i(7), IN1(6) 
                           => A_i(6), IN1(5) => A_i(5), IN1(4) => A_i(4), 
                           IN1(3) => A_i(3), IN1(2) => A_i(2), IN1(1) => A_i(1)
                           , IN1(0) => A_i(0), IN2(31) => sum_addr_i(31), 
                           IN2(30) => sum_addr_i(30), IN2(29) => sum_addr_i(29)
                           , IN2(28) => sum_addr_i(28), IN2(27) => 
                           sum_addr_i(27), IN2(26) => sum_addr_i(26), IN2(25) 
                           => sum_addr_i(25), IN2(24) => sum_addr_i(24), 
                           IN2(23) => sum_addr_i(23), IN2(22) => sum_addr_i(22)
                           , IN2(21) => sum_addr_i(21), IN2(20) => 
                           sum_addr_i(20), IN2(19) => sum_addr_i(19), IN2(18) 
                           => sum_addr_i(18), IN2(17) => sum_addr_i(17), 
                           IN2(16) => sum_addr_i(16), IN2(15) => sum_addr_i(15)
                           , IN2(14) => sum_addr_i(14), IN2(13) => 
                           sum_addr_i(13), IN2(12) => sum_addr_i(12), IN2(11) 
                           => sum_addr_i(11), IN2(10) => sum_addr_i(10), IN2(9)
                           => sum_addr_i(9), IN2(8) => sum_addr_i(8), IN2(7) =>
                           sum_addr_i(7), IN2(6) => sum_addr_i(6), IN2(5) => 
                           sum_addr_i(5), IN2(4) => sum_addr_i(4), IN2(3) => 
                           sum_addr_i(3), IN2(2) => sum_addr_i(2), IN2(1) => 
                           sum_addr_i(1), IN2(0) => sum_addr_i(0), IN3(31) => 
                           branch_target_i(31), IN3(30) => branch_target_i(30),
                           IN3(29) => branch_target_i(29), IN3(28) => 
                           branch_target_i(28), IN3(27) => branch_target_i(27),
                           IN3(26) => branch_target_i(26), IN3(25) => 
                           branch_target_i(25), IN3(24) => branch_target_i(24),
                           IN3(23) => branch_target_i(23), IN3(22) => 
                           branch_target_i(22), IN3(21) => branch_target_i(21),
                           IN3(20) => branch_target_i(20), IN3(19) => 
                           branch_target_i(19), IN3(18) => branch_target_i(18),
                           IN3(17) => branch_target_i(17), IN3(16) => 
                           branch_target_i(16), IN3(15) => branch_target_i(15),
                           IN3(14) => branch_target_i(14), IN3(13) => 
                           branch_target_i(13), IN3(12) => branch_target_i(12),
                           IN3(11) => branch_target_i(11), IN3(10) => 
                           branch_target_i(10), IN3(9) => branch_target_i(9), 
                           IN3(8) => branch_target_i(8), IN3(7) => 
                           branch_target_i(7), IN3(6) => branch_target_i(6), 
                           IN3(5) => branch_target_i(5), IN3(4) => 
                           branch_target_i(4), IN3(3) => branch_target_i(3), 
                           IN3(2) => branch_target_i(2), IN3(1) => 
                           branch_target_i(1), IN3(0) => branch_target_i(0), 
                           CTRL(1) => S_MUX_PC_BUS_i(1), CTRL(0) => 
                           S_MUX_PC_BUS_i(0), OUT1(31) => 
                           PC_BUS_pre_BTB_31_port, OUT1(30) => 
                           PC_BUS_pre_BTB_30_port, OUT1(29) => 
                           PC_BUS_pre_BTB_29_port, OUT1(28) => 
                           PC_BUS_pre_BTB_28_port, OUT1(27) => 
                           PC_BUS_pre_BTB_27_port, OUT1(26) => 
                           PC_BUS_pre_BTB_26_port, OUT1(25) => 
                           PC_BUS_pre_BTB_25_port, OUT1(24) => 
                           PC_BUS_pre_BTB_24_port, OUT1(23) => 
                           PC_BUS_pre_BTB_23_port, OUT1(22) => 
                           PC_BUS_pre_BTB_22_port, OUT1(21) => 
                           PC_BUS_pre_BTB_21_port, OUT1(20) => 
                           PC_BUS_pre_BTB_20_port, OUT1(19) => 
                           PC_BUS_pre_BTB_19_port, OUT1(18) => 
                           PC_BUS_pre_BTB_18_port, OUT1(17) => 
                           PC_BUS_pre_BTB_17_port, OUT1(16) => 
                           PC_BUS_pre_BTB_16_port, OUT1(15) => 
                           PC_BUS_pre_BTB_15_port, OUT1(14) => 
                           PC_BUS_pre_BTB_14_port, OUT1(13) => 
                           PC_BUS_pre_BTB_13_port, OUT1(12) => 
                           PC_BUS_pre_BTB_12_port, OUT1(11) => 
                           PC_BUS_pre_BTB_11_port, OUT1(10) => 
                           PC_BUS_pre_BTB_10_port, OUT1(9) => 
                           PC_BUS_pre_BTB_9_port, OUT1(8) => 
                           PC_BUS_pre_BTB_8_port, OUT1(7) => 
                           PC_BUS_pre_BTB_7_port, OUT1(6) => 
                           PC_BUS_pre_BTB_6_port, OUT1(5) => 
                           PC_BUS_pre_BTB_5_port, OUT1(4) => 
                           PC_BUS_pre_BTB_4_port, OUT1(3) => 
                           PC_BUS_pre_BTB_3_port, OUT1(2) => 
                           PC_BUS_pre_BTB_2_port, OUT1(1) => 
                           PC_BUS_pre_BTB_1_port, OUT1(0) => 
                           PC_BUS_pre_BTB_0_port);
   MUXPREDICTION : mux41_1 port map( IN0(31) => PC4_o_31_port, IN0(30) => 
                           PC4_o_30_port, IN0(29) => PC4_o_29_port, IN0(28) => 
                           PC4_o_28_port, IN0(27) => PC4_o_27_port, IN0(26) => 
                           PC4_o_26_port, IN0(25) => PC4_o_25_port, IN0(24) => 
                           PC4_o_24_port, IN0(23) => PC4_o_23_port, IN0(22) => 
                           PC4_o_22_port, IN0(21) => PC4_o_21_port, IN0(20) => 
                           PC4_o_20_port, IN0(19) => PC4_o_19_port, IN0(18) => 
                           PC4_o_18_port, IN0(17) => PC4_o_17_port, IN0(16) => 
                           PC4_o_16_port, IN0(15) => PC4_o_15_port, IN0(14) => 
                           PC4_o_14_port, IN0(13) => PC4_o_13_port, IN0(12) => 
                           PC4_o_12_port, IN0(11) => PC4_o_11_port, IN0(10) => 
                           PC4_o_10_port, IN0(9) => PC4_o_9_port, IN0(8) => 
                           PC4_o_8_port, IN0(7) => PC4_o_7_port, IN0(6) => 
                           PC4_o_6_port, IN0(5) => PC4_o_5_port, IN0(4) => 
                           PC4_o_4_port, IN0(3) => PC4_o_3_port, IN0(2) => 
                           PC4_o_2_port, IN0(1) => PC4_o_1_port, IN0(0) => 
                           PC4_o_0_port, IN1(31) => predicted_PC(31), IN1(30) 
                           => predicted_PC(30), IN1(29) => predicted_PC(29), 
                           IN1(28) => predicted_PC(28), IN1(27) => 
                           predicted_PC(27), IN1(26) => predicted_PC(26), 
                           IN1(25) => predicted_PC(25), IN1(24) => 
                           predicted_PC(24), IN1(23) => predicted_PC(23), 
                           IN1(22) => predicted_PC(22), IN1(21) => 
                           predicted_PC(21), IN1(20) => predicted_PC(20), 
                           IN1(19) => predicted_PC(19), IN1(18) => 
                           predicted_PC(18), IN1(17) => predicted_PC(17), 
                           IN1(16) => predicted_PC(16), IN1(15) => 
                           predicted_PC(15), IN1(14) => predicted_PC(14), 
                           IN1(13) => predicted_PC(13), IN1(12) => 
                           predicted_PC(12), IN1(11) => predicted_PC(11), 
                           IN1(10) => predicted_PC(10), IN1(9) => 
                           predicted_PC(9), IN1(8) => predicted_PC(8), IN1(7) 
                           => predicted_PC(7), IN1(6) => predicted_PC(6), 
                           IN1(5) => predicted_PC(5), IN1(4) => predicted_PC(4)
                           , IN1(3) => predicted_PC(3), IN1(2) => 
                           predicted_PC(2), IN1(1) => predicted_PC(1), IN1(0) 
                           => predicted_PC(0), IN2(31) => 
                           PC_BUS_pre_BTB_31_port, IN2(30) => 
                           PC_BUS_pre_BTB_30_port, IN2(29) => 
                           PC_BUS_pre_BTB_29_port, IN2(28) => 
                           PC_BUS_pre_BTB_28_port, IN2(27) => 
                           PC_BUS_pre_BTB_27_port, IN2(26) => 
                           PC_BUS_pre_BTB_26_port, IN2(25) => 
                           PC_BUS_pre_BTB_25_port, IN2(24) => 
                           PC_BUS_pre_BTB_24_port, IN2(23) => 
                           PC_BUS_pre_BTB_23_port, IN2(22) => 
                           PC_BUS_pre_BTB_22_port, IN2(21) => 
                           PC_BUS_pre_BTB_21_port, IN2(20) => n1, IN2(19) => 
                           PC_BUS_pre_BTB_19_port, IN2(18) => 
                           PC_BUS_pre_BTB_18_port, IN2(17) => 
                           PC_BUS_pre_BTB_17_port, IN2(16) => 
                           PC_BUS_pre_BTB_16_port, IN2(15) => 
                           PC_BUS_pre_BTB_15_port, IN2(14) => 
                           PC_BUS_pre_BTB_14_port, IN2(13) => 
                           PC_BUS_pre_BTB_13_port, IN2(12) => 
                           PC_BUS_pre_BTB_12_port, IN2(11) => 
                           PC_BUS_pre_BTB_11_port, IN2(10) => 
                           PC_BUS_pre_BTB_10_port, IN2(9) => 
                           PC_BUS_pre_BTB_9_port, IN2(8) => 
                           PC_BUS_pre_BTB_8_port, IN2(7) => 
                           PC_BUS_pre_BTB_7_port, IN2(6) => 
                           PC_BUS_pre_BTB_6_port, IN2(5) => 
                           PC_BUS_pre_BTB_5_port, IN2(4) => 
                           PC_BUS_pre_BTB_4_port, IN2(3) => 
                           PC_BUS_pre_BTB_3_port, IN2(2) => 
                           PC_BUS_pre_BTB_2_port, IN2(1) => 
                           PC_BUS_pre_BTB_1_port, IN2(0) => 
                           PC_BUS_pre_BTB_0_port, IN3(31) => 
                           PC_BUS_pre_BTB_31_port, IN3(30) => 
                           PC_BUS_pre_BTB_30_port, IN3(29) => 
                           PC_BUS_pre_BTB_29_port, IN3(28) => 
                           PC_BUS_pre_BTB_28_port, IN3(27) => 
                           PC_BUS_pre_BTB_27_port, IN3(26) => 
                           PC_BUS_pre_BTB_26_port, IN3(25) => 
                           PC_BUS_pre_BTB_25_port, IN3(24) => 
                           PC_BUS_pre_BTB_24_port, IN3(23) => 
                           PC_BUS_pre_BTB_23_port, IN3(22) => 
                           PC_BUS_pre_BTB_22_port, IN3(21) => 
                           PC_BUS_pre_BTB_21_port, IN3(20) => n1, IN3(19) => 
                           PC_BUS_pre_BTB_19_port, IN3(18) => 
                           PC_BUS_pre_BTB_18_port, IN3(17) => 
                           PC_BUS_pre_BTB_17_port, IN3(16) => 
                           PC_BUS_pre_BTB_16_port, IN3(15) => 
                           PC_BUS_pre_BTB_15_port, IN3(14) => 
                           PC_BUS_pre_BTB_14_port, IN3(13) => 
                           PC_BUS_pre_BTB_13_port, IN3(12) => 
                           PC_BUS_pre_BTB_12_port, IN3(11) => 
                           PC_BUS_pre_BTB_11_port, IN3(10) => 
                           PC_BUS_pre_BTB_10_port, IN3(9) => 
                           PC_BUS_pre_BTB_9_port, IN3(8) => 
                           PC_BUS_pre_BTB_8_port, IN3(7) => 
                           PC_BUS_pre_BTB_7_port, IN3(6) => 
                           PC_BUS_pre_BTB_6_port, IN3(5) => 
                           PC_BUS_pre_BTB_5_port, IN3(4) => 
                           PC_BUS_pre_BTB_4_port, IN3(3) => 
                           PC_BUS_pre_BTB_3_port, IN3(2) => 
                           PC_BUS_pre_BTB_2_port, IN3(1) => 
                           PC_BUS_pre_BTB_1_port, IN3(0) => 
                           PC_BUS_pre_BTB_0_port, CTRL(1) => mispredict_i, 
                           CTRL(0) => take_prediction_i, OUT1(31) => 
                           PC_BUS_31_port, OUT1(30) => PC_BUS_30_port, OUT1(29)
                           => PC_BUS_29_port, OUT1(28) => PC_BUS_28_port, 
                           OUT1(27) => PC_BUS_27_port, OUT1(26) => 
                           PC_BUS_26_port, OUT1(25) => PC_BUS_25_port, OUT1(24)
                           => PC_BUS_24_port, OUT1(23) => PC_BUS_23_port, 
                           OUT1(22) => PC_BUS_22_port, OUT1(21) => 
                           PC_BUS_21_port, OUT1(20) => PC_BUS_20_port, OUT1(19)
                           => PC_BUS_19_port, OUT1(18) => PC_BUS_18_port, 
                           OUT1(17) => PC_BUS_17_port, OUT1(16) => 
                           PC_BUS_16_port, OUT1(15) => PC_BUS_15_port, OUT1(14)
                           => PC_BUS_14_port, OUT1(13) => PC_BUS_13_port, 
                           OUT1(12) => PC_BUS_12_port, OUT1(11) => 
                           PC_BUS_11_port, OUT1(10) => PC_BUS_10_port, OUT1(9) 
                           => PC_BUS_9_port, OUT1(8) => PC_BUS_8_port, OUT1(7) 
                           => PC_BUS_7_port, OUT1(6) => PC_BUS_6_port, OUT1(5) 
                           => PC_BUS_5_port, OUT1(4) => PC_BUS_4_port, OUT1(3) 
                           => PC_BUS_3_port, OUT1(2) => PC_BUS_2_port, OUT1(1) 
                           => PC_BUS_1_port, OUT1(0) => PC_BUS_0_port);
   U1 : INV_X1 port map( A => stall_i, ZN => en_IR);
   U2 : CLKBUF_X1 port map( A => PC_BUS_pre_BTB_20_port, Z => n1);

end SYN_Struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity top_level is

   port( clock, rst : in std_logic;  IRAM_Addr_o : out std_logic_vector (31 
         downto 0);  IRAM_Dout_i : in std_logic_vector (31 downto 0);  
         DRAM_Enable_o, DRAM_WR_o : out std_logic;  DRAM_Din_o, DRAM_Addr_o : 
         out std_logic_vector (31 downto 0);  DRAM_Dout_i : in std_logic_vector
         (31 downto 0));

end top_level;

architecture SYN_arch of top_level is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component fw_logic
      port( D1_i, rAdec_i, D2_i, D3_i, rA_i, rB_i : in std_logic_vector (4 
            downto 0);  S_mem_W, S_wb_W, S_exe_W : in std_logic;  S_FWAdec, 
            S_FWA, S_FWB : out std_logic_vector (1 downto 0);  S_mem_LOAD_BAR :
            in std_logic);
   end component;
   
   component mem_block
      port( X_i, LOAD_i : in std_logic_vector (31 downto 0);  W_o : out 
            std_logic_vector (31 downto 0);  S_MUX_MEM_i_BAR : in std_logic);
   end component;
   
   component mem_regs
      port( W_i : in std_logic_vector (31 downto 0);  D3_i : in 
            std_logic_vector (4 downto 0);  W_o : out std_logic_vector (31 
            downto 0);  D3_o : out std_logic_vector (4 downto 0);  clk, rst : 
            in std_logic);
   end component;
   
   component execute_block
      port( IMM_i, A_i : in std_logic_vector (31 downto 0);  rB_i, rC_i : in 
            std_logic_vector (4 downto 0);  MUXED_B_i : in std_logic_vector (31
            downto 0);  S_MUX_ALUIN_i : in std_logic;  FW_X_i, FW_W_i : in 
            std_logic_vector (31 downto 0);  S_FW_A_i, S_FW_B_i : in 
            std_logic_vector (1 downto 0);  muxed_dest : out std_logic_vector 
            (4 downto 0);  muxed_B : out std_logic_vector (31 downto 0);  
            S_MUX_DEST_i : in std_logic_vector (1 downto 0);  OP : in 
            std_logic_vector (0 to 4);  ALUW_i : in std_logic_vector (12 downto
            0);  DOUT : out std_logic_vector (31 downto 0);  stall_o : out 
            std_logic;  Clock, Reset : in std_logic);
   end component;
   
   component execute_regs
      port( X_i, S_i : in std_logic_vector (31 downto 0);  D2_i : in 
            std_logic_vector (4 downto 0);  X_o, S_o : out std_logic_vector (31
            downto 0);  D2_o : out std_logic_vector (4 downto 0);  stall_i, clk
            , rst : in std_logic);
   end component;
   
   component decode_regs
      port( A_i, B_i : in std_logic_vector (31 downto 0);  rA_i, rB_i, rC_i : 
            in std_logic_vector (4 downto 0);  IMM_i : in std_logic_vector (31 
            downto 0);  ALUW_i : in std_logic_vector (12 downto 0);  A_o, B_o :
            out std_logic_vector (31 downto 0);  rA_o, rB_o, rC_o : out 
            std_logic_vector (4 downto 0);  IMM_o : out std_logic_vector (31 
            downto 0);  ALUW_o : out std_logic_vector (12 downto 0);  stall_i, 
            clk, rst : in std_logic);
   end component;
   
   component dlx_regfile
      port( Clk, Rst, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, 
            ADD_RD2 : in std_logic_vector (4 downto 0);  DATAIN : in 
            std_logic_vector (31 downto 0);  OUT1, OUT2 : out std_logic_vector 
            (31 downto 0));
   end component;
   
   component 
      dlx_cu_MICROCODE_MEM_SIZE64_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE13
      port( Clk, Rst : in std_logic;  IR_IN : in std_logic_vector (31 downto 0)
            ;  stall_exe_i, mispredict_i : in std_logic;  D1_i, D2_i : in 
            std_logic_vector (4 downto 0);  S1_LATCH_EN, S2_LATCH_EN, 
            S3_LATCH_EN : out std_logic;  S_MUX_PC_BUS : out std_logic_vector 
            (1 downto 0);  S_EXT, S_EXT_SIGN, S_EQ_NEQ : out std_logic;  
            S_MUX_DEST : out std_logic_vector (1 downto 0);  S_MUX_LINK, 
            S_MEM_W_R, S_MEM_EN, S_RF_W_wb, S_RF_W_mem, S_RF_W_exe, S_MUX_ALUIN
            , stall_exe_o, stall_dec_o, stall_fetch_o, stall_btb_o, 
            was_branch_o, was_jmp_o : out std_logic;  ALU_WORD_o : out 
            std_logic_vector (12 downto 0);  ALU_OPCODE : out std_logic_vector 
            (0 to 4);  S_MUX_MEM_BAR : out std_logic);
   end component;
   
   component jump_logic
      port( NPCF_i, IR_i, A_i : in std_logic_vector (31 downto 0);  A_o : out 
            std_logic_vector (31 downto 0);  rA_o, rB_o, rC_o : out 
            std_logic_vector (4 downto 0);  branch_target_o, sum_addr_o, 
            extended_imm : out std_logic_vector (31 downto 0);  taken_o : out 
            std_logic;  FW_X_i, FW_W_i : in std_logic_vector (31 downto 0);  
            S_FW_Adec_i : in std_logic_vector (1 downto 0);  S_EXT_i, 
            S_EXT_SIGN_i, S_MUX_LINK_i, S_EQ_NEQ_i : in std_logic);
   end component;
   
   component fetch_regs
      port( NPCF_i, IR_i : in std_logic_vector (31 downto 0);  NPCF_o, IR_o : 
            out std_logic_vector (31 downto 0);  stall_i, clk, rst : in 
            std_logic);
   end component;
   
   component btb_N_LINES4_SIZE32
      port( clock, reset, stall_i : in std_logic;  TAG_i : in std_logic_vector 
            (3 downto 0);  target_PC_i : in std_logic_vector (31 downto 0);  
            was_taken_i : in std_logic;  predicted_next_PC_o : out 
            std_logic_vector (31 downto 0);  taken_o, mispredict_o : out 
            std_logic);
   end component;
   
   component fetch_block
      port( branch_target_i, sum_addr_i, A_i, NPC4_i : in std_logic_vector (31 
            downto 0);  S_MUX_PC_BUS_i : in std_logic_vector (1 downto 0);  
            PC_o, PC4_o, PC_BUS_pre_BTB : out std_logic_vector (31 downto 0);  
            stall_i, take_prediction_i, mispredict_i : in std_logic;  
            predicted_PC : in std_logic_vector (31 downto 0);  clk, rst : in 
            std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, IRAM_Addr_o_31_port, 
      IRAM_Addr_o_30_port, IRAM_Addr_o_29_port, IRAM_Addr_o_28_port, 
      IRAM_Addr_o_27_port, IRAM_Addr_o_26_port, IRAM_Addr_o_25_port, 
      IRAM_Addr_o_24_port, IRAM_Addr_o_23_port, IRAM_Addr_o_22_port, 
      IRAM_Addr_o_21_port, IRAM_Addr_o_20_port, IRAM_Addr_o_19_port, 
      IRAM_Addr_o_18_port, IRAM_Addr_o_17_port, IRAM_Addr_o_16_port, 
      IRAM_Addr_o_15_port, IRAM_Addr_o_14_port, IRAM_Addr_o_13_port, 
      IRAM_Addr_o_12_port, IRAM_Addr_o_11_port, IRAM_Addr_o_10_port, 
      IRAM_Addr_o_9_port, IRAM_Addr_o_8_port, IRAM_Addr_o_7_port, 
      IRAM_Addr_o_6_port, IRAM_Addr_o_5_port, IRAM_Addr_o_4_port, 
      IRAM_Addr_o_3_port, IRAM_Addr_o_2_port, IRAM_Addr_o_1_port, 
      IRAM_Addr_o_0_port, DRAM_Addr_o_31_port, DRAM_Addr_o_30_port, 
      DRAM_Addr_o_29_port, DRAM_Addr_o_28_port, DRAM_Addr_o_27_port, 
      DRAM_Addr_o_26_port, DRAM_Addr_o_25_port, DRAM_Addr_o_24_port, 
      DRAM_Addr_o_23_port, DRAM_Addr_o_22_port, DRAM_Addr_o_21_port, 
      DRAM_Addr_o_20_port, DRAM_Addr_o_19_port, DRAM_Addr_o_18_port, 
      DRAM_Addr_o_17_port, DRAM_Addr_o_16_port, DRAM_Addr_o_15_port, 
      DRAM_Addr_o_14_port, DRAM_Addr_o_13_port, DRAM_Addr_o_12_port, 
      DRAM_Addr_o_11_port, DRAM_Addr_o_10_port, DRAM_Addr_o_9_port, 
      DRAM_Addr_o_8_port, DRAM_Addr_o_7_port, DRAM_Addr_o_6_port, 
      DRAM_Addr_o_5_port, DRAM_Addr_o_4_port, DRAM_Addr_o_3_port, 
      DRAM_Addr_o_2_port, DRAM_Addr_o_1_port, DRAM_Addr_o_0_port, 
      was_taken_from_jl, was_branch, was_jmp, was_taken, 
      dummy_branch_target_31_port, dummy_branch_target_30_port, 
      dummy_branch_target_29_port, dummy_branch_target_28_port, 
      dummy_branch_target_27_port, dummy_branch_target_26_port, 
      dummy_branch_target_25_port, dummy_branch_target_24_port, 
      dummy_branch_target_23_port, dummy_branch_target_22_port, 
      dummy_branch_target_21_port, dummy_branch_target_20_port, 
      dummy_branch_target_19_port, dummy_branch_target_18_port, 
      dummy_branch_target_17_port, dummy_branch_target_16_port, 
      dummy_branch_target_15_port, dummy_branch_target_14_port, 
      dummy_branch_target_13_port, dummy_branch_target_12_port, 
      dummy_branch_target_11_port, dummy_branch_target_10_port, 
      dummy_branch_target_9_port, dummy_branch_target_8_port, 
      dummy_branch_target_7_port, dummy_branch_target_6_port, 
      dummy_branch_target_5_port, dummy_branch_target_4_port, 
      dummy_branch_target_3_port, dummy_branch_target_2_port, 
      dummy_branch_target_1_port, dummy_branch_target_0_port, 
      dummy_sum_addr_31_port, dummy_sum_addr_30_port, dummy_sum_addr_29_port, 
      dummy_sum_addr_28_port, dummy_sum_addr_27_port, dummy_sum_addr_26_port, 
      dummy_sum_addr_25_port, dummy_sum_addr_24_port, dummy_sum_addr_23_port, 
      dummy_sum_addr_22_port, dummy_sum_addr_21_port, dummy_sum_addr_20_port, 
      dummy_sum_addr_19_port, dummy_sum_addr_18_port, dummy_sum_addr_17_port, 
      dummy_sum_addr_16_port, dummy_sum_addr_15_port, dummy_sum_addr_14_port, 
      dummy_sum_addr_13_port, dummy_sum_addr_12_port, dummy_sum_addr_11_port, 
      dummy_sum_addr_10_port, dummy_sum_addr_9_port, dummy_sum_addr_8_port, 
      dummy_sum_addr_7_port, dummy_sum_addr_6_port, dummy_sum_addr_5_port, 
      dummy_sum_addr_4_port, dummy_sum_addr_3_port, dummy_sum_addr_2_port, 
      dummy_sum_addr_1_port, dummy_sum_addr_0_port, dummy_A_31_port, 
      dummy_A_30_port, dummy_A_29_port, dummy_A_28_port, dummy_A_27_port, 
      dummy_A_26_port, dummy_A_25_port, dummy_A_24_port, dummy_A_23_port, 
      dummy_A_22_port, dummy_A_21_port, dummy_A_20_port, dummy_A_19_port, 
      dummy_A_18_port, dummy_A_17_port, dummy_A_16_port, dummy_A_15_port, 
      dummy_A_14_port, dummy_A_13_port, dummy_A_12_port, dummy_A_11_port, 
      dummy_A_10_port, dummy_A_9_port, dummy_A_8_port, dummy_A_7_port, 
      dummy_A_6_port, dummy_A_5_port, dummy_A_4_port, dummy_A_3_port, 
      dummy_A_2_port, dummy_A_1_port, dummy_A_0_port, NPCF_31_port, 
      NPCF_30_port, NPCF_29_port, NPCF_28_port, NPCF_27_port, NPCF_26_port, 
      NPCF_25_port, NPCF_24_port, NPCF_23_port, NPCF_22_port, NPCF_21_port, 
      NPCF_20_port, NPCF_19_port, NPCF_18_port, NPCF_17_port, NPCF_16_port, 
      NPCF_15_port, NPCF_14_port, NPCF_13_port, NPCF_12_port, NPCF_11_port, 
      NPCF_10_port, NPCF_9_port, NPCF_8_port, NPCF_7_port, NPCF_6_port, 
      NPCF_5_port, NPCF_4_port, NPCF_3_port, NPCF_2_port, NPCF_1_port, 
      NPCF_0_port, dummy_S_MUX_PC_BUS_1_port, dummy_S_MUX_PC_BUS_0_port, 
      PC4_31_port, PC4_30_port, PC4_29_port, PC4_28_port, PC4_27_port, 
      PC4_26_port, PC4_25_port, PC4_24_port, PC4_23_port, PC4_22_port, 
      PC4_21_port, PC4_20_port, PC4_19_port, PC4_18_port, PC4_17_port, 
      PC4_16_port, PC4_15_port, PC4_14_port, PC4_13_port, PC4_12_port, 
      PC4_11_port, PC4_10_port, PC4_9_port, PC4_8_port, PC4_7_port, PC4_6_port,
      PC4_5_port, PC4_4_port, PC4_3_port, PC4_2_port, PC4_1_port, PC4_0_port, 
      TARGET_PC_31_port, TARGET_PC_30_port, TARGET_PC_28_port, 
      TARGET_PC_27_port, TARGET_PC_26_port, TARGET_PC_25_port, 
      TARGET_PC_24_port, TARGET_PC_23_port, TARGET_PC_22_port, 
      TARGET_PC_21_port, TARGET_PC_20_port, TARGET_PC_19_port, 
      TARGET_PC_18_port, TARGET_PC_17_port, TARGET_PC_16_port, 
      TARGET_PC_15_port, TARGET_PC_14_port, TARGET_PC_13_port, 
      TARGET_PC_12_port, TARGET_PC_11_port, TARGET_PC_10_port, TARGET_PC_9_port
      , TARGET_PC_8_port, TARGET_PC_7_port, TARGET_PC_6_port, TARGET_PC_5_port,
      TARGET_PC_4_port, TARGET_PC_3_port, TARGET_PC_2_port, TARGET_PC_1_port, 
      TARGET_PC_0_port, stall_fetch, mispredict, take_prediction, 
      predicted_PC_31_port, predicted_PC_30_port, predicted_PC_29_port, 
      predicted_PC_28_port, predicted_PC_27_port, predicted_PC_26_port, 
      predicted_PC_25_port, predicted_PC_24_port, predicted_PC_23_port, 
      predicted_PC_22_port, predicted_PC_21_port, predicted_PC_20_port, 
      predicted_PC_19_port, predicted_PC_18_port, predicted_PC_17_port, 
      predicted_PC_16_port, predicted_PC_15_port, predicted_PC_14_port, 
      predicted_PC_13_port, predicted_PC_12_port, predicted_PC_11_port, 
      predicted_PC_10_port, predicted_PC_9_port, predicted_PC_8_port, 
      predicted_PC_7_port, predicted_PC_6_port, predicted_PC_5_port, 
      predicted_PC_4_port, predicted_PC_3_port, predicted_PC_2_port, 
      predicted_PC_1_port, predicted_PC_0_port, stall_btb, IR_31_port, 
      IR_30_port, IR_29_port, IR_28_port, IR_27_port, IR_26_port, IR_25_port, 
      IR_24_port, IR_23_port, IR_22_port, IR_21_port, IR_20_port, IR_19_port, 
      IR_18_port, IR_17_port, IR_16_port, IR_15_port, IR_14_port, IR_13_port, 
      IR_12_port, IR_11_port, IR_10_port, IR_9_port, IR_8_port, IR_7_port, 
      IR_6_port, IR_5_port, IR_4_port, IR_3_port, IR_2_port, IR_1_port, 
      IR_0_port, stall_decode, AtoComp_31_port, AtoComp_30_port, 
      AtoComp_29_port, AtoComp_28_port, AtoComp_27_port, AtoComp_26_port, 
      AtoComp_25_port, AtoComp_24_port, AtoComp_23_port, AtoComp_22_port, 
      AtoComp_21_port, AtoComp_20_port, AtoComp_19_port, AtoComp_18_port, 
      AtoComp_17_port, AtoComp_16_port, AtoComp_15_port, AtoComp_14_port, 
      AtoComp_13_port, AtoComp_12_port, AtoComp_11_port, AtoComp_10_port, 
      AtoComp_9_port, AtoComp_8_port, AtoComp_7_port, AtoComp_6_port, 
      AtoComp_5_port, AtoComp_4_port, AtoComp_3_port, AtoComp_2_port, 
      AtoComp_1_port, AtoComp_0_port, rA2reg_4_port, rA2reg_3_port, 
      rA2reg_2_port, rA2reg_1_port, rA2reg_0_port, rB2reg_4_port, rB2reg_3_port
      , rB2reg_2_port, rB2reg_1_port, rB2reg_0_port, rC2reg_4_port, 
      rC2reg_3_port, rC2reg_2_port, rC2reg_1_port, rC2reg_0_port, 
      help_IMM_31_port, help_IMM_30_port, help_IMM_29_port, help_IMM_28_port, 
      help_IMM_27_port, help_IMM_26_port, help_IMM_25_port, help_IMM_24_port, 
      help_IMM_23_port, help_IMM_22_port, help_IMM_21_port, help_IMM_20_port, 
      help_IMM_19_port, help_IMM_18_port, help_IMM_17_port, help_IMM_16_port, 
      help_IMM_15_port, help_IMM_14_port, help_IMM_13_port, help_IMM_12_port, 
      help_IMM_11_port, help_IMM_10_port, help_IMM_9_port, help_IMM_8_port, 
      help_IMM_7_port, help_IMM_6_port, help_IMM_5_port, help_IMM_4_port, 
      help_IMM_3_port, help_IMM_2_port, help_IMM_1_port, help_IMM_0_port, 
      wb2reg_31_port, wb2reg_30_port, wb2reg_29_port, wb2reg_28_port, 
      wb2reg_27_port, wb2reg_26_port, wb2reg_25_port, wb2reg_24_port, 
      wb2reg_23_port, wb2reg_22_port, wb2reg_21_port, wb2reg_20_port, 
      wb2reg_19_port, wb2reg_18_port, wb2reg_17_port, wb2reg_16_port, 
      wb2reg_15_port, wb2reg_14_port, wb2reg_13_port, wb2reg_12_port, 
      wb2reg_11_port, wb2reg_10_port, wb2reg_9_port, wb2reg_8_port, 
      wb2reg_7_port, wb2reg_6_port, wb2reg_5_port, wb2reg_4_port, wb2reg_3_port
      , wb2reg_2_port, wb2reg_1_port, wb2reg_0_port, dummy_S_FWAdec_1_port, 
      dummy_S_FWAdec_0_port, dummy_S_EXT, dummy_S_EXT_SIGN, dummy_S_EQ_NEQ, 
      exe_stall_cu, muxed_dest2exe_4_port, muxed_dest2exe_3_port, 
      muxed_dest2exe_2_port, muxed_dest2exe_1_port, muxed_dest2exe_0_port, 
      D22D3_4_port, D22D3_3_port, D22D3_1_port, D22D3_0_port, 
      dummy_S_MUX_DEST_1_port, dummy_S_MUX_DEST_0_port, dummy_S_MUX_MEM, 
      dummy_S_RF_W_wb, dummy_S_RF_W_mem, dummy_S_MUX_ALUIN, stall_exe, 
      ALUW_dec_12_port, ALUW_dec_11_port, ALUW_dec_10_port, ALUW_dec_9_port, 
      ALUW_dec_8_port, ALUW_dec_7_port, ALUW_dec_6_port, ALUW_dec_5_port, 
      ALUW_dec_4_port, ALUW_dec_3_port, ALUW_dec_2_port, ALUW_dec_1_port, 
      ALUW_dec_0_port, enable_regfile, W2wb_31_port, W2wb_30_port, W2wb_29_port
      , W2wb_28_port, W2wb_27_port, W2wb_26_port, W2wb_25_port, W2wb_24_port, 
      W2wb_23_port, W2wb_22_port, W2wb_21_port, W2wb_20_port, W2wb_19_port, 
      W2wb_18_port, W2wb_17_port, W2wb_16_port, W2wb_15_port, W2wb_14_port, 
      W2wb_13_port, W2wb_12_port, W2wb_11_port, W2wb_10_port, W2wb_9_port, 
      W2wb_8_port, W2wb_7_port, W2wb_6_port, W2wb_5_port, W2wb_4_port, 
      W2wb_3_port, W2wb_2_port, W2wb_1_port, W2wb_0_port, dummy_B_31_port, 
      dummy_B_30_port, dummy_B_29_port, dummy_B_28_port, dummy_B_27_port, 
      dummy_B_26_port, dummy_B_25_port, dummy_B_24_port, dummy_B_23_port, 
      dummy_B_22_port, dummy_B_21_port, dummy_B_20_port, dummy_B_19_port, 
      dummy_B_18_port, dummy_B_17_port, dummy_B_16_port, dummy_B_15_port, 
      dummy_B_14_port, dummy_B_13_port, dummy_B_12_port, dummy_B_11_port, 
      dummy_B_10_port, dummy_B_9_port, dummy_B_8_port, dummy_B_7_port, 
      dummy_B_6_port, dummy_B_5_port, dummy_B_4_port, dummy_B_3_port, 
      dummy_B_2_port, dummy_B_1_port, dummy_B_0_port, A2exe_31_port, 
      A2exe_30_port, A2exe_29_port, A2exe_28_port, A2exe_27_port, A2exe_26_port
      , A2exe_25_port, A2exe_24_port, A2exe_23_port, A2exe_22_port, 
      A2exe_21_port, A2exe_20_port, A2exe_19_port, A2exe_18_port, A2exe_17_port
      , A2exe_16_port, A2exe_15_port, A2exe_14_port, A2exe_13_port, 
      A2exe_12_port, A2exe_11_port, A2exe_10_port, A2exe_9_port, A2exe_8_port, 
      A2exe_7_port, A2exe_6_port, A2exe_5_port, A2exe_4_port, A2exe_3_port, 
      A2exe_2_port, A2exe_1_port, A2exe_0_port, B2exe_31_port, B2exe_30_port, 
      B2exe_29_port, B2exe_28_port, B2exe_27_port, B2exe_26_port, B2exe_25_port
      , B2exe_24_port, B2exe_23_port, B2exe_22_port, B2exe_21_port, 
      B2exe_20_port, B2exe_19_port, B2exe_18_port, B2exe_17_port, B2exe_16_port
      , B2exe_15_port, B2exe_14_port, B2exe_13_port, B2exe_12_port, 
      B2exe_11_port, B2exe_10_port, B2exe_9_port, B2exe_8_port, B2exe_7_port, 
      B2exe_6_port, B2exe_5_port, B2exe_4_port, B2exe_3_port, B2exe_2_port, 
      B2exe_1_port, B2exe_0_port, rA2fw_4_port, rA2fw_3_port, rA2fw_2_port, 
      rA2fw_1_port, rA2fw_0_port, rB2mux_4_port, rB2mux_3_port, rB2mux_2_port, 
      rB2mux_1_port, rB2mux_0_port, rC2mux_4_port, rC2mux_3_port, rC2mux_2_port
      , rC2mux_1_port, rC2mux_0_port, IMM2exe_31_port, IMM2exe_30_port, 
      IMM2exe_29_port, IMM2exe_28_port, IMM2exe_27_port, IMM2exe_26_port, 
      IMM2exe_25_port, IMM2exe_24_port, IMM2exe_23_port, IMM2exe_22_port, 
      IMM2exe_21_port, IMM2exe_20_port, IMM2exe_19_port, IMM2exe_18_port, 
      IMM2exe_17_port, IMM2exe_16_port, IMM2exe_15_port, IMM2exe_14_port, 
      IMM2exe_13_port, IMM2exe_12_port, IMM2exe_11_port, IMM2exe_10_port, 
      IMM2exe_9_port, IMM2exe_8_port, IMM2exe_7_port, IMM2exe_6_port, 
      IMM2exe_5_port, IMM2exe_4_port, IMM2exe_3_port, IMM2exe_2_port, 
      IMM2exe_1_port, IMM2exe_0_port, ALUW_12_port, ALUW_11_port, ALUW_10_port,
      ALUW_9_port, ALUW_8_port, ALUW_7_port, ALUW_6_port, ALUW_5_port, 
      ALUW_4_port, ALUW_3_port, ALUW_2_port, ALUW_1_port, ALUW_0_port, 
      X2mem_31_port, X2mem_30_port, X2mem_29_port, X2mem_28_port, X2mem_27_port
      , X2mem_26_port, X2mem_25_port, X2mem_24_port, X2mem_23_port, 
      X2mem_22_port, X2mem_21_port, X2mem_20_port, X2mem_19_port, X2mem_18_port
      , X2mem_17_port, X2mem_16_port, X2mem_15_port, X2mem_14_port, 
      X2mem_13_port, X2mem_12_port, X2mem_11_port, X2mem_10_port, X2mem_9_port,
      X2mem_8_port, X2mem_7_port, X2mem_6_port, X2mem_5_port, X2mem_4_port, 
      X2mem_3_port, X2mem_2_port, X2mem_1_port, X2mem_0_port, S2mem_31_port, 
      S2mem_30_port, S2mem_29_port, S2mem_28_port, S2mem_27_port, S2mem_26_port
      , S2mem_25_port, S2mem_24_port, S2mem_23_port, S2mem_22_port, 
      S2mem_21_port, S2mem_20_port, S2mem_19_port, S2mem_18_port, S2mem_17_port
      , S2mem_16_port, S2mem_15_port, S2mem_14_port, S2mem_13_port, 
      S2mem_12_port, S2mem_11_port, S2mem_10_port, S2mem_9_port, S2mem_8_port, 
      S2mem_7_port, S2mem_6_port, S2mem_5_port, S2mem_4_port, S2mem_3_port, 
      S2mem_2_port, S2mem_0_port, dummy_S_FWA2exe_1_port, 
      dummy_S_FWA2exe_0_port, dummy_S_FWB2exe_1_port, dummy_S_FWB2exe_0_port, 
      D32reg_4_port, D32reg_3_port, D32reg_2_port, D32reg_1_port, D32reg_0_port
      , n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18
      , n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, 
      n33, n34, n35, net47162, net47163, net47164, net47165, net47166, net47167
      , net47168, net47169, net47170 : std_logic;

begin
   IRAM_Addr_o <= ( IRAM_Addr_o_31_port, IRAM_Addr_o_30_port, 
      IRAM_Addr_o_29_port, IRAM_Addr_o_28_port, IRAM_Addr_o_27_port, 
      IRAM_Addr_o_26_port, IRAM_Addr_o_25_port, IRAM_Addr_o_24_port, 
      IRAM_Addr_o_23_port, IRAM_Addr_o_22_port, IRAM_Addr_o_21_port, 
      IRAM_Addr_o_20_port, IRAM_Addr_o_19_port, IRAM_Addr_o_18_port, 
      IRAM_Addr_o_17_port, IRAM_Addr_o_16_port, IRAM_Addr_o_15_port, 
      IRAM_Addr_o_14_port, IRAM_Addr_o_13_port, IRAM_Addr_o_12_port, 
      IRAM_Addr_o_11_port, IRAM_Addr_o_10_port, IRAM_Addr_o_9_port, 
      IRAM_Addr_o_8_port, IRAM_Addr_o_7_port, IRAM_Addr_o_6_port, 
      IRAM_Addr_o_5_port, IRAM_Addr_o_4_port, IRAM_Addr_o_3_port, 
      IRAM_Addr_o_2_port, IRAM_Addr_o_1_port, IRAM_Addr_o_0_port );
   DRAM_Addr_o <= ( DRAM_Addr_o_31_port, DRAM_Addr_o_30_port, 
      DRAM_Addr_o_29_port, DRAM_Addr_o_28_port, DRAM_Addr_o_27_port, 
      DRAM_Addr_o_26_port, DRAM_Addr_o_25_port, DRAM_Addr_o_24_port, 
      DRAM_Addr_o_23_port, DRAM_Addr_o_22_port, DRAM_Addr_o_21_port, 
      DRAM_Addr_o_20_port, DRAM_Addr_o_19_port, DRAM_Addr_o_18_port, 
      DRAM_Addr_o_17_port, DRAM_Addr_o_16_port, DRAM_Addr_o_15_port, 
      DRAM_Addr_o_14_port, DRAM_Addr_o_13_port, DRAM_Addr_o_12_port, 
      DRAM_Addr_o_11_port, DRAM_Addr_o_10_port, DRAM_Addr_o_9_port, 
      DRAM_Addr_o_8_port, DRAM_Addr_o_7_port, DRAM_Addr_o_6_port, 
      DRAM_Addr_o_5_port, DRAM_Addr_o_4_port, DRAM_Addr_o_3_port, 
      DRAM_Addr_o_2_port, DRAM_Addr_o_1_port, DRAM_Addr_o_0_port );
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   UFETCH_BLOCK : fetch_block port map( branch_target_i(31) => 
                           dummy_branch_target_31_port, branch_target_i(30) => 
                           dummy_branch_target_30_port, branch_target_i(29) => 
                           dummy_branch_target_29_port, branch_target_i(28) => 
                           dummy_branch_target_28_port, branch_target_i(27) => 
                           dummy_branch_target_27_port, branch_target_i(26) => 
                           dummy_branch_target_26_port, branch_target_i(25) => 
                           dummy_branch_target_25_port, branch_target_i(24) => 
                           dummy_branch_target_24_port, branch_target_i(23) => 
                           dummy_branch_target_23_port, branch_target_i(22) => 
                           dummy_branch_target_22_port, branch_target_i(21) => 
                           dummy_branch_target_21_port, branch_target_i(20) => 
                           dummy_branch_target_20_port, branch_target_i(19) => 
                           dummy_branch_target_19_port, branch_target_i(18) => 
                           dummy_branch_target_18_port, branch_target_i(17) => 
                           dummy_branch_target_17_port, branch_target_i(16) => 
                           dummy_branch_target_16_port, branch_target_i(15) => 
                           dummy_branch_target_15_port, branch_target_i(14) => 
                           dummy_branch_target_14_port, branch_target_i(13) => 
                           dummy_branch_target_13_port, branch_target_i(12) => 
                           dummy_branch_target_12_port, branch_target_i(11) => 
                           dummy_branch_target_11_port, branch_target_i(10) => 
                           dummy_branch_target_10_port, branch_target_i(9) => 
                           dummy_branch_target_9_port, branch_target_i(8) => 
                           dummy_branch_target_8_port, branch_target_i(7) => 
                           dummy_branch_target_7_port, branch_target_i(6) => 
                           dummy_branch_target_6_port, branch_target_i(5) => 
                           dummy_branch_target_5_port, branch_target_i(4) => 
                           dummy_branch_target_4_port, branch_target_i(3) => 
                           dummy_branch_target_3_port, branch_target_i(2) => 
                           dummy_branch_target_2_port, branch_target_i(1) => 
                           dummy_branch_target_1_port, branch_target_i(0) => 
                           dummy_branch_target_0_port, sum_addr_i(31) => 
                           dummy_sum_addr_31_port, sum_addr_i(30) => 
                           dummy_sum_addr_30_port, sum_addr_i(29) => 
                           dummy_sum_addr_29_port, sum_addr_i(28) => 
                           dummy_sum_addr_28_port, sum_addr_i(27) => 
                           dummy_sum_addr_27_port, sum_addr_i(26) => 
                           dummy_sum_addr_26_port, sum_addr_i(25) => 
                           dummy_sum_addr_25_port, sum_addr_i(24) => 
                           dummy_sum_addr_24_port, sum_addr_i(23) => 
                           dummy_sum_addr_23_port, sum_addr_i(22) => 
                           dummy_sum_addr_22_port, sum_addr_i(21) => 
                           dummy_sum_addr_21_port, sum_addr_i(20) => 
                           dummy_sum_addr_20_port, sum_addr_i(19) => 
                           dummy_sum_addr_19_port, sum_addr_i(18) => 
                           dummy_sum_addr_18_port, sum_addr_i(17) => 
                           dummy_sum_addr_17_port, sum_addr_i(16) => 
                           dummy_sum_addr_16_port, sum_addr_i(15) => 
                           dummy_sum_addr_15_port, sum_addr_i(14) => 
                           dummy_sum_addr_14_port, sum_addr_i(13) => 
                           dummy_sum_addr_13_port, sum_addr_i(12) => 
                           dummy_sum_addr_12_port, sum_addr_i(11) => 
                           dummy_sum_addr_11_port, sum_addr_i(10) => 
                           dummy_sum_addr_10_port, sum_addr_i(9) => 
                           dummy_sum_addr_9_port, sum_addr_i(8) => 
                           dummy_sum_addr_8_port, sum_addr_i(7) => 
                           dummy_sum_addr_7_port, sum_addr_i(6) => 
                           dummy_sum_addr_6_port, sum_addr_i(5) => 
                           dummy_sum_addr_5_port, sum_addr_i(4) => 
                           dummy_sum_addr_4_port, sum_addr_i(3) => 
                           dummy_sum_addr_3_port, sum_addr_i(2) => 
                           dummy_sum_addr_2_port, sum_addr_i(1) => 
                           dummy_sum_addr_1_port, sum_addr_i(0) => 
                           dummy_sum_addr_0_port, A_i(31) => dummy_A_31_port, 
                           A_i(30) => dummy_A_30_port, A_i(29) => 
                           dummy_A_29_port, A_i(28) => dummy_A_28_port, A_i(27)
                           => dummy_A_27_port, A_i(26) => dummy_A_26_port, 
                           A_i(25) => dummy_A_25_port, A_i(24) => 
                           dummy_A_24_port, A_i(23) => dummy_A_23_port, A_i(22)
                           => dummy_A_22_port, A_i(21) => dummy_A_21_port, 
                           A_i(20) => dummy_A_20_port, A_i(19) => 
                           dummy_A_19_port, A_i(18) => dummy_A_18_port, A_i(17)
                           => dummy_A_17_port, A_i(16) => dummy_A_16_port, 
                           A_i(15) => dummy_A_15_port, A_i(14) => 
                           dummy_A_14_port, A_i(13) => dummy_A_13_port, A_i(12)
                           => dummy_A_12_port, A_i(11) => dummy_A_11_port, 
                           A_i(10) => dummy_A_10_port, A_i(9) => dummy_A_9_port
                           , A_i(8) => dummy_A_8_port, A_i(7) => dummy_A_7_port
                           , A_i(6) => dummy_A_6_port, A_i(5) => dummy_A_5_port
                           , A_i(4) => dummy_A_4_port, A_i(3) => dummy_A_3_port
                           , A_i(2) => dummy_A_2_port, A_i(1) => dummy_A_1_port
                           , A_i(0) => dummy_A_0_port, NPC4_i(31) => 
                           NPCF_31_port, NPC4_i(30) => NPCF_30_port, NPC4_i(29)
                           => NPCF_29_port, NPC4_i(28) => NPCF_28_port, 
                           NPC4_i(27) => NPCF_27_port, NPC4_i(26) => 
                           NPCF_26_port, NPC4_i(25) => NPCF_25_port, NPC4_i(24)
                           => NPCF_24_port, NPC4_i(23) => NPCF_23_port, 
                           NPC4_i(22) => NPCF_22_port, NPC4_i(21) => 
                           NPCF_21_port, NPC4_i(20) => NPCF_20_port, NPC4_i(19)
                           => NPCF_19_port, NPC4_i(18) => NPCF_18_port, 
                           NPC4_i(17) => NPCF_17_port, NPC4_i(16) => 
                           NPCF_16_port, NPC4_i(15) => NPCF_15_port, NPC4_i(14)
                           => NPCF_14_port, NPC4_i(13) => NPCF_13_port, 
                           NPC4_i(12) => NPCF_12_port, NPC4_i(11) => 
                           NPCF_11_port, NPC4_i(10) => NPCF_10_port, NPC4_i(9) 
                           => NPCF_9_port, NPC4_i(8) => NPCF_8_port, NPC4_i(7) 
                           => NPCF_7_port, NPC4_i(6) => NPCF_6_port, NPC4_i(5) 
                           => NPCF_5_port, NPC4_i(4) => NPCF_4_port, NPC4_i(3) 
                           => NPCF_3_port, NPC4_i(2) => NPCF_2_port, NPC4_i(1) 
                           => NPCF_1_port, NPC4_i(0) => NPCF_0_port, 
                           S_MUX_PC_BUS_i(1) => dummy_S_MUX_PC_BUS_1_port, 
                           S_MUX_PC_BUS_i(0) => dummy_S_MUX_PC_BUS_0_port, 
                           PC_o(31) => IRAM_Addr_o_31_port, PC_o(30) => 
                           IRAM_Addr_o_30_port, PC_o(29) => IRAM_Addr_o_29_port
                           , PC_o(28) => IRAM_Addr_o_28_port, PC_o(27) => 
                           IRAM_Addr_o_27_port, PC_o(26) => IRAM_Addr_o_26_port
                           , PC_o(25) => IRAM_Addr_o_25_port, PC_o(24) => 
                           IRAM_Addr_o_24_port, PC_o(23) => IRAM_Addr_o_23_port
                           , PC_o(22) => IRAM_Addr_o_22_port, PC_o(21) => 
                           IRAM_Addr_o_21_port, PC_o(20) => IRAM_Addr_o_20_port
                           , PC_o(19) => IRAM_Addr_o_19_port, PC_o(18) => 
                           IRAM_Addr_o_18_port, PC_o(17) => IRAM_Addr_o_17_port
                           , PC_o(16) => IRAM_Addr_o_16_port, PC_o(15) => 
                           IRAM_Addr_o_15_port, PC_o(14) => IRAM_Addr_o_14_port
                           , PC_o(13) => IRAM_Addr_o_13_port, PC_o(12) => 
                           IRAM_Addr_o_12_port, PC_o(11) => IRAM_Addr_o_11_port
                           , PC_o(10) => IRAM_Addr_o_10_port, PC_o(9) => 
                           IRAM_Addr_o_9_port, PC_o(8) => IRAM_Addr_o_8_port, 
                           PC_o(7) => IRAM_Addr_o_7_port, PC_o(6) => 
                           IRAM_Addr_o_6_port, PC_o(5) => IRAM_Addr_o_5_port, 
                           PC_o(4) => IRAM_Addr_o_4_port, PC_o(3) => 
                           IRAM_Addr_o_3_port, PC_o(2) => IRAM_Addr_o_2_port, 
                           PC_o(1) => IRAM_Addr_o_1_port, PC_o(0) => 
                           IRAM_Addr_o_0_port, PC4_o(31) => PC4_31_port, 
                           PC4_o(30) => PC4_30_port, PC4_o(29) => PC4_29_port, 
                           PC4_o(28) => PC4_28_port, PC4_o(27) => PC4_27_port, 
                           PC4_o(26) => PC4_26_port, PC4_o(25) => PC4_25_port, 
                           PC4_o(24) => PC4_24_port, PC4_o(23) => PC4_23_port, 
                           PC4_o(22) => PC4_22_port, PC4_o(21) => PC4_21_port, 
                           PC4_o(20) => PC4_20_port, PC4_o(19) => PC4_19_port, 
                           PC4_o(18) => PC4_18_port, PC4_o(17) => PC4_17_port, 
                           PC4_o(16) => PC4_16_port, PC4_o(15) => PC4_15_port, 
                           PC4_o(14) => PC4_14_port, PC4_o(13) => PC4_13_port, 
                           PC4_o(12) => PC4_12_port, PC4_o(11) => PC4_11_port, 
                           PC4_o(10) => PC4_10_port, PC4_o(9) => PC4_9_port, 
                           PC4_o(8) => PC4_8_port, PC4_o(7) => PC4_7_port, 
                           PC4_o(6) => PC4_6_port, PC4_o(5) => PC4_5_port, 
                           PC4_o(4) => PC4_4_port, PC4_o(3) => PC4_3_port, 
                           PC4_o(2) => PC4_2_port, PC4_o(1) => PC4_1_port, 
                           PC4_o(0) => PC4_0_port, PC_BUS_pre_BTB(31) => 
                           TARGET_PC_31_port, PC_BUS_pre_BTB(30) => 
                           TARGET_PC_30_port, PC_BUS_pre_BTB(29) => n5, 
                           PC_BUS_pre_BTB(28) => TARGET_PC_28_port, 
                           PC_BUS_pre_BTB(27) => TARGET_PC_27_port, 
                           PC_BUS_pre_BTB(26) => TARGET_PC_26_port, 
                           PC_BUS_pre_BTB(25) => TARGET_PC_25_port, 
                           PC_BUS_pre_BTB(24) => TARGET_PC_24_port, 
                           PC_BUS_pre_BTB(23) => TARGET_PC_23_port, 
                           PC_BUS_pre_BTB(22) => TARGET_PC_22_port, 
                           PC_BUS_pre_BTB(21) => TARGET_PC_21_port, 
                           PC_BUS_pre_BTB(20) => TARGET_PC_20_port, 
                           PC_BUS_pre_BTB(19) => TARGET_PC_19_port, 
                           PC_BUS_pre_BTB(18) => TARGET_PC_18_port, 
                           PC_BUS_pre_BTB(17) => TARGET_PC_17_port, 
                           PC_BUS_pre_BTB(16) => TARGET_PC_16_port, 
                           PC_BUS_pre_BTB(15) => TARGET_PC_15_port, 
                           PC_BUS_pre_BTB(14) => TARGET_PC_14_port, 
                           PC_BUS_pre_BTB(13) => TARGET_PC_13_port, 
                           PC_BUS_pre_BTB(12) => TARGET_PC_12_port, 
                           PC_BUS_pre_BTB(11) => TARGET_PC_11_port, 
                           PC_BUS_pre_BTB(10) => TARGET_PC_10_port, 
                           PC_BUS_pre_BTB(9) => TARGET_PC_9_port, 
                           PC_BUS_pre_BTB(8) => TARGET_PC_8_port, 
                           PC_BUS_pre_BTB(7) => TARGET_PC_7_port, 
                           PC_BUS_pre_BTB(6) => TARGET_PC_6_port, 
                           PC_BUS_pre_BTB(5) => TARGET_PC_5_port, 
                           PC_BUS_pre_BTB(4) => TARGET_PC_4_port, 
                           PC_BUS_pre_BTB(3) => TARGET_PC_3_port, 
                           PC_BUS_pre_BTB(2) => TARGET_PC_2_port, 
                           PC_BUS_pre_BTB(1) => TARGET_PC_1_port, 
                           PC_BUS_pre_BTB(0) => TARGET_PC_0_port, stall_i => 
                           stall_fetch, take_prediction_i => take_prediction, 
                           mispredict_i => mispredict, predicted_PC(31) => 
                           predicted_PC_31_port, predicted_PC(30) => 
                           predicted_PC_30_port, predicted_PC(29) => 
                           predicted_PC_29_port, predicted_PC(28) => 
                           predicted_PC_28_port, predicted_PC(27) => 
                           predicted_PC_27_port, predicted_PC(26) => 
                           predicted_PC_26_port, predicted_PC(25) => 
                           predicted_PC_25_port, predicted_PC(24) => 
                           predicted_PC_24_port, predicted_PC(23) => 
                           predicted_PC_23_port, predicted_PC(22) => 
                           predicted_PC_22_port, predicted_PC(21) => 
                           predicted_PC_21_port, predicted_PC(20) => 
                           predicted_PC_20_port, predicted_PC(19) => 
                           predicted_PC_19_port, predicted_PC(18) => 
                           predicted_PC_18_port, predicted_PC(17) => 
                           predicted_PC_17_port, predicted_PC(16) => 
                           predicted_PC_16_port, predicted_PC(15) => 
                           predicted_PC_15_port, predicted_PC(14) => 
                           predicted_PC_14_port, predicted_PC(13) => 
                           predicted_PC_13_port, predicted_PC(12) => 
                           predicted_PC_12_port, predicted_PC(11) => 
                           predicted_PC_11_port, predicted_PC(10) => 
                           predicted_PC_10_port, predicted_PC(9) => 
                           predicted_PC_9_port, predicted_PC(8) => 
                           predicted_PC_8_port, predicted_PC(7) => 
                           predicted_PC_7_port, predicted_PC(6) => 
                           predicted_PC_6_port, predicted_PC(5) => 
                           predicted_PC_5_port, predicted_PC(4) => 
                           predicted_PC_4_port, predicted_PC(3) => 
                           predicted_PC_3_port, predicted_PC(2) => 
                           predicted_PC_2_port, predicted_PC(1) => 
                           predicted_PC_1_port, predicted_PC(0) => 
                           predicted_PC_0_port, clk => clock, rst => rst);
   UBTB : btb_N_LINES4_SIZE32 port map( clock => clock, reset => rst, stall_i 
                           => stall_btb, TAG_i(3) => IRAM_Addr_o_5_port, 
                           TAG_i(2) => IRAM_Addr_o_4_port, TAG_i(1) => 
                           IRAM_Addr_o_3_port, TAG_i(0) => IRAM_Addr_o_2_port, 
                           target_PC_i(31) => TARGET_PC_31_port, 
                           target_PC_i(30) => TARGET_PC_30_port, 
                           target_PC_i(29) => n5, target_PC_i(28) => 
                           TARGET_PC_28_port, target_PC_i(27) => 
                           TARGET_PC_27_port, target_PC_i(26) => 
                           TARGET_PC_26_port, target_PC_i(25) => 
                           TARGET_PC_25_port, target_PC_i(24) => 
                           TARGET_PC_24_port, target_PC_i(23) => 
                           TARGET_PC_23_port, target_PC_i(22) => 
                           TARGET_PC_22_port, target_PC_i(21) => 
                           TARGET_PC_21_port, target_PC_i(20) => 
                           TARGET_PC_20_port, target_PC_i(19) => 
                           TARGET_PC_19_port, target_PC_i(18) => 
                           TARGET_PC_18_port, target_PC_i(17) => 
                           TARGET_PC_17_port, target_PC_i(16) => 
                           TARGET_PC_16_port, target_PC_i(15) => 
                           TARGET_PC_15_port, target_PC_i(14) => 
                           TARGET_PC_14_port, target_PC_i(13) => 
                           TARGET_PC_13_port, target_PC_i(12) => 
                           TARGET_PC_12_port, target_PC_i(11) => 
                           TARGET_PC_11_port, target_PC_i(10) => 
                           TARGET_PC_10_port, target_PC_i(9) => 
                           TARGET_PC_9_port, target_PC_i(8) => TARGET_PC_8_port
                           , target_PC_i(7) => TARGET_PC_7_port, target_PC_i(6)
                           => TARGET_PC_6_port, target_PC_i(5) => 
                           TARGET_PC_5_port, target_PC_i(4) => TARGET_PC_4_port
                           , target_PC_i(3) => TARGET_PC_3_port, target_PC_i(2)
                           => TARGET_PC_2_port, target_PC_i(1) => 
                           TARGET_PC_1_port, target_PC_i(0) => TARGET_PC_0_port
                           , was_taken_i => was_taken, predicted_next_PC_o(31) 
                           => predicted_PC_31_port, predicted_next_PC_o(30) => 
                           predicted_PC_30_port, predicted_next_PC_o(29) => 
                           predicted_PC_29_port, predicted_next_PC_o(28) => 
                           predicted_PC_28_port, predicted_next_PC_o(27) => 
                           predicted_PC_27_port, predicted_next_PC_o(26) => 
                           predicted_PC_26_port, predicted_next_PC_o(25) => 
                           predicted_PC_25_port, predicted_next_PC_o(24) => 
                           predicted_PC_24_port, predicted_next_PC_o(23) => 
                           predicted_PC_23_port, predicted_next_PC_o(22) => 
                           predicted_PC_22_port, predicted_next_PC_o(21) => 
                           predicted_PC_21_port, predicted_next_PC_o(20) => 
                           predicted_PC_20_port, predicted_next_PC_o(19) => 
                           predicted_PC_19_port, predicted_next_PC_o(18) => 
                           predicted_PC_18_port, predicted_next_PC_o(17) => 
                           predicted_PC_17_port, predicted_next_PC_o(16) => 
                           predicted_PC_16_port, predicted_next_PC_o(15) => 
                           predicted_PC_15_port, predicted_next_PC_o(14) => 
                           predicted_PC_14_port, predicted_next_PC_o(13) => 
                           predicted_PC_13_port, predicted_next_PC_o(12) => 
                           predicted_PC_12_port, predicted_next_PC_o(11) => 
                           predicted_PC_11_port, predicted_next_PC_o(10) => 
                           predicted_PC_10_port, predicted_next_PC_o(9) => 
                           predicted_PC_9_port, predicted_next_PC_o(8) => 
                           predicted_PC_8_port, predicted_next_PC_o(7) => 
                           predicted_PC_7_port, predicted_next_PC_o(6) => 
                           predicted_PC_6_port, predicted_next_PC_o(5) => 
                           predicted_PC_5_port, predicted_next_PC_o(4) => 
                           predicted_PC_4_port, predicted_next_PC_o(3) => 
                           predicted_PC_3_port, predicted_next_PC_o(2) => 
                           predicted_PC_2_port, predicted_next_PC_o(1) => 
                           predicted_PC_1_port, predicted_next_PC_o(0) => 
                           predicted_PC_0_port, taken_o => take_prediction, 
                           mispredict_o => mispredict);
   UFEETCH_REGS : fetch_regs port map( NPCF_i(31) => PC4_31_port, NPCF_i(30) =>
                           PC4_30_port, NPCF_i(29) => PC4_29_port, NPCF_i(28) 
                           => PC4_28_port, NPCF_i(27) => PC4_27_port, 
                           NPCF_i(26) => PC4_26_port, NPCF_i(25) => PC4_25_port
                           , NPCF_i(24) => PC4_24_port, NPCF_i(23) => 
                           PC4_23_port, NPCF_i(22) => PC4_22_port, NPCF_i(21) 
                           => PC4_21_port, NPCF_i(20) => PC4_20_port, 
                           NPCF_i(19) => PC4_19_port, NPCF_i(18) => PC4_18_port
                           , NPCF_i(17) => PC4_17_port, NPCF_i(16) => 
                           PC4_16_port, NPCF_i(15) => PC4_15_port, NPCF_i(14) 
                           => PC4_14_port, NPCF_i(13) => PC4_13_port, 
                           NPCF_i(12) => PC4_12_port, NPCF_i(11) => PC4_11_port
                           , NPCF_i(10) => PC4_10_port, NPCF_i(9) => PC4_9_port
                           , NPCF_i(8) => PC4_8_port, NPCF_i(7) => PC4_7_port, 
                           NPCF_i(6) => PC4_6_port, NPCF_i(5) => PC4_5_port, 
                           NPCF_i(4) => PC4_4_port, NPCF_i(3) => PC4_3_port, 
                           NPCF_i(2) => PC4_2_port, NPCF_i(1) => PC4_1_port, 
                           NPCF_i(0) => PC4_0_port, IR_i(31) => IRAM_Dout_i(31)
                           , IR_i(30) => IRAM_Dout_i(30), IR_i(29) => 
                           IRAM_Dout_i(29), IR_i(28) => IRAM_Dout_i(28), 
                           IR_i(27) => IRAM_Dout_i(27), IR_i(26) => 
                           IRAM_Dout_i(26), IR_i(25) => IRAM_Dout_i(25), 
                           IR_i(24) => IRAM_Dout_i(24), IR_i(23) => 
                           IRAM_Dout_i(23), IR_i(22) => IRAM_Dout_i(22), 
                           IR_i(21) => IRAM_Dout_i(21), IR_i(20) => 
                           IRAM_Dout_i(20), IR_i(19) => IRAM_Dout_i(19), 
                           IR_i(18) => IRAM_Dout_i(18), IR_i(17) => 
                           IRAM_Dout_i(17), IR_i(16) => IRAM_Dout_i(16), 
                           IR_i(15) => IRAM_Dout_i(15), IR_i(14) => 
                           IRAM_Dout_i(14), IR_i(13) => IRAM_Dout_i(13), 
                           IR_i(12) => IRAM_Dout_i(12), IR_i(11) => 
                           IRAM_Dout_i(11), IR_i(10) => IRAM_Dout_i(10), 
                           IR_i(9) => IRAM_Dout_i(9), IR_i(8) => IRAM_Dout_i(8)
                           , IR_i(7) => IRAM_Dout_i(7), IR_i(6) => 
                           IRAM_Dout_i(6), IR_i(5) => IRAM_Dout_i(5), IR_i(4) 
                           => IRAM_Dout_i(4), IR_i(3) => IRAM_Dout_i(3), 
                           IR_i(2) => IRAM_Dout_i(2), IR_i(1) => IRAM_Dout_i(1)
                           , IR_i(0) => IRAM_Dout_i(0), NPCF_o(31) => 
                           NPCF_31_port, NPCF_o(30) => NPCF_30_port, NPCF_o(29)
                           => NPCF_29_port, NPCF_o(28) => NPCF_28_port, 
                           NPCF_o(27) => NPCF_27_port, NPCF_o(26) => 
                           NPCF_26_port, NPCF_o(25) => NPCF_25_port, NPCF_o(24)
                           => NPCF_24_port, NPCF_o(23) => NPCF_23_port, 
                           NPCF_o(22) => NPCF_22_port, NPCF_o(21) => 
                           NPCF_21_port, NPCF_o(20) => NPCF_20_port, NPCF_o(19)
                           => NPCF_19_port, NPCF_o(18) => NPCF_18_port, 
                           NPCF_o(17) => NPCF_17_port, NPCF_o(16) => 
                           NPCF_16_port, NPCF_o(15) => NPCF_15_port, NPCF_o(14)
                           => NPCF_14_port, NPCF_o(13) => NPCF_13_port, 
                           NPCF_o(12) => NPCF_12_port, NPCF_o(11) => 
                           NPCF_11_port, NPCF_o(10) => NPCF_10_port, NPCF_o(9) 
                           => NPCF_9_port, NPCF_o(8) => NPCF_8_port, NPCF_o(7) 
                           => NPCF_7_port, NPCF_o(6) => NPCF_6_port, NPCF_o(5) 
                           => NPCF_5_port, NPCF_o(4) => NPCF_4_port, NPCF_o(3) 
                           => NPCF_3_port, NPCF_o(2) => NPCF_2_port, NPCF_o(1) 
                           => NPCF_1_port, NPCF_o(0) => NPCF_0_port, IR_o(31) 
                           => IR_31_port, IR_o(30) => IR_30_port, IR_o(29) => 
                           IR_29_port, IR_o(28) => IR_28_port, IR_o(27) => 
                           IR_27_port, IR_o(26) => IR_26_port, IR_o(25) => 
                           IR_25_port, IR_o(24) => IR_24_port, IR_o(23) => 
                           IR_23_port, IR_o(22) => IR_22_port, IR_o(21) => 
                           IR_21_port, IR_o(20) => IR_20_port, IR_o(19) => 
                           IR_19_port, IR_o(18) => IR_18_port, IR_o(17) => 
                           IR_17_port, IR_o(16) => IR_16_port, IR_o(15) => 
                           IR_15_port, IR_o(14) => IR_14_port, IR_o(13) => 
                           IR_13_port, IR_o(12) => IR_12_port, IR_o(11) => 
                           IR_11_port, IR_o(10) => IR_10_port, IR_o(9) => 
                           IR_9_port, IR_o(8) => IR_8_port, IR_o(7) => 
                           IR_7_port, IR_o(6) => IR_6_port, IR_o(5) => 
                           IR_5_port, IR_o(4) => IR_4_port, IR_o(3) => 
                           IR_3_port, IR_o(2) => IR_2_port, IR_o(1) => 
                           IR_1_port, IR_o(0) => IR_0_port, stall_i => 
                           stall_decode, clk => clock, rst => rst);
   UJUMP_LOGIC : jump_logic port map( NPCF_i(31) => NPCF_31_port, NPCF_i(30) =>
                           NPCF_30_port, NPCF_i(29) => NPCF_29_port, NPCF_i(28)
                           => NPCF_28_port, NPCF_i(27) => NPCF_27_port, 
                           NPCF_i(26) => NPCF_26_port, NPCF_i(25) => 
                           NPCF_25_port, NPCF_i(24) => NPCF_24_port, NPCF_i(23)
                           => NPCF_23_port, NPCF_i(22) => NPCF_22_port, 
                           NPCF_i(21) => NPCF_21_port, NPCF_i(20) => 
                           NPCF_20_port, NPCF_i(19) => NPCF_19_port, NPCF_i(18)
                           => NPCF_18_port, NPCF_i(17) => NPCF_17_port, 
                           NPCF_i(16) => NPCF_16_port, NPCF_i(15) => 
                           NPCF_15_port, NPCF_i(14) => NPCF_14_port, NPCF_i(13)
                           => NPCF_13_port, NPCF_i(12) => NPCF_12_port, 
                           NPCF_i(11) => NPCF_11_port, NPCF_i(10) => 
                           NPCF_10_port, NPCF_i(9) => NPCF_9_port, NPCF_i(8) =>
                           NPCF_8_port, NPCF_i(7) => NPCF_7_port, NPCF_i(6) => 
                           NPCF_6_port, NPCF_i(5) => NPCF_5_port, NPCF_i(4) => 
                           NPCF_4_port, NPCF_i(3) => NPCF_3_port, NPCF_i(2) => 
                           NPCF_2_port, NPCF_i(1) => NPCF_1_port, NPCF_i(0) => 
                           NPCF_0_port, IR_i(31) => n14, IR_i(30) => n15, 
                           IR_i(29) => n16, IR_i(28) => n17, IR_i(27) => n18, 
                           IR_i(26) => n19, IR_i(25) => IR_25_port, IR_i(24) =>
                           IR_24_port, IR_i(23) => IR_23_port, IR_i(22) => 
                           IR_22_port, IR_i(21) => IR_21_port, IR_i(20) => 
                           IR_20_port, IR_i(19) => IR_19_port, IR_i(18) => 
                           IR_18_port, IR_i(17) => IR_17_port, IR_i(16) => 
                           IR_16_port, IR_i(15) => IR_15_port, IR_i(14) => 
                           IR_14_port, IR_i(13) => IR_13_port, IR_i(12) => 
                           IR_12_port, IR_i(11) => IR_11_port, IR_i(10) => 
                           IR_10_port, IR_i(9) => IR_9_port, IR_i(8) => 
                           IR_8_port, IR_i(7) => IR_7_port, IR_i(6) => 
                           IR_6_port, IR_i(5) => IR_5_port, IR_i(4) => 
                           IR_4_port, IR_i(3) => IR_3_port, IR_i(2) => 
                           IR_2_port, IR_i(1) => IR_1_port, IR_i(0) => 
                           IR_0_port, A_i(31) => AtoComp_31_port, A_i(30) => 
                           AtoComp_30_port, A_i(29) => AtoComp_29_port, A_i(28)
                           => AtoComp_28_port, A_i(27) => AtoComp_27_port, 
                           A_i(26) => AtoComp_26_port, A_i(25) => 
                           AtoComp_25_port, A_i(24) => AtoComp_24_port, A_i(23)
                           => AtoComp_23_port, A_i(22) => AtoComp_22_port, 
                           A_i(21) => AtoComp_21_port, A_i(20) => 
                           AtoComp_20_port, A_i(19) => AtoComp_19_port, A_i(18)
                           => AtoComp_18_port, A_i(17) => AtoComp_17_port, 
                           A_i(16) => AtoComp_16_port, A_i(15) => 
                           AtoComp_15_port, A_i(14) => AtoComp_14_port, A_i(13)
                           => AtoComp_13_port, A_i(12) => AtoComp_12_port, 
                           A_i(11) => AtoComp_11_port, A_i(10) => 
                           AtoComp_10_port, A_i(9) => AtoComp_9_port, A_i(8) =>
                           AtoComp_8_port, A_i(7) => AtoComp_7_port, A_i(6) => 
                           AtoComp_6_port, A_i(5) => AtoComp_5_port, A_i(4) => 
                           AtoComp_4_port, A_i(3) => AtoComp_3_port, A_i(2) => 
                           AtoComp_2_port, A_i(1) => AtoComp_1_port, A_i(0) => 
                           AtoComp_0_port, A_o(31) => dummy_A_31_port, A_o(30) 
                           => dummy_A_30_port, A_o(29) => dummy_A_29_port, 
                           A_o(28) => dummy_A_28_port, A_o(27) => 
                           dummy_A_27_port, A_o(26) => dummy_A_26_port, A_o(25)
                           => dummy_A_25_port, A_o(24) => dummy_A_24_port, 
                           A_o(23) => dummy_A_23_port, A_o(22) => 
                           dummy_A_22_port, A_o(21) => dummy_A_21_port, A_o(20)
                           => dummy_A_20_port, A_o(19) => dummy_A_19_port, 
                           A_o(18) => dummy_A_18_port, A_o(17) => 
                           dummy_A_17_port, A_o(16) => dummy_A_16_port, A_o(15)
                           => dummy_A_15_port, A_o(14) => dummy_A_14_port, 
                           A_o(13) => dummy_A_13_port, A_o(12) => 
                           dummy_A_12_port, A_o(11) => dummy_A_11_port, A_o(10)
                           => dummy_A_10_port, A_o(9) => dummy_A_9_port, A_o(8)
                           => dummy_A_8_port, A_o(7) => dummy_A_7_port, A_o(6) 
                           => dummy_A_6_port, A_o(5) => dummy_A_5_port, A_o(4) 
                           => dummy_A_4_port, A_o(3) => dummy_A_3_port, A_o(2) 
                           => dummy_A_2_port, A_o(1) => dummy_A_1_port, A_o(0) 
                           => dummy_A_0_port, rA_o(4) => rA2reg_4_port, rA_o(3)
                           => rA2reg_3_port, rA_o(2) => rA2reg_2_port, rA_o(1) 
                           => rA2reg_1_port, rA_o(0) => rA2reg_0_port, rB_o(4) 
                           => rB2reg_4_port, rB_o(3) => rB2reg_3_port, rB_o(2) 
                           => rB2reg_2_port, rB_o(1) => rB2reg_1_port, rB_o(0) 
                           => rB2reg_0_port, rC_o(4) => rC2reg_4_port, rC_o(3) 
                           => rC2reg_3_port, rC_o(2) => rC2reg_2_port, rC_o(1) 
                           => rC2reg_1_port, rC_o(0) => rC2reg_0_port, 
                           branch_target_o(31) => dummy_branch_target_31_port, 
                           branch_target_o(30) => dummy_branch_target_30_port, 
                           branch_target_o(29) => dummy_branch_target_29_port, 
                           branch_target_o(28) => dummy_branch_target_28_port, 
                           branch_target_o(27) => dummy_branch_target_27_port, 
                           branch_target_o(26) => dummy_branch_target_26_port, 
                           branch_target_o(25) => dummy_branch_target_25_port, 
                           branch_target_o(24) => dummy_branch_target_24_port, 
                           branch_target_o(23) => dummy_branch_target_23_port, 
                           branch_target_o(22) => dummy_branch_target_22_port, 
                           branch_target_o(21) => dummy_branch_target_21_port, 
                           branch_target_o(20) => dummy_branch_target_20_port, 
                           branch_target_o(19) => dummy_branch_target_19_port, 
                           branch_target_o(18) => dummy_branch_target_18_port, 
                           branch_target_o(17) => dummy_branch_target_17_port, 
                           branch_target_o(16) => dummy_branch_target_16_port, 
                           branch_target_o(15) => dummy_branch_target_15_port, 
                           branch_target_o(14) => dummy_branch_target_14_port, 
                           branch_target_o(13) => dummy_branch_target_13_port, 
                           branch_target_o(12) => dummy_branch_target_12_port, 
                           branch_target_o(11) => dummy_branch_target_11_port, 
                           branch_target_o(10) => dummy_branch_target_10_port, 
                           branch_target_o(9) => dummy_branch_target_9_port, 
                           branch_target_o(8) => dummy_branch_target_8_port, 
                           branch_target_o(7) => dummy_branch_target_7_port, 
                           branch_target_o(6) => dummy_branch_target_6_port, 
                           branch_target_o(5) => dummy_branch_target_5_port, 
                           branch_target_o(4) => dummy_branch_target_4_port, 
                           branch_target_o(3) => dummy_branch_target_3_port, 
                           branch_target_o(2) => dummy_branch_target_2_port, 
                           branch_target_o(1) => dummy_branch_target_1_port, 
                           branch_target_o(0) => dummy_branch_target_0_port, 
                           sum_addr_o(31) => dummy_sum_addr_31_port, 
                           sum_addr_o(30) => dummy_sum_addr_30_port, 
                           sum_addr_o(29) => dummy_sum_addr_29_port, 
                           sum_addr_o(28) => dummy_sum_addr_28_port, 
                           sum_addr_o(27) => dummy_sum_addr_27_port, 
                           sum_addr_o(26) => dummy_sum_addr_26_port, 
                           sum_addr_o(25) => dummy_sum_addr_25_port, 
                           sum_addr_o(24) => dummy_sum_addr_24_port, 
                           sum_addr_o(23) => dummy_sum_addr_23_port, 
                           sum_addr_o(22) => dummy_sum_addr_22_port, 
                           sum_addr_o(21) => dummy_sum_addr_21_port, 
                           sum_addr_o(20) => dummy_sum_addr_20_port, 
                           sum_addr_o(19) => dummy_sum_addr_19_port, 
                           sum_addr_o(18) => dummy_sum_addr_18_port, 
                           sum_addr_o(17) => dummy_sum_addr_17_port, 
                           sum_addr_o(16) => dummy_sum_addr_16_port, 
                           sum_addr_o(15) => dummy_sum_addr_15_port, 
                           sum_addr_o(14) => dummy_sum_addr_14_port, 
                           sum_addr_o(13) => dummy_sum_addr_13_port, 
                           sum_addr_o(12) => dummy_sum_addr_12_port, 
                           sum_addr_o(11) => dummy_sum_addr_11_port, 
                           sum_addr_o(10) => dummy_sum_addr_10_port, 
                           sum_addr_o(9) => dummy_sum_addr_9_port, 
                           sum_addr_o(8) => dummy_sum_addr_8_port, 
                           sum_addr_o(7) => dummy_sum_addr_7_port, 
                           sum_addr_o(6) => dummy_sum_addr_6_port, 
                           sum_addr_o(5) => dummy_sum_addr_5_port, 
                           sum_addr_o(4) => dummy_sum_addr_4_port, 
                           sum_addr_o(3) => dummy_sum_addr_3_port, 
                           sum_addr_o(2) => dummy_sum_addr_2_port, 
                           sum_addr_o(1) => dummy_sum_addr_1_port, 
                           sum_addr_o(0) => dummy_sum_addr_0_port, 
                           extended_imm(31) => help_IMM_31_port, 
                           extended_imm(30) => help_IMM_30_port, 
                           extended_imm(29) => help_IMM_29_port, 
                           extended_imm(28) => help_IMM_28_port, 
                           extended_imm(27) => help_IMM_27_port, 
                           extended_imm(26) => help_IMM_26_port, 
                           extended_imm(25) => help_IMM_25_port, 
                           extended_imm(24) => help_IMM_24_port, 
                           extended_imm(23) => help_IMM_23_port, 
                           extended_imm(22) => help_IMM_22_port, 
                           extended_imm(21) => help_IMM_21_port, 
                           extended_imm(20) => help_IMM_20_port, 
                           extended_imm(19) => help_IMM_19_port, 
                           extended_imm(18) => help_IMM_18_port, 
                           extended_imm(17) => help_IMM_17_port, 
                           extended_imm(16) => help_IMM_16_port, 
                           extended_imm(15) => help_IMM_15_port, 
                           extended_imm(14) => help_IMM_14_port, 
                           extended_imm(13) => help_IMM_13_port, 
                           extended_imm(12) => help_IMM_12_port, 
                           extended_imm(11) => help_IMM_11_port, 
                           extended_imm(10) => help_IMM_10_port, 
                           extended_imm(9) => help_IMM_9_port, extended_imm(8) 
                           => help_IMM_8_port, extended_imm(7) => 
                           help_IMM_7_port, extended_imm(6) => help_IMM_6_port,
                           extended_imm(5) => help_IMM_5_port, extended_imm(4) 
                           => help_IMM_4_port, extended_imm(3) => 
                           help_IMM_3_port, extended_imm(2) => help_IMM_2_port,
                           extended_imm(1) => help_IMM_1_port, extended_imm(0) 
                           => help_IMM_0_port, taken_o => was_taken_from_jl, 
                           FW_X_i(31) => DRAM_Addr_o_31_port, FW_X_i(30) => 
                           DRAM_Addr_o_30_port, FW_X_i(29) => 
                           DRAM_Addr_o_29_port, FW_X_i(28) => 
                           DRAM_Addr_o_28_port, FW_X_i(27) => 
                           DRAM_Addr_o_27_port, FW_X_i(26) => 
                           DRAM_Addr_o_26_port, FW_X_i(25) => 
                           DRAM_Addr_o_25_port, FW_X_i(24) => 
                           DRAM_Addr_o_24_port, FW_X_i(23) => 
                           DRAM_Addr_o_23_port, FW_X_i(22) => 
                           DRAM_Addr_o_22_port, FW_X_i(21) => 
                           DRAM_Addr_o_21_port, FW_X_i(20) => 
                           DRAM_Addr_o_20_port, FW_X_i(19) => 
                           DRAM_Addr_o_19_port, FW_X_i(18) => 
                           DRAM_Addr_o_18_port, FW_X_i(17) => 
                           DRAM_Addr_o_17_port, FW_X_i(16) => 
                           DRAM_Addr_o_16_port, FW_X_i(15) => 
                           DRAM_Addr_o_15_port, FW_X_i(14) => 
                           DRAM_Addr_o_14_port, FW_X_i(13) => 
                           DRAM_Addr_o_13_port, FW_X_i(12) => 
                           DRAM_Addr_o_12_port, FW_X_i(11) => 
                           DRAM_Addr_o_11_port, FW_X_i(10) => 
                           DRAM_Addr_o_10_port, FW_X_i(9) => DRAM_Addr_o_9_port
                           , FW_X_i(8) => DRAM_Addr_o_8_port, FW_X_i(7) => 
                           DRAM_Addr_o_7_port, FW_X_i(6) => DRAM_Addr_o_6_port,
                           FW_X_i(5) => DRAM_Addr_o_5_port, FW_X_i(4) => 
                           DRAM_Addr_o_4_port, FW_X_i(3) => DRAM_Addr_o_3_port,
                           FW_X_i(2) => DRAM_Addr_o_2_port, FW_X_i(1) => 
                           DRAM_Addr_o_1_port, FW_X_i(0) => DRAM_Addr_o_0_port,
                           FW_W_i(31) => wb2reg_31_port, FW_W_i(30) => 
                           wb2reg_30_port, FW_W_i(29) => wb2reg_29_port, 
                           FW_W_i(28) => wb2reg_28_port, FW_W_i(27) => 
                           wb2reg_27_port, FW_W_i(26) => wb2reg_26_port, 
                           FW_W_i(25) => wb2reg_25_port, FW_W_i(24) => 
                           wb2reg_24_port, FW_W_i(23) => wb2reg_23_port, 
                           FW_W_i(22) => wb2reg_22_port, FW_W_i(21) => 
                           wb2reg_21_port, FW_W_i(20) => wb2reg_20_port, 
                           FW_W_i(19) => wb2reg_19_port, FW_W_i(18) => 
                           wb2reg_18_port, FW_W_i(17) => wb2reg_17_port, 
                           FW_W_i(16) => wb2reg_16_port, FW_W_i(15) => 
                           wb2reg_15_port, FW_W_i(14) => wb2reg_14_port, 
                           FW_W_i(13) => wb2reg_13_port, FW_W_i(12) => 
                           wb2reg_12_port, FW_W_i(11) => wb2reg_11_port, 
                           FW_W_i(10) => wb2reg_10_port, FW_W_i(9) => 
                           wb2reg_9_port, FW_W_i(8) => wb2reg_8_port, FW_W_i(7)
                           => wb2reg_7_port, FW_W_i(6) => wb2reg_6_port, 
                           FW_W_i(5) => wb2reg_5_port, FW_W_i(4) => 
                           wb2reg_4_port, FW_W_i(3) => wb2reg_3_port, FW_W_i(2)
                           => wb2reg_2_port, FW_W_i(1) => wb2reg_1_port, 
                           FW_W_i(0) => wb2reg_0_port, S_FW_Adec_i(1) => 
                           dummy_S_FWAdec_1_port, S_FW_Adec_i(0) => 
                           dummy_S_FWAdec_0_port, S_EXT_i => dummy_S_EXT, 
                           S_EXT_SIGN_i => dummy_S_EXT_SIGN, S_MUX_LINK_i => n6
                           , S_EQ_NEQ_i => dummy_S_EQ_NEQ);
   UCU : 
                           dlx_cu_MICROCODE_MEM_SIZE64_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE13 
                           port map( Clk => clock, Rst => rst, IR_IN(31) => 
                           IR_31_port, IR_IN(30) => IR_30_port, IR_IN(29) => 
                           IR_29_port, IR_IN(28) => IR_28_port, IR_IN(27) => 
                           IR_27_port, IR_IN(26) => IR_26_port, IR_IN(25) => 
                           IR_25_port, IR_IN(24) => IR_24_port, IR_IN(23) => 
                           IR_23_port, IR_IN(22) => IR_22_port, IR_IN(21) => 
                           IR_21_port, IR_IN(20) => IR_20_port, IR_IN(19) => 
                           IR_19_port, IR_IN(18) => IR_18_port, IR_IN(17) => 
                           IR_17_port, IR_IN(16) => IR_16_port, IR_IN(15) => 
                           n20, IR_IN(14) => n21, IR_IN(13) => n22, IR_IN(12) 
                           => n23, IR_IN(11) => n24, IR_IN(10) => IR_10_port, 
                           IR_IN(9) => IR_9_port, IR_IN(8) => IR_8_port, 
                           IR_IN(7) => IR_7_port, IR_IN(6) => IR_6_port, 
                           IR_IN(5) => IR_5_port, IR_IN(4) => IR_4_port, 
                           IR_IN(3) => IR_3_port, IR_IN(2) => IR_2_port, 
                           IR_IN(1) => IR_1_port, IR_IN(0) => IR_0_port, 
                           stall_exe_i => exe_stall_cu, mispredict_i => n4, 
                           D1_i(4) => muxed_dest2exe_4_port, D1_i(3) => 
                           muxed_dest2exe_3_port, D1_i(2) => 
                           muxed_dest2exe_2_port, D1_i(1) => 
                           muxed_dest2exe_1_port, D1_i(0) => 
                           muxed_dest2exe_0_port, D2_i(4) => n10, D2_i(3) => 
                           n12, D2_i(2) => n9, D2_i(1) => n13, D2_i(0) => n11, 
                           S1_LATCH_EN => net47162, S2_LATCH_EN => net47163, 
                           S3_LATCH_EN => net47164, S_MUX_PC_BUS(1) => 
                           dummy_S_MUX_PC_BUS_1_port, S_MUX_PC_BUS(0) => 
                           dummy_S_MUX_PC_BUS_0_port, S_EXT => dummy_S_EXT, 
                           S_EXT_SIGN => dummy_S_EXT_SIGN, S_EQ_NEQ => 
                           dummy_S_EQ_NEQ, S_MUX_DEST(1) => 
                           dummy_S_MUX_DEST_1_port, S_MUX_DEST(0) => 
                           dummy_S_MUX_DEST_0_port, S_MUX_LINK => n6, S_MEM_W_R
                           => DRAM_WR_o, S_MEM_EN => DRAM_Enable_o, S_RF_W_wb 
                           => dummy_S_RF_W_wb, S_RF_W_mem => dummy_S_RF_W_mem, 
                           S_RF_W_exe => net47165, S_MUX_ALUIN => 
                           dummy_S_MUX_ALUIN, stall_exe_o => stall_exe, 
                           stall_dec_o => stall_decode, stall_fetch_o => 
                           stall_fetch, stall_btb_o => stall_btb, was_branch_o 
                           => was_branch, was_jmp_o => was_jmp, ALU_WORD_o(12) 
                           => ALUW_dec_12_port, ALU_WORD_o(11) => 
                           ALUW_dec_11_port, ALU_WORD_o(10) => ALUW_dec_10_port
                           , ALU_WORD_o(9) => ALUW_dec_9_port, ALU_WORD_o(8) =>
                           ALUW_dec_8_port, ALU_WORD_o(7) => ALUW_dec_7_port, 
                           ALU_WORD_o(6) => ALUW_dec_6_port, ALU_WORD_o(5) => 
                           ALUW_dec_5_port, ALU_WORD_o(4) => ALUW_dec_4_port, 
                           ALU_WORD_o(3) => ALUW_dec_3_port, ALU_WORD_o(2) => 
                           ALUW_dec_2_port, ALU_WORD_o(1) => ALUW_dec_1_port, 
                           ALU_WORD_o(0) => ALUW_dec_0_port, ALU_OPCODE(0) => 
                           net47166, ALU_OPCODE(1) => net47167, ALU_OPCODE(2) 
                           => net47168, ALU_OPCODE(3) => net47169, 
                           ALU_OPCODE(4) => net47170, S_MUX_MEM_BAR => 
                           dummy_S_MUX_MEM);
   RF : dlx_regfile port map( Clk => clock, Rst => rst, ENABLE => 
                           enable_regfile, RD1 => X_Logic1_port, RD2 => 
                           X_Logic1_port, WR => dummy_S_RF_W_mem, ADD_WR(4) => 
                           n10, ADD_WR(3) => n12, ADD_WR(2) => n9, ADD_WR(1) =>
                           n13, ADD_WR(0) => n11, ADD_RD1(4) => IRAM_Dout_i(25)
                           , ADD_RD1(3) => IRAM_Dout_i(24), ADD_RD1(2) => 
                           IRAM_Dout_i(23), ADD_RD1(1) => IRAM_Dout_i(22), 
                           ADD_RD1(0) => IRAM_Dout_i(21), ADD_RD2(4) => 
                           IRAM_Dout_i(20), ADD_RD2(3) => IRAM_Dout_i(19), 
                           ADD_RD2(2) => IRAM_Dout_i(18), ADD_RD2(1) => 
                           IRAM_Dout_i(17), ADD_RD2(0) => IRAM_Dout_i(16), 
                           DATAIN(31) => W2wb_31_port, DATAIN(30) => 
                           W2wb_30_port, DATAIN(29) => W2wb_29_port, DATAIN(28)
                           => W2wb_28_port, DATAIN(27) => W2wb_27_port, 
                           DATAIN(26) => W2wb_26_port, DATAIN(25) => 
                           W2wb_25_port, DATAIN(24) => W2wb_24_port, DATAIN(23)
                           => W2wb_23_port, DATAIN(22) => W2wb_22_port, 
                           DATAIN(21) => W2wb_21_port, DATAIN(20) => 
                           W2wb_20_port, DATAIN(19) => W2wb_19_port, DATAIN(18)
                           => W2wb_18_port, DATAIN(17) => W2wb_17_port, 
                           DATAIN(16) => W2wb_16_port, DATAIN(15) => 
                           W2wb_15_port, DATAIN(14) => W2wb_14_port, DATAIN(13)
                           => W2wb_13_port, DATAIN(12) => W2wb_12_port, 
                           DATAIN(11) => W2wb_11_port, DATAIN(10) => 
                           W2wb_10_port, DATAIN(9) => W2wb_9_port, DATAIN(8) =>
                           W2wb_8_port, DATAIN(7) => W2wb_7_port, DATAIN(6) => 
                           W2wb_6_port, DATAIN(5) => W2wb_5_port, DATAIN(4) => 
                           W2wb_4_port, DATAIN(3) => W2wb_3_port, DATAIN(2) => 
                           W2wb_2_port, DATAIN(1) => W2wb_1_port, DATAIN(0) => 
                           W2wb_0_port, OUT1(31) => AtoComp_31_port, OUT1(30) 
                           => AtoComp_30_port, OUT1(29) => AtoComp_29_port, 
                           OUT1(28) => AtoComp_28_port, OUT1(27) => 
                           AtoComp_27_port, OUT1(26) => AtoComp_26_port, 
                           OUT1(25) => AtoComp_25_port, OUT1(24) => 
                           AtoComp_24_port, OUT1(23) => AtoComp_23_port, 
                           OUT1(22) => AtoComp_22_port, OUT1(21) => 
                           AtoComp_21_port, OUT1(20) => AtoComp_20_port, 
                           OUT1(19) => AtoComp_19_port, OUT1(18) => 
                           AtoComp_18_port, OUT1(17) => AtoComp_17_port, 
                           OUT1(16) => AtoComp_16_port, OUT1(15) => 
                           AtoComp_15_port, OUT1(14) => AtoComp_14_port, 
                           OUT1(13) => AtoComp_13_port, OUT1(12) => 
                           AtoComp_12_port, OUT1(11) => AtoComp_11_port, 
                           OUT1(10) => AtoComp_10_port, OUT1(9) => 
                           AtoComp_9_port, OUT1(8) => AtoComp_8_port, OUT1(7) 
                           => AtoComp_7_port, OUT1(6) => AtoComp_6_port, 
                           OUT1(5) => AtoComp_5_port, OUT1(4) => AtoComp_4_port
                           , OUT1(3) => AtoComp_3_port, OUT1(2) => 
                           AtoComp_2_port, OUT1(1) => AtoComp_1_port, OUT1(0) 
                           => AtoComp_0_port, OUT2(31) => dummy_B_31_port, 
                           OUT2(30) => dummy_B_30_port, OUT2(29) => 
                           dummy_B_29_port, OUT2(28) => dummy_B_28_port, 
                           OUT2(27) => dummy_B_27_port, OUT2(26) => 
                           dummy_B_26_port, OUT2(25) => dummy_B_25_port, 
                           OUT2(24) => dummy_B_24_port, OUT2(23) => 
                           dummy_B_23_port, OUT2(22) => dummy_B_22_port, 
                           OUT2(21) => dummy_B_21_port, OUT2(20) => 
                           dummy_B_20_port, OUT2(19) => dummy_B_19_port, 
                           OUT2(18) => dummy_B_18_port, OUT2(17) => 
                           dummy_B_17_port, OUT2(16) => dummy_B_16_port, 
                           OUT2(15) => dummy_B_15_port, OUT2(14) => 
                           dummy_B_14_port, OUT2(13) => dummy_B_13_port, 
                           OUT2(12) => dummy_B_12_port, OUT2(11) => 
                           dummy_B_11_port, OUT2(10) => dummy_B_10_port, 
                           OUT2(9) => dummy_B_9_port, OUT2(8) => dummy_B_8_port
                           , OUT2(7) => dummy_B_7_port, OUT2(6) => 
                           dummy_B_6_port, OUT2(5) => dummy_B_5_port, OUT2(4) 
                           => dummy_B_4_port, OUT2(3) => dummy_B_3_port, 
                           OUT2(2) => dummy_B_2_port, OUT2(1) => dummy_B_1_port
                           , OUT2(0) => dummy_B_0_port);
   UDECODE_REGS : decode_regs port map( A_i(31) => AtoComp_31_port, A_i(30) => 
                           AtoComp_30_port, A_i(29) => AtoComp_29_port, A_i(28)
                           => AtoComp_28_port, A_i(27) => AtoComp_27_port, 
                           A_i(26) => AtoComp_26_port, A_i(25) => 
                           AtoComp_25_port, A_i(24) => AtoComp_24_port, A_i(23)
                           => AtoComp_23_port, A_i(22) => AtoComp_22_port, 
                           A_i(21) => AtoComp_21_port, A_i(20) => 
                           AtoComp_20_port, A_i(19) => AtoComp_19_port, A_i(18)
                           => AtoComp_18_port, A_i(17) => AtoComp_17_port, 
                           A_i(16) => AtoComp_16_port, A_i(15) => 
                           AtoComp_15_port, A_i(14) => AtoComp_14_port, A_i(13)
                           => AtoComp_13_port, A_i(12) => AtoComp_12_port, 
                           A_i(11) => AtoComp_11_port, A_i(10) => 
                           AtoComp_10_port, A_i(9) => AtoComp_9_port, A_i(8) =>
                           AtoComp_8_port, A_i(7) => AtoComp_7_port, A_i(6) => 
                           AtoComp_6_port, A_i(5) => AtoComp_5_port, A_i(4) => 
                           AtoComp_4_port, A_i(3) => AtoComp_3_port, A_i(2) => 
                           AtoComp_2_port, A_i(1) => AtoComp_1_port, A_i(0) => 
                           AtoComp_0_port, B_i(31) => dummy_B_31_port, B_i(30) 
                           => dummy_B_30_port, B_i(29) => dummy_B_29_port, 
                           B_i(28) => dummy_B_28_port, B_i(27) => 
                           dummy_B_27_port, B_i(26) => dummy_B_26_port, B_i(25)
                           => dummy_B_25_port, B_i(24) => dummy_B_24_port, 
                           B_i(23) => dummy_B_23_port, B_i(22) => 
                           dummy_B_22_port, B_i(21) => dummy_B_21_port, B_i(20)
                           => dummy_B_20_port, B_i(19) => dummy_B_19_port, 
                           B_i(18) => dummy_B_18_port, B_i(17) => 
                           dummy_B_17_port, B_i(16) => dummy_B_16_port, B_i(15)
                           => dummy_B_15_port, B_i(14) => dummy_B_14_port, 
                           B_i(13) => dummy_B_13_port, B_i(12) => 
                           dummy_B_12_port, B_i(11) => dummy_B_11_port, B_i(10)
                           => dummy_B_10_port, B_i(9) => dummy_B_9_port, B_i(8)
                           => dummy_B_8_port, B_i(7) => dummy_B_7_port, B_i(6) 
                           => dummy_B_6_port, B_i(5) => dummy_B_5_port, B_i(4) 
                           => dummy_B_4_port, B_i(3) => dummy_B_3_port, B_i(2) 
                           => dummy_B_2_port, B_i(1) => dummy_B_1_port, B_i(0) 
                           => dummy_B_0_port, rA_i(4) => rA2reg_4_port, rA_i(3)
                           => rA2reg_3_port, rA_i(2) => rA2reg_2_port, rA_i(1) 
                           => rA2reg_1_port, rA_i(0) => rA2reg_0_port, rB_i(4) 
                           => rB2reg_4_port, rB_i(3) => rB2reg_3_port, rB_i(2) 
                           => rB2reg_2_port, rB_i(1) => rB2reg_1_port, rB_i(0) 
                           => rB2reg_0_port, rC_i(4) => rC2reg_4_port, rC_i(3) 
                           => rC2reg_3_port, rC_i(2) => rC2reg_2_port, rC_i(1) 
                           => rC2reg_1_port, rC_i(0) => rC2reg_0_port, 
                           IMM_i(31) => help_IMM_31_port, IMM_i(30) => 
                           help_IMM_30_port, IMM_i(29) => help_IMM_29_port, 
                           IMM_i(28) => help_IMM_28_port, IMM_i(27) => 
                           help_IMM_27_port, IMM_i(26) => help_IMM_26_port, 
                           IMM_i(25) => help_IMM_25_port, IMM_i(24) => 
                           help_IMM_24_port, IMM_i(23) => help_IMM_23_port, 
                           IMM_i(22) => help_IMM_22_port, IMM_i(21) => 
                           help_IMM_21_port, IMM_i(20) => help_IMM_20_port, 
                           IMM_i(19) => help_IMM_19_port, IMM_i(18) => 
                           help_IMM_18_port, IMM_i(17) => help_IMM_17_port, 
                           IMM_i(16) => help_IMM_16_port, IMM_i(15) => 
                           help_IMM_15_port, IMM_i(14) => help_IMM_14_port, 
                           IMM_i(13) => help_IMM_13_port, IMM_i(12) => 
                           help_IMM_12_port, IMM_i(11) => help_IMM_11_port, 
                           IMM_i(10) => help_IMM_10_port, IMM_i(9) => 
                           help_IMM_9_port, IMM_i(8) => help_IMM_8_port, 
                           IMM_i(7) => help_IMM_7_port, IMM_i(6) => 
                           help_IMM_6_port, IMM_i(5) => help_IMM_5_port, 
                           IMM_i(4) => help_IMM_4_port, IMM_i(3) => 
                           help_IMM_3_port, IMM_i(2) => help_IMM_2_port, 
                           IMM_i(1) => help_IMM_1_port, IMM_i(0) => 
                           help_IMM_0_port, ALUW_i(12) => ALUW_dec_12_port, 
                           ALUW_i(11) => ALUW_dec_11_port, ALUW_i(10) => 
                           ALUW_dec_10_port, ALUW_i(9) => ALUW_dec_9_port, 
                           ALUW_i(8) => ALUW_dec_8_port, ALUW_i(7) => 
                           ALUW_dec_7_port, ALUW_i(6) => ALUW_dec_6_port, 
                           ALUW_i(5) => ALUW_dec_5_port, ALUW_i(4) => 
                           ALUW_dec_4_port, ALUW_i(3) => ALUW_dec_3_port, 
                           ALUW_i(2) => ALUW_dec_2_port, ALUW_i(1) => 
                           ALUW_dec_1_port, ALUW_i(0) => ALUW_dec_0_port, 
                           A_o(31) => A2exe_31_port, A_o(30) => A2exe_30_port, 
                           A_o(29) => A2exe_29_port, A_o(28) => A2exe_28_port, 
                           A_o(27) => A2exe_27_port, A_o(26) => A2exe_26_port, 
                           A_o(25) => A2exe_25_port, A_o(24) => A2exe_24_port, 
                           A_o(23) => A2exe_23_port, A_o(22) => A2exe_22_port, 
                           A_o(21) => A2exe_21_port, A_o(20) => A2exe_20_port, 
                           A_o(19) => A2exe_19_port, A_o(18) => A2exe_18_port, 
                           A_o(17) => A2exe_17_port, A_o(16) => A2exe_16_port, 
                           A_o(15) => A2exe_15_port, A_o(14) => A2exe_14_port, 
                           A_o(13) => A2exe_13_port, A_o(12) => A2exe_12_port, 
                           A_o(11) => A2exe_11_port, A_o(10) => A2exe_10_port, 
                           A_o(9) => A2exe_9_port, A_o(8) => A2exe_8_port, 
                           A_o(7) => A2exe_7_port, A_o(6) => A2exe_6_port, 
                           A_o(5) => A2exe_5_port, A_o(4) => A2exe_4_port, 
                           A_o(3) => A2exe_3_port, A_o(2) => A2exe_2_port, 
                           A_o(1) => A2exe_1_port, A_o(0) => A2exe_0_port, 
                           B_o(31) => B2exe_31_port, B_o(30) => B2exe_30_port, 
                           B_o(29) => B2exe_29_port, B_o(28) => B2exe_28_port, 
                           B_o(27) => B2exe_27_port, B_o(26) => B2exe_26_port, 
                           B_o(25) => B2exe_25_port, B_o(24) => B2exe_24_port, 
                           B_o(23) => B2exe_23_port, B_o(22) => B2exe_22_port, 
                           B_o(21) => B2exe_21_port, B_o(20) => B2exe_20_port, 
                           B_o(19) => B2exe_19_port, B_o(18) => B2exe_18_port, 
                           B_o(17) => B2exe_17_port, B_o(16) => B2exe_16_port, 
                           B_o(15) => B2exe_15_port, B_o(14) => B2exe_14_port, 
                           B_o(13) => B2exe_13_port, B_o(12) => B2exe_12_port, 
                           B_o(11) => B2exe_11_port, B_o(10) => B2exe_10_port, 
                           B_o(9) => B2exe_9_port, B_o(8) => B2exe_8_port, 
                           B_o(7) => B2exe_7_port, B_o(6) => B2exe_6_port, 
                           B_o(5) => B2exe_5_port, B_o(4) => B2exe_4_port, 
                           B_o(3) => B2exe_3_port, B_o(2) => B2exe_2_port, 
                           B_o(1) => B2exe_1_port, B_o(0) => B2exe_0_port, 
                           rA_o(4) => rA2fw_4_port, rA_o(3) => rA2fw_3_port, 
                           rA_o(2) => rA2fw_2_port, rA_o(1) => rA2fw_1_port, 
                           rA_o(0) => rA2fw_0_port, rB_o(4) => rB2mux_4_port, 
                           rB_o(3) => rB2mux_3_port, rB_o(2) => rB2mux_2_port, 
                           rB_o(1) => rB2mux_1_port, rB_o(0) => rB2mux_0_port, 
                           rC_o(4) => rC2mux_4_port, rC_o(3) => rC2mux_3_port, 
                           rC_o(2) => rC2mux_2_port, rC_o(1) => rC2mux_1_port, 
                           rC_o(0) => rC2mux_0_port, IMM_o(31) => 
                           IMM2exe_31_port, IMM_o(30) => IMM2exe_30_port, 
                           IMM_o(29) => IMM2exe_29_port, IMM_o(28) => 
                           IMM2exe_28_port, IMM_o(27) => IMM2exe_27_port, 
                           IMM_o(26) => IMM2exe_26_port, IMM_o(25) => 
                           IMM2exe_25_port, IMM_o(24) => IMM2exe_24_port, 
                           IMM_o(23) => IMM2exe_23_port, IMM_o(22) => 
                           IMM2exe_22_port, IMM_o(21) => IMM2exe_21_port, 
                           IMM_o(20) => IMM2exe_20_port, IMM_o(19) => 
                           IMM2exe_19_port, IMM_o(18) => IMM2exe_18_port, 
                           IMM_o(17) => IMM2exe_17_port, IMM_o(16) => 
                           IMM2exe_16_port, IMM_o(15) => IMM2exe_15_port, 
                           IMM_o(14) => IMM2exe_14_port, IMM_o(13) => 
                           IMM2exe_13_port, IMM_o(12) => IMM2exe_12_port, 
                           IMM_o(11) => IMM2exe_11_port, IMM_o(10) => 
                           IMM2exe_10_port, IMM_o(9) => IMM2exe_9_port, 
                           IMM_o(8) => IMM2exe_8_port, IMM_o(7) => 
                           IMM2exe_7_port, IMM_o(6) => IMM2exe_6_port, IMM_o(5)
                           => IMM2exe_5_port, IMM_o(4) => IMM2exe_4_port, 
                           IMM_o(3) => IMM2exe_3_port, IMM_o(2) => 
                           IMM2exe_2_port, IMM_o(1) => IMM2exe_1_port, IMM_o(0)
                           => IMM2exe_0_port, ALUW_o(12) => ALUW_12_port, 
                           ALUW_o(11) => ALUW_11_port, ALUW_o(10) => 
                           ALUW_10_port, ALUW_o(9) => ALUW_9_port, ALUW_o(8) =>
                           ALUW_8_port, ALUW_o(7) => ALUW_7_port, ALUW_o(6) => 
                           ALUW_6_port, ALUW_o(5) => ALUW_5_port, ALUW_o(4) => 
                           ALUW_4_port, ALUW_o(3) => ALUW_3_port, ALUW_o(2) => 
                           ALUW_2_port, ALUW_o(1) => ALUW_1_port, ALUW_o(0) => 
                           ALUW_0_port, stall_i => stall_exe, clk => clock, rst
                           => rst);
   UEXECUTE_REGS : execute_regs port map( X_i(31) => X2mem_31_port, X_i(30) => 
                           X2mem_30_port, X_i(29) => X2mem_29_port, X_i(28) => 
                           X2mem_28_port, X_i(27) => X2mem_27_port, X_i(26) => 
                           X2mem_26_port, X_i(25) => X2mem_25_port, X_i(24) => 
                           X2mem_24_port, X_i(23) => X2mem_23_port, X_i(22) => 
                           X2mem_22_port, X_i(21) => X2mem_21_port, X_i(20) => 
                           X2mem_20_port, X_i(19) => X2mem_19_port, X_i(18) => 
                           X2mem_18_port, X_i(17) => X2mem_17_port, X_i(16) => 
                           X2mem_16_port, X_i(15) => X2mem_15_port, X_i(14) => 
                           X2mem_14_port, X_i(13) => X2mem_13_port, X_i(12) => 
                           X2mem_12_port, X_i(11) => X2mem_11_port, X_i(10) => 
                           X2mem_10_port, X_i(9) => X2mem_9_port, X_i(8) => 
                           X2mem_8_port, X_i(7) => X2mem_7_port, X_i(6) => 
                           X2mem_6_port, X_i(5) => X2mem_5_port, X_i(4) => 
                           X2mem_4_port, X_i(3) => X2mem_3_port, X_i(2) => 
                           X2mem_2_port, X_i(1) => X2mem_1_port, X_i(0) => 
                           X2mem_0_port, S_i(31) => S2mem_31_port, S_i(30) => 
                           S2mem_30_port, S_i(29) => S2mem_29_port, S_i(28) => 
                           S2mem_28_port, S_i(27) => S2mem_27_port, S_i(26) => 
                           S2mem_26_port, S_i(25) => S2mem_25_port, S_i(24) => 
                           S2mem_24_port, S_i(23) => S2mem_23_port, S_i(22) => 
                           S2mem_22_port, S_i(21) => S2mem_21_port, S_i(20) => 
                           S2mem_20_port, S_i(19) => S2mem_19_port, S_i(18) => 
                           S2mem_18_port, S_i(17) => S2mem_17_port, S_i(16) => 
                           S2mem_16_port, S_i(15) => S2mem_15_port, S_i(14) => 
                           S2mem_14_port, S_i(13) => S2mem_13_port, S_i(12) => 
                           S2mem_12_port, S_i(11) => S2mem_11_port, S_i(10) => 
                           S2mem_10_port, S_i(9) => S2mem_9_port, S_i(8) => 
                           S2mem_8_port, S_i(7) => S2mem_7_port, S_i(6) => 
                           S2mem_6_port, S_i(5) => S2mem_5_port, S_i(4) => 
                           S2mem_4_port, S_i(3) => S2mem_3_port, S_i(2) => 
                           S2mem_2_port, S_i(1) => n7, S_i(0) => S2mem_0_port, 
                           D2_i(4) => muxed_dest2exe_4_port, D2_i(3) => 
                           muxed_dest2exe_3_port, D2_i(2) => 
                           muxed_dest2exe_2_port, D2_i(1) => 
                           muxed_dest2exe_1_port, D2_i(0) => 
                           muxed_dest2exe_0_port, X_o(31) => 
                           DRAM_Addr_o_31_port, X_o(30) => DRAM_Addr_o_30_port,
                           X_o(29) => DRAM_Addr_o_29_port, X_o(28) => 
                           DRAM_Addr_o_28_port, X_o(27) => DRAM_Addr_o_27_port,
                           X_o(26) => DRAM_Addr_o_26_port, X_o(25) => 
                           DRAM_Addr_o_25_port, X_o(24) => DRAM_Addr_o_24_port,
                           X_o(23) => DRAM_Addr_o_23_port, X_o(22) => 
                           DRAM_Addr_o_22_port, X_o(21) => DRAM_Addr_o_21_port,
                           X_o(20) => DRAM_Addr_o_20_port, X_o(19) => 
                           DRAM_Addr_o_19_port, X_o(18) => DRAM_Addr_o_18_port,
                           X_o(17) => DRAM_Addr_o_17_port, X_o(16) => 
                           DRAM_Addr_o_16_port, X_o(15) => DRAM_Addr_o_15_port,
                           X_o(14) => DRAM_Addr_o_14_port, X_o(13) => 
                           DRAM_Addr_o_13_port, X_o(12) => DRAM_Addr_o_12_port,
                           X_o(11) => DRAM_Addr_o_11_port, X_o(10) => 
                           DRAM_Addr_o_10_port, X_o(9) => DRAM_Addr_o_9_port, 
                           X_o(8) => DRAM_Addr_o_8_port, X_o(7) => 
                           DRAM_Addr_o_7_port, X_o(6) => DRAM_Addr_o_6_port, 
                           X_o(5) => DRAM_Addr_o_5_port, X_o(4) => 
                           DRAM_Addr_o_4_port, X_o(3) => DRAM_Addr_o_3_port, 
                           X_o(2) => DRAM_Addr_o_2_port, X_o(1) => 
                           DRAM_Addr_o_1_port, X_o(0) => DRAM_Addr_o_0_port, 
                           S_o(31) => DRAM_Din_o(31), S_o(30) => DRAM_Din_o(30)
                           , S_o(29) => DRAM_Din_o(29), S_o(28) => 
                           DRAM_Din_o(28), S_o(27) => DRAM_Din_o(27), S_o(26) 
                           => DRAM_Din_o(26), S_o(25) => DRAM_Din_o(25), 
                           S_o(24) => DRAM_Din_o(24), S_o(23) => DRAM_Din_o(23)
                           , S_o(22) => DRAM_Din_o(22), S_o(21) => 
                           DRAM_Din_o(21), S_o(20) => DRAM_Din_o(20), S_o(19) 
                           => DRAM_Din_o(19), S_o(18) => DRAM_Din_o(18), 
                           S_o(17) => DRAM_Din_o(17), S_o(16) => DRAM_Din_o(16)
                           , S_o(15) => DRAM_Din_o(15), S_o(14) => 
                           DRAM_Din_o(14), S_o(13) => DRAM_Din_o(13), S_o(12) 
                           => DRAM_Din_o(12), S_o(11) => DRAM_Din_o(11), 
                           S_o(10) => DRAM_Din_o(10), S_o(9) => DRAM_Din_o(9), 
                           S_o(8) => DRAM_Din_o(8), S_o(7) => DRAM_Din_o(7), 
                           S_o(6) => DRAM_Din_o(6), S_o(5) => DRAM_Din_o(5), 
                           S_o(4) => DRAM_Din_o(4), S_o(3) => DRAM_Din_o(3), 
                           S_o(2) => DRAM_Din_o(2), S_o(1) => DRAM_Din_o(1), 
                           S_o(0) => DRAM_Din_o(0), D2_o(4) => D22D3_4_port, 
                           D2_o(3) => D22D3_3_port, D2_o(2) => n8, D2_o(1) => 
                           D22D3_1_port, D2_o(0) => D22D3_0_port, stall_i => 
                           X_Logic0_port, clk => clock, rst => rst);
   UEXECUTE_BLOCK : execute_block port map( IMM_i(31) => IMM2exe_31_port, 
                           IMM_i(30) => IMM2exe_30_port, IMM_i(29) => 
                           IMM2exe_29_port, IMM_i(28) => IMM2exe_28_port, 
                           IMM_i(27) => IMM2exe_27_port, IMM_i(26) => 
                           IMM2exe_26_port, IMM_i(25) => IMM2exe_25_port, 
                           IMM_i(24) => IMM2exe_24_port, IMM_i(23) => 
                           IMM2exe_23_port, IMM_i(22) => IMM2exe_22_port, 
                           IMM_i(21) => IMM2exe_21_port, IMM_i(20) => 
                           IMM2exe_20_port, IMM_i(19) => IMM2exe_19_port, 
                           IMM_i(18) => IMM2exe_18_port, IMM_i(17) => 
                           IMM2exe_17_port, IMM_i(16) => IMM2exe_16_port, 
                           IMM_i(15) => IMM2exe_15_port, IMM_i(14) => 
                           IMM2exe_14_port, IMM_i(13) => IMM2exe_13_port, 
                           IMM_i(12) => IMM2exe_12_port, IMM_i(11) => 
                           IMM2exe_11_port, IMM_i(10) => IMM2exe_10_port, 
                           IMM_i(9) => IMM2exe_9_port, IMM_i(8) => 
                           IMM2exe_8_port, IMM_i(7) => IMM2exe_7_port, IMM_i(6)
                           => IMM2exe_6_port, IMM_i(5) => IMM2exe_5_port, 
                           IMM_i(4) => IMM2exe_4_port, IMM_i(3) => 
                           IMM2exe_3_port, IMM_i(2) => IMM2exe_2_port, IMM_i(1)
                           => IMM2exe_1_port, IMM_i(0) => IMM2exe_0_port, 
                           A_i(31) => A2exe_31_port, A_i(30) => A2exe_30_port, 
                           A_i(29) => A2exe_29_port, A_i(28) => A2exe_28_port, 
                           A_i(27) => A2exe_27_port, A_i(26) => A2exe_26_port, 
                           A_i(25) => A2exe_25_port, A_i(24) => A2exe_24_port, 
                           A_i(23) => A2exe_23_port, A_i(22) => A2exe_22_port, 
                           A_i(21) => A2exe_21_port, A_i(20) => A2exe_20_port, 
                           A_i(19) => A2exe_19_port, A_i(18) => A2exe_18_port, 
                           A_i(17) => A2exe_17_port, A_i(16) => A2exe_16_port, 
                           A_i(15) => A2exe_15_port, A_i(14) => A2exe_14_port, 
                           A_i(13) => A2exe_13_port, A_i(12) => A2exe_12_port, 
                           A_i(11) => A2exe_11_port, A_i(10) => A2exe_10_port, 
                           A_i(9) => A2exe_9_port, A_i(8) => A2exe_8_port, 
                           A_i(7) => A2exe_7_port, A_i(6) => A2exe_6_port, 
                           A_i(5) => A2exe_5_port, A_i(4) => A2exe_4_port, 
                           A_i(3) => A2exe_3_port, A_i(2) => A2exe_2_port, 
                           A_i(1) => A2exe_1_port, A_i(0) => A2exe_0_port, 
                           rB_i(4) => rB2mux_4_port, rB_i(3) => rB2mux_3_port, 
                           rB_i(2) => rB2mux_2_port, rB_i(1) => rB2mux_1_port, 
                           rB_i(0) => rB2mux_0_port, rC_i(4) => rC2mux_4_port, 
                           rC_i(3) => rC2mux_3_port, rC_i(2) => rC2mux_2_port, 
                           rC_i(1) => rC2mux_1_port, rC_i(0) => rC2mux_0_port, 
                           MUXED_B_i(31) => B2exe_31_port, MUXED_B_i(30) => 
                           B2exe_30_port, MUXED_B_i(29) => B2exe_29_port, 
                           MUXED_B_i(28) => B2exe_28_port, MUXED_B_i(27) => 
                           B2exe_27_port, MUXED_B_i(26) => B2exe_26_port, 
                           MUXED_B_i(25) => B2exe_25_port, MUXED_B_i(24) => 
                           B2exe_24_port, MUXED_B_i(23) => B2exe_23_port, 
                           MUXED_B_i(22) => B2exe_22_port, MUXED_B_i(21) => 
                           B2exe_21_port, MUXED_B_i(20) => B2exe_20_port, 
                           MUXED_B_i(19) => B2exe_19_port, MUXED_B_i(18) => 
                           B2exe_18_port, MUXED_B_i(17) => B2exe_17_port, 
                           MUXED_B_i(16) => B2exe_16_port, MUXED_B_i(15) => 
                           B2exe_15_port, MUXED_B_i(14) => B2exe_14_port, 
                           MUXED_B_i(13) => B2exe_13_port, MUXED_B_i(12) => 
                           B2exe_12_port, MUXED_B_i(11) => B2exe_11_port, 
                           MUXED_B_i(10) => B2exe_10_port, MUXED_B_i(9) => 
                           B2exe_9_port, MUXED_B_i(8) => B2exe_8_port, 
                           MUXED_B_i(7) => B2exe_7_port, MUXED_B_i(6) => 
                           B2exe_6_port, MUXED_B_i(5) => B2exe_5_port, 
                           MUXED_B_i(4) => B2exe_4_port, MUXED_B_i(3) => 
                           B2exe_3_port, MUXED_B_i(2) => B2exe_2_port, 
                           MUXED_B_i(1) => B2exe_1_port, MUXED_B_i(0) => 
                           B2exe_0_port, S_MUX_ALUIN_i => dummy_S_MUX_ALUIN, 
                           FW_X_i(31) => DRAM_Addr_o_31_port, FW_X_i(30) => 
                           DRAM_Addr_o_30_port, FW_X_i(29) => 
                           DRAM_Addr_o_29_port, FW_X_i(28) => 
                           DRAM_Addr_o_28_port, FW_X_i(27) => 
                           DRAM_Addr_o_27_port, FW_X_i(26) => 
                           DRAM_Addr_o_26_port, FW_X_i(25) => 
                           DRAM_Addr_o_25_port, FW_X_i(24) => 
                           DRAM_Addr_o_24_port, FW_X_i(23) => 
                           DRAM_Addr_o_23_port, FW_X_i(22) => 
                           DRAM_Addr_o_22_port, FW_X_i(21) => 
                           DRAM_Addr_o_21_port, FW_X_i(20) => 
                           DRAM_Addr_o_20_port, FW_X_i(19) => 
                           DRAM_Addr_o_19_port, FW_X_i(18) => 
                           DRAM_Addr_o_18_port, FW_X_i(17) => 
                           DRAM_Addr_o_17_port, FW_X_i(16) => 
                           DRAM_Addr_o_16_port, FW_X_i(15) => 
                           DRAM_Addr_o_15_port, FW_X_i(14) => 
                           DRAM_Addr_o_14_port, FW_X_i(13) => 
                           DRAM_Addr_o_13_port, FW_X_i(12) => 
                           DRAM_Addr_o_12_port, FW_X_i(11) => 
                           DRAM_Addr_o_11_port, FW_X_i(10) => 
                           DRAM_Addr_o_10_port, FW_X_i(9) => DRAM_Addr_o_9_port
                           , FW_X_i(8) => DRAM_Addr_o_8_port, FW_X_i(7) => 
                           DRAM_Addr_o_7_port, FW_X_i(6) => DRAM_Addr_o_6_port,
                           FW_X_i(5) => DRAM_Addr_o_5_port, FW_X_i(4) => 
                           DRAM_Addr_o_4_port, FW_X_i(3) => DRAM_Addr_o_3_port,
                           FW_X_i(2) => DRAM_Addr_o_2_port, FW_X_i(1) => 
                           DRAM_Addr_o_1_port, FW_X_i(0) => DRAM_Addr_o_0_port,
                           FW_W_i(31) => wb2reg_31_port, FW_W_i(30) => 
                           wb2reg_30_port, FW_W_i(29) => wb2reg_29_port, 
                           FW_W_i(28) => wb2reg_28_port, FW_W_i(27) => 
                           wb2reg_27_port, FW_W_i(26) => wb2reg_26_port, 
                           FW_W_i(25) => wb2reg_25_port, FW_W_i(24) => 
                           wb2reg_24_port, FW_W_i(23) => wb2reg_23_port, 
                           FW_W_i(22) => wb2reg_22_port, FW_W_i(21) => 
                           wb2reg_21_port, FW_W_i(20) => wb2reg_20_port, 
                           FW_W_i(19) => wb2reg_19_port, FW_W_i(18) => 
                           wb2reg_18_port, FW_W_i(17) => wb2reg_17_port, 
                           FW_W_i(16) => wb2reg_16_port, FW_W_i(15) => 
                           wb2reg_15_port, FW_W_i(14) => wb2reg_14_port, 
                           FW_W_i(13) => wb2reg_13_port, FW_W_i(12) => 
                           wb2reg_12_port, FW_W_i(11) => wb2reg_11_port, 
                           FW_W_i(10) => wb2reg_10_port, FW_W_i(9) => 
                           wb2reg_9_port, FW_W_i(8) => wb2reg_8_port, FW_W_i(7)
                           => wb2reg_7_port, FW_W_i(6) => wb2reg_6_port, 
                           FW_W_i(5) => wb2reg_5_port, FW_W_i(4) => 
                           wb2reg_4_port, FW_W_i(3) => wb2reg_3_port, FW_W_i(2)
                           => wb2reg_2_port, FW_W_i(1) => wb2reg_1_port, 
                           FW_W_i(0) => wb2reg_0_port, S_FW_A_i(1) => 
                           dummy_S_FWA2exe_1_port, S_FW_A_i(0) => 
                           dummy_S_FWA2exe_0_port, S_FW_B_i(1) => 
                           dummy_S_FWB2exe_1_port, S_FW_B_i(0) => 
                           dummy_S_FWB2exe_0_port, muxed_dest(4) => 
                           muxed_dest2exe_4_port, muxed_dest(3) => 
                           muxed_dest2exe_3_port, muxed_dest(2) => 
                           muxed_dest2exe_2_port, muxed_dest(1) => 
                           muxed_dest2exe_1_port, muxed_dest(0) => 
                           muxed_dest2exe_0_port, muxed_B(31) => S2mem_31_port,
                           muxed_B(30) => S2mem_30_port, muxed_B(29) => 
                           S2mem_29_port, muxed_B(28) => S2mem_28_port, 
                           muxed_B(27) => S2mem_27_port, muxed_B(26) => 
                           S2mem_26_port, muxed_B(25) => S2mem_25_port, 
                           muxed_B(24) => S2mem_24_port, muxed_B(23) => 
                           S2mem_23_port, muxed_B(22) => S2mem_22_port, 
                           muxed_B(21) => S2mem_21_port, muxed_B(20) => 
                           S2mem_20_port, muxed_B(19) => S2mem_19_port, 
                           muxed_B(18) => S2mem_18_port, muxed_B(17) => 
                           S2mem_17_port, muxed_B(16) => S2mem_16_port, 
                           muxed_B(15) => S2mem_15_port, muxed_B(14) => 
                           S2mem_14_port, muxed_B(13) => S2mem_13_port, 
                           muxed_B(12) => S2mem_12_port, muxed_B(11) => 
                           S2mem_11_port, muxed_B(10) => S2mem_10_port, 
                           muxed_B(9) => S2mem_9_port, muxed_B(8) => 
                           S2mem_8_port, muxed_B(7) => S2mem_7_port, muxed_B(6)
                           => S2mem_6_port, muxed_B(5) => S2mem_5_port, 
                           muxed_B(4) => S2mem_4_port, muxed_B(3) => 
                           S2mem_3_port, muxed_B(2) => S2mem_2_port, muxed_B(1)
                           => n7, muxed_B(0) => S2mem_0_port, S_MUX_DEST_i(1) 
                           => dummy_S_MUX_DEST_1_port, S_MUX_DEST_i(0) => 
                           dummy_S_MUX_DEST_0_port, OP(0) => n25, OP(1) => n26,
                           OP(2) => n27, OP(3) => n28, OP(4) => n29, ALUW_i(12)
                           => ALUW_12_port, ALUW_i(11) => ALUW_11_port, 
                           ALUW_i(10) => ALUW_10_port, ALUW_i(9) => ALUW_9_port
                           , ALUW_i(8) => ALUW_8_port, ALUW_i(7) => ALUW_7_port
                           , ALUW_i(6) => ALUW_6_port, ALUW_i(5) => ALUW_5_port
                           , ALUW_i(4) => ALUW_4_port, ALUW_i(3) => ALUW_3_port
                           , ALUW_i(2) => ALUW_2_port, ALUW_i(1) => ALUW_1_port
                           , ALUW_i(0) => ALUW_0_port, DOUT(31) => 
                           X2mem_31_port, DOUT(30) => X2mem_30_port, DOUT(29) 
                           => X2mem_29_port, DOUT(28) => X2mem_28_port, 
                           DOUT(27) => X2mem_27_port, DOUT(26) => X2mem_26_port
                           , DOUT(25) => X2mem_25_port, DOUT(24) => 
                           X2mem_24_port, DOUT(23) => X2mem_23_port, DOUT(22) 
                           => X2mem_22_port, DOUT(21) => X2mem_21_port, 
                           DOUT(20) => X2mem_20_port, DOUT(19) => X2mem_19_port
                           , DOUT(18) => X2mem_18_port, DOUT(17) => 
                           X2mem_17_port, DOUT(16) => X2mem_16_port, DOUT(15) 
                           => X2mem_15_port, DOUT(14) => X2mem_14_port, 
                           DOUT(13) => X2mem_13_port, DOUT(12) => X2mem_12_port
                           , DOUT(11) => X2mem_11_port, DOUT(10) => 
                           X2mem_10_port, DOUT(9) => X2mem_9_port, DOUT(8) => 
                           X2mem_8_port, DOUT(7) => X2mem_7_port, DOUT(6) => 
                           X2mem_6_port, DOUT(5) => X2mem_5_port, DOUT(4) => 
                           X2mem_4_port, DOUT(3) => X2mem_3_port, DOUT(2) => 
                           X2mem_2_port, DOUT(1) => X2mem_1_port, DOUT(0) => 
                           X2mem_0_port, stall_o => exe_stall_cu, Clock => 
                           clock, Reset => rst);
   UMEM_REGS : mem_regs port map( W_i(31) => W2wb_31_port, W_i(30) => 
                           W2wb_30_port, W_i(29) => W2wb_29_port, W_i(28) => 
                           W2wb_28_port, W_i(27) => W2wb_27_port, W_i(26) => 
                           W2wb_26_port, W_i(25) => W2wb_25_port, W_i(24) => 
                           W2wb_24_port, W_i(23) => W2wb_23_port, W_i(22) => 
                           W2wb_22_port, W_i(21) => W2wb_21_port, W_i(20) => 
                           W2wb_20_port, W_i(19) => W2wb_19_port, W_i(18) => 
                           W2wb_18_port, W_i(17) => W2wb_17_port, W_i(16) => 
                           W2wb_16_port, W_i(15) => W2wb_15_port, W_i(14) => 
                           W2wb_14_port, W_i(13) => W2wb_13_port, W_i(12) => 
                           W2wb_12_port, W_i(11) => W2wb_11_port, W_i(10) => 
                           W2wb_10_port, W_i(9) => W2wb_9_port, W_i(8) => 
                           W2wb_8_port, W_i(7) => W2wb_7_port, W_i(6) => 
                           W2wb_6_port, W_i(5) => W2wb_5_port, W_i(4) => 
                           W2wb_4_port, W_i(3) => W2wb_3_port, W_i(2) => 
                           W2wb_2_port, W_i(1) => W2wb_1_port, W_i(0) => 
                           W2wb_0_port, D3_i(4) => n10, D3_i(3) => n12, D3_i(2)
                           => n9, D3_i(1) => n13, D3_i(0) => n11, W_o(31) => 
                           wb2reg_31_port, W_o(30) => wb2reg_30_port, W_o(29) 
                           => wb2reg_29_port, W_o(28) => wb2reg_28_port, 
                           W_o(27) => wb2reg_27_port, W_o(26) => wb2reg_26_port
                           , W_o(25) => wb2reg_25_port, W_o(24) => 
                           wb2reg_24_port, W_o(23) => wb2reg_23_port, W_o(22) 
                           => wb2reg_22_port, W_o(21) => wb2reg_21_port, 
                           W_o(20) => wb2reg_20_port, W_o(19) => wb2reg_19_port
                           , W_o(18) => wb2reg_18_port, W_o(17) => 
                           wb2reg_17_port, W_o(16) => wb2reg_16_port, W_o(15) 
                           => wb2reg_15_port, W_o(14) => wb2reg_14_port, 
                           W_o(13) => wb2reg_13_port, W_o(12) => wb2reg_12_port
                           , W_o(11) => wb2reg_11_port, W_o(10) => 
                           wb2reg_10_port, W_o(9) => wb2reg_9_port, W_o(8) => 
                           wb2reg_8_port, W_o(7) => wb2reg_7_port, W_o(6) => 
                           wb2reg_6_port, W_o(5) => wb2reg_5_port, W_o(4) => 
                           wb2reg_4_port, W_o(3) => wb2reg_3_port, W_o(2) => 
                           wb2reg_2_port, W_o(1) => wb2reg_1_port, W_o(0) => 
                           wb2reg_0_port, D3_o(4) => D32reg_4_port, D3_o(3) => 
                           D32reg_3_port, D3_o(2) => D32reg_2_port, D3_o(1) => 
                           D32reg_1_port, D3_o(0) => D32reg_0_port, clk => 
                           clock, rst => rst);
   UMEM_BLOCK : mem_block port map( X_i(31) => DRAM_Addr_o_31_port, X_i(30) => 
                           DRAM_Addr_o_30_port, X_i(29) => DRAM_Addr_o_29_port,
                           X_i(28) => DRAM_Addr_o_28_port, X_i(27) => 
                           DRAM_Addr_o_27_port, X_i(26) => DRAM_Addr_o_26_port,
                           X_i(25) => DRAM_Addr_o_25_port, X_i(24) => 
                           DRAM_Addr_o_24_port, X_i(23) => DRAM_Addr_o_23_port,
                           X_i(22) => DRAM_Addr_o_22_port, X_i(21) => 
                           DRAM_Addr_o_21_port, X_i(20) => DRAM_Addr_o_20_port,
                           X_i(19) => DRAM_Addr_o_19_port, X_i(18) => 
                           DRAM_Addr_o_18_port, X_i(17) => DRAM_Addr_o_17_port,
                           X_i(16) => DRAM_Addr_o_16_port, X_i(15) => 
                           DRAM_Addr_o_15_port, X_i(14) => DRAM_Addr_o_14_port,
                           X_i(13) => DRAM_Addr_o_13_port, X_i(12) => 
                           DRAM_Addr_o_12_port, X_i(11) => DRAM_Addr_o_11_port,
                           X_i(10) => DRAM_Addr_o_10_port, X_i(9) => 
                           DRAM_Addr_o_9_port, X_i(8) => DRAM_Addr_o_8_port, 
                           X_i(7) => DRAM_Addr_o_7_port, X_i(6) => 
                           DRAM_Addr_o_6_port, X_i(5) => DRAM_Addr_o_5_port, 
                           X_i(4) => DRAM_Addr_o_4_port, X_i(3) => 
                           DRAM_Addr_o_3_port, X_i(2) => DRAM_Addr_o_2_port, 
                           X_i(1) => DRAM_Addr_o_1_port, X_i(0) => 
                           DRAM_Addr_o_0_port, LOAD_i(31) => DRAM_Dout_i(31), 
                           LOAD_i(30) => DRAM_Dout_i(30), LOAD_i(29) => 
                           DRAM_Dout_i(29), LOAD_i(28) => DRAM_Dout_i(28), 
                           LOAD_i(27) => DRAM_Dout_i(27), LOAD_i(26) => 
                           DRAM_Dout_i(26), LOAD_i(25) => DRAM_Dout_i(25), 
                           LOAD_i(24) => DRAM_Dout_i(24), LOAD_i(23) => 
                           DRAM_Dout_i(23), LOAD_i(22) => DRAM_Dout_i(22), 
                           LOAD_i(21) => DRAM_Dout_i(21), LOAD_i(20) => 
                           DRAM_Dout_i(20), LOAD_i(19) => DRAM_Dout_i(19), 
                           LOAD_i(18) => DRAM_Dout_i(18), LOAD_i(17) => 
                           DRAM_Dout_i(17), LOAD_i(16) => DRAM_Dout_i(16), 
                           LOAD_i(15) => DRAM_Dout_i(15), LOAD_i(14) => 
                           DRAM_Dout_i(14), LOAD_i(13) => DRAM_Dout_i(13), 
                           LOAD_i(12) => DRAM_Dout_i(12), LOAD_i(11) => 
                           DRAM_Dout_i(11), LOAD_i(10) => DRAM_Dout_i(10), 
                           LOAD_i(9) => DRAM_Dout_i(9), LOAD_i(8) => 
                           DRAM_Dout_i(8), LOAD_i(7) => DRAM_Dout_i(7), 
                           LOAD_i(6) => DRAM_Dout_i(6), LOAD_i(5) => 
                           DRAM_Dout_i(5), LOAD_i(4) => DRAM_Dout_i(4), 
                           LOAD_i(3) => DRAM_Dout_i(3), LOAD_i(2) => 
                           DRAM_Dout_i(2), LOAD_i(1) => DRAM_Dout_i(1), 
                           LOAD_i(0) => DRAM_Dout_i(0), W_o(31) => W2wb_31_port
                           , W_o(30) => W2wb_30_port, W_o(29) => W2wb_29_port, 
                           W_o(28) => W2wb_28_port, W_o(27) => W2wb_27_port, 
                           W_o(26) => W2wb_26_port, W_o(25) => W2wb_25_port, 
                           W_o(24) => W2wb_24_port, W_o(23) => W2wb_23_port, 
                           W_o(22) => W2wb_22_port, W_o(21) => W2wb_21_port, 
                           W_o(20) => W2wb_20_port, W_o(19) => W2wb_19_port, 
                           W_o(18) => W2wb_18_port, W_o(17) => W2wb_17_port, 
                           W_o(16) => W2wb_16_port, W_o(15) => W2wb_15_port, 
                           W_o(14) => W2wb_14_port, W_o(13) => W2wb_13_port, 
                           W_o(12) => W2wb_12_port, W_o(11) => W2wb_11_port, 
                           W_o(10) => W2wb_10_port, W_o(9) => W2wb_9_port, 
                           W_o(8) => W2wb_8_port, W_o(7) => W2wb_7_port, W_o(6)
                           => W2wb_6_port, W_o(5) => W2wb_5_port, W_o(4) => 
                           W2wb_4_port, W_o(3) => W2wb_3_port, W_o(2) => 
                           W2wb_2_port, W_o(1) => W2wb_1_port, W_o(0) => 
                           W2wb_0_port, S_MUX_MEM_i_BAR => dummy_S_MUX_MEM);
   UFW_LOGIC : fw_logic port map( D1_i(4) => n30, D1_i(3) => n31, D1_i(2) => 
                           n32, D1_i(1) => n33, D1_i(0) => n34, rAdec_i(4) => 
                           IR_25_port, rAdec_i(3) => IR_24_port, rAdec_i(2) => 
                           IR_23_port, rAdec_i(1) => IR_22_port, rAdec_i(0) => 
                           IR_21_port, D2_i(4) => D22D3_4_port, D2_i(3) => 
                           D22D3_3_port, D2_i(2) => n8, D2_i(1) => D22D3_1_port
                           , D2_i(0) => D22D3_0_port, D3_i(4) => D32reg_4_port,
                           D3_i(3) => D32reg_3_port, D3_i(2) => D32reg_2_port, 
                           D3_i(1) => D32reg_1_port, D3_i(0) => D32reg_0_port, 
                           rA_i(4) => rA2fw_4_port, rA_i(3) => rA2fw_3_port, 
                           rA_i(2) => rA2fw_2_port, rA_i(1) => rA2fw_1_port, 
                           rA_i(0) => rA2fw_0_port, rB_i(4) => rB2mux_4_port, 
                           rB_i(3) => rB2mux_3_port, rB_i(2) => rB2mux_2_port, 
                           rB_i(1) => rB2mux_1_port, rB_i(0) => rB2mux_0_port, 
                           S_mem_W => dummy_S_RF_W_mem, S_wb_W => 
                           dummy_S_RF_W_wb, S_exe_W => n35, S_FWAdec(1) => 
                           dummy_S_FWAdec_1_port, S_FWAdec(0) => 
                           dummy_S_FWAdec_0_port, S_FWA(1) => 
                           dummy_S_FWA2exe_1_port, S_FWA(0) => 
                           dummy_S_FWA2exe_0_port, S_FWB(1) => 
                           dummy_S_FWB2exe_1_port, S_FWB(0) => 
                           dummy_S_FWB2exe_0_port, S_mem_LOAD_BAR => 
                           dummy_S_MUX_MEM);
   U5 : INV_X1 port map( A => stall_decode, ZN => enable_regfile);
   U6 : CLKBUF_X1 port map( A => mispredict, Z => n4);
   U7 : CLKBUF_X1 port map( A => D22D3_1_port, Z => n13);
   U8 : BUF_X1 port map( A => D22D3_4_port, Z => n10);
   U9 : BUF_X1 port map( A => n8, Z => n9);
   U10 : BUF_X1 port map( A => D22D3_0_port, Z => n11);
   U11 : BUF_X1 port map( A => D22D3_3_port, Z => n12);
   U12 : INV_X2 port map( A => n3, ZN => was_taken);
   U13 : AOI21_X1 port map( B1 => was_taken_from_jl, B2 => was_branch, A => 
                           was_jmp, ZN => n3);
   n14 <= '0';
   n15 <= '0';
   n16 <= '0';
   n17 <= '0';
   n18 <= '0';
   n19 <= '0';
   n20 <= '0';
   n21 <= '0';
   n22 <= '0';
   n23 <= '0';
   n24 <= '0';
   n25 <= '0';
   n26 <= '0';
   n27 <= '0';
   n28 <= '0';
   n29 <= '0';
   n30 <= '0';
   n31 <= '0';
   n32 <= '0';
   n33 <= '0';
   n34 <= '0';
   n35 <= '0';

end SYN_arch;
