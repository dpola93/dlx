
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_top_level is

-- define attributes
attribute ENUM_ENCODING : STRING;

-- define any necessary types
type aluOp is (NOP, SLLS, SRLS, SRAS, ADDS, ADDUS, SUBS, SUBUS, ANDS, ORS, 
   XORS, SEQS, SNES, SLTS, SGTS, SLES, SGES, MOVI2SS, MOVS2IS, MOVFS, MOVDS, 
   MOVFP2IS, MOVI2FP, MOVI2TS, MOVT2IS, SLTUS, SGTUS, SLEUS, SGEUS, MULTU, 
   MULTS);
attribute ENUM_ENCODING of aluOp : type is 
   "00000 00001 00010 00011 00100 00101 00110 00111 01000 01001 01010 01011 01100 01101 01110 01111 10000 10001 10010 10011 10100 10101 10110 10111 11000 11001 11010 11011 11100 11101 11110";
type UNSIGNED is array (INTEGER range <>) of std_logic;
   
   -- Declarations for conversion functions.
   function std_logic_vector_to_aluOp(arg : in std_logic_vector( 1 to 5 )) 
               return aluOp;
   function aluOp_to_std_logic_vector(arg : in aluOp) return std_logic_vector;

end CONV_PACK_top_level;

package body CONV_PACK_top_level is
   
   -- std_logic_vector to enum type function
   function std_logic_vector_to_aluOp(arg : in std_logic_vector( 1 to 5 )) 
   return aluOp is
   -- synopsys built_in SYN_FEED_THRU;
   begin
      case arg is
         when "00000" => return NOP;
         when "00001" => return SLLS;
         when "00010" => return SRLS;
         when "00011" => return SRAS;
         when "00100" => return ADDS;
         when "00101" => return ADDUS;
         when "00110" => return SUBS;
         when "00111" => return SUBUS;
         when "01000" => return ANDS;
         when "01001" => return ORS;
         when "01010" => return XORS;
         when "01011" => return SEQS;
         when "01100" => return SNES;
         when "01101" => return SLTS;
         when "01110" => return SGTS;
         when "01111" => return SLES;
         when "10000" => return SGES;
         when "10001" => return MOVI2SS;
         when "10010" => return MOVS2IS;
         when "10011" => return MOVFS;
         when "10100" => return MOVDS;
         when "10101" => return MOVFP2IS;
         when "10110" => return MOVI2FP;
         when "10111" => return MOVI2TS;
         when "11000" => return MOVT2IS;
         when "11001" => return SLTUS;
         when "11010" => return SGTUS;
         when "11011" => return SLEUS;
         when "11100" => return SGEUS;
         when "11101" => return MULTU;
         when "11110" => return MULTS;
         when others => assert FALSE -- this should not happen.
               report "un-convertible value"
               severity warning;
               return NOP;
      end case;
   end;
   
   -- enum type to std_logic_vector function
   function aluOp_to_std_logic_vector(arg : in aluOp) return std_logic_vector 
   is
   -- synopsys built_in SYN_FEED_THRU;
   begin
      case arg is
         when NOP => return "00000";
         when SLLS => return "00001";
         when SRLS => return "00010";
         when SRAS => return "00011";
         when ADDS => return "00100";
         when ADDUS => return "00101";
         when SUBS => return "00110";
         when SUBUS => return "00111";
         when ANDS => return "01000";
         when ORS => return "01001";
         when XORS => return "01010";
         when SEQS => return "01011";
         when SNES => return "01100";
         when SLTS => return "01101";
         when SGTS => return "01110";
         when SLES => return "01111";
         when SGES => return "10000";
         when MOVI2SS => return "10001";
         when MOVS2IS => return "10010";
         when MOVFS => return "10011";
         when MOVDS => return "10100";
         when MOVFP2IS => return "10101";
         when MOVI2FP => return "10110";
         when MOVI2TS => return "10111";
         when MOVT2IS => return "11000";
         when SLTUS => return "11001";
         when SGTUS => return "11010";
         when SLEUS => return "11011";
         when SGEUS => return "11100";
         when MULTU => return "11101";
         when MULTS => return "11110";
         when others => assert FALSE -- this should not happen.
               report "un-convertible value"
               severity warning;
               return "00000";
      end case;
   end;

end CONV_PACK_top_level;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_16 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_16;

architecture SYN_USE_DEFA_ARCH_NAME of 
   SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_16 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net199627 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net199627);
   main_gate : AND2_X1 port map( A1 => net199627, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_15 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_15;

architecture SYN_USE_DEFA_ARCH_NAME of 
   SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_15 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net199627 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net199627);
   main_gate : AND2_X1 port map( A1 => net199627, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_14 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_14;

architecture SYN_USE_DEFA_ARCH_NAME of 
   SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_14 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net199627 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net199627);
   main_gate : AND2_X1 port map( A1 => net199627, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_13 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_13;

architecture SYN_USE_DEFA_ARCH_NAME of 
   SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_13 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net199627 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net199627);
   main_gate : AND2_X1 port map( A1 => net199627, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_12 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_12;

architecture SYN_USE_DEFA_ARCH_NAME of 
   SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_12 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net199627 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net199627);
   main_gate : AND2_X1 port map( A1 => net199627, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_11 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_11;

architecture SYN_USE_DEFA_ARCH_NAME of 
   SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_11 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net199627 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net199627);
   main_gate : AND2_X1 port map( A1 => net199627, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_10 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_10;

architecture SYN_USE_DEFA_ARCH_NAME of 
   SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_10 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net199627 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net199627);
   main_gate : AND2_X1 port map( A1 => net199627, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_9 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_9;

architecture SYN_USE_DEFA_ARCH_NAME of 
   SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_9 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net199627 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net199627);
   main_gate : AND2_X1 port map( A1 => net199627, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_8 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_8;

architecture SYN_USE_DEFA_ARCH_NAME of 
   SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_8 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net199627 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net199627);
   main_gate : AND2_X1 port map( A1 => net199627, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_7 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_7;

architecture SYN_USE_DEFA_ARCH_NAME of 
   SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_7 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net199627 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net199627);
   main_gate : AND2_X1 port map( A1 => net199627, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_6 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_6;

architecture SYN_USE_DEFA_ARCH_NAME of 
   SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_6 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net199627 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net199627);
   main_gate : AND2_X1 port map( A1 => net199627, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_5 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_5;

architecture SYN_USE_DEFA_ARCH_NAME of 
   SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_5 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net199627 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net199627);
   main_gate : AND2_X1 port map( A1 => net199627, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_4 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_4;

architecture SYN_USE_DEFA_ARCH_NAME of 
   SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_4 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net199627 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net199627);
   main_gate : AND2_X1 port map( A1 => net199627, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_3 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_3;

architecture SYN_USE_DEFA_ARCH_NAME of 
   SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_3 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net199627 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net199627);
   main_gate : AND2_X1 port map( A1 => net199627, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_2 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_2;

architecture SYN_USE_DEFA_ARCH_NAME of 
   SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_2 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net199627 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net199627);
   main_gate : AND2_X1 port map( A1 => net199627, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_1 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_1;

architecture SYN_USE_DEFA_ARCH_NAME of 
   SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_1 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net199627 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net199627);
   main_gate : AND2_X1 port map( A1 => net199627, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_ff32_en_1 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_ff32_en_1;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_ff32_en_1 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net199612 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net199612);
   main_gate : AND2_X1 port map( A1 => net199612, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_dlx_regfile_33 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_dlx_regfile_33;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_dlx_regfile_33 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net199397 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net199397);
   main_gate : AND2_X1 port map( A1 => net199397, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_dlx_regfile_32 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_dlx_regfile_32;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_dlx_regfile_32 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net199397 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net199397);
   main_gate : AND2_X1 port map( A1 => net199397, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_dlx_regfile_31 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_dlx_regfile_31;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_dlx_regfile_31 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net199397 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net199397);
   main_gate : AND2_X1 port map( A1 => net199397, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_dlx_regfile_30 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_dlx_regfile_30;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_dlx_regfile_30 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net199397 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net199397);
   main_gate : AND2_X1 port map( A1 => net199397, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_dlx_regfile_29 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_dlx_regfile_29;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_dlx_regfile_29 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net199397 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net199397);
   main_gate : AND2_X1 port map( A1 => net199397, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_dlx_regfile_28 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_dlx_regfile_28;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_dlx_regfile_28 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net199397 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net199397);
   main_gate : AND2_X1 port map( A1 => net199397, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_dlx_regfile_27 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_dlx_regfile_27;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_dlx_regfile_27 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net199397 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net199397);
   main_gate : AND2_X1 port map( A1 => net199397, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_dlx_regfile_26 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_dlx_regfile_26;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_dlx_regfile_26 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net199397 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net199397);
   main_gate : AND2_X1 port map( A1 => net199397, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_dlx_regfile_25 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_dlx_regfile_25;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_dlx_regfile_25 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net199397 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net199397);
   main_gate : AND2_X1 port map( A1 => net199397, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_dlx_regfile_24 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_dlx_regfile_24;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_dlx_regfile_24 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net199397 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net199397);
   main_gate : AND2_X1 port map( A1 => net199397, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_dlx_regfile_23 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_dlx_regfile_23;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_dlx_regfile_23 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net199397 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net199397);
   main_gate : AND2_X1 port map( A1 => net199397, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_dlx_regfile_22 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_dlx_regfile_22;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_dlx_regfile_22 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net199397 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net199397);
   main_gate : AND2_X1 port map( A1 => net199397, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_dlx_regfile_21 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_dlx_regfile_21;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_dlx_regfile_21 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net199397 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net199397);
   main_gate : AND2_X1 port map( A1 => net199397, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_dlx_regfile_20 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_dlx_regfile_20;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_dlx_regfile_20 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net199397 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net199397);
   main_gate : AND2_X1 port map( A1 => net199397, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_dlx_regfile_19 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_dlx_regfile_19;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_dlx_regfile_19 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net199397 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net199397);
   main_gate : AND2_X1 port map( A1 => net199397, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_dlx_regfile_18 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_dlx_regfile_18;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_dlx_regfile_18 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net199397 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net199397);
   main_gate : AND2_X1 port map( A1 => net199397, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_dlx_regfile_17 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_dlx_regfile_17;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_dlx_regfile_17 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net199397 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net199397);
   main_gate : AND2_X1 port map( A1 => net199397, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_dlx_regfile_16 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_dlx_regfile_16;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_dlx_regfile_16 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net199397 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net199397);
   main_gate : AND2_X1 port map( A1 => net199397, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_dlx_regfile_15 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_dlx_regfile_15;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_dlx_regfile_15 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net199397 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net199397);
   main_gate : AND2_X1 port map( A1 => net199397, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_dlx_regfile_14 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_dlx_regfile_14;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_dlx_regfile_14 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net199397 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net199397);
   main_gate : AND2_X1 port map( A1 => net199397, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_dlx_regfile_13 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_dlx_regfile_13;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_dlx_regfile_13 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net199397 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net199397);
   main_gate : AND2_X1 port map( A1 => net199397, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_dlx_regfile_12 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_dlx_regfile_12;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_dlx_regfile_12 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net199397 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net199397);
   main_gate : AND2_X1 port map( A1 => net199397, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_dlx_regfile_11 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_dlx_regfile_11;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_dlx_regfile_11 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net199397 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net199397);
   main_gate : AND2_X1 port map( A1 => net199397, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_dlx_regfile_10 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_dlx_regfile_10;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_dlx_regfile_10 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net199397 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net199397);
   main_gate : AND2_X1 port map( A1 => net199397, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_dlx_regfile_9 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_dlx_regfile_9;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_dlx_regfile_9 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net199397 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net199397);
   main_gate : AND2_X1 port map( A1 => net199397, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_dlx_regfile_8 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_dlx_regfile_8;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_dlx_regfile_8 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net199397 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net199397);
   main_gate : AND2_X1 port map( A1 => net199397, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_dlx_regfile_7 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_dlx_regfile_7;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_dlx_regfile_7 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net199397 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net199397);
   main_gate : AND2_X1 port map( A1 => net199397, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_dlx_regfile_6 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_dlx_regfile_6;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_dlx_regfile_6 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net199397 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net199397);
   main_gate : AND2_X1 port map( A1 => net199397, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_dlx_regfile_5 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_dlx_regfile_5;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_dlx_regfile_5 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net199397 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net199397);
   main_gate : AND2_X1 port map( A1 => net199397, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_dlx_regfile_4 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_dlx_regfile_4;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_dlx_regfile_4 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net199397 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net199397);
   main_gate : AND2_X1 port map( A1 => net199397, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_dlx_regfile_3 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_dlx_regfile_3;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_dlx_regfile_3 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net199397 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net199397);
   main_gate : AND2_X1 port map( A1 => net199397, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_dlx_regfile_2 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_dlx_regfile_2;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_dlx_regfile_2 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net199397 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net199397);
   main_gate : AND2_X1 port map( A1 => net199397, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_dlx_regfile_1 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_dlx_regfile_1;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_dlx_regfile_1 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net199397 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net199397);
   main_gate : AND2_X1 port map( A1 => net199397, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_ff32_en_SIZE5_3 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_ff32_en_SIZE5_3;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_ff32_en_SIZE5_3 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net199367 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net199367);
   main_gate : AND2_X1 port map( A1 => net199367, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_ff32_en_SIZE5_2 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_ff32_en_SIZE5_2;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_ff32_en_SIZE5_2 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net199367 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net199367);
   main_gate : AND2_X1 port map( A1 => net199367, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_ff32_en_SIZE32_5 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_ff32_en_SIZE32_5;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_ff32_en_SIZE32_5 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net199352 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net199352);
   main_gate : AND2_X1 port map( A1 => net199352, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_ff32_en_SIZE32_4 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_ff32_en_SIZE32_4;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_ff32_en_SIZE32_4 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net199352 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net199352);
   main_gate : AND2_X1 port map( A1 => net199352, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_ff32_en_SIZE32_1 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_ff32_en_SIZE32_1;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_ff32_en_SIZE32_1 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net199352 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net199352);
   main_gate : AND2_X1 port map( A1 => net199352, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_127 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_127;

architecture SYN_BEHAVIORAL of FA_127 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U5 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => B, A2 => Ci, ZN => n4);
   U3 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U1 : XNOR2_X1 port map( A => n6, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_126 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_126;

architecture SYN_BEHAVIORAL of FA_126 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U5 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => B, A2 => Ci, ZN => n4);
   U3 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U1 : XNOR2_X1 port map( A => n6, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_125 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_125;

architecture SYN_BEHAVIORAL of FA_125 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n2);
   U1 : XNOR2_X1 port map( A => n2, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_120 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_120;

architecture SYN_BEHAVIORAL of FA_120 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => S);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_119 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_119;

architecture SYN_BEHAVIORAL of FA_119 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U1 : XNOR2_X1 port map( A => n6, B => B, ZN => S);
   U5 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => B, A2 => Ci, ZN => n4);
   U3 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_118 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_118;

architecture SYN_BEHAVIORAL of FA_118 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U1 : XNOR2_X1 port map( A => n6, B => B, ZN => S);
   U5 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => B, A2 => Ci, ZN => n4);
   U3 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_117 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_117;

architecture SYN_BEHAVIORAL of FA_117 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n2);
   U1 : XNOR2_X1 port map( A => n2, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_116 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_116;

architecture SYN_BEHAVIORAL of FA_116 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => A, A2 => B, ZN => Co);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_115 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_115;

architecture SYN_BEHAVIORAL of FA_115 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U1 : XNOR2_X1 port map( A => n6, B => B, ZN => S);
   U5 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => B, A2 => Ci, ZN => n4);
   U3 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_114 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_114;

architecture SYN_BEHAVIORAL of FA_114 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U1 : XNOR2_X1 port map( A => n6, B => B, ZN => S);
   U5 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => B, A2 => Ci, ZN => n4);
   U3 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_113 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_113;

architecture SYN_BEHAVIORAL of FA_113 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n2);
   U1 : XNOR2_X1 port map( A => n2, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_112 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_112;

architecture SYN_BEHAVIORAL of FA_112 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => S);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_111 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_111;

architecture SYN_BEHAVIORAL of FA_111 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U1 : XNOR2_X1 port map( A => n6, B => B, ZN => S);
   U5 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => B, A2 => Ci, ZN => n4);
   U3 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_110 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_110;

architecture SYN_BEHAVIORAL of FA_110 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U1 : XNOR2_X1 port map( A => n6, B => B, ZN => S);
   U5 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => B, A2 => Ci, ZN => n4);
   U3 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_109 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_109;

architecture SYN_BEHAVIORAL of FA_109 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n2);
   U1 : XNOR2_X1 port map( A => n2, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_108 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_108;

architecture SYN_BEHAVIORAL of FA_108 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => A, A2 => B, ZN => Co);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_107 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_107;

architecture SYN_BEHAVIORAL of FA_107 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U1 : XNOR2_X1 port map( A => n6, B => B, ZN => S);
   U5 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => B, A2 => Ci, ZN => n4);
   U3 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_106 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_106;

architecture SYN_BEHAVIORAL of FA_106 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U1 : XNOR2_X1 port map( A => n6, B => B, ZN => S);
   U5 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => B, A2 => Ci, ZN => n4);
   U3 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_105 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_105;

architecture SYN_BEHAVIORAL of FA_105 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n2);
   U1 : XNOR2_X1 port map( A => n2, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_104 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_104;

architecture SYN_BEHAVIORAL of FA_104 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => S);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_103 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_103;

architecture SYN_BEHAVIORAL of FA_103 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U5 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => B, A2 => Ci, ZN => n4);
   U3 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U1 : XNOR2_X1 port map( A => n6, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_102 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_102;

architecture SYN_BEHAVIORAL of FA_102 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U1 : XNOR2_X1 port map( A => n6, B => B, ZN => S);
   U5 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => B, A2 => Ci, ZN => n4);
   U3 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_101 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_101;

architecture SYN_BEHAVIORAL of FA_101 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n2);
   U1 : XNOR2_X1 port map( A => n2, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_100 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_100;

architecture SYN_BEHAVIORAL of FA_100 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => A, A2 => B, ZN => Co);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_99 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_99;

architecture SYN_BEHAVIORAL of FA_99 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U5 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => B, A2 => Ci, ZN => n4);
   U3 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U1 : XNOR2_X1 port map( A => n6, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_98 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_98;

architecture SYN_BEHAVIORAL of FA_98 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U1 : XNOR2_X1 port map( A => n6, B => B, ZN => S);
   U5 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => B, A2 => Ci, ZN => n4);
   U3 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_97 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_97;

architecture SYN_BEHAVIORAL of FA_97 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n2);
   U1 : XNOR2_X1 port map( A => n2, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_96 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_96;

architecture SYN_BEHAVIORAL of FA_96 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => S);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_95 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_95;

architecture SYN_BEHAVIORAL of FA_95 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n5);
   U1 : XNOR2_X1 port map( A => n5, B => B, ZN => S);
   U3 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n3);
   U4 : NAND2_X1 port map( A1 => n3, A2 => n4, ZN => Co);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => B, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_94 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_94;

architecture SYN_BEHAVIORAL of FA_94 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n4 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n4);
   U1 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n2);
   U3 : NAND2_X1 port map( A1 => n2, A2 => n3, ZN => Co);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => B, ZN => n3);
   U5 : XNOR2_X1 port map( A => n4, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_93 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_93;

architecture SYN_BEHAVIORAL of FA_93 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal net246211 : std_logic;

begin
   
   U1 : FA_X1 port map( A => B, B => A, CI => Ci, CO => net246211, S => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_92 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_92;

architecture SYN_BEHAVIORAL of FA_92 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => S);
   U2 : OR2_X1 port map( A1 => B, A2 => A, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_91 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_91;

architecture SYN_BEHAVIORAL of FA_91 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n5);
   U1 : XNOR2_X1 port map( A => n5, B => B, ZN => S);
   U3 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n3);
   U4 : NAND2_X1 port map( A1 => n3, A2 => n4, ZN => Co);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => B, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_90 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_90;

architecture SYN_BEHAVIORAL of FA_90 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n4 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n4);
   U1 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n2);
   U3 : NAND2_X1 port map( A1 => n2, A2 => n3, ZN => Co);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => B, ZN => n3);
   U5 : XNOR2_X1 port map( A => n4, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_89 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_89;

architecture SYN_BEHAVIORAL of FA_89 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal net246210 : std_logic;

begin
   
   U1 : FA_X1 port map( A => B, B => A, CI => Ci, CO => net246210, S => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_88 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_88;

architecture SYN_BEHAVIORAL of FA_88 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n2, B => B, ZN => S);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => Co);
   U3 : INV_X1 port map( A => A, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_87 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_87;

architecture SYN_BEHAVIORAL of FA_87 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n4 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n4);
   U1 : XNOR2_X1 port map( A => n4, B => B, ZN => S);
   U3 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n2);
   U4 : NAND2_X1 port map( A1 => n2, A2 => n3, ZN => Co);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => B, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_86 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_86;

architecture SYN_BEHAVIORAL of FA_86 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n4 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n4);
   U1 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n2);
   U3 : NAND2_X1 port map( A1 => n2, A2 => n3, ZN => Co);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => B, ZN => n3);
   U5 : XNOR2_X1 port map( A => n4, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_85 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_85;

architecture SYN_BEHAVIORAL of FA_85 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => Ci, ZN => n2);
   U2 : XNOR2_X1 port map( A => n2, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_84 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_84;

architecture SYN_BEHAVIORAL of FA_84 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => S);
   U2 : OR2_X1 port map( A1 => B, A2 => A, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_83 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_83;

architecture SYN_BEHAVIORAL of FA_83 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n4 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n4);
   U1 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n2);
   U3 : NAND2_X1 port map( A1 => n2, A2 => n3, ZN => Co);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => B, ZN => n3);
   U5 : XNOR2_X1 port map( A => n4, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_82 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_82;

architecture SYN_BEHAVIORAL of FA_82 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n4 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n4);
   U1 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n2);
   U3 : NAND2_X1 port map( A1 => n2, A2 => n3, ZN => Co);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => B, ZN => n3);
   U5 : XNOR2_X1 port map( A => n4, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_81 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_81;

architecture SYN_BEHAVIORAL of FA_81 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal net246209 : std_logic;

begin
   
   U1 : FA_X1 port map( A => B, B => A, CI => Ci, CO => net246209, S => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_80 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_80;

architecture SYN_BEHAVIORAL of FA_80 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => S);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_79 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_79;

architecture SYN_BEHAVIORAL of FA_79 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n6, n7 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n7);
   U1 : XNOR2_X1 port map( A => n7, B => B, ZN => S);
   U3 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => Co);
   U4 : NAND2_X1 port map( A1 => B, A2 => Ci, ZN => n5);
   U5 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_78 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_78;

architecture SYN_BEHAVIORAL of FA_78 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n6, B => B, ZN => S);
   U3 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U4 : NAND2_X1 port map( A1 => B, A2 => Ci, ZN => n4);
   U5 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_77 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_77;

architecture SYN_BEHAVIORAL of FA_77 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal net246208 : std_logic;

begin
   
   U1 : FA_X1 port map( A => B, B => A, CI => Ci, CO => net246208, S => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_76 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_76;

architecture SYN_BEHAVIORAL of FA_76 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => A, A2 => B, ZN => Co);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_75 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_75;

architecture SYN_BEHAVIORAL of FA_75 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n6, n7 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n7, B => B, ZN => S);
   U3 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => Co);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n7);
   U4 : NAND2_X1 port map( A1 => B, A2 => Ci, ZN => n5);
   U5 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_74 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_74;

architecture SYN_BEHAVIORAL of FA_74 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n6, B => B, ZN => S);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U3 : NAND2_X1 port map( A1 => B, A2 => Ci, ZN => n4);
   U4 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n5);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_73 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_73;

architecture SYN_BEHAVIORAL of FA_73 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => Ci, ZN => n3);
   U2 : XNOR2_X1 port map( A => n3, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_72 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_72;

architecture SYN_BEHAVIORAL of FA_72 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Co);
   U2 : INV_X1 port map( A => A, ZN => n3);
   U3 : XNOR2_X1 port map( A => n3, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_71 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_71;

architecture SYN_BEHAVIORAL of FA_71 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n6, n7 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n7);
   U5 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n6);
   U4 : NAND2_X1 port map( A1 => B, A2 => Ci, ZN => n5);
   U3 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => Co);
   U1 : XNOR2_X1 port map( A => n7, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_70 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_70;

architecture SYN_BEHAVIORAL of FA_70 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n4 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n4);
   U1 : XNOR2_X1 port map( A => n4, B => B, ZN => S);
   U3 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n2);
   U4 : NAND2_X1 port map( A1 => n2, A2 => n3, ZN => Co);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => B, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_69 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_69;

architecture SYN_BEHAVIORAL of FA_69 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal net246207 : std_logic;

begin
   
   U1 : FA_X1 port map( A => B, B => A, CI => Ci, CO => net246207, S => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_68 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_68;

architecture SYN_BEHAVIORAL of FA_68 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => S);
   U2 : OR2_X1 port map( A1 => B, A2 => A, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_67 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_67;

architecture SYN_BEHAVIORAL of FA_67 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n5);
   U1 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n3);
   U3 : NAND2_X1 port map( A1 => n3, A2 => n4, ZN => Co);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => B, ZN => n4);
   U5 : XNOR2_X1 port map( A => n5, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_66 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_66;

architecture SYN_BEHAVIORAL of FA_66 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n4 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n4);
   U1 : XNOR2_X1 port map( A => n4, B => B, ZN => S);
   U3 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n2);
   U4 : NAND2_X1 port map( A1 => n2, A2 => n3, ZN => Co);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => B, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_65 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_65;

architecture SYN_BEHAVIORAL of FA_65 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n2);
   U1 : XNOR2_X1 port map( A => n2, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_64 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_64;

architecture SYN_BEHAVIORAL of FA_64 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n3);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => Co);
   U3 : XNOR2_X1 port map( A => n3, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_63 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_63;

architecture SYN_BEHAVIORAL of FA_63 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n6, n7 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n7);
   U3 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => Co);
   U1 : XNOR2_X1 port map( A => n7, B => B, ZN => S);
   U4 : NAND2_X1 port map( A1 => B, A2 => Ci, ZN => n5);
   U5 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_62 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_62;

architecture SYN_BEHAVIORAL of FA_62 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U3 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U1 : XNOR2_X1 port map( A => n6, B => B, ZN => S);
   U4 : NAND2_X1 port map( A1 => B, A2 => Ci, ZN => n4);
   U5 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_61 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_61;

architecture SYN_BEHAVIORAL of FA_61 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n2);
   U1 : XNOR2_X1 port map( A => n2, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_60 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_60;

architecture SYN_BEHAVIORAL of FA_60 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => A, A2 => B, ZN => Co);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_59 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_59;

architecture SYN_BEHAVIORAL of FA_59 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n6, n7 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n7);
   U3 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => Co);
   U1 : XNOR2_X1 port map( A => n7, B => B, ZN => S);
   U4 : NAND2_X1 port map( A1 => B, A2 => Ci, ZN => n5);
   U5 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_58 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_58;

architecture SYN_BEHAVIORAL of FA_58 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U3 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U1 : XNOR2_X1 port map( A => n6, B => B, ZN => S);
   U4 : NAND2_X1 port map( A1 => B, A2 => Ci, ZN => n4);
   U5 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_57 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_57;

architecture SYN_BEHAVIORAL of FA_57 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n2);
   U1 : XNOR2_X1 port map( A => n2, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_56 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_56;

architecture SYN_BEHAVIORAL of FA_56 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => S);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_55 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_55;

architecture SYN_BEHAVIORAL of FA_55 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U1 : XNOR2_X1 port map( A => n6, B => B, ZN => S);
   U4 : NAND2_X1 port map( A1 => B, A2 => Ci, ZN => n4);
   U5 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_54 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_54;

architecture SYN_BEHAVIORAL of FA_54 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U1 : XNOR2_X1 port map( A => n6, B => B, ZN => S);
   U4 : NAND2_X1 port map( A1 => B, A2 => Ci, ZN => n4);
   U5 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_53 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_53;

architecture SYN_BEHAVIORAL of FA_53 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n2);
   U1 : XNOR2_X1 port map( A => n2, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_52 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_52;

architecture SYN_BEHAVIORAL of FA_52 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => A, A2 => B, ZN => Co);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_51 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_51;

architecture SYN_BEHAVIORAL of FA_51 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U1 : XNOR2_X1 port map( A => n6, B => B, ZN => S);
   U4 : NAND2_X1 port map( A1 => B, A2 => Ci, ZN => n4);
   U5 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_50 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_50;

architecture SYN_BEHAVIORAL of FA_50 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U1 : XNOR2_X1 port map( A => n6, B => B, ZN => S);
   U4 : NAND2_X1 port map( A1 => B, A2 => Ci, ZN => n4);
   U5 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_49 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_49;

architecture SYN_BEHAVIORAL of FA_49 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n2);
   U1 : XNOR2_X1 port map( A => n2, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_48 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_48;

architecture SYN_BEHAVIORAL of FA_48 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => S);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_47 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_47;

architecture SYN_BEHAVIORAL of FA_47 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U1 : XNOR2_X1 port map( A => n6, B => B, ZN => S);
   U4 : NAND2_X1 port map( A1 => B, A2 => Ci, ZN => n4);
   U5 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_46 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_46;

architecture SYN_BEHAVIORAL of FA_46 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n3, net246206 : std_logic;

begin
   
   U5 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n3);
   U4 : NAND2_X1 port map( A1 => B, A2 => Ci, ZN => n1);
   U3 : NAND2_X1 port map( A1 => n3, A2 => n1, ZN => Co);
   U1 : FA_X1 port map( A => B, B => A, CI => Ci, CO => net246206, S => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_45 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_45;

architecture SYN_BEHAVIORAL of FA_45 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U2 : XOR2_X1 port map( A => B, B => n2, Z => n1);
   U3 : XNOR2_X1 port map( A => Ci, B => n1, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_44 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_44;

architecture SYN_BEHAVIORAL of FA_44 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => A, A2 => B, ZN => Co);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_43 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_43;

architecture SYN_BEHAVIORAL of FA_43 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U1 : XNOR2_X1 port map( A => n6, B => B, ZN => S);
   U4 : NAND2_X1 port map( A1 => B, A2 => Ci, ZN => n4);
   U5 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_42 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_42;

architecture SYN_BEHAVIORAL of FA_42 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U5 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => B, A2 => Ci, ZN => n4);
   U3 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U1 : XNOR2_X1 port map( A => n6, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_41 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_41;

architecture SYN_BEHAVIORAL of FA_41 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U2 : XOR2_X1 port map( A => B, B => n2, Z => n1);
   U3 : XNOR2_X1 port map( A => Ci, B => n1, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_40 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_40;

architecture SYN_BEHAVIORAL of FA_40 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => S);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_39 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_39;

architecture SYN_BEHAVIORAL of FA_39 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U1 : XNOR2_X1 port map( A => n6, B => B, ZN => S);
   U4 : NAND2_X1 port map( A1 => B, A2 => Ci, ZN => n4);
   U5 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_38 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_38;

architecture SYN_BEHAVIORAL of FA_38 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U1 : XNOR2_X1 port map( A => n6, B => B, ZN => S);
   U4 : NAND2_X1 port map( A1 => B, A2 => Ci, ZN => n4);
   U5 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_37 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_37;

architecture SYN_BEHAVIORAL of FA_37 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n2);
   U1 : XNOR2_X1 port map( A => n2, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_36 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_36;

architecture SYN_BEHAVIORAL of FA_36 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => S);
   U2 : OR2_X1 port map( A1 => A, A2 => B, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_35 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_35;

architecture SYN_BEHAVIORAL of FA_35 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U1 : XNOR2_X1 port map( A => n6, B => B, ZN => S);
   U4 : NAND2_X1 port map( A1 => B, A2 => Ci, ZN => n4);
   U5 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_34 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_34;

architecture SYN_BEHAVIORAL of FA_34 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U1 : XNOR2_X1 port map( A => n6, B => B, ZN => S);
   U4 : NAND2_X1 port map( A1 => B, A2 => Ci, ZN => n4);
   U5 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_33 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_33;

architecture SYN_BEHAVIORAL of FA_33 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n2);
   U1 : XNOR2_X1 port map( A => n2, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_32 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_32;

architecture SYN_BEHAVIORAL of FA_32 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => S);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_31 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_31;

architecture SYN_BEHAVIORAL of FA_31 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U1 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U3 : XNOR2_X1 port map( A => n6, B => B, ZN => S);
   U4 : NAND2_X1 port map( A1 => B, A2 => Ci, ZN => n4);
   U5 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_30 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_30;

architecture SYN_BEHAVIORAL of FA_30 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U3 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U1 : XNOR2_X1 port map( A => n6, B => B, ZN => S);
   U4 : NAND2_X1 port map( A1 => B, A2 => Ci, ZN => n4);
   U5 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_29 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_29;

architecture SYN_BEHAVIORAL of FA_29 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n2);
   U1 : XNOR2_X1 port map( A => n2, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_28 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_28;

architecture SYN_BEHAVIORAL of FA_28 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : OR2_X1 port map( A1 => A, A2 => B, ZN => Co);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_27 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_27;

architecture SYN_BEHAVIORAL of FA_27 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U1 : XNOR2_X1 port map( A => n6, B => B, ZN => S);
   U4 : NAND2_X1 port map( A1 => B, A2 => Ci, ZN => n4);
   U5 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_26 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_26;

architecture SYN_BEHAVIORAL of FA_26 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U3 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U1 : XNOR2_X1 port map( A => n6, B => B, ZN => S);
   U4 : NAND2_X1 port map( A1 => B, A2 => Ci, ZN => n4);
   U5 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_25 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_25;

architecture SYN_BEHAVIORAL of FA_25 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n2);
   U1 : XNOR2_X1 port map( A => n2, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_24 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_24;

architecture SYN_BEHAVIORAL of FA_24 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n3, B => B, ZN => S);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => Co);
   U3 : INV_X1 port map( A => A, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_23 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_23;

architecture SYN_BEHAVIORAL of FA_23 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U1 : XNOR2_X1 port map( A => n6, B => B, ZN => S);
   U4 : NAND2_X1 port map( A1 => B, A2 => Ci, ZN => n4);
   U5 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_22 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_22;

architecture SYN_BEHAVIORAL of FA_22 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U1 : XNOR2_X1 port map( A => n6, B => B, ZN => S);
   U4 : NAND2_X1 port map( A1 => B, A2 => Ci, ZN => n4);
   U5 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_21 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_21;

architecture SYN_BEHAVIORAL of FA_21 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n2);
   U1 : XNOR2_X1 port map( A => n2, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_20 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_20;

architecture SYN_BEHAVIORAL of FA_20 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => S);
   U2 : OR2_X1 port map( A1 => A, A2 => B, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_19 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_19;

architecture SYN_BEHAVIORAL of FA_19 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U1 : XNOR2_X1 port map( A => n6, B => B, ZN => S);
   U4 : NAND2_X1 port map( A1 => B, A2 => Ci, ZN => n4);
   U5 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_18 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_18;

architecture SYN_BEHAVIORAL of FA_18 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U1 : XNOR2_X1 port map( A => n6, B => B, ZN => S);
   U4 : NAND2_X1 port map( A1 => B, A2 => Ci, ZN => n4);
   U5 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_17 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_17;

architecture SYN_BEHAVIORAL of FA_17 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n2);
   U1 : XNOR2_X1 port map( A => n2, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_16 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_16;

architecture SYN_BEHAVIORAL of FA_16 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n3, B => B, ZN => S);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => Co);
   U3 : INV_X1 port map( A => A, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_15 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_15;

architecture SYN_BEHAVIORAL of FA_15 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U1 : XNOR2_X1 port map( A => n6, B => B, ZN => S);
   U4 : NAND2_X1 port map( A1 => B, A2 => Ci, ZN => n4);
   U5 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_14 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_14;

architecture SYN_BEHAVIORAL of FA_14 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U5 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => B, A2 => Ci, ZN => n4);
   U3 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U1 : XNOR2_X1 port map( A => n6, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_13 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_13;

architecture SYN_BEHAVIORAL of FA_13 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n2);
   U1 : XNOR2_X1 port map( A => n2, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_12 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_12;

architecture SYN_BEHAVIORAL of FA_12 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => S);
   U2 : OR2_X1 port map( A1 => A, A2 => B, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_11 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_11;

architecture SYN_BEHAVIORAL of FA_11 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U3 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U1 : XNOR2_X1 port map( A => n6, B => B, ZN => S);
   U4 : NAND2_X1 port map( A1 => B, A2 => Ci, ZN => n4);
   U5 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_10 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_10;

architecture SYN_BEHAVIORAL of FA_10 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U5 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => B, A2 => Ci, ZN => n4);
   U3 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U1 : XNOR2_X1 port map( A => n6, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_9 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_9;

architecture SYN_BEHAVIORAL of FA_9 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n2);
   U1 : XNOR2_X1 port map( A => n2, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_8 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_8;

architecture SYN_BEHAVIORAL of FA_8 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n3, B => B, ZN => S);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => Co);
   U3 : INV_X1 port map( A => A, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_7 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_7;

architecture SYN_BEHAVIORAL of FA_7 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U1 : XNOR2_X1 port map( A => n6, B => B, ZN => S);
   U5 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n5);
   U3 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U4 : NAND2_X1 port map( A1 => B, A2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_6 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_6;

architecture SYN_BEHAVIORAL of FA_6 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U1 : XNOR2_X1 port map( A => n6, B => B, ZN => S);
   U5 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => B, A2 => Ci, ZN => n4);
   U3 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_5 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_5;

architecture SYN_BEHAVIORAL of FA_5 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n2, B => B, ZN => S);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_4 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_4;

architecture SYN_BEHAVIORAL of FA_4 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => S);
   U2 : OR2_X1 port map( A1 => A, A2 => B, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_3 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_3;

architecture SYN_BEHAVIORAL of FA_3 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U1 : XNOR2_X1 port map( A => n6, B => B, ZN => S);
   U5 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => B, A2 => Ci, ZN => n4);
   U3 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_2 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_2;

architecture SYN_BEHAVIORAL of FA_2 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U1 : XNOR2_X1 port map( A => n6, B => B, ZN => S);
   U5 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => B, A2 => Ci, ZN => n4);
   U3 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_1 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1;

architecture SYN_BEHAVIORAL of FA_1 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n2);
   U1 : XNOR2_X1 port map( A => n2, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity mux21_SIZE4_15 is

   port( IN0, IN1 : in std_logic_vector (3 downto 0);  CTRL : in std_logic;  
         OUT1 : out std_logic_vector (3 downto 0));

end mux21_SIZE4_15;

architecture SYN_Bhe of mux21_SIZE4_15 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => IN0(3), B => IN1(3), S => CTRL, Z => OUT1(3));
   U2 : MUX2_X1 port map( A => IN0(2), B => IN1(2), S => CTRL, Z => OUT1(2));
   U3 : MUX2_X1 port map( A => IN0(1), B => IN1(1), S => CTRL, Z => OUT1(1));
   U4 : MUX2_X1 port map( A => IN0(0), B => IN1(0), S => CTRL, Z => OUT1(0));

end SYN_Bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity mux21_SIZE4_14 is

   port( IN0, IN1 : in std_logic_vector (3 downto 0);  CTRL : in std_logic;  
         OUT1 : out std_logic_vector (3 downto 0));

end mux21_SIZE4_14;

architecture SYN_Bhe of mux21_SIZE4_14 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => IN0(3), B => IN1(3), S => CTRL, Z => OUT1(3));
   U2 : MUX2_X1 port map( A => IN0(2), B => IN1(2), S => CTRL, Z => OUT1(2));
   U3 : MUX2_X1 port map( A => IN0(1), B => IN1(1), S => CTRL, Z => OUT1(1));
   U4 : MUX2_X1 port map( A => IN0(0), B => IN1(0), S => CTRL, Z => OUT1(0));

end SYN_Bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity mux21_SIZE4_13 is

   port( IN0, IN1 : in std_logic_vector (3 downto 0);  CTRL : in std_logic;  
         OUT1 : out std_logic_vector (3 downto 0));

end mux21_SIZE4_13;

architecture SYN_Bhe of mux21_SIZE4_13 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => IN0(3), B => IN1(3), S => CTRL, Z => OUT1(3));
   U2 : MUX2_X1 port map( A => IN0(2), B => IN1(2), S => CTRL, Z => OUT1(2));
   U3 : MUX2_X1 port map( A => IN0(1), B => IN1(1), S => CTRL, Z => OUT1(1));
   U4 : MUX2_X1 port map( A => IN0(0), B => IN1(0), S => CTRL, Z => OUT1(0));

end SYN_Bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity mux21_SIZE4_12 is

   port( IN0, IN1 : in std_logic_vector (3 downto 0);  CTRL : in std_logic;  
         OUT1 : out std_logic_vector (3 downto 0));

end mux21_SIZE4_12;

architecture SYN_Bhe of mux21_SIZE4_12 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U2 : MUX2_X1 port map( A => IN0(2), B => IN1(2), S => CTRL, Z => OUT1(2));
   U3 : MUX2_X1 port map( A => IN0(1), B => IN1(1), S => CTRL, Z => OUT1(1));
   U4 : MUX2_X1 port map( A => IN0(0), B => IN1(0), S => CTRL, Z => OUT1(0));
   U1 : INV_X1 port map( A => CTRL, ZN => n3);
   U5 : NAND2_X1 port map( A1 => IN0(3), A2 => n3, ZN => n1);
   U6 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => OUT1(3));
   U7 : NAND2_X1 port map( A1 => IN1(3), A2 => CTRL, ZN => n2);

end SYN_Bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity mux21_SIZE4_11 is

   port( IN0, IN1 : in std_logic_vector (3 downto 0);  CTRL : in std_logic;  
         OUT1 : out std_logic_vector (3 downto 0));

end mux21_SIZE4_11;

architecture SYN_Bhe of mux21_SIZE4_11 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U2 : MUX2_X1 port map( A => IN0(2), B => IN1(2), S => CTRL, Z => OUT1(2));
   U4 : MUX2_X1 port map( A => IN0(0), B => IN1(0), S => CTRL, Z => OUT1(0));
   U1 : MUX2_X1 port map( A => IN0(1), B => IN1(1), S => CTRL, Z => OUT1(1));
   U3 : INV_X1 port map( A => CTRL, ZN => n3);
   U5 : NAND2_X1 port map( A1 => IN0(3), A2 => n3, ZN => n1);
   U6 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => OUT1(3));
   U7 : NAND2_X1 port map( A1 => IN1(3), A2 => CTRL, ZN => n2);

end SYN_Bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity mux21_SIZE4_10 is

   port( IN0, IN1 : in std_logic_vector (3 downto 0);  CTRL : in std_logic;  
         OUT1 : out std_logic_vector (3 downto 0));

end mux21_SIZE4_10;

architecture SYN_Bhe of mux21_SIZE4_10 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : MUX2_X1 port map( A => IN0(2), B => IN1(2), S => CTRL, Z => OUT1(2));
   U1 : MUX2_X1 port map( A => IN0(3), B => IN1(3), S => CTRL, Z => OUT1(3));
   U3 : MUX2_X1 port map( A => IN0(0), B => IN1(0), S => CTRL, Z => OUT1(0));
   U4 : MUX2_X1 port map( A => IN0(1), B => IN1(1), S => CTRL, Z => OUT1(1));

end SYN_Bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity mux21_SIZE4_9 is

   port( IN0, IN1 : in std_logic_vector (3 downto 0);  CTRL : in std_logic;  
         OUT1 : out std_logic_vector (3 downto 0));

end mux21_SIZE4_9;

architecture SYN_Bhe of mux21_SIZE4_9 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => IN0(3), B => IN1(3), S => CTRL, Z => OUT1(3));
   U2 : MUX2_X1 port map( A => IN0(2), B => IN1(2), S => CTRL, Z => OUT1(2));
   U3 : MUX2_X1 port map( A => IN0(1), B => IN1(1), S => CTRL, Z => OUT1(1));
   U4 : MUX2_X1 port map( A => IN0(0), B => IN1(0), S => CTRL, Z => OUT1(0));

end SYN_Bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity mux21_SIZE4_8 is

   port( IN0, IN1 : in std_logic_vector (3 downto 0);  CTRL : in std_logic;  
         OUT1 : out std_logic_vector (3 downto 0));

end mux21_SIZE4_8;

architecture SYN_Bhe of mux21_SIZE4_8 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => IN0(3), B => IN1(3), S => CTRL, Z => OUT1(3));
   U2 : MUX2_X1 port map( A => IN0(2), B => IN1(2), S => CTRL, Z => OUT1(2));
   U3 : MUX2_X1 port map( A => IN0(1), B => IN1(1), S => CTRL, Z => OUT1(1));
   U4 : MUX2_X1 port map( A => IN0(0), B => IN1(0), S => CTRL, Z => OUT1(0));

end SYN_Bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity mux21_SIZE4_7 is

   port( IN0, IN1 : in std_logic_vector (3 downto 0);  CTRL : in std_logic;  
         OUT1 : out std_logic_vector (3 downto 0));

end mux21_SIZE4_7;

architecture SYN_Bhe of mux21_SIZE4_7 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => IN0(3), B => IN1(3), S => CTRL, Z => OUT1(3));
   U2 : MUX2_X1 port map( A => IN0(2), B => IN1(2), S => CTRL, Z => OUT1(2));
   U3 : MUX2_X1 port map( A => IN0(1), B => IN1(1), S => CTRL, Z => OUT1(1));
   U4 : MUX2_X1 port map( A => IN0(0), B => IN1(0), S => CTRL, Z => OUT1(0));

end SYN_Bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity mux21_SIZE4_6 is

   port( IN0, IN1 : in std_logic_vector (3 downto 0);  CTRL : in std_logic;  
         OUT1 : out std_logic_vector (3 downto 0));

end mux21_SIZE4_6;

architecture SYN_Bhe of mux21_SIZE4_6 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U3 : MUX2_X1 port map( A => IN0(1), B => IN1(1), S => CTRL, Z => OUT1(1));
   U1 : MUX2_X1 port map( A => IN0(3), B => IN1(3), S => CTRL, Z => OUT1(3));
   U2 : MUX2_X1 port map( A => IN0(2), B => IN1(2), S => CTRL, Z => OUT1(2));
   U4 : MUX2_X1 port map( A => IN0(0), B => IN1(0), S => CTRL, Z => OUT1(0));

end SYN_Bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity mux21_SIZE4_5 is

   port( IN0, IN1 : in std_logic_vector (3 downto 0);  CTRL : in std_logic;  
         OUT1 : out std_logic_vector (3 downto 0));

end mux21_SIZE4_5;

architecture SYN_Bhe of mux21_SIZE4_5 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => IN0(3), B => IN1(3), S => CTRL, Z => OUT1(3));
   U2 : MUX2_X1 port map( A => IN0(2), B => IN1(2), S => CTRL, Z => OUT1(2));
   U3 : MUX2_X1 port map( A => IN0(1), B => IN1(1), S => CTRL, Z => OUT1(1));
   U4 : MUX2_X1 port map( A => IN0(0), B => IN1(0), S => CTRL, Z => OUT1(0));

end SYN_Bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity mux21_SIZE4_4 is

   port( IN0, IN1 : in std_logic_vector (3 downto 0);  CTRL : in std_logic;  
         OUT1 : out std_logic_vector (3 downto 0));

end mux21_SIZE4_4;

architecture SYN_Bhe of mux21_SIZE4_4 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => IN0(3), B => IN1(3), S => CTRL, Z => OUT1(3));
   U2 : MUX2_X1 port map( A => IN0(2), B => IN1(2), S => CTRL, Z => OUT1(2));
   U3 : MUX2_X1 port map( A => IN0(1), B => IN1(1), S => CTRL, Z => OUT1(1));
   U4 : MUX2_X1 port map( A => IN0(0), B => IN1(0), S => CTRL, Z => OUT1(0));

end SYN_Bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity mux21_SIZE4_3 is

   port( IN0, IN1 : in std_logic_vector (3 downto 0);  CTRL : in std_logic;  
         OUT1 : out std_logic_vector (3 downto 0));

end mux21_SIZE4_3;

architecture SYN_Bhe of mux21_SIZE4_3 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => IN0(3), B => IN1(3), S => CTRL, Z => OUT1(3));
   U2 : MUX2_X1 port map( A => IN0(2), B => IN1(2), S => CTRL, Z => OUT1(2));
   U3 : MUX2_X1 port map( A => IN0(0), B => IN1(0), S => CTRL, Z => OUT1(0));
   U4 : MUX2_X1 port map( A => IN0(1), B => IN1(1), S => CTRL, Z => OUT1(1));

end SYN_Bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity mux21_SIZE4_2 is

   port( IN0, IN1 : in std_logic_vector (3 downto 0);  CTRL : in std_logic;  
         OUT1 : out std_logic_vector (3 downto 0));

end mux21_SIZE4_2;

architecture SYN_Bhe of mux21_SIZE4_2 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => IN0(3), B => IN1(3), S => CTRL, Z => OUT1(3));
   U2 : MUX2_X1 port map( A => IN0(2), B => IN1(2), S => CTRL, Z => OUT1(2));
   U3 : MUX2_X1 port map( A => IN0(1), B => IN1(1), S => CTRL, Z => OUT1(1));
   U4 : MUX2_X1 port map( A => IN0(0), B => IN1(0), S => CTRL, Z => OUT1(0));

end SYN_Bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity mux21_SIZE4_1 is

   port( IN0, IN1 : in std_logic_vector (3 downto 0);  CTRL : in std_logic;  
         OUT1 : out std_logic_vector (3 downto 0));

end mux21_SIZE4_1;

architecture SYN_Bhe of mux21_SIZE4_1 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : MUX2_X1 port map( A => IN0(2), B => IN1(2), S => CTRL, Z => OUT1(2));
   U3 : MUX2_X1 port map( A => IN0(1), B => IN1(1), S => CTRL, Z => OUT1(1));
   U4 : MUX2_X1 port map( A => IN0(0), B => IN1(0), S => CTRL, Z => OUT1(0));
   U1 : MUX2_X1 port map( A => IN0(3), B => IN1(3), S => CTRL, Z => OUT1(3));

end SYN_Bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity RCA_N4_30 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_30;

architecture SYN_STRUCTURAL of RCA_N4_30 is

   component FA_117
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_118
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_119
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_120
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal n1, CTMP_3_port, CTMP_2_port, CTMP_1_port, net246205 : std_logic;

begin
   
   FAI_1 : FA_120 port map( A => A(0), B => B(0), Ci => n1, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_119 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_118 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_117 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => net246205);
   n1 <= '0';

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity RCA_N4_29 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_29;

architecture SYN_STRUCTURAL of RCA_N4_29 is

   component FA_113
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_114
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_115
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_116
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal n1, CTMP_3_port, CTMP_2_port, CTMP_1_port, net246204 : std_logic;

begin
   
   FAI_1 : FA_116 port map( A => A(0), B => B(0), Ci => n1, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_115 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_114 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_113 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => net246204);
   n1 <= '1';

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity RCA_N4_28 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_28;

architecture SYN_STRUCTURAL of RCA_N4_28 is

   component FA_109
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_110
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_111
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_112
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal n1, CTMP_3_port, CTMP_2_port, CTMP_1_port, net246203 : std_logic;

begin
   
   FAI_1 : FA_112 port map( A => A(0), B => B(0), Ci => n1, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_111 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_110 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_109 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => net246203);
   n1 <= '0';

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity RCA_N4_27 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_27;

architecture SYN_STRUCTURAL of RCA_N4_27 is

   component FA_105
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_106
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_107
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_108
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal n1, CTMP_3_port, CTMP_2_port, CTMP_1_port, net246202 : std_logic;

begin
   
   FAI_1 : FA_108 port map( A => A(0), B => B(0), Ci => n1, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_107 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_106 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_105 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => net246202);
   n1 <= '1';

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity RCA_N4_26 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_26;

architecture SYN_STRUCTURAL of RCA_N4_26 is

   component FA_101
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_102
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_103
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_104
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal n1, CTMP_3_port, CTMP_2_port, CTMP_1_port, net246201 : std_logic;

begin
   
   FAI_1 : FA_104 port map( A => A(0), B => B(0), Ci => n1, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_103 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_102 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_101 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => net246201);
   n1 <= '0';

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity RCA_N4_25 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_25;

architecture SYN_STRUCTURAL of RCA_N4_25 is

   component FA_97
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_98
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_99
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_100
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal n1, CTMP_3_port, CTMP_2_port, CTMP_1_port, net246200 : std_logic;

begin
   
   FAI_1 : FA_100 port map( A => A(0), B => B(0), Ci => n1, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_99 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_98 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_97 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => net246200);
   n1 <= '1';

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity RCA_N4_24 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_24;

architecture SYN_STRUCTURAL of RCA_N4_24 is

   component FA_93
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_94
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_95
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_96
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal n2, CTMP_3_port, CTMP_2_port, CTMP_1_port, net246199 : std_logic;

begin
   
   FAI_1 : FA_96 port map( A => A(0), B => B(0), Ci => n2, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_95 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_94 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_93 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => net246199);
   n2 <= '0';

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity RCA_N4_23 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_23;

architecture SYN_STRUCTURAL of RCA_N4_23 is

   component FA_89
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_90
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_91
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_92
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal n2, CTMP_3_port, CTMP_2_port, CTMP_1_port, net246198 : std_logic;

begin
   
   FAI_1 : FA_92 port map( A => A(0), B => B(0), Ci => n2, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_91 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_90 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_89 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => net246198);
   n2 <= '1';

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity RCA_N4_22 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_22;

architecture SYN_STRUCTURAL of RCA_N4_22 is

   component FA_85
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_86
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_87
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_88
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal n1, CTMP_3_port, CTMP_2_port, CTMP_1_port, net246197 : std_logic;

begin
   
   FAI_1 : FA_88 port map( A => A(0), B => B(0), Ci => n1, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_87 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_86 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_85 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => net246197);
   n1 <= '0';

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity RCA_N4_21 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_21;

architecture SYN_STRUCTURAL of RCA_N4_21 is

   component FA_81
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_82
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_83
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_84
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal n1, CTMP_3_port, CTMP_2_port, CTMP_1_port, net246196 : std_logic;

begin
   
   FAI_1 : FA_84 port map( A => A(0), B => B(0), Ci => n1, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_83 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_82 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_81 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => net246196);
   n1 <= '1';

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity RCA_N4_20 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_20;

architecture SYN_STRUCTURAL of RCA_N4_20 is

   component FA_77
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_78
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_79
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_80
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal n3, CTMP_3_port, CTMP_2_port, CTMP_1_port, net246195 : std_logic;

begin
   
   FAI_1 : FA_80 port map( A => A(0), B => B(0), Ci => n3, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_79 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_78 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_77 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => net246195);
   n3 <= '0';

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity RCA_N4_19 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_19;

architecture SYN_STRUCTURAL of RCA_N4_19 is

   component FA_73
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_74
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_75
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_76
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal n3, CTMP_3_port, CTMP_2_port, CTMP_1_port, net246194 : std_logic;

begin
   
   FAI_1 : FA_76 port map( A => A(0), B => B(0), Ci => n3, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_75 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_74 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_73 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => net246194);
   n3 <= '1';

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity RCA_N4_18 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_18;

architecture SYN_STRUCTURAL of RCA_N4_18 is

   component FA_69
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_70
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_71
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_72
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal n2, CTMP_3_port, CTMP_2_port, CTMP_1_port, net246193 : std_logic;

begin
   
   FAI_1 : FA_72 port map( A => A(0), B => B(0), Ci => n2, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_71 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_70 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_69 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => net246193);
   n2 <= '0';

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity RCA_N4_17 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_17;

architecture SYN_STRUCTURAL of RCA_N4_17 is

   component FA_65
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_66
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_67
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_68
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal n2, CTMP_3_port, CTMP_2_port, CTMP_1_port, net246192 : std_logic;

begin
   
   FAI_1 : FA_68 port map( A => A(0), B => B(0), Ci => n2, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_67 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_66 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_65 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => net246192);
   n2 <= '1';

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity RCA_N4_16 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_16;

architecture SYN_STRUCTURAL of RCA_N4_16 is

   component FA_61
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_62
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_63
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_64
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal n2, CTMP_3_port, CTMP_2_port, CTMP_1_port, net246191 : std_logic;

begin
   
   FAI_1 : FA_64 port map( A => A(0), B => B(0), Ci => n2, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_63 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_62 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_61 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => net246191);
   n2 <= '0';

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity RCA_N4_15 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_15;

architecture SYN_STRUCTURAL of RCA_N4_15 is

   component FA_57
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_58
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_59
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_60
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal n2, CTMP_3_port, CTMP_2_port, CTMP_1_port, net246190 : std_logic;

begin
   
   FAI_1 : FA_60 port map( A => A(0), B => B(0), Ci => n2, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_59 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_58 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_57 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => net246190);
   n2 <= '1';

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity RCA_N4_14 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_14;

architecture SYN_STRUCTURAL of RCA_N4_14 is

   component FA_53
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_54
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_55
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_56
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal n1, CTMP_3_port, CTMP_2_port, CTMP_1_port, net246189 : std_logic;

begin
   
   FAI_1 : FA_56 port map( A => A(0), B => B(0), Ci => n1, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_55 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_54 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_53 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => net246189);
   n1 <= '0';

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity RCA_N4_13 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_13;

architecture SYN_STRUCTURAL of RCA_N4_13 is

   component FA_49
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_50
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_51
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_52
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal n1, CTMP_3_port, CTMP_2_port, CTMP_1_port, net246188 : std_logic;

begin
   
   FAI_1 : FA_52 port map( A => A(0), B => B(0), Ci => n1, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_51 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_50 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_49 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => net246188);
   n1 <= '1';

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity RCA_N4_12 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_12;

architecture SYN_STRUCTURAL of RCA_N4_12 is

   component FA_45
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_46
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_47
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_48
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal n1, CTMP_3_port, CTMP_2_port, CTMP_1_port, net246187 : std_logic;

begin
   
   FAI_1 : FA_48 port map( A => A(0), B => B(0), Ci => n1, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_47 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_46 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_45 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => net246187);
   n1 <= '0';

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity RCA_N4_11 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_11;

architecture SYN_STRUCTURAL of RCA_N4_11 is

   component FA_41
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_42
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_43
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_44
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal n1, CTMP_3_port, CTMP_2_port, CTMP_1_port, net246186 : std_logic;

begin
   
   FAI_1 : FA_44 port map( A => A(0), B => B(0), Ci => n1, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_43 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_42 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_41 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => net246186);
   n1 <= '1';

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity RCA_N4_10 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_10;

architecture SYN_STRUCTURAL of RCA_N4_10 is

   component FA_37
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_38
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_39
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_40
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal n1, CTMP_3_port, CTMP_2_port, CTMP_1_port, net246185 : std_logic;

begin
   
   FAI_1 : FA_40 port map( A => A(0), B => B(0), Ci => n1, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_39 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_38 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_37 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => net246185);
   n1 <= '0';

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity RCA_N4_9 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_9;

architecture SYN_STRUCTURAL of RCA_N4_9 is

   component FA_33
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_34
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_35
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_36
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal n1, CTMP_3_port, CTMP_2_port, CTMP_1_port, net246184 : std_logic;

begin
   
   FAI_1 : FA_36 port map( A => A(0), B => B(0), Ci => n1, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_35 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_34 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_33 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => net246184);
   n1 <= '1';

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity RCA_N4_8 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_8;

architecture SYN_STRUCTURAL of RCA_N4_8 is

   component FA_29
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_30
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_31
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_32
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal n1, CTMP_3_port, CTMP_2_port, CTMP_1_port, net246183 : std_logic;

begin
   
   FAI_1 : FA_32 port map( A => A(0), B => B(0), Ci => n1, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_31 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_30 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_29 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => net246183);
   n1 <= '0';

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity RCA_N4_7 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_7;

architecture SYN_STRUCTURAL of RCA_N4_7 is

   component FA_25
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_26
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_27
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_28
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal n1, CTMP_3_port, CTMP_2_port, CTMP_1_port, net246182 : std_logic;

begin
   
   FAI_1 : FA_28 port map( A => A(0), B => B(0), Ci => n1, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_27 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_26 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_25 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => net246182);
   n1 <= '1';

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity RCA_N4_6 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_6;

architecture SYN_STRUCTURAL of RCA_N4_6 is

   component FA_21
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_22
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_23
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_24
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal n1, CTMP_3_port, CTMP_2_port, CTMP_1_port, net246181 : std_logic;

begin
   
   FAI_1 : FA_24 port map( A => A(0), B => B(0), Ci => n1, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_23 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_22 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_21 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => net246181);
   n1 <= '0';

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity RCA_N4_5 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_5;

architecture SYN_STRUCTURAL of RCA_N4_5 is

   component FA_17
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_18
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_19
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_20
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal n1, CTMP_3_port, CTMP_2_port, CTMP_1_port, net246180 : std_logic;

begin
   
   FAI_1 : FA_20 port map( A => A(0), B => B(0), Ci => n1, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_19 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_18 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_17 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => net246180);
   n1 <= '1';

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity RCA_N4_4 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_4;

architecture SYN_STRUCTURAL of RCA_N4_4 is

   component FA_13
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_14
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_15
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_16
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal n1, CTMP_3_port, CTMP_2_port, CTMP_1_port, net246179 : std_logic;

begin
   
   FAI_1 : FA_16 port map( A => A(0), B => B(0), Ci => n1, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_15 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_14 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_13 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => net246179);
   n1 <= '0';

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity RCA_N4_3 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_3;

architecture SYN_STRUCTURAL of RCA_N4_3 is

   component FA_9
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_10
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_11
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_12
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal n1, CTMP_3_port, CTMP_2_port, CTMP_1_port, net246178 : std_logic;

begin
   
   FAI_1 : FA_12 port map( A => A(0), B => B(0), Ci => n1, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_11 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_10 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_9 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => net246178);
   n1 <= '1';

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity RCA_N4_2 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_2;

architecture SYN_STRUCTURAL of RCA_N4_2 is

   component FA_5
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_6
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_7
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_8
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal n1, CTMP_3_port, CTMP_2_port, CTMP_1_port, net246177 : std_logic;

begin
   
   FAI_1 : FA_8 port map( A => A(0), B => B(0), Ci => n1, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_7 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_6 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_5 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => net246177);
   n1 <= '0';

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity RCA_N4_1 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_1;

architecture SYN_STRUCTURAL of RCA_N4_1 is

   component FA_1
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_2
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_3
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_4
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal n1, CTMP_3_port, CTMP_2_port, CTMP_1_port, net246176 : std_logic;

begin
   
   FAI_1 : FA_4 port map( A => A(0), B => B(0), Ci => n1, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_3 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_2 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_1 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => net246176);
   n1 <= '1';

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity shift_N9_2 is

   port( Clock, ALOAD : in std_logic;  D : in std_logic_vector (8 downto 0);  
         SO : out std_logic);

end shift_N9_2;

architecture SYN_archi of shift_N9_2 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component SDFF_X1
      port( D, SI, SE, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal tmp_8_port, tmp_7_port, tmp_6_port, tmp_5_port, tmp_4_port, 
      tmp_3_port, tmp_2_port, tmp_1_port, N11, n1, n10, n11_port, n12, n13, n14
      , n15, n16, n17 : std_logic;

begin
   
   tmp_reg_8_inst : DFF_X1 port map( D => N11, CK => Clock, Q => tmp_8_port, QN
                           => n1);
   tmp_reg_7_inst : SDFF_X1 port map( D => tmp_8_port, SI => D(7), SE => ALOAD,
                           CK => Clock, Q => tmp_7_port, QN => n10);
   tmp_reg_6_inst : SDFF_X1 port map( D => tmp_7_port, SI => D(6), SE => ALOAD,
                           CK => Clock, Q => tmp_6_port, QN => n11_port);
   tmp_reg_5_inst : SDFF_X1 port map( D => tmp_6_port, SI => D(5), SE => ALOAD,
                           CK => Clock, Q => tmp_5_port, QN => n12);
   tmp_reg_4_inst : SDFF_X1 port map( D => tmp_5_port, SI => D(4), SE => ALOAD,
                           CK => Clock, Q => tmp_4_port, QN => n13);
   tmp_reg_3_inst : SDFF_X1 port map( D => tmp_4_port, SI => D(3), SE => ALOAD,
                           CK => Clock, Q => tmp_3_port, QN => n14);
   tmp_reg_2_inst : SDFF_X1 port map( D => tmp_3_port, SI => D(2), SE => ALOAD,
                           CK => Clock, Q => tmp_2_port, QN => n15);
   tmp_reg_1_inst : SDFF_X1 port map( D => tmp_2_port, SI => D(1), SE => ALOAD,
                           CK => Clock, Q => tmp_1_port, QN => n16);
   tmp_reg_0_inst : SDFF_X1 port map( D => tmp_1_port, SI => D(0), SE => ALOAD,
                           CK => Clock, Q => SO, QN => n17);
   U3 : AND2_X1 port map( A1 => ALOAD, A2 => D(8), ZN => N11);

end SYN_archi;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity shift_N9_1 is

   port( Clock, ALOAD : in std_logic;  D : in std_logic_vector (8 downto 0);  
         SO : out std_logic);

end shift_N9_1;

architecture SYN_archi of shift_N9_1 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component SDFF_X2
      port( D, SI, SE, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component SDFF_X1
      port( D, SI, SE, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal tmp_8_port, tmp_7_port, tmp_6_port, tmp_5_port, tmp_4_port, 
      tmp_3_port, tmp_2_port, tmp_1_port, N11, n1, n2, n10, n11_port, n12, n13,
      n14, n15, n16 : std_logic;

begin
   
   tmp_reg_8_inst : DFF_X1 port map( D => N11, CK => Clock, Q => tmp_8_port, QN
                           => n2);
   tmp_reg_7_inst : SDFF_X1 port map( D => tmp_8_port, SI => D(7), SE => ALOAD,
                           CK => Clock, Q => tmp_7_port, QN => n10);
   tmp_reg_6_inst : SDFF_X1 port map( D => tmp_7_port, SI => D(6), SE => ALOAD,
                           CK => Clock, Q => tmp_6_port, QN => n11_port);
   tmp_reg_5_inst : SDFF_X1 port map( D => tmp_6_port, SI => D(5), SE => ALOAD,
                           CK => Clock, Q => tmp_5_port, QN => n12);
   tmp_reg_4_inst : SDFF_X1 port map( D => tmp_5_port, SI => D(4), SE => ALOAD,
                           CK => Clock, Q => tmp_4_port, QN => n13);
   tmp_reg_3_inst : SDFF_X1 port map( D => tmp_4_port, SI => D(3), SE => ALOAD,
                           CK => Clock, Q => tmp_3_port, QN => n14);
   tmp_reg_2_inst : SDFF_X1 port map( D => tmp_3_port, SI => D(2), SE => ALOAD,
                           CK => Clock, Q => tmp_2_port, QN => n15);
   tmp_reg_1_inst : SDFF_X1 port map( D => tmp_2_port, SI => D(1), SE => ALOAD,
                           CK => Clock, Q => tmp_1_port, QN => n16);
   tmp_reg_0_inst : SDFF_X2 port map( D => tmp_1_port, SI => D(0), SE => ALOAD,
                           CK => Clock, Q => SO, QN => n1);
   U3 : AND2_X1 port map( A1 => ALOAD, A2 => D(8), ZN => N11);

end SYN_archi;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity booth_encoder_8 is

   port( B_in : in std_logic_vector (2 downto 0);  A_out : out std_logic_vector
         (2 downto 0));

end booth_encoder_8;

architecture SYN_bhe of booth_encoder_8 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI33_X1
      port( A1, A2, A3, B1, B2, B3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n5, n6, n7 : std_logic;

begin
   
   U6 : OAI33_X1 port map( A1 => B_in(0), A2 => B_in(1), A3 => n1, B1 => n7, B2
                           => n6, B3 => B_in(2), ZN => A_out(0));
   U4 : NAND2_X1 port map( A1 => B_in(2), A2 => n7, ZN => n5);
   U9 : INV_X1 port map( A => B_in(2), ZN => n1);
   U3 : INV_X1 port map( A => B_in(0), ZN => n7);
   U5 : INV_X1 port map( A => B_in(1), ZN => n6);
   U7 : OAI221_X1 port map( B1 => B_in(1), B2 => n7, C1 => n6, C2 => B_in(2), A
                           => n5, ZN => A_out(2));
   U8 : AOI21_X1 port map( B1 => B_in(0), B2 => B_in(1), A => n1, ZN => 
                           A_out(1));

end SYN_bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity booth_encoder_7 is

   port( B_in : in std_logic_vector (2 downto 0);  A_out : out std_logic_vector
         (2 downto 0));

end booth_encoder_7;

architecture SYN_bhe of booth_encoder_7 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI33_X1
      port( A1, A2, A3, B1, B2, B3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n5, n6, n7 : std_logic;

begin
   
   U6 : OAI33_X1 port map( A1 => B_in(0), A2 => B_in(1), A3 => n1, B1 => n7, B2
                           => n6, B3 => B_in(2), ZN => A_out(0));
   U8 : INV_X1 port map( A => B_in(0), ZN => n7);
   U3 : INV_X1 port map( A => B_in(2), ZN => n1);
   U4 : INV_X1 port map( A => B_in(1), ZN => n6);
   U5 : AOI21_X1 port map( B1 => B_in(0), B2 => B_in(1), A => n1, ZN => 
                           A_out(1));
   U7 : OAI221_X1 port map( B1 => B_in(1), B2 => n7, C1 => n6, C2 => B_in(2), A
                           => n5, ZN => A_out(2));
   U9 : NAND2_X1 port map( A1 => B_in(2), A2 => n7, ZN => n5);

end SYN_bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity booth_encoder_6 is

   port( B_in : in std_logic_vector (2 downto 0);  A_out : out std_logic_vector
         (2 downto 0));

end booth_encoder_6;

architecture SYN_bhe of booth_encoder_6 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI33_X1
      port( A1, A2, A3, B1, B2, B3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n5, n6, n7 : std_logic;

begin
   
   U6 : OAI33_X1 port map( A1 => B_in(0), A2 => B_in(1), A3 => n1, B1 => n7, B2
                           => n6, B3 => B_in(2), ZN => A_out(0));
   U3 : INV_X1 port map( A => B_in(2), ZN => n1);
   U4 : INV_X1 port map( A => B_in(0), ZN => n7);
   U5 : INV_X1 port map( A => B_in(1), ZN => n6);
   U7 : NAND2_X1 port map( A1 => B_in(2), A2 => n7, ZN => n5);
   U8 : OAI221_X1 port map( B1 => B_in(1), B2 => n7, C1 => n6, C2 => B_in(2), A
                           => n5, ZN => A_out(2));
   U9 : AOI21_X1 port map( B1 => B_in(0), B2 => B_in(1), A => n1, ZN => 
                           A_out(1));

end SYN_bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity booth_encoder_5 is

   port( B_in : in std_logic_vector (2 downto 0);  A_out : out std_logic_vector
         (2 downto 0));

end booth_encoder_5;

architecture SYN_bhe of booth_encoder_5 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI33_X1
      port( A1, A2, A3, B1, B2, B3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n5, n6, n7 : std_logic;

begin
   
   U6 : OAI33_X1 port map( A1 => B_in(0), A2 => B_in(1), A3 => n1, B1 => n7, B2
                           => n6, B3 => B_in(2), ZN => A_out(0));
   U7 : INV_X1 port map( A => B_in(1), ZN => n6);
   U3 : INV_X1 port map( A => B_in(0), ZN => n7);
   U4 : INV_X1 port map( A => B_in(2), ZN => n1);
   U5 : OAI221_X1 port map( B1 => B_in(1), B2 => n7, C1 => n6, C2 => B_in(2), A
                           => n5, ZN => A_out(2));
   U8 : NAND2_X1 port map( A1 => B_in(2), A2 => n7, ZN => n5);
   U9 : AOI21_X1 port map( B1 => B_in(0), B2 => B_in(1), A => n1, ZN => 
                           A_out(1));

end SYN_bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity booth_encoder_4 is

   port( B_in : in std_logic_vector (2 downto 0);  A_out : out std_logic_vector
         (2 downto 0));

end booth_encoder_4;

architecture SYN_bhe of booth_encoder_4 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI33_X1
      port( A1, A2, A3, B1, B2, B3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n5, n6, n7 : std_logic;

begin
   
   U6 : OAI33_X1 port map( A1 => B_in(0), A2 => B_in(1), A3 => n1, B1 => n7, B2
                           => n6, B3 => B_in(2), ZN => A_out(0));
   U3 : INV_X1 port map( A => B_in(0), ZN => n7);
   U4 : INV_X1 port map( A => B_in(1), ZN => n6);
   U5 : INV_X1 port map( A => B_in(2), ZN => n1);
   U7 : AOI21_X1 port map( B1 => B_in(0), B2 => B_in(1), A => n1, ZN => 
                           A_out(1));
   U8 : OAI221_X1 port map( B1 => B_in(1), B2 => n7, C1 => n6, C2 => B_in(2), A
                           => n5, ZN => A_out(2));
   U9 : NAND2_X1 port map( A1 => B_in(2), A2 => n7, ZN => n5);

end SYN_bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity booth_encoder_3 is

   port( B_in : in std_logic_vector (2 downto 0);  A_out : out std_logic_vector
         (2 downto 0));

end booth_encoder_3;

architecture SYN_bhe of booth_encoder_3 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI33_X1
      port( A1, A2, A3, B1, B2, B3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n5, n6, n7 : std_logic;

begin
   
   U6 : OAI33_X1 port map( A1 => B_in(0), A2 => B_in(1), A3 => n1, B1 => n7, B2
                           => n6, B3 => B_in(2), ZN => A_out(0));
   U7 : INV_X1 port map( A => B_in(1), ZN => n6);
   U3 : INV_X1 port map( A => B_in(2), ZN => n1);
   U4 : INV_X1 port map( A => B_in(0), ZN => n7);
   U5 : NAND2_X1 port map( A1 => B_in(2), A2 => n7, ZN => n5);
   U8 : OAI221_X1 port map( B1 => B_in(1), B2 => n7, C1 => n6, C2 => B_in(2), A
                           => n5, ZN => A_out(2));
   U9 : AOI21_X1 port map( B1 => B_in(0), B2 => B_in(1), A => n1, ZN => 
                           A_out(1));

end SYN_bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity booth_encoder_2 is

   port( B_in : in std_logic_vector (2 downto 0);  A_out : out std_logic_vector
         (2 downto 0));

end booth_encoder_2;

architecture SYN_bhe of booth_encoder_2 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI33_X1
      port( A1, A2, A3, B1, B2, B3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n5, n6, n7 : std_logic;

begin
   
   U6 : OAI33_X1 port map( A1 => B_in(0), A2 => B_in(1), A3 => n1, B1 => n7, B2
                           => n6, B3 => B_in(2), ZN => A_out(0));
   U3 : INV_X1 port map( A => B_in(1), ZN => n6);
   U4 : INV_X1 port map( A => B_in(0), ZN => n7);
   U5 : INV_X1 port map( A => B_in(2), ZN => n1);
   U7 : AOI21_X1 port map( B1 => B_in(0), B2 => B_in(1), A => n1, ZN => 
                           A_out(1));
   U8 : OAI221_X1 port map( B1 => B_in(1), B2 => n7, C1 => n6, C2 => B_in(2), A
                           => n5, ZN => A_out(2));
   U9 : NAND2_X1 port map( A1 => B_in(2), A2 => n7, ZN => n5);

end SYN_bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity booth_encoder_1 is

   port( B_in : in std_logic_vector (2 downto 0);  A_out : out std_logic_vector
         (2 downto 0));

end booth_encoder_1;

architecture SYN_bhe of booth_encoder_1 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI33_X1
      port( A1, A2, A3, B1, B2, B3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4, n5 : std_logic;

begin
   
   U6 : OAI33_X1 port map( A1 => B_in(0), A2 => B_in(1), A3 => n4, B1 => n5, B2
                           => n4, B3 => B_in(2), ZN => A_out(0));
   U4 : NAND2_X1 port map( A1 => B_in(2), A2 => n5, ZN => n1);
   U3 : OAI221_X1 port map( B1 => B_in(1), B2 => n5, C1 => n4, C2 => B_in(2), A
                           => n1, ZN => A_out(2));
   U5 : INV_X1 port map( A => B_in(1), ZN => n4);
   U7 : INV_X1 port map( A => B_in(0), ZN => n5);
   U8 : AOI21_X1 port map( B1 => B_in(0), B2 => B_in(1), A => n4, ZN => 
                           A_out(1));

end SYN_bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity carry_sel_gen_N4_15 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end carry_sel_gen_N4_15;

architecture SYN_STRUCTURAL of carry_sel_gen_N4_15 is

   component mux21_SIZE4_15
      port( IN0, IN1 : in std_logic_vector (3 downto 0);  CTRL : in std_logic; 
            OUT1 : out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_N4_29
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_30
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, nocarry_sum_to_mux_3_port, 
      nocarry_sum_to_mux_2_port, nocarry_sum_to_mux_1_port, 
      nocarry_sum_to_mux_0_port, carry_sum_to_mux_3_port, 
      carry_sum_to_mux_2_port, carry_sum_to_mux_1_port, carry_sum_to_mux_0_port
      , net246174, net246175 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   rca_nocarry : RCA_N4_30 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           nocarry_sum_to_mux_3_port, S(2) => 
                           nocarry_sum_to_mux_2_port, S(1) => 
                           nocarry_sum_to_mux_1_port, S(0) => 
                           nocarry_sum_to_mux_0_port, Co => net246175);
   rca_carry : RCA_N4_29 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           carry_sum_to_mux_3_port, S(2) => 
                           carry_sum_to_mux_2_port, S(1) => 
                           carry_sum_to_mux_1_port, S(0) => 
                           carry_sum_to_mux_0_port, Co => net246174);
   outmux : mux21_SIZE4_15 port map( IN0(3) => nocarry_sum_to_mux_3_port, 
                           IN0(2) => nocarry_sum_to_mux_2_port, IN0(1) => 
                           nocarry_sum_to_mux_1_port, IN0(0) => 
                           nocarry_sum_to_mux_0_port, IN1(3) => 
                           carry_sum_to_mux_3_port, IN1(2) => 
                           carry_sum_to_mux_2_port, IN1(1) => 
                           carry_sum_to_mux_1_port, IN1(0) => 
                           carry_sum_to_mux_0_port, CTRL => Ci, OUT1(3) => S(3)
                           , OUT1(2) => S(2), OUT1(1) => S(1), OUT1(0) => S(0))
                           ;

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity carry_sel_gen_N4_14 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end carry_sel_gen_N4_14;

architecture SYN_STRUCTURAL of carry_sel_gen_N4_14 is

   component mux21_SIZE4_14
      port( IN0, IN1 : in std_logic_vector (3 downto 0);  CTRL : in std_logic; 
            OUT1 : out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_N4_27
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_28
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, nocarry_sum_to_mux_3_port, 
      nocarry_sum_to_mux_2_port, nocarry_sum_to_mux_1_port, 
      nocarry_sum_to_mux_0_port, carry_sum_to_mux_3_port, 
      carry_sum_to_mux_2_port, carry_sum_to_mux_1_port, carry_sum_to_mux_0_port
      , net246172, net246173 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   rca_nocarry : RCA_N4_28 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           nocarry_sum_to_mux_3_port, S(2) => 
                           nocarry_sum_to_mux_2_port, S(1) => 
                           nocarry_sum_to_mux_1_port, S(0) => 
                           nocarry_sum_to_mux_0_port, Co => net246173);
   rca_carry : RCA_N4_27 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           carry_sum_to_mux_3_port, S(2) => 
                           carry_sum_to_mux_2_port, S(1) => 
                           carry_sum_to_mux_1_port, S(0) => 
                           carry_sum_to_mux_0_port, Co => net246172);
   outmux : mux21_SIZE4_14 port map( IN0(3) => nocarry_sum_to_mux_3_port, 
                           IN0(2) => nocarry_sum_to_mux_2_port, IN0(1) => 
                           nocarry_sum_to_mux_1_port, IN0(0) => 
                           nocarry_sum_to_mux_0_port, IN1(3) => 
                           carry_sum_to_mux_3_port, IN1(2) => 
                           carry_sum_to_mux_2_port, IN1(1) => 
                           carry_sum_to_mux_1_port, IN1(0) => 
                           carry_sum_to_mux_0_port, CTRL => Ci, OUT1(3) => S(3)
                           , OUT1(2) => S(2), OUT1(1) => S(1), OUT1(0) => S(0))
                           ;

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity carry_sel_gen_N4_13 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end carry_sel_gen_N4_13;

architecture SYN_STRUCTURAL of carry_sel_gen_N4_13 is

   component mux21_SIZE4_13
      port( IN0, IN1 : in std_logic_vector (3 downto 0);  CTRL : in std_logic; 
            OUT1 : out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_N4_25
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_26
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, nocarry_sum_to_mux_3_port, 
      nocarry_sum_to_mux_2_port, nocarry_sum_to_mux_1_port, 
      nocarry_sum_to_mux_0_port, carry_sum_to_mux_3_port, 
      carry_sum_to_mux_2_port, carry_sum_to_mux_1_port, carry_sum_to_mux_0_port
      , net246170, net246171 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   rca_nocarry : RCA_N4_26 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           nocarry_sum_to_mux_3_port, S(2) => 
                           nocarry_sum_to_mux_2_port, S(1) => 
                           nocarry_sum_to_mux_1_port, S(0) => 
                           nocarry_sum_to_mux_0_port, Co => net246171);
   rca_carry : RCA_N4_25 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           carry_sum_to_mux_3_port, S(2) => 
                           carry_sum_to_mux_2_port, S(1) => 
                           carry_sum_to_mux_1_port, S(0) => 
                           carry_sum_to_mux_0_port, Co => net246170);
   outmux : mux21_SIZE4_13 port map( IN0(3) => nocarry_sum_to_mux_3_port, 
                           IN0(2) => nocarry_sum_to_mux_2_port, IN0(1) => 
                           nocarry_sum_to_mux_1_port, IN0(0) => 
                           nocarry_sum_to_mux_0_port, IN1(3) => 
                           carry_sum_to_mux_3_port, IN1(2) => 
                           carry_sum_to_mux_2_port, IN1(1) => 
                           carry_sum_to_mux_1_port, IN1(0) => 
                           carry_sum_to_mux_0_port, CTRL => Ci, OUT1(3) => S(3)
                           , OUT1(2) => S(2), OUT1(1) => S(1), OUT1(0) => S(0))
                           ;

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity carry_sel_gen_N4_12 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end carry_sel_gen_N4_12;

architecture SYN_STRUCTURAL of carry_sel_gen_N4_12 is

   component mux21_SIZE4_12
      port( IN0, IN1 : in std_logic_vector (3 downto 0);  CTRL : in std_logic; 
            OUT1 : out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_N4_23
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_24
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, nocarry_sum_to_mux_3_port, 
      nocarry_sum_to_mux_2_port, nocarry_sum_to_mux_1_port, 
      nocarry_sum_to_mux_0_port, carry_sum_to_mux_3_port, 
      carry_sum_to_mux_2_port, carry_sum_to_mux_1_port, carry_sum_to_mux_0_port
      , net246168, net246169 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   rca_nocarry : RCA_N4_24 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           nocarry_sum_to_mux_3_port, S(2) => 
                           nocarry_sum_to_mux_2_port, S(1) => 
                           nocarry_sum_to_mux_1_port, S(0) => 
                           nocarry_sum_to_mux_0_port, Co => net246169);
   rca_carry : RCA_N4_23 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           carry_sum_to_mux_3_port, S(2) => 
                           carry_sum_to_mux_2_port, S(1) => 
                           carry_sum_to_mux_1_port, S(0) => 
                           carry_sum_to_mux_0_port, Co => net246168);
   outmux : mux21_SIZE4_12 port map( IN0(3) => nocarry_sum_to_mux_3_port, 
                           IN0(2) => nocarry_sum_to_mux_2_port, IN0(1) => 
                           nocarry_sum_to_mux_1_port, IN0(0) => 
                           nocarry_sum_to_mux_0_port, IN1(3) => 
                           carry_sum_to_mux_3_port, IN1(2) => 
                           carry_sum_to_mux_2_port, IN1(1) => 
                           carry_sum_to_mux_1_port, IN1(0) => 
                           carry_sum_to_mux_0_port, CTRL => Ci, OUT1(3) => S(3)
                           , OUT1(2) => S(2), OUT1(1) => S(1), OUT1(0) => S(0))
                           ;

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity carry_sel_gen_N4_11 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end carry_sel_gen_N4_11;

architecture SYN_STRUCTURAL of carry_sel_gen_N4_11 is

   component mux21_SIZE4_11
      port( IN0, IN1 : in std_logic_vector (3 downto 0);  CTRL : in std_logic; 
            OUT1 : out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_N4_21
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_22
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, nocarry_sum_to_mux_3_port, 
      nocarry_sum_to_mux_2_port, nocarry_sum_to_mux_1_port, 
      nocarry_sum_to_mux_0_port, carry_sum_to_mux_3_port, 
      carry_sum_to_mux_2_port, carry_sum_to_mux_1_port, carry_sum_to_mux_0_port
      , net246166, net246167 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   rca_nocarry : RCA_N4_22 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           nocarry_sum_to_mux_3_port, S(2) => 
                           nocarry_sum_to_mux_2_port, S(1) => 
                           nocarry_sum_to_mux_1_port, S(0) => 
                           nocarry_sum_to_mux_0_port, Co => net246167);
   rca_carry : RCA_N4_21 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           carry_sum_to_mux_3_port, S(2) => 
                           carry_sum_to_mux_2_port, S(1) => 
                           carry_sum_to_mux_1_port, S(0) => 
                           carry_sum_to_mux_0_port, Co => net246166);
   outmux : mux21_SIZE4_11 port map( IN0(3) => nocarry_sum_to_mux_3_port, 
                           IN0(2) => nocarry_sum_to_mux_2_port, IN0(1) => 
                           nocarry_sum_to_mux_1_port, IN0(0) => 
                           nocarry_sum_to_mux_0_port, IN1(3) => 
                           carry_sum_to_mux_3_port, IN1(2) => 
                           carry_sum_to_mux_2_port, IN1(1) => 
                           carry_sum_to_mux_1_port, IN1(0) => 
                           carry_sum_to_mux_0_port, CTRL => Ci, OUT1(3) => S(3)
                           , OUT1(2) => S(2), OUT1(1) => S(1), OUT1(0) => S(0))
                           ;

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity carry_sel_gen_N4_10 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end carry_sel_gen_N4_10;

architecture SYN_STRUCTURAL of carry_sel_gen_N4_10 is

   component mux21_SIZE4_10
      port( IN0, IN1 : in std_logic_vector (3 downto 0);  CTRL : in std_logic; 
            OUT1 : out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_N4_19
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_20
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, nocarry_sum_to_mux_3_port, 
      nocarry_sum_to_mux_2_port, nocarry_sum_to_mux_1_port, 
      nocarry_sum_to_mux_0_port, carry_sum_to_mux_3_port, 
      carry_sum_to_mux_2_port, carry_sum_to_mux_1_port, carry_sum_to_mux_0_port
      , net246164, net246165 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   rca_nocarry : RCA_N4_20 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           nocarry_sum_to_mux_3_port, S(2) => 
                           nocarry_sum_to_mux_2_port, S(1) => 
                           nocarry_sum_to_mux_1_port, S(0) => 
                           nocarry_sum_to_mux_0_port, Co => net246165);
   rca_carry : RCA_N4_19 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           carry_sum_to_mux_3_port, S(2) => 
                           carry_sum_to_mux_2_port, S(1) => 
                           carry_sum_to_mux_1_port, S(0) => 
                           carry_sum_to_mux_0_port, Co => net246164);
   outmux : mux21_SIZE4_10 port map( IN0(3) => nocarry_sum_to_mux_3_port, 
                           IN0(2) => nocarry_sum_to_mux_2_port, IN0(1) => 
                           nocarry_sum_to_mux_1_port, IN0(0) => 
                           nocarry_sum_to_mux_0_port, IN1(3) => 
                           carry_sum_to_mux_3_port, IN1(2) => 
                           carry_sum_to_mux_2_port, IN1(1) => 
                           carry_sum_to_mux_1_port, IN1(0) => 
                           carry_sum_to_mux_0_port, CTRL => Ci, OUT1(3) => S(3)
                           , OUT1(2) => S(2), OUT1(1) => S(1), OUT1(0) => S(0))
                           ;

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity carry_sel_gen_N4_9 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end carry_sel_gen_N4_9;

architecture SYN_STRUCTURAL of carry_sel_gen_N4_9 is

   component mux21_SIZE4_9
      port( IN0, IN1 : in std_logic_vector (3 downto 0);  CTRL : in std_logic; 
            OUT1 : out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_N4_17
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_18
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, nocarry_sum_to_mux_3_port, 
      nocarry_sum_to_mux_2_port, nocarry_sum_to_mux_1_port, 
      nocarry_sum_to_mux_0_port, carry_sum_to_mux_3_port, 
      carry_sum_to_mux_2_port, carry_sum_to_mux_1_port, carry_sum_to_mux_0_port
      , net246162, net246163 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   rca_nocarry : RCA_N4_18 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           nocarry_sum_to_mux_3_port, S(2) => 
                           nocarry_sum_to_mux_2_port, S(1) => 
                           nocarry_sum_to_mux_1_port, S(0) => 
                           nocarry_sum_to_mux_0_port, Co => net246163);
   rca_carry : RCA_N4_17 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           carry_sum_to_mux_3_port, S(2) => 
                           carry_sum_to_mux_2_port, S(1) => 
                           carry_sum_to_mux_1_port, S(0) => 
                           carry_sum_to_mux_0_port, Co => net246162);
   outmux : mux21_SIZE4_9 port map( IN0(3) => nocarry_sum_to_mux_3_port, IN0(2)
                           => nocarry_sum_to_mux_2_port, IN0(1) => 
                           nocarry_sum_to_mux_1_port, IN0(0) => 
                           nocarry_sum_to_mux_0_port, IN1(3) => 
                           carry_sum_to_mux_3_port, IN1(2) => 
                           carry_sum_to_mux_2_port, IN1(1) => 
                           carry_sum_to_mux_1_port, IN1(0) => 
                           carry_sum_to_mux_0_port, CTRL => Ci, OUT1(3) => S(3)
                           , OUT1(2) => S(2), OUT1(1) => S(1), OUT1(0) => S(0))
                           ;

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity carry_sel_gen_N4_8 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end carry_sel_gen_N4_8;

architecture SYN_STRUCTURAL of carry_sel_gen_N4_8 is

   component mux21_SIZE4_8
      port( IN0, IN1 : in std_logic_vector (3 downto 0);  CTRL : in std_logic; 
            OUT1 : out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_N4_15
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_16
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, nocarry_sum_to_mux_3_port, 
      nocarry_sum_to_mux_2_port, nocarry_sum_to_mux_1_port, 
      nocarry_sum_to_mux_0_port, carry_sum_to_mux_3_port, 
      carry_sum_to_mux_2_port, carry_sum_to_mux_1_port, carry_sum_to_mux_0_port
      , net246160, net246161 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   rca_nocarry : RCA_N4_16 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           nocarry_sum_to_mux_3_port, S(2) => 
                           nocarry_sum_to_mux_2_port, S(1) => 
                           nocarry_sum_to_mux_1_port, S(0) => 
                           nocarry_sum_to_mux_0_port, Co => net246161);
   rca_carry : RCA_N4_15 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           carry_sum_to_mux_3_port, S(2) => 
                           carry_sum_to_mux_2_port, S(1) => 
                           carry_sum_to_mux_1_port, S(0) => 
                           carry_sum_to_mux_0_port, Co => net246160);
   outmux : mux21_SIZE4_8 port map( IN0(3) => nocarry_sum_to_mux_3_port, IN0(2)
                           => nocarry_sum_to_mux_2_port, IN0(1) => 
                           nocarry_sum_to_mux_1_port, IN0(0) => 
                           nocarry_sum_to_mux_0_port, IN1(3) => 
                           carry_sum_to_mux_3_port, IN1(2) => 
                           carry_sum_to_mux_2_port, IN1(1) => 
                           carry_sum_to_mux_1_port, IN1(0) => 
                           carry_sum_to_mux_0_port, CTRL => Ci, OUT1(3) => S(3)
                           , OUT1(2) => S(2), OUT1(1) => S(1), OUT1(0) => S(0))
                           ;

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity carry_sel_gen_N4_7 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end carry_sel_gen_N4_7;

architecture SYN_STRUCTURAL of carry_sel_gen_N4_7 is

   component mux21_SIZE4_7
      port( IN0, IN1 : in std_logic_vector (3 downto 0);  CTRL : in std_logic; 
            OUT1 : out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_N4_13
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_14
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, nocarry_sum_to_mux_3_port, 
      nocarry_sum_to_mux_2_port, nocarry_sum_to_mux_1_port, 
      nocarry_sum_to_mux_0_port, carry_sum_to_mux_3_port, 
      carry_sum_to_mux_2_port, carry_sum_to_mux_1_port, carry_sum_to_mux_0_port
      , net246158, net246159 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   rca_nocarry : RCA_N4_14 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           nocarry_sum_to_mux_3_port, S(2) => 
                           nocarry_sum_to_mux_2_port, S(1) => 
                           nocarry_sum_to_mux_1_port, S(0) => 
                           nocarry_sum_to_mux_0_port, Co => net246159);
   rca_carry : RCA_N4_13 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           carry_sum_to_mux_3_port, S(2) => 
                           carry_sum_to_mux_2_port, S(1) => 
                           carry_sum_to_mux_1_port, S(0) => 
                           carry_sum_to_mux_0_port, Co => net246158);
   outmux : mux21_SIZE4_7 port map( IN0(3) => nocarry_sum_to_mux_3_port, IN0(2)
                           => nocarry_sum_to_mux_2_port, IN0(1) => 
                           nocarry_sum_to_mux_1_port, IN0(0) => 
                           nocarry_sum_to_mux_0_port, IN1(3) => 
                           carry_sum_to_mux_3_port, IN1(2) => 
                           carry_sum_to_mux_2_port, IN1(1) => 
                           carry_sum_to_mux_1_port, IN1(0) => 
                           carry_sum_to_mux_0_port, CTRL => Ci, OUT1(3) => S(3)
                           , OUT1(2) => S(2), OUT1(1) => S(1), OUT1(0) => S(0))
                           ;

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity carry_sel_gen_N4_6 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end carry_sel_gen_N4_6;

architecture SYN_STRUCTURAL of carry_sel_gen_N4_6 is

   component mux21_SIZE4_6
      port( IN0, IN1 : in std_logic_vector (3 downto 0);  CTRL : in std_logic; 
            OUT1 : out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_N4_11
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_12
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, nocarry_sum_to_mux_3_port, 
      nocarry_sum_to_mux_2_port, nocarry_sum_to_mux_1_port, 
      nocarry_sum_to_mux_0_port, carry_sum_to_mux_3_port, 
      carry_sum_to_mux_2_port, carry_sum_to_mux_1_port, carry_sum_to_mux_0_port
      , net246156, net246157 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   rca_nocarry : RCA_N4_12 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           nocarry_sum_to_mux_3_port, S(2) => 
                           nocarry_sum_to_mux_2_port, S(1) => 
                           nocarry_sum_to_mux_1_port, S(0) => 
                           nocarry_sum_to_mux_0_port, Co => net246157);
   rca_carry : RCA_N4_11 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           carry_sum_to_mux_3_port, S(2) => 
                           carry_sum_to_mux_2_port, S(1) => 
                           carry_sum_to_mux_1_port, S(0) => 
                           carry_sum_to_mux_0_port, Co => net246156);
   outmux : mux21_SIZE4_6 port map( IN0(3) => nocarry_sum_to_mux_3_port, IN0(2)
                           => nocarry_sum_to_mux_2_port, IN0(1) => 
                           nocarry_sum_to_mux_1_port, IN0(0) => 
                           nocarry_sum_to_mux_0_port, IN1(3) => 
                           carry_sum_to_mux_3_port, IN1(2) => 
                           carry_sum_to_mux_2_port, IN1(1) => 
                           carry_sum_to_mux_1_port, IN1(0) => 
                           carry_sum_to_mux_0_port, CTRL => Ci, OUT1(3) => S(3)
                           , OUT1(2) => S(2), OUT1(1) => S(1), OUT1(0) => S(0))
                           ;

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity carry_sel_gen_N4_5 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end carry_sel_gen_N4_5;

architecture SYN_STRUCTURAL of carry_sel_gen_N4_5 is

   component mux21_SIZE4_5
      port( IN0, IN1 : in std_logic_vector (3 downto 0);  CTRL : in std_logic; 
            OUT1 : out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_N4_9
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_10
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, nocarry_sum_to_mux_3_port, 
      nocarry_sum_to_mux_2_port, nocarry_sum_to_mux_1_port, 
      nocarry_sum_to_mux_0_port, carry_sum_to_mux_3_port, 
      carry_sum_to_mux_2_port, carry_sum_to_mux_1_port, carry_sum_to_mux_0_port
      , net246154, net246155 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   rca_nocarry : RCA_N4_10 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           nocarry_sum_to_mux_3_port, S(2) => 
                           nocarry_sum_to_mux_2_port, S(1) => 
                           nocarry_sum_to_mux_1_port, S(0) => 
                           nocarry_sum_to_mux_0_port, Co => net246155);
   rca_carry : RCA_N4_9 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           carry_sum_to_mux_3_port, S(2) => 
                           carry_sum_to_mux_2_port, S(1) => 
                           carry_sum_to_mux_1_port, S(0) => 
                           carry_sum_to_mux_0_port, Co => net246154);
   outmux : mux21_SIZE4_5 port map( IN0(3) => nocarry_sum_to_mux_3_port, IN0(2)
                           => nocarry_sum_to_mux_2_port, IN0(1) => 
                           nocarry_sum_to_mux_1_port, IN0(0) => 
                           nocarry_sum_to_mux_0_port, IN1(3) => 
                           carry_sum_to_mux_3_port, IN1(2) => 
                           carry_sum_to_mux_2_port, IN1(1) => 
                           carry_sum_to_mux_1_port, IN1(0) => 
                           carry_sum_to_mux_0_port, CTRL => Ci, OUT1(3) => S(3)
                           , OUT1(2) => S(2), OUT1(1) => S(1), OUT1(0) => S(0))
                           ;

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity carry_sel_gen_N4_4 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end carry_sel_gen_N4_4;

architecture SYN_STRUCTURAL of carry_sel_gen_N4_4 is

   component mux21_SIZE4_4
      port( IN0, IN1 : in std_logic_vector (3 downto 0);  CTRL : in std_logic; 
            OUT1 : out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_N4_7
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_8
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, nocarry_sum_to_mux_3_port, 
      nocarry_sum_to_mux_2_port, nocarry_sum_to_mux_1_port, 
      nocarry_sum_to_mux_0_port, carry_sum_to_mux_3_port, 
      carry_sum_to_mux_2_port, carry_sum_to_mux_1_port, carry_sum_to_mux_0_port
      , net246152, net246153 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   rca_nocarry : RCA_N4_8 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           nocarry_sum_to_mux_3_port, S(2) => 
                           nocarry_sum_to_mux_2_port, S(1) => 
                           nocarry_sum_to_mux_1_port, S(0) => 
                           nocarry_sum_to_mux_0_port, Co => net246153);
   rca_carry : RCA_N4_7 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           carry_sum_to_mux_3_port, S(2) => 
                           carry_sum_to_mux_2_port, S(1) => 
                           carry_sum_to_mux_1_port, S(0) => 
                           carry_sum_to_mux_0_port, Co => net246152);
   outmux : mux21_SIZE4_4 port map( IN0(3) => nocarry_sum_to_mux_3_port, IN0(2)
                           => nocarry_sum_to_mux_2_port, IN0(1) => 
                           nocarry_sum_to_mux_1_port, IN0(0) => 
                           nocarry_sum_to_mux_0_port, IN1(3) => 
                           carry_sum_to_mux_3_port, IN1(2) => 
                           carry_sum_to_mux_2_port, IN1(1) => 
                           carry_sum_to_mux_1_port, IN1(0) => 
                           carry_sum_to_mux_0_port, CTRL => Ci, OUT1(3) => S(3)
                           , OUT1(2) => S(2), OUT1(1) => S(1), OUT1(0) => S(0))
                           ;

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity carry_sel_gen_N4_3 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end carry_sel_gen_N4_3;

architecture SYN_STRUCTURAL of carry_sel_gen_N4_3 is

   component mux21_SIZE4_3
      port( IN0, IN1 : in std_logic_vector (3 downto 0);  CTRL : in std_logic; 
            OUT1 : out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_N4_5
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_6
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, nocarry_sum_to_mux_3_port, 
      nocarry_sum_to_mux_2_port, nocarry_sum_to_mux_1_port, 
      nocarry_sum_to_mux_0_port, carry_sum_to_mux_3_port, 
      carry_sum_to_mux_2_port, carry_sum_to_mux_1_port, carry_sum_to_mux_0_port
      , net246150, net246151 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   rca_nocarry : RCA_N4_6 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           nocarry_sum_to_mux_3_port, S(2) => 
                           nocarry_sum_to_mux_2_port, S(1) => 
                           nocarry_sum_to_mux_1_port, S(0) => 
                           nocarry_sum_to_mux_0_port, Co => net246151);
   rca_carry : RCA_N4_5 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           carry_sum_to_mux_3_port, S(2) => 
                           carry_sum_to_mux_2_port, S(1) => 
                           carry_sum_to_mux_1_port, S(0) => 
                           carry_sum_to_mux_0_port, Co => net246150);
   outmux : mux21_SIZE4_3 port map( IN0(3) => nocarry_sum_to_mux_3_port, IN0(2)
                           => nocarry_sum_to_mux_2_port, IN0(1) => 
                           nocarry_sum_to_mux_1_port, IN0(0) => 
                           nocarry_sum_to_mux_0_port, IN1(3) => 
                           carry_sum_to_mux_3_port, IN1(2) => 
                           carry_sum_to_mux_2_port, IN1(1) => 
                           carry_sum_to_mux_1_port, IN1(0) => 
                           carry_sum_to_mux_0_port, CTRL => Ci, OUT1(3) => S(3)
                           , OUT1(2) => S(2), OUT1(1) => S(1), OUT1(0) => S(0))
                           ;

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity carry_sel_gen_N4_2 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end carry_sel_gen_N4_2;

architecture SYN_STRUCTURAL of carry_sel_gen_N4_2 is

   component mux21_SIZE4_2
      port( IN0, IN1 : in std_logic_vector (3 downto 0);  CTRL : in std_logic; 
            OUT1 : out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_N4_3
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_4
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, nocarry_sum_to_mux_3_port, 
      nocarry_sum_to_mux_2_port, nocarry_sum_to_mux_1_port, 
      nocarry_sum_to_mux_0_port, carry_sum_to_mux_3_port, 
      carry_sum_to_mux_2_port, carry_sum_to_mux_1_port, carry_sum_to_mux_0_port
      , net246148, net246149 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   rca_nocarry : RCA_N4_4 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           nocarry_sum_to_mux_3_port, S(2) => 
                           nocarry_sum_to_mux_2_port, S(1) => 
                           nocarry_sum_to_mux_1_port, S(0) => 
                           nocarry_sum_to_mux_0_port, Co => net246149);
   rca_carry : RCA_N4_3 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           carry_sum_to_mux_3_port, S(2) => 
                           carry_sum_to_mux_2_port, S(1) => 
                           carry_sum_to_mux_1_port, S(0) => 
                           carry_sum_to_mux_0_port, Co => net246148);
   outmux : mux21_SIZE4_2 port map( IN0(3) => nocarry_sum_to_mux_3_port, IN0(2)
                           => nocarry_sum_to_mux_2_port, IN0(1) => 
                           nocarry_sum_to_mux_1_port, IN0(0) => 
                           nocarry_sum_to_mux_0_port, IN1(3) => 
                           carry_sum_to_mux_3_port, IN1(2) => 
                           carry_sum_to_mux_2_port, IN1(1) => 
                           carry_sum_to_mux_1_port, IN1(0) => 
                           carry_sum_to_mux_0_port, CTRL => Ci, OUT1(3) => S(3)
                           , OUT1(2) => S(2), OUT1(1) => S(1), OUT1(0) => S(0))
                           ;

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity carry_sel_gen_N4_1 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end carry_sel_gen_N4_1;

architecture SYN_STRUCTURAL of carry_sel_gen_N4_1 is

   component mux21_SIZE4_1
      port( IN0, IN1 : in std_logic_vector (3 downto 0);  CTRL : in std_logic; 
            OUT1 : out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_N4_1
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_2
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, nocarry_sum_to_mux_3_port, 
      nocarry_sum_to_mux_2_port, nocarry_sum_to_mux_1_port, 
      nocarry_sum_to_mux_0_port, carry_sum_to_mux_3_port, 
      carry_sum_to_mux_2_port, carry_sum_to_mux_1_port, carry_sum_to_mux_0_port
      , net246146, net246147 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   rca_nocarry : RCA_N4_2 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           nocarry_sum_to_mux_3_port, S(2) => 
                           nocarry_sum_to_mux_2_port, S(1) => 
                           nocarry_sum_to_mux_1_port, S(0) => 
                           nocarry_sum_to_mux_0_port, Co => net246147);
   rca_carry : RCA_N4_1 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           carry_sum_to_mux_3_port, S(2) => 
                           carry_sum_to_mux_2_port, S(1) => 
                           carry_sum_to_mux_1_port, S(0) => 
                           carry_sum_to_mux_0_port, Co => net246146);
   outmux : mux21_SIZE4_1 port map( IN0(3) => nocarry_sum_to_mux_3_port, IN0(2)
                           => nocarry_sum_to_mux_2_port, IN0(1) => 
                           nocarry_sum_to_mux_1_port, IN0(0) => 
                           nocarry_sum_to_mux_0_port, IN1(3) => 
                           carry_sum_to_mux_3_port, IN1(2) => 
                           carry_sum_to_mux_2_port, IN1(1) => 
                           carry_sum_to_mux_1_port, IN1(0) => 
                           carry_sum_to_mux_0_port, CTRL => Ci, OUT1(3) => S(3)
                           , OUT1(2) => S(2), OUT1(1) => S(1), OUT1(0) => S(0))
                           ;

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_53 is

   port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic);

end pg_53;

architecture SYN_beh of pg_53 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U3 : AOI21_X1 port map( B1 => g_prec, B2 => p, A => g, ZN => n1);
   U1 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);
   U2 : INV_X1 port map( A => n1, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_52 is

   port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic);

end pg_52;

architecture SYN_beh of pg_52 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U3 : AOI21_X1 port map( B1 => g_prec, B2 => p, A => g, ZN => n1);
   U1 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);
   U2 : INV_X1 port map( A => n1, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_51 is

   port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic);

end pg_51;

architecture SYN_beh of pg_51 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U3 : AOI21_X1 port map( B1 => g_prec, B2 => p, A => g, ZN => n1);
   U1 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);
   U2 : INV_X1 port map( A => n1, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_50 is

   port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic);

end pg_50;

architecture SYN_beh of pg_50 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U3 : AOI21_X1 port map( B1 => g_prec, B2 => p, A => g, ZN => n1);
   U1 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);
   U2 : INV_X1 port map( A => n1, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_49 is

   port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic);

end pg_49;

architecture SYN_beh of pg_49 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U3 : AOI21_X1 port map( B1 => g_prec, B2 => p, A => g, ZN => n1);
   U1 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);
   U2 : INV_X1 port map( A => n1, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_48 is

   port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic);

end pg_48;

architecture SYN_beh of pg_48 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U3 : AOI21_X1 port map( B1 => g_prec, B2 => p, A => g, ZN => n1);
   U1 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);
   U2 : INV_X1 port map( A => n1, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_47 is

   port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic);

end pg_47;

architecture SYN_beh of pg_47 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);
   U2 : INV_X1 port map( A => g, ZN => n2);
   U3 : NAND2_X1 port map( A1 => g_prec, A2 => p, ZN => n1);
   U4 : NAND2_X1 port map( A1 => n1, A2 => n2, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_46 is

   port( g, p, g_prec, p_prec : in std_logic;  p_out, g_out_BAR : out std_logic
         );

end pg_46;

architecture SYN_beh of pg_46 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);
   U2 : AOI21_X1 port map( B1 => g_prec, B2 => p, A => g, ZN => g_out_BAR);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_45 is

   port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic);

end pg_45;

architecture SYN_beh of pg_45 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => g, ZN => n2);
   U2 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);
   U3 : NAND2_X1 port map( A1 => p, A2 => g_prec, ZN => n1);
   U4 : NAND2_X1 port map( A1 => n1, A2 => n2, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_44 is

   port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic);

end pg_44;

architecture SYN_beh of pg_44 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => p, B2 => g_prec, A => g, ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => g_out);
   U3 : AND2_X1 port map( A1 => p_prec, A2 => p, ZN => p_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_43 is

   port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic);

end pg_43;

architecture SYN_beh of pg_43 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => g_out);
   U2 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);
   U3 : AOI21_X1 port map( B1 => g_prec, B2 => p, A => g, ZN => n1);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_42 is

   port( g, p, g_prec, p_prec : in std_logic;  p_out, g_out_BAR : out std_logic
         );

end pg_42;

architecture SYN_beh of pg_42 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);
   U2 : AOI21_X1 port map( B1 => p, B2 => g_prec, A => g, ZN => g_out_BAR);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_39 is

   port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic);

end pg_39;

architecture SYN_beh of pg_39 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U3 : AOI21_X1 port map( B1 => g_prec, B2 => p, A => g, ZN => n1);
   U1 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);
   U2 : INV_X1 port map( A => n1, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_38 is

   port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic);

end pg_38;

architecture SYN_beh of pg_38 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U3 : AOI21_X1 port map( B1 => g_prec, B2 => p, A => g, ZN => n1);
   U1 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);
   U2 : INV_X1 port map( A => n1, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_37 is

   port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic);

end pg_37;

architecture SYN_beh of pg_37 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U3 : AOI21_X1 port map( B1 => g_prec, B2 => p, A => g, ZN => n1);
   U1 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);
   U2 : INV_X1 port map( A => n1, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_36 is

   port( p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic;  
         g_BAR : in std_logic);

end pg_36;

architecture SYN_beh of pg_36 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);
   U2 : NAND2_X1 port map( A1 => n1, A2 => g_BAR, ZN => g_out);
   U3 : NAND2_X1 port map( A1 => g_prec, A2 => p, ZN => n1);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_35 is

   port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic);

end pg_35;

architecture SYN_beh of pg_35 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);
   U2 : INV_X1 port map( A => g, ZN => n2);
   U3 : NAND2_X1 port map( A1 => g_prec, A2 => p, ZN => n1);
   U4 : NAND2_X1 port map( A1 => n1, A2 => n2, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_34 is

   port( p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic;  
         g_BAR : in std_logic);

end pg_34;

architecture SYN_beh of pg_34 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);
   U2 : NAND2_X1 port map( A1 => g_BAR, A2 => n1, ZN => g_out);
   U3 : NAND2_X1 port map( A1 => g_prec, A2 => p, ZN => n1);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_32 is

   port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic);

end pg_32;

architecture SYN_beh of pg_32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U3 : AOI21_X1 port map( B1 => g_prec, B2 => p, A => g, ZN => n1);
   U1 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);
   U2 : INV_X1 port map( A => n1, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_31 is

   port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic);

end pg_31;

architecture SYN_beh of pg_31 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);
   U2 : INV_X1 port map( A => n1, ZN => g_out);
   U3 : AOI21_X1 port map( B1 => g_prec, B2 => p, A => g, ZN => n1);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_29 is

   port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic);

end pg_29;

architecture SYN_beh of pg_29 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);
   U2 : INV_X1 port map( A => g, ZN => n2);
   U3 : NAND2_X1 port map( A1 => g_prec, A2 => p, ZN => n1);
   U4 : NAND2_X1 port map( A1 => n1, A2 => n2, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_27 is

   port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic);

end pg_27;

architecture SYN_beh of pg_27 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => g, ZN => n2);
   U2 : AND2_X1 port map( A1 => p_prec, A2 => p, ZN => p_out);
   U3 : NAND2_X1 port map( A1 => p, A2 => g_prec, ZN => n1);
   U4 : NAND2_X1 port map( A1 => n1, A2 => n2, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_26 is

   port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic);

end pg_26;

architecture SYN_beh of pg_26 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);
   U2 : INV_X1 port map( A => n1, ZN => g_out);
   U3 : AOI21_X1 port map( B1 => g_prec, B2 => p, A => g, ZN => n1);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_25 is

   port( g, p, g_prec, p_prec : in std_logic;  p_out, g_out_BAR : out std_logic
         );

end pg_25;

architecture SYN_beh of pg_25 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);
   U2 : AOI21_X1 port map( B1 => g_prec, B2 => p, A => g, ZN => g_out_BAR);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_24 is

   port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic);

end pg_24;

architecture SYN_beh of pg_24 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => g, ZN => n2);
   U2 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);
   U3 : NAND2_X1 port map( A1 => g_prec, A2 => p, ZN => n1);
   U4 : NAND2_X1 port map( A1 => n1, A2 => n2, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_23 is

   port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic);

end pg_23;

architecture SYN_beh of pg_23 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => g_out);
   U2 : AND2_X1 port map( A1 => p_prec, A2 => p, ZN => p_out);
   U3 : AOI21_X1 port map( B1 => g_prec, B2 => p, A => g, ZN => n1);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_22 is

   port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic);

end pg_22;

architecture SYN_beh of pg_22 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p_prec, A2 => p, ZN => p_out);
   U2 : INV_X1 port map( A => n1, ZN => g_out);
   U3 : AOI21_X1 port map( B1 => g_prec, B2 => p, A => g, ZN => n1);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_21 is

   port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic);

end pg_21;

architecture SYN_beh of pg_21 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => g_prec, B2 => p, A => g, ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => g_out);
   U3 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_20 is

   port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic);

end pg_20;

architecture SYN_beh of pg_20 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);
   U2 : INV_X1 port map( A => n1, ZN => g_out);
   U3 : AOI21_X1 port map( B1 => g_prec, B2 => p, A => g, ZN => n1);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_19 is

   port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic);

end pg_19;

architecture SYN_beh of pg_19 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U3 : AOI21_X1 port map( B1 => g_prec, B2 => p, A => g, ZN => n1);
   U1 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);
   U2 : INV_X1 port map( A => n1, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_18 is

   port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic);

end pg_18;

architecture SYN_beh of pg_18 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U3 : AOI21_X1 port map( B1 => g_prec, B2 => p, A => g, ZN => n1);
   U1 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);
   U2 : INV_X1 port map( A => n1, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_17 is

   port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic);

end pg_17;

architecture SYN_beh of pg_17 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => g_out);
   U2 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);
   U3 : AOI21_X1 port map( B1 => g_prec, B2 => p, A => g, ZN => n1);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_16 is

   port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic);

end pg_16;

architecture SYN_beh of pg_16 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => g_out);
   U2 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);
   U3 : AOI21_X1 port map( B1 => g_prec, B2 => p, A => g, ZN => n1);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_15 is

   port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic);

end pg_15;

architecture SYN_beh of pg_15 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U3 : AOI21_X1 port map( B1 => g_prec, B2 => p, A => g, ZN => n1);
   U1 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);
   U2 : INV_X1 port map( A => n1, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_14 is

   port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic);

end pg_14;

architecture SYN_beh of pg_14 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U3 : AOI21_X1 port map( B1 => g_prec, B2 => p, A => g, ZN => n1);
   U1 : INV_X1 port map( A => n1, ZN => g_out);
   U2 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_13 is

   port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic);

end pg_13;

architecture SYN_beh of pg_13 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => g_prec, B2 => p, A => g, ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => g_out);
   U3 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_12 is

   port( p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic;  
         g_BAR : in std_logic);

end pg_12;

architecture SYN_beh of pg_12 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);
   U2 : NAND2_X1 port map( A1 => g_prec, A2 => p, ZN => n1);
   U3 : NAND2_X1 port map( A1 => n1, A2 => g_BAR, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_11 is

   port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic);

end pg_11;

architecture SYN_beh of pg_11 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);
   U2 : INV_X1 port map( A => n1, ZN => g_out);
   U3 : AOI21_X1 port map( B1 => g_prec, B2 => p, A => g, ZN => n1);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_10 is

   port( g, p, g_prec, p_prec : in std_logic;  p_out, g_out_BAR : out std_logic
         );

end pg_10;

architecture SYN_beh of pg_10 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p_prec, A2 => p, ZN => p_out);
   U2 : AOI21_X1 port map( B1 => g_prec, B2 => p, A => g, ZN => g_out_BAR);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_9 is

   port( g, p, g_prec, p_prec : in std_logic;  p_out, g_out_BAR : out std_logic
         );

end pg_9;

architecture SYN_beh of pg_9 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U3 : AOI21_X1 port map( B1 => g_prec, B2 => p, A => g, ZN => g_out_BAR);
   U1 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_8 is

   port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic);

end pg_8;

architecture SYN_beh of pg_8 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);
   U2 : INV_X1 port map( A => n1, ZN => g_out);
   U3 : AOI21_X1 port map( B1 => g_prec, B2 => p, A => g, ZN => n1);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_7 is

   port( g, p, g_prec, p_prec : in std_logic;  p_out, g_out_BAR : out std_logic
         );

end pg_7;

architecture SYN_beh of pg_7 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U3 : AOI21_X1 port map( B1 => g_prec, B2 => p, A => g, ZN => g_out_BAR);
   U1 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_6 is

   port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic);

end pg_6;

architecture SYN_beh of pg_6 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => g_prec, B2 => p, A => g, ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => g_out);
   U3 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_5 is

   port( p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic;  
         g_BAR : in std_logic);

end pg_5;

architecture SYN_beh of pg_5 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);
   U2 : NAND2_X1 port map( A1 => g_prec, A2 => p, ZN => n1);
   U3 : NAND2_X1 port map( A1 => n1, A2 => g_BAR, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_4 is

   port( g, p, p_prec : in std_logic;  g_out, p_out : out std_logic;  
         g_prec_BAR : in std_logic);

end pg_4;

architecture SYN_beh of pg_4 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);
   U2 : INV_X1 port map( A => g_prec_BAR, ZN => n1);
   U3 : INV_X1 port map( A => n3, ZN => g_out);
   U4 : AOI21_X1 port map( B1 => n1, B2 => p, A => g, ZN => n3);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_3 is

   port( g, p, p_prec : in std_logic;  g_out, p_out : out std_logic;  
         g_prec_BAR : in std_logic);

end pg_3;

architecture SYN_beh of pg_3 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : OAI21_X1 port map( B1 => g_prec_BAR, B2 => n1, A => n2, ZN => g_out);
   U2 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);
   U3 : INV_X1 port map( A => p, ZN => n1);
   U4 : INV_X1 port map( A => g, ZN => n2);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_2 is

   port( p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic;  
         g_BAR : in std_logic);

end pg_2;

architecture SYN_beh of pg_2 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);
   U2 : NAND2_X1 port map( A1 => g_prec, A2 => p, ZN => n1);
   U3 : NAND2_X1 port map( A1 => n1, A2 => g_BAR, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_1 is

   port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic);

end pg_1;

architecture SYN_beh of pg_1 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => g_prec, B2 => p, A => g, ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => g_out);
   U3 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity g_19 is

   port( g, p, g_prec : in std_logic;  g_out : out std_logic);

end g_19;

architecture SYN_beh of g_19 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U2 : AOI21_X1 port map( B1 => p, B2 => g_prec, A => g, ZN => n1);
   U1 : INV_X1 port map( A => n1, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity g_18 is

   port( g, p, g_prec : in std_logic;  g_out : out std_logic);

end g_18;

architecture SYN_beh of g_18 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U2 : AOI21_X1 port map( B1 => p, B2 => g_prec, A => g, ZN => n1);
   U1 : INV_X1 port map( A => n1, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity g_17 is

   port( g, p, g_prec : in std_logic;  g_out : out std_logic);

end g_17;

architecture SYN_beh of g_17 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U2 : AOI21_X1 port map( B1 => p, B2 => g_prec, A => g, ZN => n1);
   U1 : INV_X1 port map( A => n1, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity g_16 is

   port( g, p, g_prec : in std_logic;  g_out : out std_logic);

end g_16;

architecture SYN_beh of g_16 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U2 : AOI21_X1 port map( B1 => p, B2 => g_prec, A => g, ZN => n1);
   U1 : INV_X1 port map( A => n1, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity g_15 is

   port( g, p, g_prec : in std_logic;  g_out : out std_logic);

end g_15;

architecture SYN_beh of g_15 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U2 : AOI21_X1 port map( B1 => p, B2 => g_prec, A => g, ZN => n1);
   U1 : INV_X1 port map( A => n1, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity g_14 is

   port( g, p, g_prec : in std_logic;  g_out : out std_logic);

end g_14;

architecture SYN_beh of g_14 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => g_out);
   U2 : AOI21_X1 port map( B1 => p, B2 => g_prec, A => g, ZN => n1);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity g_13 is

   port( g, p, g_prec : in std_logic;  g_out : out std_logic);

end g_13;

architecture SYN_beh of g_13 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => p, B2 => g_prec, A => g, ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity g_12 is

   port( g, p, g_prec : in std_logic;  g_out : out std_logic);

end g_12;

architecture SYN_beh of g_12 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : OR2_X1 port map( A1 => g, A2 => n1, ZN => g_out);
   U2 : AND2_X1 port map( A1 => p, A2 => g_prec, ZN => n1);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity g_10 is

   port( g, p, g_prec : in std_logic;  g_out : out std_logic);

end g_10;

architecture SYN_beh of g_10 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => g, ZN => n2);
   U2 : NAND2_X1 port map( A1 => n1, A2 => n2, ZN => g_out);
   U3 : NAND2_X1 port map( A1 => p, A2 => g_prec, ZN => n1);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity g_9 is

   port( g, p, g_prec : in std_logic;  g_out : out std_logic);

end g_9;

architecture SYN_beh of g_9 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => g, ZN => n2);
   U2 : NAND2_X1 port map( A1 => n1, A2 => n2, ZN => g_out);
   U3 : NAND2_X1 port map( A1 => g_prec, A2 => p, ZN => n1);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity g_8 is

   port( g, p, g_prec : in std_logic;  g_out : out std_logic);

end g_8;

architecture SYN_beh of g_8 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X2 port map( A => n1, ZN => g_out);
   U2 : AOI21_X1 port map( B1 => g_prec, B2 => p, A => g, ZN => n1);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity g_7 is

   port( g, p, g_prec : in std_logic;  g_out : out std_logic);

end g_7;

architecture SYN_beh of g_7 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => g_out);
   U2 : AOI21_X1 port map( B1 => g_prec, B2 => p, A => g, ZN => n1);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity g_6 is

   port( g, p, g_prec : in std_logic;  g_out : out std_logic);

end g_6;

architecture SYN_beh of g_6 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => g_out);
   U2 : AOI21_X1 port map( B1 => p, B2 => g_prec, A => g, ZN => n1);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity g_5 is

   port( g, p, g_prec : in std_logic;  g_out : out std_logic);

end g_5;

architecture SYN_beh of g_5 is

   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => p, B2 => g_prec, A => g, ZN => n1);
   U2 : INV_X2 port map( A => n1, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity g_4 is

   port( p, g_prec : in std_logic;  g_out : out std_logic;  g_BAR : in 
         std_logic);

end g_4;

architecture SYN_beh of g_4 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n1, A2 => g_BAR, ZN => g_out);
   U2 : NAND2_X1 port map( A1 => g_prec, A2 => p, ZN => n1);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity g_3 is

   port( g, p, g_prec : in std_logic;  g_out : out std_logic);

end g_3;

architecture SYN_beh of g_3 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => g_out);
   U2 : AOI21_X1 port map( B1 => p, B2 => g_prec, A => g, ZN => n1);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity g_2 is

   port( g, p, g_prec : in std_logic;  g_out : out std_logic);

end g_2;

architecture SYN_beh of g_2 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => g_out);
   U2 : AOI21_X1 port map( B1 => g_prec, B2 => p, A => g, ZN => n1);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity g_1 is

   port( g, p, g_prec : in std_logic;  g_out : out std_logic);

end g_1;

architecture SYN_beh of g_1 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => p, B2 => g_prec, A => g, ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_63 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_63;

architecture SYN_beh of pg_net_63 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_62 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_62;

architecture SYN_beh of pg_net_62 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_61 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_61;

architecture SYN_beh of pg_net_61 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_60 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_60;

architecture SYN_beh of pg_net_60 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_59 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_59;

architecture SYN_beh of pg_net_59 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_58 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_58;

architecture SYN_beh of pg_net_58 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_57 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_57;

architecture SYN_beh of pg_net_57 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_56 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_56;

architecture SYN_beh of pg_net_56 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_55 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_55;

architecture SYN_beh of pg_net_55 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_54 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_54;

architecture SYN_beh of pg_net_54 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_53 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_53;

architecture SYN_beh of pg_net_53 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_52 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_52;

architecture SYN_beh of pg_net_52 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_51 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_51;

architecture SYN_beh of pg_net_51 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_50 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_50;

architecture SYN_beh of pg_net_50 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_49 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_49;

architecture SYN_beh of pg_net_49 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_48 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_48;

architecture SYN_beh of pg_net_48 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_47 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_47;

architecture SYN_beh of pg_net_47 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_46 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_46;

architecture SYN_beh of pg_net_46 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_45 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_45;

architecture SYN_beh of pg_net_45 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_44 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_44;

architecture SYN_beh of pg_net_44 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => a, ZN => n1);
   U2 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);
   U3 : XNOR2_X1 port map( A => b, B => n1, ZN => p_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_43 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_43;

architecture SYN_beh of pg_net_43 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_42 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_42;

architecture SYN_beh of pg_net_42 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_41 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_41;

architecture SYN_beh of pg_net_41 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_40 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_40;

architecture SYN_beh of pg_net_40 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_39 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_39;

architecture SYN_beh of pg_net_39 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_38 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_38;

architecture SYN_beh of pg_net_38 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U2 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_33 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_33;

architecture SYN_beh of pg_net_33 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_32 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_32;

architecture SYN_beh of pg_net_32 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_31 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_31;

architecture SYN_beh of pg_net_31 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_30 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_30;

architecture SYN_beh of pg_net_30 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_29 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_29;

architecture SYN_beh of pg_net_29 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_28 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_28;

architecture SYN_beh of pg_net_28 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_27 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_27;

architecture SYN_beh of pg_net_27 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_26 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_26;

architecture SYN_beh of pg_net_26 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_25 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_25;

architecture SYN_beh of pg_net_25 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_24 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_24;

architecture SYN_beh of pg_net_24 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_23 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_23;

architecture SYN_beh of pg_net_23 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_22 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_22;

architecture SYN_beh of pg_net_22 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_21 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_21;

architecture SYN_beh of pg_net_21 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U2 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_20 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_20;

architecture SYN_beh of pg_net_20 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_19 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_19;

architecture SYN_beh of pg_net_19 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_18 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_18;

architecture SYN_beh of pg_net_18 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_17 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_17;

architecture SYN_beh of pg_net_17 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_16 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_16;

architecture SYN_beh of pg_net_16 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_15 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_15;

architecture SYN_beh of pg_net_15 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_14 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_14;

architecture SYN_beh of pg_net_14 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_13 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_13;

architecture SYN_beh of pg_net_13 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_12 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_12;

architecture SYN_beh of pg_net_12 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_11 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_11;

architecture SYN_beh of pg_net_11 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_10 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_10;

architecture SYN_beh of pg_net_10 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_9 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_9;

architecture SYN_beh of pg_net_9 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_8 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_8;

architecture SYN_beh of pg_net_8 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_7 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_7;

architecture SYN_beh of pg_net_7 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_6 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_6;

architecture SYN_beh of pg_net_6 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_5 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_5;

architecture SYN_beh of pg_net_5 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_4 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_4;

architecture SYN_beh of pg_net_4 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_3 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_3;

architecture SYN_beh of pg_net_3 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_2 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_2;

architecture SYN_beh of pg_net_2 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_1 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_1;

architecture SYN_beh of pg_net_1 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);
   U2 : INV_X1 port map( A => a, ZN => n1);
   U3 : XNOR2_X1 port map( A => b, B => n1, ZN => p_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity sum_gen_N32_1 is

   port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic_vector 
         (8 downto 0);  S : out std_logic_vector (31 downto 0));

end sum_gen_N32_1;

architecture SYN_STRUCTURAL of sum_gen_N32_1 is

   component carry_sel_gen_N4_1
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component carry_sel_gen_N4_2
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component carry_sel_gen_N4_3
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component carry_sel_gen_N4_4
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component carry_sel_gen_N4_5
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component carry_sel_gen_N4_6
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component carry_sel_gen_N4_7
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component carry_sel_gen_N4_8
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal net199157, net199158, net199159, net199160, net199161, net199162, 
      net199163, net199164 : std_logic;

begin
   
   csel_N_0 : carry_sel_gen_N4_8 port map( A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), Ci => Cin(0), S(3) => S(3), 
                           S(2) => S(2), S(1) => S(1), S(0) => S(0), Co => 
                           net199164);
   csel_N_1 : carry_sel_gen_N4_7 port map( A(3) => A(7), A(2) => A(6), A(1) => 
                           A(5), A(0) => A(4), B(3) => B(7), B(2) => B(6), B(1)
                           => B(5), B(0) => B(4), Ci => Cin(1), S(3) => S(7), 
                           S(2) => S(6), S(1) => S(5), S(0) => S(4), Co => 
                           net199163);
   csel_N_2 : carry_sel_gen_N4_6 port map( A(3) => A(11), A(2) => A(10), A(1) 
                           => A(9), A(0) => A(8), B(3) => B(11), B(2) => B(10),
                           B(1) => B(9), B(0) => B(8), Ci => Cin(2), S(3) => 
                           S(11), S(2) => S(10), S(1) => S(9), S(0) => S(8), Co
                           => net199162);
   csel_N_3 : carry_sel_gen_N4_5 port map( A(3) => A(15), A(2) => A(14), A(1) 
                           => A(13), A(0) => A(12), B(3) => B(15), B(2) => 
                           B(14), B(1) => B(13), B(0) => B(12), Ci => Cin(3), 
                           S(3) => S(15), S(2) => S(14), S(1) => S(13), S(0) =>
                           S(12), Co => net199161);
   csel_N_4 : carry_sel_gen_N4_4 port map( A(3) => A(19), A(2) => A(18), A(1) 
                           => A(17), A(0) => A(16), B(3) => B(19), B(2) => 
                           B(18), B(1) => B(17), B(0) => B(16), Ci => Cin(4), 
                           S(3) => S(19), S(2) => S(18), S(1) => S(17), S(0) =>
                           S(16), Co => net199160);
   csel_N_5 : carry_sel_gen_N4_3 port map( A(3) => A(23), A(2) => A(22), A(1) 
                           => A(21), A(0) => A(20), B(3) => B(23), B(2) => 
                           B(22), B(1) => B(21), B(0) => B(20), Ci => Cin(5), 
                           S(3) => S(23), S(2) => S(22), S(1) => S(21), S(0) =>
                           S(20), Co => net199159);
   csel_N_6 : carry_sel_gen_N4_2 port map( A(3) => A(27), A(2) => A(26), A(1) 
                           => A(25), A(0) => A(24), B(3) => B(27), B(2) => 
                           B(26), B(1) => B(25), B(0) => B(24), Ci => Cin(6), 
                           S(3) => S(27), S(2) => S(26), S(1) => S(25), S(0) =>
                           S(24), Co => net199158);
   csel_N_7 : carry_sel_gen_N4_1 port map( A(3) => A(31), A(2) => A(30), A(1) 
                           => A(29), A(0) => A(28), B(3) => B(31), B(2) => 
                           B(30), B(1) => B(29), B(0) => B(28), Ci => Cin(7), 
                           S(3) => S(31), S(2) => S(30), S(1) => S(29), S(0) =>
                           S(28), Co => net199157);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity carry_tree_N32_logN5_1 is

   port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  Cout :
         out std_logic_vector (7 downto 0));

end carry_tree_N32_logN5_1;

architecture SYN_arch of carry_tree_N32_logN5_1 is

   component pg_1
      port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic
            );
   end component;
   
   component pg_2
      port( p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic;  
            g_BAR : in std_logic);
   end component;
   
   component pg_3
      port( g, p, p_prec : in std_logic;  g_out, p_out : out std_logic;  
            g_prec_BAR : in std_logic);
   end component;
   
   component pg_4
      port( g, p, p_prec : in std_logic;  g_out, p_out : out std_logic;  
            g_prec_BAR : in std_logic);
   end component;
   
   component pg_5
      port( p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic;  
            g_BAR : in std_logic);
   end component;
   
   component g_1
      port( g, p, g_prec : in std_logic;  g_out : out std_logic);
   end component;
   
   component g_2
      port( g, p, g_prec : in std_logic;  g_out : out std_logic);
   end component;
   
   component g_3
      port( g, p, g_prec : in std_logic;  g_out : out std_logic);
   end component;
   
   component g_4
      port( p, g_prec : in std_logic;  g_out : out std_logic;  g_BAR : in 
            std_logic);
   end component;
   
   component g_5
      port( g, p, g_prec : in std_logic;  g_out : out std_logic);
   end component;
   
   component g_6
      port( g, p, g_prec : in std_logic;  g_out : out std_logic);
   end component;
   
   component g_7
      port( g, p, g_prec : in std_logic;  g_out : out std_logic);
   end component;
   
   component pg_6
      port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic
            );
   end component;
   
   component pg_7
      port( g, p, g_prec, p_prec : in std_logic;  p_out, g_out_BAR : out 
            std_logic);
   end component;
   
   component pg_8
      port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic
            );
   end component;
   
   component pg_9
      port( g, p, g_prec, p_prec : in std_logic;  p_out, g_out_BAR : out 
            std_logic);
   end component;
   
   component pg_10
      port( g, p, g_prec, p_prec : in std_logic;  p_out, g_out_BAR : out 
            std_logic);
   end component;
   
   component pg_11
      port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic
            );
   end component;
   
   component pg_12
      port( p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic;  
            g_BAR : in std_logic);
   end component;
   
   component g_8
      port( g, p, g_prec : in std_logic;  g_out : out std_logic);
   end component;
   
   component pg_13
      port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic
            );
   end component;
   
   component pg_14
      port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic
            );
   end component;
   
   component pg_15
      port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic
            );
   end component;
   
   component pg_16
      port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic
            );
   end component;
   
   component pg_17
      port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic
            );
   end component;
   
   component pg_18
      port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic
            );
   end component;
   
   component pg_19
      port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic
            );
   end component;
   
   component pg_20
      port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic
            );
   end component;
   
   component pg_21
      port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic
            );
   end component;
   
   component pg_22
      port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic
            );
   end component;
   
   component pg_23
      port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic
            );
   end component;
   
   component pg_24
      port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic
            );
   end component;
   
   component pg_25
      port( g, p, g_prec, p_prec : in std_logic;  p_out, g_out_BAR : out 
            std_logic);
   end component;
   
   component pg_26
      port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic
            );
   end component;
   
   component pg_27
      port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic
            );
   end component;
   
   component g_9
      port( g, p, g_prec : in std_logic;  g_out : out std_logic);
   end component;
   
   component g_10
      port( g, p, g_prec : in std_logic;  g_out : out std_logic);
   end component;
   
   component pg_net_1
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_2
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_3
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_4
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_5
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_6
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_7
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_8
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_9
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_10
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_11
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_12
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_13
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_14
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_15
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_16
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_17
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_18
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_19
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_20
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_21
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_22
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_23
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_24
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_25
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_26
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_27
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_28
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_29
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_30
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_31
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_32
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   signal Cout_7_port, Cout_6_port, Cout_5_port, Cout_4_port, Cout_3_port, 
      Cout_2_port, Cout_1_port, Cout_0_port, p_net_31_port, p_net_30_port, 
      p_net_29_port, p_net_28_port, p_net_27_port, p_net_26_port, p_net_25_port
      , p_net_24_port, p_net_23_port, p_net_22_port, p_net_21_port, 
      p_net_20_port, p_net_19_port, p_net_18_port, p_net_17_port, p_net_16_port
      , p_net_15_port, p_net_14_port, p_net_13_port, p_net_12_port, 
      p_net_11_port, p_net_10_port, p_net_9_port, p_net_8_port, p_net_7_port, 
      p_net_6_port, p_net_5_port, p_net_4_port, p_net_3_port, p_net_2_port, 
      p_net_1_port, g_net_31_port, g_net_30_port, g_net_29_port, g_net_28_port,
      g_net_27_port, g_net_26_port, g_net_25_port, g_net_24_port, g_net_23_port
      , g_net_22_port, g_net_21_port, g_net_20_port, g_net_19_port, 
      g_net_18_port, g_net_17_port, g_net_16_port, g_net_15_port, g_net_14_port
      , g_net_13_port, g_net_12_port, g_net_11_port, g_net_10_port, 
      g_net_9_port, g_net_8_port, g_net_7_port, g_net_6_port, g_net_5_port, 
      g_net_4_port, g_net_3_port, g_net_2_port, g_net_1_port, g_net_0_port, 
      magic_pro_1_port, magic_pro_0_port, pg_1_15_1_port, pg_1_15_0_port, 
      pg_1_14_1_port, pg_1_14_0_port, pg_1_13_1_port, pg_1_13_0_port, 
      pg_1_12_1_port, pg_1_12_0_port, pg_1_11_1_port, pg_1_11_0_port, 
      pg_1_10_1_port, pg_1_10_0_port, pg_1_9_1_port, pg_1_9_0_port, 
      pg_1_8_1_port, pg_1_8_0_port, pg_1_7_1_port, pg_1_7_0_port, pg_1_6_1_port
      , pg_1_6_0_port, pg_1_5_1_port, pg_1_5_0_port, pg_1_4_1_port, 
      pg_1_4_0_port, pg_1_3_1_port, pg_1_3_0_port, pg_1_2_1_port, pg_1_2_0_port
      , pg_1_1_1_port, pg_1_1_0_port, pg_1_0_0_port, pg_n_4_7_1_port, 
      pg_n_4_7_0_port, pg_n_4_6_1_port, pg_n_4_6_0_port, pg_n_3_7_1_port, 
      pg_n_3_7_0_port, pg_n_3_5_1_port, pg_n_3_5_0_port, pg_n_3_3_1_port, 
      pg_n_3_3_0_port, pg_n_2_7_1_port, pg_n_2_7_0_port, pg_n_2_6_1_port, 
      pg_n_2_6_0_port, pg_n_2_5_1_port, pg_n_2_5_0_port, pg_n_2_4_1_port, 
      pg_n_2_4_0_port, pg_n_2_3_1_port, pg_n_2_3_0_port, pg_n_2_2_1_port, 
      pg_n_2_2_0_port, pg_n_2_1_1_port, pg_n_2_1_0_port : std_logic;

begin
   Cout <= ( Cout_7_port, Cout_6_port, Cout_5_port, Cout_4_port, Cout_3_port, 
      Cout_2_port, Cout_1_port, Cout_0_port );
   
   pg_net_x_1 : pg_net_32 port map( a => A(1), b => B(1), g_out => g_net_1_port
                           , p_out => p_net_1_port);
   pg_net_x_2 : pg_net_31 port map( a => A(2), b => B(2), g_out => g_net_2_port
                           , p_out => p_net_2_port);
   pg_net_x_3 : pg_net_30 port map( a => A(3), b => B(3), g_out => g_net_3_port
                           , p_out => p_net_3_port);
   pg_net_x_4 : pg_net_29 port map( a => A(4), b => B(4), g_out => g_net_4_port
                           , p_out => p_net_4_port);
   pg_net_x_5 : pg_net_28 port map( a => A(5), b => B(5), g_out => g_net_5_port
                           , p_out => p_net_5_port);
   pg_net_x_6 : pg_net_27 port map( a => A(6), b => B(6), g_out => g_net_6_port
                           , p_out => p_net_6_port);
   pg_net_x_7 : pg_net_26 port map( a => A(7), b => B(7), g_out => g_net_7_port
                           , p_out => p_net_7_port);
   pg_net_x_8 : pg_net_25 port map( a => A(8), b => B(8), g_out => g_net_8_port
                           , p_out => p_net_8_port);
   pg_net_x_9 : pg_net_24 port map( a => A(9), b => B(9), g_out => g_net_9_port
                           , p_out => p_net_9_port);
   pg_net_x_10 : pg_net_23 port map( a => A(10), b => B(10), g_out => 
                           g_net_10_port, p_out => p_net_10_port);
   pg_net_x_11 : pg_net_22 port map( a => A(11), b => B(11), g_out => 
                           g_net_11_port, p_out => p_net_11_port);
   pg_net_x_12 : pg_net_21 port map( a => A(12), b => B(12), g_out => 
                           g_net_12_port, p_out => p_net_12_port);
   pg_net_x_13 : pg_net_20 port map( a => A(13), b => B(13), g_out => 
                           g_net_13_port, p_out => p_net_13_port);
   pg_net_x_14 : pg_net_19 port map( a => A(14), b => B(14), g_out => 
                           g_net_14_port, p_out => p_net_14_port);
   pg_net_x_15 : pg_net_18 port map( a => A(15), b => B(15), g_out => 
                           g_net_15_port, p_out => p_net_15_port);
   pg_net_x_16 : pg_net_17 port map( a => A(16), b => B(16), g_out => 
                           g_net_16_port, p_out => p_net_16_port);
   pg_net_x_17 : pg_net_16 port map( a => A(17), b => B(17), g_out => 
                           g_net_17_port, p_out => p_net_17_port);
   pg_net_x_18 : pg_net_15 port map( a => A(18), b => B(18), g_out => 
                           g_net_18_port, p_out => p_net_18_port);
   pg_net_x_19 : pg_net_14 port map( a => A(19), b => B(19), g_out => 
                           g_net_19_port, p_out => p_net_19_port);
   pg_net_x_20 : pg_net_13 port map( a => A(20), b => B(20), g_out => 
                           g_net_20_port, p_out => p_net_20_port);
   pg_net_x_21 : pg_net_12 port map( a => A(21), b => B(21), g_out => 
                           g_net_21_port, p_out => p_net_21_port);
   pg_net_x_22 : pg_net_11 port map( a => A(22), b => B(22), g_out => 
                           g_net_22_port, p_out => p_net_22_port);
   pg_net_x_23 : pg_net_10 port map( a => A(23), b => B(23), g_out => 
                           g_net_23_port, p_out => p_net_23_port);
   pg_net_x_24 : pg_net_9 port map( a => A(24), b => B(24), g_out => 
                           g_net_24_port, p_out => p_net_24_port);
   pg_net_x_25 : pg_net_8 port map( a => A(25), b => B(25), g_out => 
                           g_net_25_port, p_out => p_net_25_port);
   pg_net_x_26 : pg_net_7 port map( a => A(26), b => B(26), g_out => 
                           g_net_26_port, p_out => p_net_26_port);
   pg_net_x_27 : pg_net_6 port map( a => A(27), b => B(27), g_out => 
                           g_net_27_port, p_out => p_net_27_port);
   pg_net_x_28 : pg_net_5 port map( a => A(28), b => B(28), g_out => 
                           g_net_28_port, p_out => p_net_28_port);
   pg_net_x_29 : pg_net_4 port map( a => A(29), b => B(29), g_out => 
                           g_net_29_port, p_out => p_net_29_port);
   pg_net_x_30 : pg_net_3 port map( a => A(30), b => B(30), g_out => 
                           g_net_30_port, p_out => p_net_30_port);
   pg_net_x_31 : pg_net_2 port map( a => A(31), b => B(31), g_out => 
                           g_net_31_port, p_out => p_net_31_port);
   pg_net_0_MAGIC : pg_net_1 port map( a => A(0), b => B(0), g_out => 
                           magic_pro_0_port, p_out => magic_pro_1_port);
   xG_0_0_MAGIC : g_10 port map( g => magic_pro_0_port, p => magic_pro_1_port, 
                           g_prec => Cin, g_out => g_net_0_port);
   xG_1_0 : g_9 port map( g => g_net_1_port, p => p_net_1_port, g_prec => 
                           g_net_0_port, g_out => pg_1_0_0_port);
   xPG_1_1 : pg_27 port map( g => g_net_3_port, p => p_net_3_port, g_prec => 
                           g_net_2_port, p_prec => p_net_2_port, g_out => 
                           pg_1_1_0_port, p_out => pg_1_1_1_port);
   xPG_1_2 : pg_26 port map( g => g_net_5_port, p => p_net_5_port, g_prec => 
                           g_net_4_port, p_prec => p_net_4_port, g_out => 
                           pg_1_2_0_port, p_out => pg_1_2_1_port);
   xPG_1_3 : pg_25 port map( g => g_net_7_port, p => p_net_7_port, g_prec => 
                           g_net_6_port, p_prec => p_net_6_port, p_out => 
                           pg_1_3_1_port, g_out_BAR => pg_1_3_0_port);
   xPG_1_4 : pg_24 port map( g => g_net_9_port, p => p_net_9_port, g_prec => 
                           g_net_8_port, p_prec => p_net_8_port, g_out => 
                           pg_1_4_0_port, p_out => pg_1_4_1_port);
   xPG_1_5 : pg_23 port map( g => g_net_11_port, p => p_net_11_port, g_prec => 
                           g_net_10_port, p_prec => p_net_10_port, g_out => 
                           pg_1_5_0_port, p_out => pg_1_5_1_port);
   xPG_1_6 : pg_22 port map( g => g_net_13_port, p => p_net_13_port, g_prec => 
                           g_net_12_port, p_prec => p_net_12_port, g_out => 
                           pg_1_6_0_port, p_out => pg_1_6_1_port);
   xPG_1_7 : pg_21 port map( g => g_net_15_port, p => p_net_15_port, g_prec => 
                           g_net_14_port, p_prec => p_net_14_port, g_out => 
                           pg_1_7_0_port, p_out => pg_1_7_1_port);
   xPG_1_8 : pg_20 port map( g => g_net_17_port, p => p_net_17_port, g_prec => 
                           g_net_16_port, p_prec => p_net_16_port, g_out => 
                           pg_1_8_0_port, p_out => pg_1_8_1_port);
   xPG_1_9 : pg_19 port map( g => g_net_19_port, p => p_net_19_port, g_prec => 
                           g_net_18_port, p_prec => p_net_18_port, g_out => 
                           pg_1_9_0_port, p_out => pg_1_9_1_port);
   xPG_1_10 : pg_18 port map( g => g_net_21_port, p => p_net_21_port, g_prec =>
                           g_net_20_port, p_prec => p_net_20_port, g_out => 
                           pg_1_10_0_port, p_out => pg_1_10_1_port);
   xPG_1_11 : pg_17 port map( g => g_net_23_port, p => p_net_23_port, g_prec =>
                           g_net_22_port, p_prec => p_net_22_port, g_out => 
                           pg_1_11_0_port, p_out => pg_1_11_1_port);
   xPG_1_12 : pg_16 port map( g => g_net_25_port, p => p_net_25_port, g_prec =>
                           g_net_24_port, p_prec => p_net_24_port, g_out => 
                           pg_1_12_0_port, p_out => pg_1_12_1_port);
   xPG_1_13 : pg_15 port map( g => g_net_27_port, p => p_net_27_port, g_prec =>
                           g_net_26_port, p_prec => p_net_26_port, g_out => 
                           pg_1_13_0_port, p_out => pg_1_13_1_port);
   xPG_1_14 : pg_14 port map( g => g_net_29_port, p => p_net_29_port, g_prec =>
                           g_net_28_port, p_prec => p_net_28_port, g_out => 
                           pg_1_14_0_port, p_out => pg_1_14_1_port);
   xPG_1_15 : pg_13 port map( g => g_net_31_port, p => p_net_31_port, g_prec =>
                           g_net_30_port, p_prec => p_net_30_port, g_out => 
                           pg_1_15_0_port, p_out => pg_1_15_1_port);
   xG_2_0 : g_8 port map( g => pg_1_1_0_port, p => pg_1_1_1_port, g_prec => 
                           pg_1_0_0_port, g_out => Cout_0_port);
   xPG_2_1 : pg_12 port map( p => pg_1_3_1_port, g_prec => pg_1_2_0_port, 
                           p_prec => pg_1_2_1_port, g_out => pg_n_2_1_0_port, 
                           p_out => pg_n_2_1_1_port, g_BAR => pg_1_3_0_port);
   xPG_2_2 : pg_11 port map( g => pg_1_5_0_port, p => pg_1_5_1_port, g_prec => 
                           pg_1_4_0_port, p_prec => pg_1_4_1_port, g_out => 
                           pg_n_2_2_0_port, p_out => pg_n_2_2_1_port);
   xPG_2_3 : pg_10 port map( g => pg_1_7_0_port, p => pg_1_7_1_port, g_prec => 
                           pg_1_6_0_port, p_prec => pg_1_6_1_port, p_out => 
                           pg_n_2_3_1_port, g_out_BAR => pg_n_2_3_0_port);
   xPG_2_4 : pg_9 port map( g => pg_1_9_0_port, p => pg_1_9_1_port, g_prec => 
                           pg_1_8_0_port, p_prec => pg_1_8_1_port, p_out => 
                           pg_n_2_4_1_port, g_out_BAR => pg_n_2_4_0_port);
   xPG_2_5 : pg_8 port map( g => pg_1_11_0_port, p => pg_1_11_1_port, g_prec =>
                           pg_1_10_0_port, p_prec => pg_1_10_1_port, g_out => 
                           pg_n_2_5_0_port, p_out => pg_n_2_5_1_port);
   xPG_2_6 : pg_7 port map( g => pg_1_13_0_port, p => pg_1_13_1_port, g_prec =>
                           pg_1_12_0_port, p_prec => pg_1_12_1_port, p_out => 
                           pg_n_2_6_1_port, g_out_BAR => pg_n_2_6_0_port);
   xPG_2_7 : pg_6 port map( g => pg_1_15_0_port, p => pg_1_15_1_port, g_prec =>
                           pg_1_14_0_port, p_prec => pg_1_14_1_port, g_out => 
                           pg_n_2_7_0_port, p_out => pg_n_2_7_1_port);
   xG_3_1 : g_7 port map( g => pg_n_2_1_0_port, p => pg_n_2_1_1_port, g_prec =>
                           Cout_0_port, g_out => Cout_1_port);
   xG_4_2 : g_6 port map( g => pg_n_2_2_0_port, p => pg_n_2_2_1_port, g_prec =>
                           Cout_1_port, g_out => Cout_2_port);
   xG_4_3 : g_5 port map( g => pg_n_3_3_0_port, p => pg_n_3_3_1_port, g_prec =>
                           Cout_1_port, g_out => Cout_3_port);
   xG_5_4 : g_4 port map( p => pg_n_2_4_1_port, g_prec => Cout_3_port, g_out =>
                           Cout_4_port, g_BAR => pg_n_2_4_0_port);
   xG_5_5 : g_3 port map( g => pg_n_3_5_0_port, p => pg_n_3_5_1_port, g_prec =>
                           Cout_3_port, g_out => Cout_5_port);
   xG_5_6 : g_2 port map( g => pg_n_4_6_0_port, p => pg_n_4_6_1_port, g_prec =>
                           Cout_3_port, g_out => Cout_6_port);
   xG_5_7 : g_1 port map( g => pg_n_4_7_0_port, p => pg_n_4_7_1_port, g_prec =>
                           Cout_3_port, g_out => Cout_7_port);
   xPG_3_3 : pg_5 port map( p => pg_n_2_3_1_port, g_prec => pg_n_2_2_0_port, 
                           p_prec => pg_n_2_2_1_port, g_out => pg_n_3_3_0_port,
                           p_out => pg_n_3_3_1_port, g_BAR => pg_n_2_3_0_port);
   xPG_3_5 : pg_4 port map( g => pg_n_2_5_0_port, p => pg_n_2_5_1_port, p_prec 
                           => pg_n_2_4_1_port, g_out => pg_n_3_5_0_port, p_out 
                           => pg_n_3_5_1_port, g_prec_BAR => pg_n_2_4_0_port);
   xPG_3_7 : pg_3 port map( g => pg_n_2_7_0_port, p => pg_n_2_7_1_port, p_prec 
                           => pg_n_2_6_1_port, g_out => pg_n_3_7_0_port, p_out 
                           => pg_n_3_7_1_port, g_prec_BAR => pg_n_2_6_0_port);
   xPG_4_6 : pg_2 port map( p => pg_n_2_6_1_port, g_prec => pg_n_3_5_0_port, 
                           p_prec => pg_n_3_5_1_port, g_out => pg_n_4_6_0_port,
                           p_out => pg_n_4_6_1_port, g_BAR => pg_n_2_6_0_port);
   xPG_4_7 : pg_1 port map( g => pg_n_3_7_0_port, p => pg_n_3_7_1_port, g_prec 
                           => pg_n_3_5_0_port, p_prec => pg_n_3_5_1_port, g_out
                           => pg_n_4_7_0_port, p_out => pg_n_4_7_1_port);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity xor_gen_N32_1 is

   port( A : in std_logic_vector (31 downto 0);  B : in std_logic;  S : out 
         std_logic_vector (31 downto 0));

end xor_gen_N32_1;

architecture SYN_bhe of xor_gen_N32_1 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X2
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U4 : XOR2_X1 port map( A => B, B => A(6), Z => S(6));
   U8 : XOR2_X1 port map( A => B, B => A(31), Z => S(31));
   U9 : XOR2_X1 port map( A => B, B => A(30), Z => S(30));
   U11 : XOR2_X1 port map( A => B, B => A(29), Z => S(29));
   U12 : XOR2_X1 port map( A => B, B => A(28), Z => S(28));
   U13 : XOR2_X1 port map( A => B, B => A(27), Z => S(27));
   U14 : XOR2_X1 port map( A => B, B => A(26), Z => S(26));
   U15 : XOR2_X1 port map( A => B, B => A(25), Z => S(25));
   U16 : XOR2_X1 port map( A => B, B => A(24), Z => S(24));
   U17 : XOR2_X1 port map( A => B, B => A(23), Z => S(23));
   U18 : XOR2_X1 port map( A => B, B => A(22), Z => S(22));
   U20 : XOR2_X1 port map( A => B, B => A(20), Z => S(20));
   U22 : XOR2_X1 port map( A => B, B => A(19), Z => S(19));
   U23 : XOR2_X1 port map( A => B, B => A(18), Z => S(18));
   U26 : XOR2_X1 port map( A => B, B => A(15), Z => S(15));
   U29 : XOR2_X1 port map( A => B, B => A(12), Z => S(12));
   U30 : XOR2_X1 port map( A => A(11), B => B, Z => S(11));
   U24 : XOR2_X1 port map( A => B, B => A(17), Z => S(17));
   U1 : XOR2_X1 port map( A => B, B => A(4), Z => S(4));
   U2 : XOR2_X1 port map( A => B, B => A(2), Z => S(2));
   U3 : MUX2_X1 port map( A => B, B => n4, S => A(5), Z => S(5));
   U5 : XOR2_X1 port map( A => B, B => A(7), Z => S(7));
   U6 : XOR2_X1 port map( A => B, B => A(21), Z => S(21));
   U7 : INV_X1 port map( A => B, ZN => n4);
   U10 : XOR2_X1 port map( A => B, B => A(9), Z => S(9));
   U19 : INV_X1 port map( A => A(3), ZN => n1);
   U21 : XOR2_X2 port map( A => B, B => A(10), Z => S(10));
   U25 : XOR2_X2 port map( A => A(0), B => B, Z => S(0));
   U27 : NAND2_X1 port map( A1 => n2, A2 => n3, ZN => S(3));
   U28 : XOR2_X1 port map( A => B, B => A(16), Z => S(16));
   U31 : XOR2_X1 port map( A => A(8), B => B, Z => S(8));
   U32 : XOR2_X1 port map( A => B, B => A(14), Z => S(14));
   U33 : NAND2_X1 port map( A1 => B, A2 => n1, ZN => n2);
   U34 : NAND2_X1 port map( A1 => n4, A2 => A(3), ZN => n3);
   U35 : XOR2_X1 port map( A => B, B => A(13), Z => S(13));
   U36 : XOR2_X1 port map( A => A(1), B => B, Z => S(1));

end SYN_bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity ff32_en_SIZE5_3 is

   port( D : in std_logic_vector (4 downto 0);  en, clk, rst : in std_logic;  Q
         : out std_logic_vector (4 downto 0));

end ff32_en_SIZE5_3;

architecture SYN_behavioral of ff32_en_SIZE5_3 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_ff32_en_SIZE5_3
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   signal net199373, n1, n5, n6, n7, n8, n9, net246145 : std_logic;

begin
   
   Q_reg_4_inst : DFFR_X1 port map( D => D(4), CK => net199373, RN => n7, Q => 
                           net246145, QN => n1);
   Q_reg_3_inst : DFFR_X1 port map( D => D(3), CK => net199373, RN => n7, Q => 
                           Q(3), QN => n8);
   Q_reg_1_inst : DFFR_X1 port map( D => D(1), CK => net199373, RN => n7, Q => 
                           Q(1), QN => n9);
   clk_gate_Q_reg : SNPS_CLOCK_GATE_HIGH_ff32_en_SIZE5_3 port map( CLK => clk, 
                           EN => en, ENCLK => net199373);
   Q_reg_2_inst : DFFR_X1 port map( D => D(2), CK => net199373, RN => n7, Q => 
                           Q(2), QN => n6);
   Q_reg_0_inst : DFFR_X1 port map( D => D(0), CK => net199373, RN => n7, Q => 
                           Q(0), QN => n5);
   U2 : INV_X1 port map( A => n1, ZN => Q(4));
   U3 : INV_X1 port map( A => rst, ZN => n7);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity ff32_en_SIZE5_2 is

   port( D : in std_logic_vector (4 downto 0);  en, clk, rst : in std_logic;  Q
         : out std_logic_vector (4 downto 0));

end ff32_en_SIZE5_2;

architecture SYN_behavioral of ff32_en_SIZE5_2 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_ff32_en_SIZE5_2
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal net199373, n5, n7, n8, n9, n10, n11 : std_logic;

begin
   
   Q_reg_4_inst : DFFR_X1 port map( D => D(4), CK => net199373, RN => n5, Q => 
                           Q(4), QN => n7);
   Q_reg_3_inst : DFFR_X1 port map( D => D(3), CK => net199373, RN => n5, Q => 
                           Q(3), QN => n8);
   Q_reg_2_inst : DFFR_X1 port map( D => D(2), CK => net199373, RN => n5, Q => 
                           Q(2), QN => n9);
   Q_reg_1_inst : DFFR_X1 port map( D => D(1), CK => net199373, RN => n5, Q => 
                           Q(1), QN => n10);
   Q_reg_0_inst : DFFR_X1 port map( D => D(0), CK => net199373, RN => n5, Q => 
                           Q(0), QN => n11);
   clk_gate_Q_reg : SNPS_CLOCK_GATE_HIGH_ff32_en_SIZE5_2 port map( CLK => clk, 
                           EN => en, ENCLK => net199373);
   U2 : INV_X1 port map( A => rst, ZN => n5);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity ff32_en_SIZE5_1 is

   port( D : in std_logic_vector (4 downto 0);  en, clk, rst : in std_logic;  Q
         : out std_logic_vector (4 downto 0));

end ff32_en_SIZE5_1;

architecture SYN_behavioral of ff32_en_SIZE5_1 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n3, n4, n5, n7, net246143, net246144 : std_logic;

begin
   
   Q_reg_4_inst : DFFR_X1 port map( D => D(4), CK => clk, RN => n5, Q => Q(4), 
                           QN => n7);
   Q_reg_1_inst : DFFR_X1 port map( D => D(1), CK => clk, RN => n5, Q => Q(1), 
                           QN => net246144);
   Q_reg_0_inst : DFFR_X1 port map( D => D(0), CK => clk, RN => n5, Q => Q(0), 
                           QN => n4);
   Q_reg_2_inst : DFFR_X1 port map( D => D(2), CK => clk, RN => n5, Q => Q(2), 
                           QN => n3);
   Q_reg_3_inst : DFFR_X1 port map( D => D(3), CK => clk, RN => n5, Q => Q(3), 
                           QN => net246143);
   U2 : INV_X1 port map( A => rst, ZN => n5);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity ff32_en_SIZE32_5 is

   port( D : in std_logic_vector (31 downto 0);  en, clk, rst : in std_logic;  
         Q : out std_logic_vector (31 downto 0));

end ff32_en_SIZE32_5;

architecture SYN_behavioral of ff32_en_SIZE32_5 is

   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_ff32_en_SIZE32_5
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal net199358, n32, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44
      , n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, 
      n59, n60, n61, n62, n63, n64, n65 : std_logic;

begin
   
   Q_reg_31_inst : DFFR_X1 port map( D => D(31), CK => net199358, RN => n32, Q 
                           => Q(31), QN => n34);
   Q_reg_30_inst : DFFR_X1 port map( D => D(30), CK => net199358, RN => n32, Q 
                           => Q(30), QN => n35);
   Q_reg_29_inst : DFFR_X1 port map( D => D(29), CK => net199358, RN => n32, Q 
                           => Q(29), QN => n36);
   Q_reg_28_inst : DFFR_X1 port map( D => D(28), CK => net199358, RN => n32, Q 
                           => Q(28), QN => n37);
   Q_reg_27_inst : DFFR_X1 port map( D => D(27), CK => net199358, RN => n32, Q 
                           => Q(27), QN => n38);
   Q_reg_26_inst : DFFR_X1 port map( D => D(26), CK => net199358, RN => n32, Q 
                           => Q(26), QN => n39);
   Q_reg_25_inst : DFFR_X1 port map( D => D(25), CK => net199358, RN => n32, Q 
                           => Q(25), QN => n40);
   Q_reg_24_inst : DFFR_X1 port map( D => D(24), CK => net199358, RN => n32, Q 
                           => Q(24), QN => n41);
   Q_reg_23_inst : DFFR_X1 port map( D => D(23), CK => net199358, RN => n32, Q 
                           => Q(23), QN => n42);
   Q_reg_22_inst : DFFR_X1 port map( D => D(22), CK => net199358, RN => n32, Q 
                           => Q(22), QN => n43);
   Q_reg_21_inst : DFFR_X1 port map( D => D(21), CK => net199358, RN => n32, Q 
                           => Q(21), QN => n44);
   Q_reg_20_inst : DFFR_X1 port map( D => D(20), CK => net199358, RN => n32, Q 
                           => Q(20), QN => n45);
   Q_reg_19_inst : DFFR_X1 port map( D => D(19), CK => net199358, RN => n32, Q 
                           => Q(19), QN => n46);
   Q_reg_18_inst : DFFR_X1 port map( D => D(18), CK => net199358, RN => n32, Q 
                           => Q(18), QN => n47);
   Q_reg_17_inst : DFFR_X1 port map( D => D(17), CK => net199358, RN => n32, Q 
                           => Q(17), QN => n48);
   Q_reg_16_inst : DFFR_X1 port map( D => D(16), CK => net199358, RN => n32, Q 
                           => Q(16), QN => n49);
   Q_reg_15_inst : DFFR_X1 port map( D => D(15), CK => net199358, RN => n32, Q 
                           => Q(15), QN => n50);
   Q_reg_14_inst : DFFR_X1 port map( D => D(14), CK => net199358, RN => n32, Q 
                           => Q(14), QN => n51);
   Q_reg_13_inst : DFFR_X1 port map( D => D(13), CK => net199358, RN => n32, Q 
                           => Q(13), QN => n52);
   Q_reg_12_inst : DFFR_X1 port map( D => D(12), CK => net199358, RN => n32, Q 
                           => Q(12), QN => n53);
   Q_reg_11_inst : DFFR_X1 port map( D => D(11), CK => net199358, RN => n32, Q 
                           => Q(11), QN => n54);
   Q_reg_10_inst : DFFR_X1 port map( D => D(10), CK => net199358, RN => n32, Q 
                           => Q(10), QN => n55);
   Q_reg_9_inst : DFFR_X1 port map( D => D(9), CK => net199358, RN => n32, Q =>
                           Q(9), QN => n56);
   Q_reg_8_inst : DFFR_X1 port map( D => D(8), CK => net199358, RN => n32, Q =>
                           Q(8), QN => n57);
   Q_reg_7_inst : DFFR_X1 port map( D => D(7), CK => net199358, RN => n32, Q =>
                           Q(7), QN => n58);
   Q_reg_6_inst : DFFR_X1 port map( D => D(6), CK => net199358, RN => n32, Q =>
                           Q(6), QN => n59);
   Q_reg_5_inst : DFFR_X1 port map( D => D(5), CK => net199358, RN => n32, Q =>
                           Q(5), QN => n60);
   Q_reg_4_inst : DFFR_X1 port map( D => D(4), CK => net199358, RN => n32, Q =>
                           Q(4), QN => n61);
   Q_reg_3_inst : DFFR_X1 port map( D => D(3), CK => net199358, RN => n32, Q =>
                           Q(3), QN => n62);
   Q_reg_2_inst : DFFR_X1 port map( D => D(2), CK => net199358, RN => n32, Q =>
                           Q(2), QN => n63);
   Q_reg_1_inst : DFFR_X1 port map( D => D(1), CK => net199358, RN => n32, Q =>
                           Q(1), QN => n64);
   Q_reg_0_inst : DFFR_X1 port map( D => D(0), CK => net199358, RN => n32, Q =>
                           Q(0), QN => n65);
   clk_gate_Q_reg : SNPS_CLOCK_GATE_HIGH_ff32_en_SIZE32_5 port map( CLK => clk,
                           EN => en, ENCLK => net199358);
   U2 : INV_X2 port map( A => rst, ZN => n32);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity ff32_en_SIZE32_4 is

   port( D : in std_logic_vector (31 downto 0);  en, clk, rst : in std_logic;  
         Q : out std_logic_vector (31 downto 0));

end ff32_en_SIZE32_4;

architecture SYN_behavioral of ff32_en_SIZE32_4 is

   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_ff32_en_SIZE32_4
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal net199358, n32, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44
      , n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, 
      n59, n60, n61, n62, n63, n64, n65 : std_logic;

begin
   
   Q_reg_31_inst : DFFR_X1 port map( D => D(31), CK => net199358, RN => n32, Q 
                           => Q(31), QN => n34);
   Q_reg_30_inst : DFFR_X1 port map( D => D(30), CK => net199358, RN => n32, Q 
                           => Q(30), QN => n35);
   Q_reg_29_inst : DFFR_X1 port map( D => D(29), CK => net199358, RN => n32, Q 
                           => Q(29), QN => n36);
   Q_reg_28_inst : DFFR_X1 port map( D => D(28), CK => net199358, RN => n32, Q 
                           => Q(28), QN => n37);
   Q_reg_27_inst : DFFR_X1 port map( D => D(27), CK => net199358, RN => n32, Q 
                           => Q(27), QN => n38);
   Q_reg_26_inst : DFFR_X1 port map( D => D(26), CK => net199358, RN => n32, Q 
                           => Q(26), QN => n39);
   Q_reg_25_inst : DFFR_X1 port map( D => D(25), CK => net199358, RN => n32, Q 
                           => Q(25), QN => n40);
   Q_reg_24_inst : DFFR_X1 port map( D => D(24), CK => net199358, RN => n32, Q 
                           => Q(24), QN => n41);
   Q_reg_23_inst : DFFR_X1 port map( D => D(23), CK => net199358, RN => n32, Q 
                           => Q(23), QN => n42);
   Q_reg_22_inst : DFFR_X1 port map( D => D(22), CK => net199358, RN => n32, Q 
                           => Q(22), QN => n43);
   Q_reg_21_inst : DFFR_X1 port map( D => D(21), CK => net199358, RN => n32, Q 
                           => Q(21), QN => n44);
   Q_reg_20_inst : DFFR_X1 port map( D => D(20), CK => net199358, RN => n32, Q 
                           => Q(20), QN => n45);
   Q_reg_19_inst : DFFR_X1 port map( D => D(19), CK => net199358, RN => n32, Q 
                           => Q(19), QN => n46);
   Q_reg_18_inst : DFFR_X1 port map( D => D(18), CK => net199358, RN => n32, Q 
                           => Q(18), QN => n47);
   Q_reg_17_inst : DFFR_X1 port map( D => D(17), CK => net199358, RN => n32, Q 
                           => Q(17), QN => n48);
   Q_reg_16_inst : DFFR_X1 port map( D => D(16), CK => net199358, RN => n32, Q 
                           => Q(16), QN => n49);
   Q_reg_15_inst : DFFR_X1 port map( D => D(15), CK => net199358, RN => n32, Q 
                           => Q(15), QN => n50);
   Q_reg_14_inst : DFFR_X1 port map( D => D(14), CK => net199358, RN => n32, Q 
                           => Q(14), QN => n51);
   Q_reg_13_inst : DFFR_X1 port map( D => D(13), CK => net199358, RN => n32, Q 
                           => Q(13), QN => n52);
   Q_reg_12_inst : DFFR_X1 port map( D => D(12), CK => net199358, RN => n32, Q 
                           => Q(12), QN => n53);
   Q_reg_11_inst : DFFR_X1 port map( D => D(11), CK => net199358, RN => n32, Q 
                           => Q(11), QN => n54);
   Q_reg_10_inst : DFFR_X1 port map( D => D(10), CK => net199358, RN => n32, Q 
                           => Q(10), QN => n55);
   Q_reg_9_inst : DFFR_X1 port map( D => D(9), CK => net199358, RN => n32, Q =>
                           Q(9), QN => n56);
   Q_reg_8_inst : DFFR_X1 port map( D => D(8), CK => net199358, RN => n32, Q =>
                           Q(8), QN => n57);
   Q_reg_7_inst : DFFR_X1 port map( D => D(7), CK => net199358, RN => n32, Q =>
                           Q(7), QN => n58);
   Q_reg_6_inst : DFFR_X1 port map( D => D(6), CK => net199358, RN => n32, Q =>
                           Q(6), QN => n59);
   Q_reg_5_inst : DFFR_X1 port map( D => D(5), CK => net199358, RN => n32, Q =>
                           Q(5), QN => n60);
   Q_reg_4_inst : DFFR_X1 port map( D => D(4), CK => net199358, RN => n32, Q =>
                           Q(4), QN => n61);
   Q_reg_3_inst : DFFR_X1 port map( D => D(3), CK => net199358, RN => n32, Q =>
                           Q(3), QN => n62);
   Q_reg_2_inst : DFFR_X1 port map( D => D(2), CK => net199358, RN => n32, Q =>
                           Q(2), QN => n63);
   Q_reg_1_inst : DFFR_X1 port map( D => D(1), CK => net199358, RN => n32, Q =>
                           Q(1), QN => n64);
   Q_reg_0_inst : DFFR_X1 port map( D => D(0), CK => net199358, RN => n32, Q =>
                           Q(0), QN => n65);
   clk_gate_Q_reg : SNPS_CLOCK_GATE_HIGH_ff32_en_SIZE32_4 port map( CLK => clk,
                           EN => en, ENCLK => net199358);
   U2 : INV_X2 port map( A => rst, ZN => n32);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity ff32_en_SIZE32_3 is

   port( D : in std_logic_vector (31 downto 0);  en, clk, rst : in std_logic;  
         Q : out std_logic_vector (31 downto 0));

end ff32_en_SIZE32_3;

architecture SYN_behavioral of ff32_en_SIZE32_3 is

   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n32, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
      n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61
      , n62, n63, n64, n65 : std_logic;

begin
   
   Q_reg_31_inst : DFFR_X1 port map( D => D(31), CK => clk, RN => n32, Q => 
                           Q(31), QN => n34);
   Q_reg_30_inst : DFFR_X1 port map( D => D(30), CK => clk, RN => n32, Q => 
                           Q(30), QN => n35);
   Q_reg_29_inst : DFFR_X1 port map( D => D(29), CK => clk, RN => n32, Q => 
                           Q(29), QN => n36);
   Q_reg_28_inst : DFFR_X1 port map( D => D(28), CK => clk, RN => n32, Q => 
                           Q(28), QN => n37);
   Q_reg_27_inst : DFFR_X1 port map( D => D(27), CK => clk, RN => n32, Q => 
                           Q(27), QN => n38);
   Q_reg_26_inst : DFFR_X1 port map( D => D(26), CK => clk, RN => n32, Q => 
                           Q(26), QN => n39);
   Q_reg_25_inst : DFFR_X1 port map( D => D(25), CK => clk, RN => n32, Q => 
                           Q(25), QN => n40);
   Q_reg_24_inst : DFFR_X1 port map( D => D(24), CK => clk, RN => n32, Q => 
                           Q(24), QN => n41);
   Q_reg_23_inst : DFFR_X1 port map( D => D(23), CK => clk, RN => n32, Q => 
                           Q(23), QN => n42);
   Q_reg_22_inst : DFFR_X1 port map( D => D(22), CK => clk, RN => n32, Q => 
                           Q(22), QN => n43);
   Q_reg_21_inst : DFFR_X1 port map( D => D(21), CK => clk, RN => n32, Q => 
                           Q(21), QN => n44);
   Q_reg_20_inst : DFFR_X1 port map( D => D(20), CK => clk, RN => n32, Q => 
                           Q(20), QN => n45);
   Q_reg_19_inst : DFFR_X1 port map( D => D(19), CK => clk, RN => n32, Q => 
                           Q(19), QN => n46);
   Q_reg_18_inst : DFFR_X1 port map( D => D(18), CK => clk, RN => n32, Q => 
                           Q(18), QN => n47);
   Q_reg_17_inst : DFFR_X1 port map( D => D(17), CK => clk, RN => n32, Q => 
                           Q(17), QN => n48);
   Q_reg_16_inst : DFFR_X1 port map( D => D(16), CK => clk, RN => n32, Q => 
                           Q(16), QN => n49);
   Q_reg_15_inst : DFFR_X1 port map( D => D(15), CK => clk, RN => n32, Q => 
                           Q(15), QN => n50);
   Q_reg_14_inst : DFFR_X1 port map( D => D(14), CK => clk, RN => n32, Q => 
                           Q(14), QN => n51);
   Q_reg_13_inst : DFFR_X1 port map( D => D(13), CK => clk, RN => n32, Q => 
                           Q(13), QN => n52);
   Q_reg_12_inst : DFFR_X1 port map( D => D(12), CK => clk, RN => n32, Q => 
                           Q(12), QN => n53);
   Q_reg_11_inst : DFFR_X1 port map( D => D(11), CK => clk, RN => n32, Q => 
                           Q(11), QN => n54);
   Q_reg_10_inst : DFFR_X1 port map( D => D(10), CK => clk, RN => n32, Q => 
                           Q(10), QN => n55);
   Q_reg_9_inst : DFFR_X1 port map( D => D(9), CK => clk, RN => n32, Q => Q(9),
                           QN => n56);
   Q_reg_8_inst : DFFR_X1 port map( D => D(8), CK => clk, RN => n32, Q => Q(8),
                           QN => n57);
   Q_reg_7_inst : DFFR_X1 port map( D => D(7), CK => clk, RN => n32, Q => Q(7),
                           QN => n58);
   Q_reg_6_inst : DFFR_X1 port map( D => D(6), CK => clk, RN => n32, Q => Q(6),
                           QN => n59);
   Q_reg_5_inst : DFFR_X1 port map( D => D(5), CK => clk, RN => n32, Q => Q(5),
                           QN => n60);
   Q_reg_4_inst : DFFR_X1 port map( D => D(4), CK => clk, RN => n32, Q => Q(4),
                           QN => n61);
   Q_reg_3_inst : DFFR_X1 port map( D => D(3), CK => clk, RN => n32, Q => Q(3),
                           QN => n62);
   Q_reg_2_inst : DFFR_X1 port map( D => D(2), CK => clk, RN => n32, Q => Q(2),
                           QN => n63);
   Q_reg_1_inst : DFFR_X1 port map( D => D(1), CK => clk, RN => n32, Q => Q(1),
                           QN => n64);
   Q_reg_0_inst : DFFR_X1 port map( D => D(0), CK => clk, RN => n32, Q => Q(0),
                           QN => n65);
   U2 : INV_X2 port map( A => rst, ZN => n32);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity ff32_en_SIZE32_2 is

   port( D : in std_logic_vector (31 downto 0);  en, clk, rst : in std_logic;  
         Q : out std_logic_vector (31 downto 0));

end ff32_en_SIZE32_2;

architecture SYN_behavioral of ff32_en_SIZE32_2 is

   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
      n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62
      , n63, n64, n65, n66 : std_logic;

begin
   
   Q_reg_31_inst : DFFR_X1 port map( D => D(31), CK => clk, RN => n34, Q => 
                           Q(31), QN => n35);
   Q_reg_30_inst : DFFR_X1 port map( D => D(30), CK => clk, RN => n34, Q => 
                           Q(30), QN => n36);
   Q_reg_29_inst : DFFR_X1 port map( D => D(29), CK => clk, RN => n34, Q => 
                           Q(29), QN => n37);
   Q_reg_28_inst : DFFR_X1 port map( D => D(28), CK => clk, RN => n34, Q => 
                           Q(28), QN => n38);
   Q_reg_27_inst : DFFR_X1 port map( D => D(27), CK => clk, RN => n34, Q => 
                           Q(27), QN => n39);
   Q_reg_26_inst : DFFR_X1 port map( D => D(26), CK => clk, RN => n34, Q => 
                           Q(26), QN => n40);
   Q_reg_25_inst : DFFR_X1 port map( D => D(25), CK => clk, RN => n34, Q => 
                           Q(25), QN => n41);
   Q_reg_24_inst : DFFR_X1 port map( D => D(24), CK => clk, RN => n34, Q => 
                           Q(24), QN => n42);
   Q_reg_23_inst : DFFR_X1 port map( D => D(23), CK => clk, RN => n34, Q => 
                           Q(23), QN => n43);
   Q_reg_22_inst : DFFR_X1 port map( D => D(22), CK => clk, RN => n34, Q => 
                           Q(22), QN => n44);
   Q_reg_21_inst : DFFR_X1 port map( D => D(21), CK => clk, RN => n34, Q => 
                           Q(21), QN => n45);
   Q_reg_20_inst : DFFR_X1 port map( D => D(20), CK => clk, RN => n34, Q => 
                           Q(20), QN => n46);
   Q_reg_19_inst : DFFR_X1 port map( D => D(19), CK => clk, RN => n34, Q => 
                           Q(19), QN => n47);
   Q_reg_18_inst : DFFR_X1 port map( D => D(18), CK => clk, RN => n34, Q => 
                           Q(18), QN => n48);
   Q_reg_17_inst : DFFR_X1 port map( D => D(17), CK => clk, RN => n34, Q => 
                           Q(17), QN => n49);
   Q_reg_16_inst : DFFR_X1 port map( D => D(16), CK => clk, RN => n34, Q => 
                           Q(16), QN => n50);
   Q_reg_15_inst : DFFR_X1 port map( D => D(15), CK => clk, RN => n34, Q => 
                           Q(15), QN => n51);
   Q_reg_14_inst : DFFR_X1 port map( D => D(14), CK => clk, RN => n34, Q => 
                           Q(14), QN => n52);
   Q_reg_13_inst : DFFR_X1 port map( D => D(13), CK => clk, RN => n34, Q => 
                           Q(13), QN => n53);
   Q_reg_12_inst : DFFR_X1 port map( D => D(12), CK => clk, RN => n34, Q => 
                           Q(12), QN => n54);
   Q_reg_11_inst : DFFR_X1 port map( D => D(11), CK => clk, RN => n34, Q => 
                           Q(11), QN => n55);
   Q_reg_10_inst : DFFR_X1 port map( D => D(10), CK => clk, RN => n34, Q => 
                           Q(10), QN => n56);
   Q_reg_9_inst : DFFR_X1 port map( D => D(9), CK => clk, RN => n34, Q => Q(9),
                           QN => n57);
   Q_reg_8_inst : DFFR_X1 port map( D => D(8), CK => clk, RN => n34, Q => Q(8),
                           QN => n58);
   Q_reg_7_inst : DFFR_X1 port map( D => D(7), CK => clk, RN => n34, Q => Q(7),
                           QN => n59);
   Q_reg_6_inst : DFFR_X1 port map( D => D(6), CK => clk, RN => n34, Q => Q(6),
                           QN => n60);
   Q_reg_5_inst : DFFR_X1 port map( D => D(5), CK => clk, RN => n34, Q => Q(5),
                           QN => n61);
   Q_reg_4_inst : DFFR_X1 port map( D => D(4), CK => clk, RN => n34, Q => Q(4),
                           QN => n62);
   Q_reg_3_inst : DFFR_X1 port map( D => D(3), CK => clk, RN => n34, Q => Q(3),
                           QN => n63);
   Q_reg_2_inst : DFFR_X1 port map( D => D(2), CK => clk, RN => n34, Q => Q(2),
                           QN => n64);
   Q_reg_1_inst : DFFR_X1 port map( D => D(1), CK => clk, RN => n34, Q => Q(1),
                           QN => n65);
   Q_reg_0_inst : DFFR_X1 port map( D => D(0), CK => clk, RN => n34, Q => Q(0),
                           QN => n66);
   U2 : INV_X2 port map( A => rst, ZN => n34);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity ff32_en_SIZE32_1 is

   port( D : in std_logic_vector (31 downto 0);  en, clk, rst : in std_logic;  
         Q : out std_logic_vector (31 downto 0));

end ff32_en_SIZE32_1;

architecture SYN_behavioral of ff32_en_SIZE32_1 is

   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_ff32_en_SIZE32_1
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal net199358, n32, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44
      , n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, 
      n59, n60, n61, n62, n63, n64, n65 : std_logic;

begin
   
   Q_reg_31_inst : DFFR_X1 port map( D => D(31), CK => net199358, RN => n32, Q 
                           => Q(31), QN => n34);
   Q_reg_30_inst : DFFR_X1 port map( D => D(30), CK => net199358, RN => n32, Q 
                           => Q(30), QN => n35);
   Q_reg_29_inst : DFFR_X1 port map( D => D(29), CK => net199358, RN => n32, Q 
                           => Q(29), QN => n36);
   Q_reg_28_inst : DFFR_X1 port map( D => D(28), CK => net199358, RN => n32, Q 
                           => Q(28), QN => n37);
   Q_reg_27_inst : DFFR_X1 port map( D => D(27), CK => net199358, RN => n32, Q 
                           => Q(27), QN => n38);
   Q_reg_26_inst : DFFR_X1 port map( D => D(26), CK => net199358, RN => n32, Q 
                           => Q(26), QN => n39);
   Q_reg_25_inst : DFFR_X1 port map( D => D(25), CK => net199358, RN => n32, Q 
                           => Q(25), QN => n40);
   Q_reg_24_inst : DFFR_X1 port map( D => D(24), CK => net199358, RN => n32, Q 
                           => Q(24), QN => n41);
   Q_reg_23_inst : DFFR_X1 port map( D => D(23), CK => net199358, RN => n32, Q 
                           => Q(23), QN => n42);
   Q_reg_22_inst : DFFR_X1 port map( D => D(22), CK => net199358, RN => n32, Q 
                           => Q(22), QN => n43);
   Q_reg_21_inst : DFFR_X1 port map( D => D(21), CK => net199358, RN => n32, Q 
                           => Q(21), QN => n44);
   Q_reg_20_inst : DFFR_X1 port map( D => D(20), CK => net199358, RN => n32, Q 
                           => Q(20), QN => n45);
   Q_reg_19_inst : DFFR_X1 port map( D => D(19), CK => net199358, RN => n32, Q 
                           => Q(19), QN => n46);
   Q_reg_18_inst : DFFR_X1 port map( D => D(18), CK => net199358, RN => n32, Q 
                           => Q(18), QN => n47);
   Q_reg_17_inst : DFFR_X1 port map( D => D(17), CK => net199358, RN => n32, Q 
                           => Q(17), QN => n48);
   Q_reg_16_inst : DFFR_X1 port map( D => D(16), CK => net199358, RN => n32, Q 
                           => Q(16), QN => n49);
   Q_reg_15_inst : DFFR_X1 port map( D => D(15), CK => net199358, RN => n32, Q 
                           => Q(15), QN => n50);
   Q_reg_14_inst : DFFR_X1 port map( D => D(14), CK => net199358, RN => n32, Q 
                           => Q(14), QN => n51);
   Q_reg_13_inst : DFFR_X1 port map( D => D(13), CK => net199358, RN => n32, Q 
                           => Q(13), QN => n52);
   Q_reg_12_inst : DFFR_X1 port map( D => D(12), CK => net199358, RN => n32, Q 
                           => Q(12), QN => n53);
   Q_reg_11_inst : DFFR_X1 port map( D => D(11), CK => net199358, RN => n32, Q 
                           => Q(11), QN => n54);
   Q_reg_10_inst : DFFR_X1 port map( D => D(10), CK => net199358, RN => n32, Q 
                           => Q(10), QN => n55);
   Q_reg_9_inst : DFFR_X1 port map( D => D(9), CK => net199358, RN => n32, Q =>
                           Q(9), QN => n56);
   Q_reg_8_inst : DFFR_X1 port map( D => D(8), CK => net199358, RN => n32, Q =>
                           Q(8), QN => n57);
   Q_reg_7_inst : DFFR_X1 port map( D => D(7), CK => net199358, RN => n32, Q =>
                           Q(7), QN => n58);
   Q_reg_6_inst : DFFR_X1 port map( D => D(6), CK => net199358, RN => n32, Q =>
                           Q(6), QN => n59);
   Q_reg_5_inst : DFFR_X1 port map( D => D(5), CK => net199358, RN => n32, Q =>
                           Q(5), QN => n60);
   Q_reg_4_inst : DFFR_X1 port map( D => D(4), CK => net199358, RN => n32, Q =>
                           Q(4), QN => n61);
   Q_reg_3_inst : DFFR_X1 port map( D => D(3), CK => net199358, RN => n32, Q =>
                           Q(3), QN => n62);
   Q_reg_2_inst : DFFR_X1 port map( D => D(2), CK => net199358, RN => n32, Q =>
                           Q(2), QN => n63);
   Q_reg_1_inst : DFFR_X1 port map( D => D(1), CK => net199358, RN => n32, Q =>
                           Q(1), QN => n64);
   Q_reg_0_inst : DFFR_X1 port map( D => D(0), CK => net199358, RN => n32, Q =>
                           Q(0), QN => n65);
   clk_gate_Q_reg : SNPS_CLOCK_GATE_HIGH_ff32_en_SIZE32_1 port map( CLK => clk,
                           EN => en, ENCLK => net199358);
   U2 : INV_X2 port map( A => rst, ZN => n32);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity mux41_MUX_SIZE32_2 is

   port( IN0, IN1, IN2, IN3 : in std_logic_vector (31 downto 0);  CTRL : in 
         std_logic_vector (1 downto 0);  OUT1 : out std_logic_vector (31 downto
         0));

end mux41_MUX_SIZE32_2;

architecture SYN_bhe of mux41_MUX_SIZE32_2 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n69, n70, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, 
      n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96
      , n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142 : std_logic;

begin
   
   U51 : AOI22_X1 port map( A1 => n74, A2 => IN1(23), B1 => n72, B2 => IN0(23),
                           ZN => n106);
   U50 : AOI22_X1 port map( A1 => n75, A2 => IN3(23), B1 => n1, B2 => IN2(23), 
                           ZN => n105);
   U49 : NAND2_X1 port map( A1 => n106, A2 => n105, ZN => OUT1(23));
   U60 : AOI22_X1 port map( A1 => n74, A2 => IN1(20), B1 => n72, B2 => IN0(20),
                           ZN => n100);
   U59 : AOI22_X1 port map( A1 => n75, A2 => IN3(20), B1 => n1, B2 => IN2(20), 
                           ZN => n99);
   U58 : NAND2_X1 port map( A1 => n100, A2 => n99, ZN => OUT1(20));
   U57 : AOI22_X1 port map( A1 => n74, A2 => IN1(21), B1 => n72, B2 => IN0(21),
                           ZN => n102);
   U56 : AOI22_X1 port map( A1 => n75, A2 => IN3(21), B1 => n1, B2 => IN2(21), 
                           ZN => n101);
   U55 : NAND2_X1 port map( A1 => n102, A2 => n101, ZN => OUT1(21));
   U54 : AOI22_X1 port map( A1 => n74, A2 => IN1(22), B1 => n72, B2 => IN0(22),
                           ZN => n104);
   U53 : AOI22_X1 port map( A1 => n75, A2 => IN3(22), B1 => n1, B2 => IN2(22), 
                           ZN => n103);
   U52 : NAND2_X1 port map( A1 => n104, A2 => n103, ZN => OUT1(22));
   U78 : AOI22_X1 port map( A1 => n73, A2 => IN1(15), B1 => n137, B2 => IN0(15)
                           , ZN => n88);
   U81 : AOI22_X1 port map( A1 => n73, A2 => IN1(14), B1 => n137, B2 => IN0(14)
                           , ZN => n86);
   U79 : NAND2_X1 port map( A1 => n86, A2 => n85, ZN => OUT1(14));
   U84 : AOI22_X1 port map( A1 => n73, A2 => IN1(13), B1 => n137, B2 => IN0(13)
                           , ZN => n84);
   U82 : NAND2_X1 port map( A1 => n84, A2 => n83, ZN => OUT1(13));
   U87 : AOI22_X1 port map( A1 => n73, A2 => IN1(12), B1 => n137, B2 => IN0(12)
                           , ZN => n82);
   U93 : AOI22_X1 port map( A1 => n73, A2 => IN1(10), B1 => n137, B2 => IN0(10)
                           , ZN => n78);
   U91 : NAND2_X1 port map( A1 => n78, A2 => n77, ZN => OUT1(10));
   U90 : AOI22_X1 port map( A1 => n73, A2 => IN1(11), B1 => n137, B2 => IN0(11)
                           , ZN => n80);
   U88 : NAND2_X1 port map( A1 => n80, A2 => n79, ZN => OUT1(11));
   U3 : AOI22_X1 port map( A1 => n74, A2 => IN1(9), B1 => n72, B2 => IN0(9), ZN
                           => n142);
   U2 : AOI22_X1 port map( A1 => n140, A2 => IN3(9), B1 => n1, B2 => IN2(9), ZN
                           => n141);
   U6 : AOI22_X1 port map( A1 => n74, A2 => IN1(8), B1 => n72, B2 => IN0(8), ZN
                           => n136);
   U5 : AOI22_X1 port map( A1 => n140, A2 => IN3(8), B1 => n1, B2 => IN2(8), ZN
                           => n135);
   U63 : AOI22_X1 port map( A1 => n73, A2 => IN1(1), B1 => n72, B2 => IN0(1), 
                           ZN => n98);
   U30 : AOI22_X1 port map( A1 => n74, A2 => IN1(2), B1 => n72, B2 => IN0(2), 
                           ZN => n120);
   U29 : AOI22_X1 port map( A1 => n75, A2 => IN3(2), B1 => n1, B2 => IN2(2), ZN
                           => n119);
   U21 : AOI22_X1 port map( A1 => n74, A2 => IN1(3), B1 => n72, B2 => IN0(3), 
                           ZN => n126);
   U20 : AOI22_X1 port map( A1 => n140, A2 => IN3(3), B1 => n1, B2 => IN2(3), 
                           ZN => n125);
   U9 : AOI22_X1 port map( A1 => n74, A2 => IN1(7), B1 => n72, B2 => IN0(7), ZN
                           => n134);
   U8 : AOI22_X1 port map( A1 => n140, A2 => IN3(7), B1 => n1, B2 => IN2(7), ZN
                           => n133);
   U12 : AOI22_X1 port map( A1 => n74, A2 => IN1(6), B1 => n72, B2 => IN0(6), 
                           ZN => n132);
   U11 : AOI22_X1 port map( A1 => n140, A2 => IN3(6), B1 => n1, B2 => IN2(6), 
                           ZN => n131);
   U15 : AOI22_X1 port map( A1 => n74, A2 => IN1(5), B1 => n72, B2 => IN0(5), 
                           ZN => n130);
   U14 : AOI22_X1 port map( A1 => n140, A2 => IN3(5), B1 => n1, B2 => IN2(5), 
                           ZN => n129);
   U18 : AOI22_X1 port map( A1 => n74, A2 => IN1(4), B1 => n72, B2 => IN0(4), 
                           ZN => n128);
   U17 : AOI22_X1 port map( A1 => n140, A2 => IN3(4), B1 => n1, B2 => IN2(4), 
                           ZN => n127);
   U66 : AOI22_X1 port map( A1 => n73, A2 => IN1(19), B1 => n137, B2 => IN0(19)
                           , ZN => n96);
   U64 : NAND2_X1 port map( A1 => n96, A2 => n95, ZN => OUT1(19));
   U69 : AOI22_X1 port map( A1 => n73, A2 => IN1(18), B1 => n137, B2 => IN0(18)
                           , ZN => n94);
   U67 : NAND2_X1 port map( A1 => n94, A2 => n93, ZN => OUT1(18));
   U72 : AOI22_X1 port map( A1 => n73, A2 => IN1(17), B1 => n137, B2 => IN0(17)
                           , ZN => n92);
   U70 : NAND2_X1 port map( A1 => n92, A2 => n91, ZN => OUT1(17));
   U75 : AOI22_X1 port map( A1 => n73, A2 => IN1(16), B1 => n137, B2 => IN0(16)
                           , ZN => n90);
   U73 : NAND2_X1 port map( A1 => n90, A2 => n89, ZN => OUT1(16));
   U39 : AOI22_X1 port map( A1 => n74, A2 => IN1(27), B1 => n72, B2 => IN0(27),
                           ZN => n114);
   U38 : AOI22_X1 port map( A1 => n75, A2 => IN3(27), B1 => n1, B2 => IN2(27), 
                           ZN => n113);
   U37 : NAND2_X1 port map( A1 => n114, A2 => n113, ZN => OUT1(27));
   U48 : AOI22_X1 port map( A1 => n74, A2 => IN1(24), B1 => n72, B2 => IN0(24),
                           ZN => n108);
   U47 : AOI22_X1 port map( A1 => n75, A2 => IN3(24), B1 => n1, B2 => IN2(24), 
                           ZN => n107);
   U46 : NAND2_X1 port map( A1 => n108, A2 => n107, ZN => OUT1(24));
   U45 : AOI22_X1 port map( A1 => n74, A2 => IN1(25), B1 => n137, B2 => IN0(25)
                           , ZN => n110);
   U44 : AOI22_X1 port map( A1 => n75, A2 => IN3(25), B1 => n1, B2 => IN2(25), 
                           ZN => n109);
   U43 : NAND2_X1 port map( A1 => n110, A2 => n109, ZN => OUT1(25));
   U42 : AOI22_X1 port map( A1 => n74, A2 => IN1(26), B1 => n72, B2 => IN0(26),
                           ZN => n112);
   U41 : AOI22_X1 port map( A1 => n75, A2 => IN3(26), B1 => n1, B2 => IN2(26), 
                           ZN => n111);
   U40 : NAND2_X1 port map( A1 => n112, A2 => n111, ZN => OUT1(26));
   U33 : AOI22_X1 port map( A1 => n74, A2 => IN1(29), B1 => n72, B2 => IN0(29),
                           ZN => n118);
   U32 : AOI22_X1 port map( A1 => n75, A2 => IN3(29), B1 => n1, B2 => IN2(29), 
                           ZN => n117);
   U31 : NAND2_X1 port map( A1 => n118, A2 => n117, ZN => OUT1(29));
   U36 : AOI22_X1 port map( A1 => n74, A2 => IN1(28), B1 => n72, B2 => IN0(28),
                           ZN => n116);
   U35 : AOI22_X1 port map( A1 => n75, A2 => IN3(28), B1 => n1, B2 => IN2(28), 
                           ZN => n115);
   U34 : NAND2_X1 port map( A1 => n116, A2 => n115, ZN => OUT1(28));
   U27 : AOI22_X1 port map( A1 => n74, A2 => IN1(30), B1 => n72, B2 => IN0(30),
                           ZN => n122);
   U26 : AOI22_X1 port map( A1 => n75, A2 => IN3(30), B1 => n1, B2 => IN2(30), 
                           ZN => n121);
   U25 : NAND2_X1 port map( A1 => n122, A2 => n121, ZN => OUT1(30));
   U24 : AOI22_X1 port map( A1 => n74, A2 => IN1(31), B1 => n72, B2 => IN0(31),
                           ZN => n124);
   U23 : AOI22_X1 port map( A1 => n140, A2 => IN3(31), B1 => n1, B2 => IN2(31),
                           ZN => n123);
   U85 : NAND2_X1 port map( A1 => n82, A2 => n81, ZN => OUT1(12));
   U1 : NAND2_X1 port map( A1 => n142, A2 => n141, ZN => OUT1(9));
   U4 : NAND2_X1 port map( A1 => n136, A2 => n135, ZN => OUT1(8));
   U61 : NAND2_X1 port map( A1 => n98, A2 => n97, ZN => OUT1(1));
   U28 : NAND2_X1 port map( A1 => n120, A2 => n119, ZN => OUT1(2));
   U19 : NAND2_X1 port map( A1 => n126, A2 => n125, ZN => OUT1(3));
   U7 : NAND2_X1 port map( A1 => n134, A2 => n133, ZN => OUT1(7));
   U10 : NAND2_X1 port map( A1 => n132, A2 => n131, ZN => OUT1(6));
   U13 : NAND2_X1 port map( A1 => n130, A2 => n129, ZN => OUT1(5));
   U16 : NAND2_X1 port map( A1 => n128, A2 => n127, ZN => OUT1(4));
   U76 : NAND2_X1 port map( A1 => n88, A2 => n87, ZN => OUT1(15));
   U22 : NAND2_X1 port map( A1 => n124, A2 => n123, ZN => OUT1(31));
   U62 : AND2_X1 port map( A1 => CTRL(0), A2 => CTRL(1), ZN => n140);
   U65 : NOR2_X2 port map( A1 => CTRL(0), A2 => CTRL(1), ZN => n137);
   U68 : BUF_X2 port map( A => n137, Z => n72);
   U71 : NOR2_X2 port map( A1 => CTRL(0), A2 => n76, ZN => n139);
   U74 : BUF_X2 port map( A => n139, Z => n1);
   U77 : INV_X1 port map( A => CTRL(1), ZN => n76);
   U80 : AND2_X1 port map( A1 => n76, A2 => CTRL(0), ZN => n138);
   U83 : BUF_X2 port map( A => n140, Z => n75);
   U86 : BUF_X1 port map( A => n138, Z => n74);
   U89 : BUF_X1 port map( A => n138, Z => n73);
   U92 : NAND3_X1 port map( A1 => n69, A2 => n2, A3 => n70, ZN => OUT1(0));
   U94 : NAND2_X1 port map( A1 => n73, A2 => IN1(0), ZN => n2);
   U95 : NAND2_X1 port map( A1 => n139, A2 => IN2(0), ZN => n69);
   U96 : NAND2_X1 port map( A1 => n137, A2 => IN0(0), ZN => n70);
   U97 : AOI22_X1 port map( A1 => n75, A2 => IN3(16), B1 => n139, B2 => IN2(16)
                           , ZN => n89);
   U98 : AOI22_X1 port map( A1 => n75, A2 => IN3(18), B1 => n139, B2 => IN2(18)
                           , ZN => n93);
   U99 : AOI22_X1 port map( A1 => n75, A2 => IN3(12), B1 => n139, B2 => IN2(12)
                           , ZN => n81);
   U100 : AOI22_X1 port map( A1 => n75, A2 => IN3(10), B1 => n139, B2 => 
                           IN2(10), ZN => n77);
   U101 : AOI22_X1 port map( A1 => n75, A2 => IN3(14), B1 => n139, B2 => 
                           IN2(14), ZN => n85);
   U102 : AOI22_X1 port map( A1 => n75, A2 => IN3(17), B1 => n139, B2 => 
                           IN2(17), ZN => n91);
   U103 : AOI22_X1 port map( A1 => n75, A2 => IN3(19), B1 => n139, B2 => 
                           IN2(19), ZN => n95);
   U104 : AOI22_X1 port map( A1 => n75, A2 => IN3(11), B1 => n139, B2 => 
                           IN2(11), ZN => n79);
   U105 : AOI22_X1 port map( A1 => n75, A2 => IN3(13), B1 => n139, B2 => 
                           IN2(13), ZN => n83);
   U106 : AOI22_X1 port map( A1 => n75, A2 => IN3(15), B1 => n139, B2 => 
                           IN2(15), ZN => n87);
   U107 : AOI22_X1 port map( A1 => n75, A2 => IN3(1), B1 => n1, B2 => IN2(1), 
                           ZN => n97);

end SYN_bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity mux41_MUX_SIZE32_1 is

   port( IN0, IN1, IN2, IN3 : in std_logic_vector (31 downto 0);  CTRL : in 
         std_logic_vector (1 downto 0);  OUT1 : out std_logic_vector (31 downto
         0));

end mux41_MUX_SIZE32_1;

architecture SYN_bhe of mux41_MUX_SIZE32_1 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X3
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, 
      n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94
      , n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107
      , n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
      n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, 
      n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, 
      n144, n145, n146 : std_logic;

begin
   
   U58 : NAND2_X1 port map( A1 => n106, A2 => n105, ZN => OUT1(20));
   U49 : NAND2_X1 port map( A1 => n112, A2 => n111, ZN => OUT1(23));
   U10 : NAND2_X1 port map( A1 => n138, A2 => n137, ZN => OUT1(6));
   U46 : NAND2_X1 port map( A1 => n114, A2 => n113, ZN => OUT1(24));
   U40 : NAND2_X1 port map( A1 => n118, A2 => n117, ZN => OUT1(26));
   U37 : NAND2_X1 port map( A1 => n120, A2 => n119, ZN => OUT1(27));
   U31 : NAND2_X1 port map( A1 => n124, A2 => n123, ZN => OUT1(29));
   U25 : NAND2_X1 port map( A1 => n128, A2 => n127, ZN => OUT1(30));
   U22 : NAND2_X1 port map( A1 => n130, A2 => n129, ZN => OUT1(31));
   U1 : BUF_X2 port map( A => n144, Z => n82);
   U2 : BUF_X2 port map( A => n143, Z => n79);
   U3 : AND2_X2 port map( A1 => CTRL(1), A2 => n8, ZN => n143);
   U4 : BUF_X2 port map( A => n1, Z => n2);
   U5 : BUF_X2 port map( A => n69, Z => n75);
   U6 : BUF_X2 port map( A => n69, Z => n76);
   U7 : BUF_X2 port map( A => n143, Z => n78);
   U8 : BUF_X2 port map( A => n1, Z => n73);
   U9 : CLKBUF_X3 port map( A => n144, Z => n81);
   U11 : BUF_X2 port map( A => n1, Z => n74);
   U12 : BUF_X2 port map( A => n143, Z => n77);
   U13 : INV_X1 port map( A => CTRL(0), ZN => n8);
   U14 : AND2_X1 port map( A1 => CTRL(0), A2 => CTRL(1), ZN => n144);
   U15 : NOR2_X1 port map( A1 => n8, A2 => CTRL(1), ZN => n69);
   U16 : BUF_X1 port map( A => n144, Z => n80);
   U17 : NOR2_X1 port map( A1 => CTRL(1), A2 => CTRL(0), ZN => n1);
   U18 : NAND2_X1 port map( A1 => n2, A2 => IN0(0), ZN => n71);
   U19 : AOI22_X1 port map( A1 => n75, A2 => IN1(2), B1 => n2, B2 => IN0(2), ZN
                           => n126);
   U20 : AOI22_X1 port map( A1 => n76, A2 => IN1(30), B1 => n2, B2 => IN0(30), 
                           ZN => n128);
   U21 : AOI22_X1 port map( A1 => n76, A2 => IN1(29), B1 => n2, B2 => IN0(29), 
                           ZN => n124);
   U23 : AOI22_X1 port map( A1 => n76, A2 => IN1(20), B1 => n2, B2 => IN0(20), 
                           ZN => n106);
   U24 : AOI22_X1 port map( A1 => n76, A2 => IN1(26), B1 => n2, B2 => IN0(26), 
                           ZN => n118);
   U26 : AOI22_X1 port map( A1 => n75, A2 => IN1(14), B1 => n2, B2 => IN0(14), 
                           ZN => n92);
   U27 : AOI22_X1 port map( A1 => n76, A2 => IN1(18), B1 => n2, B2 => IN0(18), 
                           ZN => n100);
   U28 : AOI22_X1 port map( A1 => n76, A2 => IN1(19), B1 => n2, B2 => IN0(19), 
                           ZN => n102);
   U29 : AOI22_X1 port map( A1 => n75, A2 => IN1(17), B1 => n2, B2 => IN0(17), 
                           ZN => n98);
   U30 : AOI22_X1 port map( A1 => n76, A2 => IN1(16), B1 => n2, B2 => IN0(16), 
                           ZN => n96);
   U32 : NAND2_X1 port map( A1 => n69, A2 => IN1(0), ZN => n70);
   U33 : AOI22_X1 port map( A1 => n75, A2 => IN1(5), B1 => n74, B2 => IN0(5), 
                           ZN => n136);
   U34 : AOI22_X1 port map( A1 => n75, A2 => IN1(9), B1 => n74, B2 => IN0(9), 
                           ZN => n146);
   U35 : AOI22_X1 port map( A1 => n76, A2 => IN1(8), B1 => n73, B2 => IN0(8), 
                           ZN => n142);
   U36 : NAND3_X1 port map( A1 => n70, A2 => n72, A3 => n71, ZN => OUT1(0));
   U38 : NAND2_X1 port map( A1 => n78, A2 => IN2(0), ZN => n72);
   U39 : AOI22_X1 port map( A1 => n76, A2 => IN1(22), B1 => n74, B2 => IN0(22),
                           ZN => n110);
   U41 : AOI22_X1 port map( A1 => n76, A2 => IN1(24), B1 => n74, B2 => IN0(24),
                           ZN => n114);
   U42 : AOI22_X1 port map( A1 => n76, A2 => IN1(27), B1 => n73, B2 => IN0(27),
                           ZN => n120);
   U43 : AOI22_X1 port map( A1 => n75, A2 => IN1(4), B1 => n74, B2 => IN0(4), 
                           ZN => n134);
   U44 : AOI22_X1 port map( A1 => n75, A2 => IN1(21), B1 => n73, B2 => IN0(21),
                           ZN => n108);
   U45 : AOI22_X1 port map( A1 => n75, A2 => IN1(7), B1 => n73, B2 => IN0(7), 
                           ZN => n140);
   U47 : AOI22_X1 port map( A1 => n75, A2 => IN1(3), B1 => n74, B2 => IN0(3), 
                           ZN => n132);
   U48 : NAND2_X1 port map( A1 => n96, A2 => n95, ZN => OUT1(16));
   U50 : NAND2_X1 port map( A1 => n122, A2 => n121, ZN => OUT1(28));
   U51 : NAND2_X1 port map( A1 => n102, A2 => n101, ZN => OUT1(19));
   U52 : NAND2_X1 port map( A1 => n116, A2 => n115, ZN => OUT1(25));
   U53 : AOI22_X1 port map( A1 => n76, A2 => IN1(31), B1 => n74, B2 => IN0(31),
                           ZN => n130);
   U54 : AOI22_X1 port map( A1 => n76, A2 => IN1(6), B1 => n73, B2 => IN0(6), 
                           ZN => n138);
   U55 : AOI22_X1 port map( A1 => n76, A2 => IN1(28), B1 => n73, B2 => IN0(28),
                           ZN => n122);
   U56 : AOI22_X1 port map( A1 => n76, A2 => IN1(25), B1 => n73, B2 => IN0(25),
                           ZN => n116);
   U57 : AOI22_X1 port map( A1 => n76, A2 => IN1(23), B1 => n74, B2 => IN0(23),
                           ZN => n112);
   U59 : NAND2_X1 port map( A1 => n92, A2 => n91, ZN => OUT1(14));
   U60 : NAND2_X1 port map( A1 => n126, A2 => n125, ZN => OUT1(2));
   U61 : NAND2_X1 port map( A1 => n88, A2 => n87, ZN => OUT1(12));
   U62 : NAND2_X1 port map( A1 => n142, A2 => n141, ZN => OUT1(8));
   U63 : NAND2_X1 port map( A1 => n86, A2 => n85, ZN => OUT1(11));
   U64 : NAND2_X1 port map( A1 => n110, A2 => n109, ZN => OUT1(22));
   U65 : NAND2_X1 port map( A1 => n140, A2 => n139, ZN => OUT1(7));
   U66 : NAND2_X1 port map( A1 => n134, A2 => n133, ZN => OUT1(4));
   U67 : NAND2_X1 port map( A1 => n94, A2 => n93, ZN => OUT1(15));
   U68 : NAND2_X1 port map( A1 => n100, A2 => n99, ZN => OUT1(18));
   U69 : NAND2_X1 port map( A1 => n135, A2 => n136, ZN => OUT1(5));
   U70 : NAND2_X1 port map( A1 => n104, A2 => n103, ZN => OUT1(1));
   U71 : NAND2_X1 port map( A1 => n84, A2 => n83, ZN => OUT1(10));
   U72 : AOI22_X1 port map( A1 => n76, A2 => IN1(12), B1 => n74, B2 => IN0(12),
                           ZN => n88);
   U73 : AOI22_X1 port map( A1 => n75, A2 => IN1(13), B1 => n74, B2 => IN0(13),
                           ZN => n90);
   U74 : AOI22_X1 port map( A1 => n76, A2 => IN1(1), B1 => n73, B2 => IN0(1), 
                           ZN => n104);
   U75 : AOI22_X1 port map( A1 => n75, A2 => IN1(11), B1 => n73, B2 => IN0(11),
                           ZN => n86);
   U76 : AOI22_X1 port map( A1 => n75, A2 => IN1(15), B1 => n73, B2 => IN0(15),
                           ZN => n94);
   U77 : AOI22_X1 port map( A1 => n76, A2 => IN1(10), B1 => n74, B2 => IN0(10),
                           ZN => n84);
   U78 : NAND2_X1 port map( A1 => n98, A2 => n97, ZN => OUT1(17));
   U79 : NAND2_X1 port map( A1 => n108, A2 => n107, ZN => OUT1(21));
   U80 : AOI22_X1 port map( A1 => n82, A2 => IN3(31), B1 => n79, B2 => IN2(31),
                           ZN => n129);
   U81 : AOI22_X1 port map( A1 => n82, A2 => IN3(8), B1 => n79, B2 => IN2(8), 
                           ZN => n141);
   U82 : AOI22_X1 port map( A1 => n82, A2 => IN3(9), B1 => n78, B2 => IN2(9), 
                           ZN => n145);
   U83 : AOI22_X1 port map( A1 => n82, A2 => IN3(4), B1 => n79, B2 => IN2(4), 
                           ZN => n133);
   U84 : AOI22_X1 port map( A1 => n82, A2 => IN3(3), B1 => n79, B2 => IN2(3), 
                           ZN => n131);
   U85 : AOI22_X1 port map( A1 => n82, A2 => IN3(5), B1 => n79, B2 => IN2(5), 
                           ZN => n135);
   U86 : AOI22_X1 port map( A1 => n82, A2 => IN3(7), B1 => n77, B2 => IN2(7), 
                           ZN => n139);
   U87 : AOI22_X1 port map( A1 => n82, A2 => IN3(6), B1 => n79, B2 => IN2(6), 
                           ZN => n137);
   U88 : NAND2_X1 port map( A1 => n89, A2 => n90, ZN => OUT1(13));
   U89 : AOI22_X1 port map( A1 => n81, A2 => IN3(30), B1 => n77, B2 => IN2(30),
                           ZN => n127);
   U90 : AOI22_X1 port map( A1 => n81, A2 => IN3(29), B1 => n77, B2 => IN2(29),
                           ZN => n123);
   U91 : AOI22_X1 port map( A1 => n81, A2 => IN3(24), B1 => n79, B2 => IN2(24),
                           ZN => n113);
   U92 : AOI22_X1 port map( A1 => n81, A2 => IN3(27), B1 => n77, B2 => IN2(27),
                           ZN => n119);
   U93 : AOI22_X1 port map( A1 => n81, A2 => IN3(26), B1 => n143, B2 => IN2(26)
                           , ZN => n117);
   U94 : AOI22_X1 port map( A1 => n81, A2 => IN3(28), B1 => n79, B2 => IN2(28),
                           ZN => n121);
   U95 : AOI22_X1 port map( A1 => n81, A2 => IN3(20), B1 => n77, B2 => IN2(20),
                           ZN => n105);
   U96 : AOI22_X1 port map( A1 => n81, A2 => IN3(25), B1 => n79, B2 => IN2(25),
                           ZN => n115);
   U97 : AOI22_X1 port map( A1 => n81, A2 => IN3(23), B1 => n77, B2 => IN2(23),
                           ZN => n111);
   U98 : AOI22_X1 port map( A1 => n81, A2 => IN3(22), B1 => n79, B2 => IN2(22),
                           ZN => n109);
   U99 : AOI22_X1 port map( A1 => n81, A2 => IN3(2), B1 => n77, B2 => IN2(2), 
                           ZN => n125);
   U100 : AOI22_X1 port map( A1 => n81, A2 => IN3(21), B1 => n79, B2 => IN2(21)
                           , ZN => n107);
   U101 : NAND2_X1 port map( A1 => n131, A2 => n132, ZN => OUT1(3));
   U102 : NAND2_X1 port map( A1 => n146, A2 => n145, ZN => OUT1(9));
   U103 : AOI22_X1 port map( A1 => n80, A2 => IN3(16), B1 => n77, B2 => IN2(16)
                           , ZN => n95);
   U104 : AOI22_X1 port map( A1 => n80, A2 => IN3(19), B1 => n79, B2 => IN2(19)
                           , ZN => n101);
   U105 : AOI22_X1 port map( A1 => n80, A2 => IN3(12), B1 => n77, B2 => IN2(12)
                           , ZN => n87);
   U106 : AOI22_X1 port map( A1 => n80, A2 => IN3(18), B1 => n77, B2 => IN2(18)
                           , ZN => n99);
   U107 : AOI22_X1 port map( A1 => n80, A2 => IN3(11), B1 => n78, B2 => IN2(11)
                           , ZN => n85);
   U108 : AOI22_X1 port map( A1 => n80, A2 => IN3(10), B1 => n79, B2 => IN2(10)
                           , ZN => n83);
   U109 : AOI22_X1 port map( A1 => n80, A2 => IN3(17), B1 => n77, B2 => IN2(17)
                           , ZN => n97);
   U110 : AOI22_X1 port map( A1 => n80, A2 => IN3(14), B1 => n77, B2 => IN2(14)
                           , ZN => n91);
   U111 : AOI22_X1 port map( A1 => n80, A2 => IN3(15), B1 => n78, B2 => IN2(15)
                           , ZN => n93);
   U112 : AOI22_X1 port map( A1 => n80, A2 => IN3(13), B1 => n77, B2 => IN2(13)
                           , ZN => n89);
   U113 : AOI22_X1 port map( A1 => n80, A2 => IN3(1), B1 => n77, B2 => IN2(1), 
                           ZN => n103);

end SYN_bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity mux21_4 is

   port( IN0, IN1 : in std_logic_vector (31 downto 0);  CTRL : in std_logic;  
         OUT1 : out std_logic_vector (31 downto 0));

end mux21_4;

architecture SYN_Bhe of mux21_4 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => IN0(9), B => IN1(9), S => CTRL, Z => OUT1(9));
   U2 : MUX2_X1 port map( A => IN0(8), B => IN1(8), S => CTRL, Z => OUT1(8));
   U3 : MUX2_X1 port map( A => IN0(7), B => IN1(7), S => CTRL, Z => OUT1(7));
   U4 : MUX2_X1 port map( A => IN0(6), B => IN1(6), S => CTRL, Z => OUT1(6));
   U5 : MUX2_X1 port map( A => IN0(5), B => IN1(5), S => CTRL, Z => OUT1(5));
   U6 : MUX2_X1 port map( A => IN0(4), B => IN1(4), S => CTRL, Z => OUT1(4));
   U7 : MUX2_X1 port map( A => IN0(3), B => IN1(3), S => CTRL, Z => OUT1(3));
   U8 : MUX2_X1 port map( A => IN0(31), B => IN1(31), S => CTRL, Z => OUT1(31))
                           ;
   U9 : MUX2_X1 port map( A => IN0(30), B => IN1(30), S => CTRL, Z => OUT1(30))
                           ;
   U10 : MUX2_X1 port map( A => IN0(2), B => IN1(2), S => CTRL, Z => OUT1(2));
   U11 : MUX2_X1 port map( A => IN0(29), B => IN1(29), S => CTRL, Z => OUT1(29)
                           );
   U12 : MUX2_X1 port map( A => IN0(28), B => IN1(28), S => CTRL, Z => OUT1(28)
                           );
   U13 : MUX2_X1 port map( A => IN0(27), B => IN1(27), S => CTRL, Z => OUT1(27)
                           );
   U14 : MUX2_X1 port map( A => IN0(26), B => IN1(26), S => CTRL, Z => OUT1(26)
                           );
   U15 : MUX2_X1 port map( A => IN0(25), B => IN1(25), S => CTRL, Z => OUT1(25)
                           );
   U16 : MUX2_X1 port map( A => IN0(24), B => IN1(24), S => CTRL, Z => OUT1(24)
                           );
   U17 : MUX2_X1 port map( A => IN0(23), B => IN1(23), S => CTRL, Z => OUT1(23)
                           );
   U18 : MUX2_X1 port map( A => IN0(22), B => IN1(22), S => CTRL, Z => OUT1(22)
                           );
   U19 : MUX2_X1 port map( A => IN0(21), B => IN1(21), S => CTRL, Z => OUT1(21)
                           );
   U20 : MUX2_X1 port map( A => IN0(20), B => IN1(20), S => CTRL, Z => OUT1(20)
                           );
   U21 : MUX2_X1 port map( A => IN0(1), B => IN1(1), S => CTRL, Z => OUT1(1));
   U22 : MUX2_X1 port map( A => IN0(19), B => IN1(19), S => CTRL, Z => OUT1(19)
                           );
   U23 : MUX2_X1 port map( A => IN0(18), B => IN1(18), S => CTRL, Z => OUT1(18)
                           );
   U24 : MUX2_X1 port map( A => IN0(17), B => IN1(17), S => CTRL, Z => OUT1(17)
                           );
   U25 : MUX2_X1 port map( A => IN0(16), B => IN1(16), S => CTRL, Z => OUT1(16)
                           );
   U26 : MUX2_X1 port map( A => IN0(15), B => IN1(15), S => CTRL, Z => OUT1(15)
                           );
   U27 : MUX2_X1 port map( A => IN0(14), B => IN1(14), S => CTRL, Z => OUT1(14)
                           );
   U28 : MUX2_X1 port map( A => IN0(13), B => IN1(13), S => CTRL, Z => OUT1(13)
                           );
   U29 : MUX2_X1 port map( A => IN0(12), B => IN1(12), S => CTRL, Z => OUT1(12)
                           );
   U30 : MUX2_X1 port map( A => IN0(11), B => IN1(11), S => CTRL, Z => OUT1(11)
                           );
   U31 : MUX2_X1 port map( A => IN0(10), B => IN1(10), S => CTRL, Z => OUT1(10)
                           );
   U32 : MUX2_X1 port map( A => IN0(0), B => IN1(0), S => CTRL, Z => OUT1(0));

end SYN_Bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity mux21_3 is

   port( IN0, IN1 : in std_logic_vector (31 downto 0);  CTRL : in std_logic;  
         OUT1 : out std_logic_vector (31 downto 0));

end mux21_3;

architecture SYN_Bhe of mux21_3 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X2
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n4, n5, n6, n7, n8 : std_logic;

begin
   
   U2 : MUX2_X1 port map( A => IN0(8), B => IN1(8), S => CTRL, Z => OUT1(8));
   U8 : MUX2_X1 port map( A => IN0(31), B => IN1(31), S => CTRL, Z => OUT1(31))
                           ;
   U9 : MUX2_X1 port map( A => IN0(30), B => IN1(30), S => CTRL, Z => OUT1(30))
                           ;
   U11 : MUX2_X1 port map( A => IN0(29), B => IN1(29), S => CTRL, Z => OUT1(29)
                           );
   U13 : MUX2_X1 port map( A => IN0(27), B => IN1(27), S => CTRL, Z => OUT1(27)
                           );
   U14 : MUX2_X1 port map( A => IN0(26), B => IN1(26), S => CTRL, Z => OUT1(26)
                           );
   U15 : MUX2_X1 port map( A => IN0(25), B => IN1(25), S => CTRL, Z => OUT1(25)
                           );
   U16 : MUX2_X1 port map( A => IN0(24), B => IN1(24), S => CTRL, Z => OUT1(24)
                           );
   U17 : MUX2_X1 port map( A => IN0(23), B => IN1(23), S => CTRL, Z => OUT1(23)
                           );
   U18 : MUX2_X1 port map( A => IN0(22), B => IN1(22), S => CTRL, Z => OUT1(22)
                           );
   U20 : MUX2_X1 port map( A => IN0(20), B => IN1(20), S => CTRL, Z => OUT1(20)
                           );
   U22 : MUX2_X1 port map( A => IN0(19), B => IN1(19), S => CTRL, Z => OUT1(19)
                           );
   U23 : MUX2_X1 port map( A => IN0(18), B => IN1(18), S => CTRL, Z => OUT1(18)
                           );
   U24 : MUX2_X1 port map( A => IN0(17), B => IN1(17), S => CTRL, Z => OUT1(17)
                           );
   U25 : MUX2_X1 port map( A => IN0(16), B => IN1(16), S => CTRL, Z => OUT1(16)
                           );
   U1 : MUX2_X1 port map( A => IN0(4), B => IN1(4), S => CTRL, Z => OUT1(4));
   U3 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => OUT1(10));
   U4 : MUX2_X1 port map( A => IN0(6), B => IN1(6), S => CTRL, Z => OUT1(6));
   U5 : NAND2_X1 port map( A1 => IN0(9), A2 => n2, ZN => n3);
   U6 : NAND2_X1 port map( A1 => IN1(9), A2 => CTRL, ZN => n4);
   U7 : NAND2_X2 port map( A1 => n3, A2 => n4, ZN => OUT1(9));
   U10 : INV_X1 port map( A => CTRL, ZN => n2);
   U12 : NAND2_X1 port map( A1 => IN0(10), A2 => n2, ZN => n5);
   U19 : NAND2_X1 port map( A1 => IN1(10), A2 => CTRL, ZN => n6);
   U21 : MUX2_X2 port map( A => IN0(2), B => IN1(2), S => CTRL, Z => OUT1(2));
   U26 : MUX2_X1 port map( A => IN0(15), B => IN1(15), S => CTRL, Z => OUT1(15)
                           );
   U27 : MUX2_X1 port map( A => IN0(11), B => IN1(11), S => CTRL, Z => OUT1(11)
                           );
   U28 : MUX2_X1 port map( A => IN0(13), B => IN1(13), S => CTRL, Z => OUT1(13)
                           );
   U29 : MUX2_X1 port map( A => IN0(28), B => IN1(28), S => CTRL, Z => OUT1(28)
                           );
   U30 : MUX2_X1 port map( A => IN0(1), B => IN1(1), S => CTRL, Z => OUT1(1));
   U31 : MUX2_X1 port map( A => IN0(12), B => IN1(12), S => CTRL, Z => OUT1(12)
                           );
   U32 : MUX2_X1 port map( A => IN0(14), B => IN1(14), S => CTRL, Z => OUT1(14)
                           );
   U33 : MUX2_X1 port map( A => IN0(21), B => IN1(21), S => CTRL, Z => OUT1(21)
                           );
   U34 : NAND2_X1 port map( A1 => n7, A2 => n8, ZN => OUT1(0));
   U35 : NAND2_X1 port map( A1 => IN1(0), A2 => CTRL, ZN => n8);
   U36 : NAND2_X1 port map( A1 => IN0(0), A2 => n2, ZN => n7);
   U37 : MUX2_X1 port map( A => IN0(5), B => IN1(5), S => CTRL, Z => OUT1(5));
   U38 : MUX2_X1 port map( A => IN0(7), B => IN1(7), S => CTRL, Z => OUT1(7));
   U39 : MUX2_X1 port map( A => IN0(3), B => IN1(3), S => CTRL, Z => OUT1(3));

end SYN_Bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity mux21_2 is

   port( IN0, IN1 : in std_logic_vector (31 downto 0);  CTRL : in std_logic;  
         OUT1 : out std_logic_vector (31 downto 0));

end mux21_2;

architecture SYN_Bhe of mux21_2 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : MUX2_X1 port map( A => IN0(9), B => IN1(9), S => n1, Z => OUT1(9));
   U2 : MUX2_X1 port map( A => IN0(8), B => IN1(8), S => n1, Z => OUT1(8));
   U3 : MUX2_X1 port map( A => IN0(7), B => IN1(7), S => n1, Z => OUT1(7));
   U4 : MUX2_X1 port map( A => IN0(6), B => IN1(6), S => n1, Z => OUT1(6));
   U5 : MUX2_X1 port map( A => IN0(5), B => IN1(5), S => n1, Z => OUT1(5));
   U6 : MUX2_X1 port map( A => IN0(4), B => IN1(4), S => n1, Z => OUT1(4));
   U7 : MUX2_X1 port map( A => IN0(3), B => IN1(3), S => n1, Z => OUT1(3));
   U8 : MUX2_X1 port map( A => IN0(31), B => IN1(31), S => n1, Z => OUT1(31));
   U9 : MUX2_X1 port map( A => IN0(30), B => IN1(30), S => n1, Z => OUT1(30));
   U10 : MUX2_X1 port map( A => IN0(2), B => IN1(2), S => n1, Z => OUT1(2));
   U11 : MUX2_X1 port map( A => IN0(29), B => IN1(29), S => n1, Z => OUT1(29));
   U12 : MUX2_X1 port map( A => IN0(28), B => IN1(28), S => n1, Z => OUT1(28));
   U13 : MUX2_X1 port map( A => IN0(27), B => IN1(27), S => n2, Z => OUT1(27));
   U14 : MUX2_X1 port map( A => IN0(26), B => IN1(26), S => n2, Z => OUT1(26));
   U15 : MUX2_X1 port map( A => IN0(25), B => IN1(25), S => n2, Z => OUT1(25));
   U16 : MUX2_X1 port map( A => IN0(24), B => IN1(24), S => n2, Z => OUT1(24));
   U17 : MUX2_X1 port map( A => IN0(23), B => IN1(23), S => n2, Z => OUT1(23));
   U18 : MUX2_X1 port map( A => IN0(22), B => IN1(22), S => n2, Z => OUT1(22));
   U19 : MUX2_X1 port map( A => IN0(21), B => IN1(21), S => n2, Z => OUT1(21));
   U20 : MUX2_X1 port map( A => IN0(20), B => IN1(20), S => n2, Z => OUT1(20));
   U21 : MUX2_X1 port map( A => IN0(1), B => IN1(1), S => n2, Z => OUT1(1));
   U22 : MUX2_X1 port map( A => IN0(19), B => IN1(19), S => n2, Z => OUT1(19));
   U23 : MUX2_X1 port map( A => IN0(18), B => IN1(18), S => n2, Z => OUT1(18));
   U24 : MUX2_X1 port map( A => IN0(17), B => IN1(17), S => n2, Z => OUT1(17));
   U25 : MUX2_X1 port map( A => IN0(16), B => IN1(16), S => CTRL, Z => OUT1(16)
                           );
   U26 : MUX2_X1 port map( A => IN0(15), B => IN1(15), S => CTRL, Z => OUT1(15)
                           );
   U27 : MUX2_X1 port map( A => IN0(14), B => IN1(14), S => CTRL, Z => OUT1(14)
                           );
   U28 : MUX2_X1 port map( A => IN0(13), B => IN1(13), S => CTRL, Z => OUT1(13)
                           );
   U29 : MUX2_X1 port map( A => IN0(12), B => IN1(12), S => CTRL, Z => OUT1(12)
                           );
   U30 : MUX2_X1 port map( A => IN0(11), B => IN1(11), S => CTRL, Z => OUT1(11)
                           );
   U31 : MUX2_X1 port map( A => IN0(10), B => IN1(10), S => CTRL, Z => OUT1(10)
                           );
   U32 : MUX2_X1 port map( A => IN0(0), B => IN1(0), S => CTRL, Z => OUT1(0));
   U33 : BUF_X1 port map( A => CTRL, Z => n1);
   U34 : BUF_X1 port map( A => CTRL, Z => n2);

end SYN_Bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity mux21_1 is

   port( IN0, IN1 : in std_logic_vector (31 downto 0);  CTRL : in std_logic;  
         OUT1 : out std_logic_vector (31 downto 0));

end mux21_1;

architecture SYN_Bhe of mux21_1 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : MUX2_X1 port map( A => IN0(9), B => IN1(9), S => CTRL, Z => OUT1(9));
   U2 : MUX2_X1 port map( A => IN0(8), B => IN1(8), S => CTRL, Z => OUT1(8));
   U4 : MUX2_X1 port map( A => IN0(6), B => IN1(6), S => CTRL, Z => OUT1(6));
   U5 : MUX2_X1 port map( A => IN0(5), B => IN1(5), S => CTRL, Z => OUT1(5));
   U6 : MUX2_X1 port map( A => IN0(4), B => IN1(4), S => CTRL, Z => OUT1(4));
   U7 : MUX2_X1 port map( A => IN0(3), B => IN1(3), S => CTRL, Z => OUT1(3));
   U8 : MUX2_X1 port map( A => IN0(31), B => IN1(31), S => CTRL, Z => OUT1(31))
                           ;
   U9 : MUX2_X1 port map( A => IN0(30), B => IN1(30), S => CTRL, Z => OUT1(30))
                           ;
   U10 : MUX2_X1 port map( A => IN0(2), B => IN1(2), S => CTRL, Z => OUT1(2));
   U11 : MUX2_X1 port map( A => IN0(29), B => IN1(29), S => CTRL, Z => OUT1(29)
                           );
   U12 : MUX2_X1 port map( A => IN0(28), B => IN1(28), S => CTRL, Z => OUT1(28)
                           );
   U13 : MUX2_X1 port map( A => IN0(27), B => IN1(27), S => CTRL, Z => OUT1(27)
                           );
   U14 : MUX2_X1 port map( A => IN0(26), B => IN1(26), S => CTRL, Z => OUT1(26)
                           );
   U15 : MUX2_X1 port map( A => IN0(25), B => IN1(25), S => CTRL, Z => OUT1(25)
                           );
   U16 : MUX2_X1 port map( A => IN0(24), B => IN1(24), S => CTRL, Z => OUT1(24)
                           );
   U17 : MUX2_X1 port map( A => IN0(23), B => IN1(23), S => CTRL, Z => OUT1(23)
                           );
   U18 : MUX2_X1 port map( A => IN0(22), B => IN1(22), S => CTRL, Z => OUT1(22)
                           );
   U20 : MUX2_X1 port map( A => IN0(20), B => IN1(20), S => CTRL, Z => OUT1(20)
                           );
   U21 : MUX2_X1 port map( A => IN0(1), B => IN1(1), S => CTRL, Z => OUT1(1));
   U22 : MUX2_X1 port map( A => IN0(19), B => IN1(19), S => CTRL, Z => OUT1(19)
                           );
   U23 : MUX2_X1 port map( A => IN0(18), B => IN1(18), S => CTRL, Z => OUT1(18)
                           );
   U24 : MUX2_X1 port map( A => IN0(17), B => IN1(17), S => CTRL, Z => OUT1(17)
                           );
   U25 : MUX2_X1 port map( A => IN0(16), B => IN1(16), S => CTRL, Z => OUT1(16)
                           );
   U26 : MUX2_X1 port map( A => IN0(15), B => IN1(15), S => CTRL, Z => OUT1(15)
                           );
   U27 : MUX2_X1 port map( A => IN0(14), B => IN1(14), S => CTRL, Z => OUT1(14)
                           );
   U28 : MUX2_X1 port map( A => IN0(13), B => IN1(13), S => CTRL, Z => OUT1(13)
                           );
   U29 : MUX2_X1 port map( A => IN0(12), B => IN1(12), S => CTRL, Z => OUT1(12)
                           );
   U30 : MUX2_X1 port map( A => IN0(11), B => IN1(11), S => CTRL, Z => OUT1(11)
                           );
   U31 : MUX2_X1 port map( A => IN0(10), B => IN1(10), S => CTRL, Z => OUT1(10)
                           );
   U3 : INV_X1 port map( A => IN0(0), ZN => n1);
   U19 : NOR2_X1 port map( A1 => CTRL, A2 => n1, ZN => OUT1(0));
   U32 : MUX2_X1 port map( A => IN0(7), B => IN1(7), S => CTRL, Z => OUT1(7));
   U33 : MUX2_X1 port map( A => IN0(21), B => IN1(21), S => CTRL, Z => OUT1(21)
                           );

end SYN_Bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity p4add_N32_logN5_1 is

   port( A, B : in std_logic_vector (31 downto 0);  Cin, sign : in std_logic;  
         S : out std_logic_vector (31 downto 0);  Cout : out std_logic);

end p4add_N32_logN5_1;

architecture SYN_STRUCTURAL of p4add_N32_logN5_1 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component sum_gen_N32_1
      port( A, B : in std_logic_vector (31 downto 0);  Cin : in 
            std_logic_vector (8 downto 0);  S : out std_logic_vector (31 downto
            0));
   end component;
   
   component carry_tree_N32_logN5_1
      port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  
            Cout : out std_logic_vector (7 downto 0));
   end component;
   
   component xor_gen_N32_1
      port( A : in std_logic_vector (31 downto 0);  B : in std_logic;  S : out 
            std_logic_vector (31 downto 0));
   end component;
   
   signal new_B_31_port, new_B_30_port, new_B_29_port, new_B_28_port, 
      new_B_27_port, new_B_26_port, new_B_25_port, new_B_24_port, new_B_23_port
      , new_B_22_port, new_B_21_port, new_B_20_port, new_B_19_port, 
      new_B_18_port, new_B_17_port, new_B_16_port, new_B_15_port, new_B_14_port
      , new_B_13_port, new_B_12_port, new_B_11_port, new_B_10_port, 
      new_B_9_port, new_B_8_port, new_B_7_port, new_B_6_port, new_B_5_port, 
      new_B_4_port, new_B_3_port, new_B_2_port, new_B_1_port, new_B_0_port, 
      carry_pro_7_port, carry_pro_6_port, carry_pro_5_port, carry_pro_4_port, 
      carry_pro_3_port, carry_pro_2_port, carry_pro_1_port, n1, n2, n3, n4, n5 
      : std_logic;

begin
   
   xor32 : xor_gen_N32_1 port map( A(31) => B(31), A(30) => B(30), A(29) => 
                           B(29), A(28) => B(28), A(27) => B(27), A(26) => 
                           B(26), A(25) => B(25), A(24) => B(24), A(23) => 
                           B(23), A(22) => B(22), A(21) => B(21), A(20) => 
                           B(20), A(19) => B(19), A(18) => B(18), A(17) => 
                           B(17), A(16) => B(16), A(15) => B(15), A(14) => 
                           B(14), A(13) => B(13), A(12) => B(12), A(11) => 
                           B(11), A(10) => B(10), A(9) => B(9), A(8) => B(8), 
                           A(7) => B(7), A(6) => B(6), A(5) => B(5), A(4) => 
                           B(4), A(3) => B(3), A(2) => B(2), A(1) => B(1), A(0)
                           => B(0), B => sign, S(31) => new_B_31_port, S(30) =>
                           new_B_30_port, S(29) => new_B_29_port, S(28) => 
                           new_B_28_port, S(27) => new_B_27_port, S(26) => 
                           new_B_26_port, S(25) => new_B_25_port, S(24) => 
                           new_B_24_port, S(23) => new_B_23_port, S(22) => 
                           new_B_22_port, S(21) => new_B_21_port, S(20) => 
                           new_B_20_port, S(19) => new_B_19_port, S(18) => 
                           new_B_18_port, S(17) => new_B_17_port, S(16) => 
                           new_B_16_port, S(15) => new_B_15_port, S(14) => 
                           new_B_14_port, S(13) => new_B_13_port, S(12) => 
                           new_B_12_port, S(11) => new_B_11_port, S(10) => 
                           new_B_10_port, S(9) => new_B_9_port, S(8) => 
                           new_B_8_port, S(7) => new_B_7_port, S(6) => 
                           new_B_6_port, S(5) => new_B_5_port, S(4) => 
                           new_B_4_port, S(3) => new_B_3_port, S(2) => 
                           new_B_2_port, S(1) => new_B_1_port, S(0) => 
                           new_B_0_port);
   ct : carry_tree_N32_logN5_1 port map( A(31) => A(31), A(30) => A(30), A(29) 
                           => A(29), A(28) => A(28), A(27) => A(27), A(26) => 
                           A(26), A(25) => A(25), A(24) => A(24), A(23) => 
                           A(23), A(22) => A(22), A(21) => A(21), A(20) => 
                           A(20), A(19) => A(19), A(18) => A(18), A(17) => 
                           A(17), A(16) => A(16), A(15) => A(15), A(14) => 
                           A(14), A(13) => A(13), A(12) => A(12), A(11) => 
                           A(11), A(10) => A(10), A(9) => A(9), A(8) => A(8), 
                           A(7) => A(7), A(6) => A(6), A(5) => A(5), A(4) => 
                           A(4), A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(31) => new_B_31_port, B(30) => 
                           new_B_30_port, B(29) => new_B_29_port, B(28) => 
                           new_B_28_port, B(27) => new_B_27_port, B(26) => 
                           new_B_26_port, B(25) => new_B_25_port, B(24) => 
                           new_B_24_port, B(23) => new_B_23_port, B(22) => 
                           new_B_22_port, B(21) => new_B_21_port, B(20) => 
                           new_B_20_port, B(19) => new_B_19_port, B(18) => 
                           new_B_18_port, B(17) => new_B_17_port, B(16) => 
                           new_B_16_port, B(15) => new_B_15_port, B(14) => 
                           new_B_14_port, B(13) => new_B_13_port, B(12) => 
                           new_B_12_port, B(11) => new_B_11_port, B(10) => 
                           new_B_10_port, B(9) => new_B_9_port, B(8) => 
                           new_B_8_port, B(7) => new_B_7_port, B(6) => 
                           new_B_6_port, B(5) => new_B_5_port, B(4) => 
                           new_B_4_port, B(3) => new_B_3_port, B(2) => 
                           new_B_2_port, B(1) => new_B_1_port, B(0) => 
                           new_B_0_port, Cin => sign, Cout(7) => Cout, Cout(6) 
                           => carry_pro_7_port, Cout(5) => carry_pro_6_port, 
                           Cout(4) => carry_pro_5_port, Cout(3) => 
                           carry_pro_4_port, Cout(2) => carry_pro_3_port, 
                           Cout(1) => carry_pro_2_port, Cout(0) => 
                           carry_pro_1_port);
   add : sum_gen_N32_1 port map( A(31) => A(31), A(30) => A(30), A(29) => A(29)
                           , A(28) => A(28), A(27) => A(27), A(26) => A(26), 
                           A(25) => A(25), A(24) => A(24), A(23) => A(23), 
                           A(22) => A(22), A(21) => A(21), A(20) => A(20), 
                           A(19) => A(19), A(18) => A(18), A(17) => A(17), 
                           A(16) => A(16), A(15) => A(15), A(14) => A(14), 
                           A(13) => A(13), A(12) => A(12), A(11) => A(11), 
                           A(10) => A(10), A(9) => A(9), A(8) => A(8), A(7) => 
                           A(7), A(6) => A(6), A(5) => A(5), A(4) => A(4), A(3)
                           => A(3), A(2) => A(2), A(1) => A(1), A(0) => A(0), 
                           B(31) => new_B_31_port, B(30) => new_B_30_port, 
                           B(29) => new_B_29_port, B(28) => new_B_28_port, 
                           B(27) => new_B_27_port, B(26) => new_B_26_port, 
                           B(25) => new_B_25_port, B(24) => new_B_24_port, 
                           B(23) => new_B_23_port, B(22) => new_B_22_port, 
                           B(21) => new_B_21_port, B(20) => new_B_20_port, 
                           B(19) => new_B_19_port, B(18) => new_B_18_port, 
                           B(17) => new_B_17_port, B(16) => new_B_16_port, 
                           B(15) => new_B_15_port, B(14) => new_B_14_port, 
                           B(13) => n1, B(12) => new_B_12_port, B(11) => 
                           new_B_11_port, B(10) => new_B_10_port, B(9) => 
                           new_B_9_port, B(8) => new_B_8_port, B(7) => 
                           new_B_7_port, B(6) => n4, B(5) => new_B_5_port, B(4)
                           => new_B_4_port, B(3) => new_B_3_port, B(2) => n2, 
                           B(1) => n3, B(0) => new_B_0_port, Cin(8) => n5, 
                           Cin(7) => carry_pro_7_port, Cin(6) => 
                           carry_pro_6_port, Cin(5) => carry_pro_5_port, Cin(4)
                           => carry_pro_4_port, Cin(3) => carry_pro_3_port, 
                           Cin(2) => carry_pro_2_port, Cin(1) => 
                           carry_pro_1_port, Cin(0) => sign, S(31) => S(31), 
                           S(30) => S(30), S(29) => S(29), S(28) => S(28), 
                           S(27) => S(27), S(26) => S(26), S(25) => S(25), 
                           S(24) => S(24), S(23) => S(23), S(22) => S(22), 
                           S(21) => S(21), S(20) => S(20), S(19) => S(19), 
                           S(18) => S(18), S(17) => S(17), S(16) => S(16), 
                           S(15) => S(15), S(14) => S(14), S(13) => S(13), 
                           S(12) => S(12), S(11) => S(11), S(10) => S(10), S(9)
                           => S(9), S(8) => S(8), S(7) => S(7), S(6) => S(6), 
                           S(5) => S(5), S(4) => S(4), S(3) => S(3), S(2) => 
                           S(2), S(1) => S(1), S(0) => S(0));
   U1 : BUF_X1 port map( A => new_B_1_port, Z => n3);
   U2 : BUF_X1 port map( A => new_B_6_port, Z => n4);
   U3 : BUF_X1 port map( A => new_B_2_port, Z => n2);
   U4 : BUF_X1 port map( A => new_B_13_port, Z => n1);
   n5 <= '0';

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity predictor_2_15 is

   port( clock, reset, enable, taken_i : in std_logic;  prediction_o : out 
         std_logic);

end predictor_2_15;

architecture SYN_bhe of predictor_2_15 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal prediction_o_port, next_STATE_1_port, next_STATE_0_port, N11, N12, n1
      , n2, n5, n7, n8, n9, n10, net246142 : std_logic;

begin
   prediction_o <= prediction_o_port;
   
   next_STATE_reg_0_inst : DLH_X1 port map( G => enable, D => N11, Q => 
                           next_STATE_0_port);
   STATE_reg_0_inst : DFFR_X1 port map( D => n7, CK => clock, RN => n2, Q => n1
                           , QN => n5);
   next_STATE_reg_1_inst : DLH_X1 port map( G => enable, D => N12, Q => 
                           next_STATE_1_port);
   STATE_reg_1_inst : DFFR_X1 port map( D => n8, CK => clock, RN => n2, Q => 
                           prediction_o_port, QN => net246142);
   U2 : MUX2_X1 port map( A => prediction_o_port, B => next_STATE_1_port, S => 
                           enable, Z => n8);
   U4 : MUX2_X1 port map( A => n1, B => next_STATE_0_port, S => enable, Z => n7
                           );
   U9 : NOR2_X1 port map( A1 => prediction_o_port, A2 => taken_i, ZN => n10);
   U7 : NAND2_X1 port map( A1 => prediction_o_port, A2 => taken_i, ZN => n9);
   U6 : OAI21_X1 port map( B1 => n10, B2 => n1, A => n9, ZN => N11);
   U5 : OAI21_X1 port map( B1 => n5, B2 => n10, A => n9, ZN => N12);
   U3 : INV_X1 port map( A => reset, ZN => n2);

end SYN_bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity predictor_2_14 is

   port( clock, reset, enable, taken_i : in std_logic;  prediction_o : out 
         std_logic);

end predictor_2_14;

architecture SYN_bhe of predictor_2_14 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal prediction_o_port, next_STATE_1_port, next_STATE_0_port, N11, N12, n1
      , n2, n5, n7, n8, n9, n10, net246141 : std_logic;

begin
   prediction_o <= prediction_o_port;
   
   next_STATE_reg_0_inst : DLH_X1 port map( G => enable, D => N11, Q => 
                           next_STATE_0_port);
   STATE_reg_0_inst : DFFR_X1 port map( D => n7, CK => clock, RN => n2, Q => n1
                           , QN => n5);
   next_STATE_reg_1_inst : DLH_X1 port map( G => enable, D => N12, Q => 
                           next_STATE_1_port);
   STATE_reg_1_inst : DFFR_X1 port map( D => n8, CK => clock, RN => n2, Q => 
                           prediction_o_port, QN => net246141);
   U2 : MUX2_X1 port map( A => prediction_o_port, B => next_STATE_1_port, S => 
                           enable, Z => n8);
   U4 : MUX2_X1 port map( A => n1, B => next_STATE_0_port, S => enable, Z => n7
                           );
   U9 : NOR2_X1 port map( A1 => prediction_o_port, A2 => taken_i, ZN => n10);
   U7 : NAND2_X1 port map( A1 => prediction_o_port, A2 => taken_i, ZN => n9);
   U6 : OAI21_X1 port map( B1 => n10, B2 => n1, A => n9, ZN => N11);
   U5 : OAI21_X1 port map( B1 => n5, B2 => n10, A => n9, ZN => N12);
   U3 : INV_X1 port map( A => reset, ZN => n2);

end SYN_bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity predictor_2_13 is

   port( clock, reset, enable, taken_i : in std_logic;  prediction_o : out 
         std_logic);

end predictor_2_13;

architecture SYN_bhe of predictor_2_13 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal prediction_o_port, next_STATE_1_port, next_STATE_0_port, N11, N12, n1
      , n2, n5, n7, n8, n9, n10, net246140 : std_logic;

begin
   prediction_o <= prediction_o_port;
   
   next_STATE_reg_0_inst : DLH_X1 port map( G => enable, D => N11, Q => 
                           next_STATE_0_port);
   STATE_reg_0_inst : DFFR_X1 port map( D => n7, CK => clock, RN => n2, Q => n1
                           , QN => n5);
   next_STATE_reg_1_inst : DLH_X1 port map( G => enable, D => N12, Q => 
                           next_STATE_1_port);
   STATE_reg_1_inst : DFFR_X1 port map( D => n8, CK => clock, RN => n2, Q => 
                           prediction_o_port, QN => net246140);
   U2 : MUX2_X1 port map( A => prediction_o_port, B => next_STATE_1_port, S => 
                           enable, Z => n8);
   U4 : MUX2_X1 port map( A => n1, B => next_STATE_0_port, S => enable, Z => n7
                           );
   U9 : NOR2_X1 port map( A1 => prediction_o_port, A2 => taken_i, ZN => n10);
   U7 : NAND2_X1 port map( A1 => prediction_o_port, A2 => taken_i, ZN => n9);
   U5 : OAI21_X1 port map( B1 => n5, B2 => n10, A => n9, ZN => N12);
   U6 : OAI21_X1 port map( B1 => n10, B2 => n1, A => n9, ZN => N11);
   U3 : INV_X1 port map( A => reset, ZN => n2);

end SYN_bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity predictor_2_12 is

   port( clock, reset, enable, taken_i : in std_logic;  prediction_o : out 
         std_logic);

end predictor_2_12;

architecture SYN_bhe of predictor_2_12 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal prediction_o_port, next_STATE_1_port, next_STATE_0_port, N11, N12, n1
      , n2, n5, n7, n8, n9, n10, net246139 : std_logic;

begin
   prediction_o <= prediction_o_port;
   
   next_STATE_reg_0_inst : DLH_X1 port map( G => enable, D => N11, Q => 
                           next_STATE_0_port);
   STATE_reg_0_inst : DFFR_X1 port map( D => n7, CK => clock, RN => n2, Q => n1
                           , QN => n5);
   next_STATE_reg_1_inst : DLH_X1 port map( G => enable, D => N12, Q => 
                           next_STATE_1_port);
   STATE_reg_1_inst : DFFR_X1 port map( D => n8, CK => clock, RN => n2, Q => 
                           prediction_o_port, QN => net246139);
   U2 : MUX2_X1 port map( A => prediction_o_port, B => next_STATE_1_port, S => 
                           enable, Z => n8);
   U4 : MUX2_X1 port map( A => n1, B => next_STATE_0_port, S => enable, Z => n7
                           );
   U9 : NOR2_X1 port map( A1 => prediction_o_port, A2 => taken_i, ZN => n10);
   U7 : NAND2_X1 port map( A1 => prediction_o_port, A2 => taken_i, ZN => n9);
   U5 : OAI21_X1 port map( B1 => n5, B2 => n10, A => n9, ZN => N12);
   U6 : OAI21_X1 port map( B1 => n10, B2 => n1, A => n9, ZN => N11);
   U3 : INV_X1 port map( A => reset, ZN => n2);

end SYN_bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity predictor_2_11 is

   port( clock, reset, enable, taken_i : in std_logic;  prediction_o : out 
         std_logic);

end predictor_2_11;

architecture SYN_bhe of predictor_2_11 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal prediction_o_port, next_STATE_1_port, next_STATE_0_port, N11, N12, n1
      , n2, n5, n7, n8, n9, n10, net246138 : std_logic;

begin
   prediction_o <= prediction_o_port;
   
   next_STATE_reg_0_inst : DLH_X1 port map( G => enable, D => N11, Q => 
                           next_STATE_0_port);
   STATE_reg_0_inst : DFFR_X1 port map( D => n7, CK => clock, RN => n2, Q => n1
                           , QN => n5);
   next_STATE_reg_1_inst : DLH_X1 port map( G => enable, D => N12, Q => 
                           next_STATE_1_port);
   STATE_reg_1_inst : DFFR_X1 port map( D => n8, CK => clock, RN => n2, Q => 
                           prediction_o_port, QN => net246138);
   U2 : MUX2_X1 port map( A => prediction_o_port, B => next_STATE_1_port, S => 
                           enable, Z => n8);
   U4 : MUX2_X1 port map( A => n1, B => next_STATE_0_port, S => enable, Z => n7
                           );
   U9 : NOR2_X1 port map( A1 => prediction_o_port, A2 => taken_i, ZN => n10);
   U7 : NAND2_X1 port map( A1 => prediction_o_port, A2 => taken_i, ZN => n9);
   U5 : OAI21_X1 port map( B1 => n5, B2 => n10, A => n9, ZN => N12);
   U6 : OAI21_X1 port map( B1 => n10, B2 => n1, A => n9, ZN => N11);
   U3 : INV_X1 port map( A => reset, ZN => n2);

end SYN_bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity predictor_2_10 is

   port( clock, reset, enable, taken_i : in std_logic;  prediction_o : out 
         std_logic);

end predictor_2_10;

architecture SYN_bhe of predictor_2_10 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal prediction_o_port, next_STATE_1_port, next_STATE_0_port, N11, N12, n1
      , n2, n5, n7, n8, n9, n10, net246137 : std_logic;

begin
   prediction_o <= prediction_o_port;
   
   next_STATE_reg_0_inst : DLH_X1 port map( G => enable, D => N11, Q => 
                           next_STATE_0_port);
   STATE_reg_0_inst : DFFR_X1 port map( D => n7, CK => clock, RN => n2, Q => n1
                           , QN => n5);
   next_STATE_reg_1_inst : DLH_X1 port map( G => enable, D => N12, Q => 
                           next_STATE_1_port);
   STATE_reg_1_inst : DFFR_X1 port map( D => n8, CK => clock, RN => n2, Q => 
                           prediction_o_port, QN => net246137);
   U2 : MUX2_X1 port map( A => prediction_o_port, B => next_STATE_1_port, S => 
                           enable, Z => n8);
   U4 : MUX2_X1 port map( A => n1, B => next_STATE_0_port, S => enable, Z => n7
                           );
   U9 : NOR2_X1 port map( A1 => prediction_o_port, A2 => taken_i, ZN => n10);
   U7 : NAND2_X1 port map( A1 => prediction_o_port, A2 => taken_i, ZN => n9);
   U6 : OAI21_X1 port map( B1 => n10, B2 => n1, A => n9, ZN => N11);
   U5 : OAI21_X1 port map( B1 => n5, B2 => n10, A => n9, ZN => N12);
   U3 : INV_X1 port map( A => reset, ZN => n2);

end SYN_bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity predictor_2_9 is

   port( clock, reset, enable, taken_i : in std_logic;  prediction_o : out 
         std_logic);

end predictor_2_9;

architecture SYN_bhe of predictor_2_9 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal prediction_o_port, next_STATE_1_port, next_STATE_0_port, N11, N12, n1
      , n2, n5, n7, n8, n9, n10, net246136 : std_logic;

begin
   prediction_o <= prediction_o_port;
   
   next_STATE_reg_0_inst : DLH_X1 port map( G => enable, D => N11, Q => 
                           next_STATE_0_port);
   STATE_reg_0_inst : DFFR_X1 port map( D => n7, CK => clock, RN => n2, Q => n1
                           , QN => n5);
   next_STATE_reg_1_inst : DLH_X1 port map( G => enable, D => N12, Q => 
                           next_STATE_1_port);
   STATE_reg_1_inst : DFFR_X1 port map( D => n8, CK => clock, RN => n2, Q => 
                           prediction_o_port, QN => net246136);
   U2 : MUX2_X1 port map( A => prediction_o_port, B => next_STATE_1_port, S => 
                           enable, Z => n8);
   U4 : MUX2_X1 port map( A => n1, B => next_STATE_0_port, S => enable, Z => n7
                           );
   U9 : NOR2_X1 port map( A1 => prediction_o_port, A2 => taken_i, ZN => n10);
   U7 : NAND2_X1 port map( A1 => prediction_o_port, A2 => taken_i, ZN => n9);
   U6 : OAI21_X1 port map( B1 => n10, B2 => n1, A => n9, ZN => N11);
   U5 : OAI21_X1 port map( B1 => n5, B2 => n10, A => n9, ZN => N12);
   U3 : INV_X1 port map( A => reset, ZN => n2);

end SYN_bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity predictor_2_8 is

   port( clock, reset, enable, taken_i : in std_logic;  prediction_o : out 
         std_logic);

end predictor_2_8;

architecture SYN_bhe of predictor_2_8 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal prediction_o_port, next_STATE_1_port, next_STATE_0_port, N11, N12, n1
      , n2, n5, n7, n8, n9, n10, net246135 : std_logic;

begin
   prediction_o <= prediction_o_port;
   
   next_STATE_reg_0_inst : DLH_X1 port map( G => enable, D => N11, Q => 
                           next_STATE_0_port);
   STATE_reg_0_inst : DFFR_X1 port map( D => n7, CK => clock, RN => n2, Q => n1
                           , QN => n5);
   next_STATE_reg_1_inst : DLH_X1 port map( G => enable, D => N12, Q => 
                           next_STATE_1_port);
   STATE_reg_1_inst : DFFR_X1 port map( D => n8, CK => clock, RN => n2, Q => 
                           prediction_o_port, QN => net246135);
   U2 : MUX2_X1 port map( A => prediction_o_port, B => next_STATE_1_port, S => 
                           enable, Z => n8);
   U4 : MUX2_X1 port map( A => n1, B => next_STATE_0_port, S => enable, Z => n7
                           );
   U9 : NOR2_X1 port map( A1 => prediction_o_port, A2 => taken_i, ZN => n10);
   U7 : NAND2_X1 port map( A1 => prediction_o_port, A2 => taken_i, ZN => n9);
   U5 : OAI21_X1 port map( B1 => n5, B2 => n10, A => n9, ZN => N12);
   U6 : OAI21_X1 port map( B1 => n10, B2 => n1, A => n9, ZN => N11);
   U3 : INV_X1 port map( A => reset, ZN => n2);

end SYN_bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity predictor_2_7 is

   port( clock, reset, enable, taken_i : in std_logic;  prediction_o : out 
         std_logic);

end predictor_2_7;

architecture SYN_bhe of predictor_2_7 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal prediction_o_port, next_STATE_1_port, next_STATE_0_port, N11, N12, n1
      , n2, n5, n7, n8, n9, n10, net246134 : std_logic;

begin
   prediction_o <= prediction_o_port;
   
   next_STATE_reg_0_inst : DLH_X1 port map( G => enable, D => N11, Q => 
                           next_STATE_0_port);
   STATE_reg_0_inst : DFFR_X1 port map( D => n7, CK => clock, RN => n2, Q => n1
                           , QN => n5);
   next_STATE_reg_1_inst : DLH_X1 port map( G => enable, D => N12, Q => 
                           next_STATE_1_port);
   STATE_reg_1_inst : DFFR_X1 port map( D => n8, CK => clock, RN => n2, Q => 
                           prediction_o_port, QN => net246134);
   U2 : MUX2_X1 port map( A => prediction_o_port, B => next_STATE_1_port, S => 
                           enable, Z => n8);
   U4 : MUX2_X1 port map( A => n1, B => next_STATE_0_port, S => enable, Z => n7
                           );
   U9 : NOR2_X1 port map( A1 => prediction_o_port, A2 => taken_i, ZN => n10);
   U7 : NAND2_X1 port map( A1 => prediction_o_port, A2 => taken_i, ZN => n9);
   U6 : OAI21_X1 port map( B1 => n10, B2 => n1, A => n9, ZN => N11);
   U5 : OAI21_X1 port map( B1 => n5, B2 => n10, A => n9, ZN => N12);
   U3 : INV_X1 port map( A => reset, ZN => n2);

end SYN_bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity predictor_2_6 is

   port( clock, reset, enable, taken_i : in std_logic;  prediction_o : out 
         std_logic);

end predictor_2_6;

architecture SYN_bhe of predictor_2_6 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal prediction_o_port, next_STATE_1_port, next_STATE_0_port, N11, N12, n1
      , n2, n5, n7, n8, n9, n10, net246133 : std_logic;

begin
   prediction_o <= prediction_o_port;
   
   next_STATE_reg_0_inst : DLH_X1 port map( G => enable, D => N11, Q => 
                           next_STATE_0_port);
   STATE_reg_0_inst : DFFR_X1 port map( D => n7, CK => clock, RN => n2, Q => n1
                           , QN => n5);
   next_STATE_reg_1_inst : DLH_X1 port map( G => enable, D => N12, Q => 
                           next_STATE_1_port);
   STATE_reg_1_inst : DFFR_X1 port map( D => n8, CK => clock, RN => n2, Q => 
                           prediction_o_port, QN => net246133);
   U2 : MUX2_X1 port map( A => prediction_o_port, B => next_STATE_1_port, S => 
                           enable, Z => n8);
   U4 : MUX2_X1 port map( A => n1, B => next_STATE_0_port, S => enable, Z => n7
                           );
   U9 : NOR2_X1 port map( A1 => prediction_o_port, A2 => taken_i, ZN => n10);
   U7 : NAND2_X1 port map( A1 => prediction_o_port, A2 => taken_i, ZN => n9);
   U5 : OAI21_X1 port map( B1 => n5, B2 => n10, A => n9, ZN => N12);
   U6 : OAI21_X1 port map( B1 => n10, B2 => n1, A => n9, ZN => N11);
   U3 : INV_X1 port map( A => reset, ZN => n2);

end SYN_bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity predictor_2_5 is

   port( clock, reset, enable, taken_i : in std_logic;  prediction_o : out 
         std_logic);

end predictor_2_5;

architecture SYN_bhe of predictor_2_5 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal prediction_o_port, next_STATE_1_port, next_STATE_0_port, N11, N12, n1
      , n2, n5, n7, n8, n9, n10, net246132 : std_logic;

begin
   prediction_o <= prediction_o_port;
   
   next_STATE_reg_0_inst : DLH_X1 port map( G => enable, D => N11, Q => 
                           next_STATE_0_port);
   STATE_reg_0_inst : DFFR_X1 port map( D => n7, CK => clock, RN => n2, Q => n1
                           , QN => n5);
   next_STATE_reg_1_inst : DLH_X1 port map( G => enable, D => N12, Q => 
                           next_STATE_1_port);
   STATE_reg_1_inst : DFFR_X1 port map( D => n8, CK => clock, RN => n2, Q => 
                           prediction_o_port, QN => net246132);
   U2 : MUX2_X1 port map( A => prediction_o_port, B => next_STATE_1_port, S => 
                           enable, Z => n8);
   U4 : MUX2_X1 port map( A => n1, B => next_STATE_0_port, S => enable, Z => n7
                           );
   U9 : NOR2_X1 port map( A1 => prediction_o_port, A2 => taken_i, ZN => n10);
   U7 : NAND2_X1 port map( A1 => prediction_o_port, A2 => taken_i, ZN => n9);
   U5 : OAI21_X1 port map( B1 => n5, B2 => n10, A => n9, ZN => N12);
   U6 : OAI21_X1 port map( B1 => n10, B2 => n1, A => n9, ZN => N11);
   U3 : INV_X1 port map( A => reset, ZN => n2);

end SYN_bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity predictor_2_4 is

   port( clock, reset, enable, taken_i : in std_logic;  prediction_o : out 
         std_logic);

end predictor_2_4;

architecture SYN_bhe of predictor_2_4 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal prediction_o_port, next_STATE_1_port, next_STATE_0_port, N11, N12, n1
      , n2, n5, n7, n8, n9, n10, net246131 : std_logic;

begin
   prediction_o <= prediction_o_port;
   
   next_STATE_reg_0_inst : DLH_X1 port map( G => enable, D => N11, Q => 
                           next_STATE_0_port);
   STATE_reg_0_inst : DFFR_X1 port map( D => n7, CK => clock, RN => n2, Q => n1
                           , QN => n5);
   next_STATE_reg_1_inst : DLH_X1 port map( G => enable, D => N12, Q => 
                           next_STATE_1_port);
   STATE_reg_1_inst : DFFR_X1 port map( D => n8, CK => clock, RN => n2, Q => 
                           prediction_o_port, QN => net246131);
   U2 : MUX2_X1 port map( A => prediction_o_port, B => next_STATE_1_port, S => 
                           enable, Z => n8);
   U4 : MUX2_X1 port map( A => n1, B => next_STATE_0_port, S => enable, Z => n7
                           );
   U9 : NOR2_X1 port map( A1 => prediction_o_port, A2 => taken_i, ZN => n10);
   U7 : NAND2_X1 port map( A1 => prediction_o_port, A2 => taken_i, ZN => n9);
   U5 : OAI21_X1 port map( B1 => n5, B2 => n10, A => n9, ZN => N12);
   U6 : OAI21_X1 port map( B1 => n10, B2 => n1, A => n9, ZN => N11);
   U3 : INV_X1 port map( A => reset, ZN => n2);

end SYN_bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity predictor_2_3 is

   port( clock, reset, enable, taken_i : in std_logic;  prediction_o : out 
         std_logic);

end predictor_2_3;

architecture SYN_bhe of predictor_2_3 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal prediction_o_port, next_STATE_1_port, next_STATE_0_port, N11, N12, n1
      , n2, n5, n7, n8, n9, n10, net246130 : std_logic;

begin
   prediction_o <= prediction_o_port;
   
   next_STATE_reg_0_inst : DLH_X1 port map( G => enable, D => N11, Q => 
                           next_STATE_0_port);
   STATE_reg_0_inst : DFFR_X1 port map( D => n7, CK => clock, RN => n2, Q => n1
                           , QN => n5);
   next_STATE_reg_1_inst : DLH_X1 port map( G => enable, D => N12, Q => 
                           next_STATE_1_port);
   STATE_reg_1_inst : DFFR_X1 port map( D => n8, CK => clock, RN => n2, Q => 
                           prediction_o_port, QN => net246130);
   U2 : MUX2_X1 port map( A => prediction_o_port, B => next_STATE_1_port, S => 
                           enable, Z => n8);
   U4 : MUX2_X1 port map( A => n1, B => next_STATE_0_port, S => enable, Z => n7
                           );
   U9 : NOR2_X1 port map( A1 => prediction_o_port, A2 => taken_i, ZN => n10);
   U7 : NAND2_X1 port map( A1 => prediction_o_port, A2 => taken_i, ZN => n9);
   U6 : OAI21_X1 port map( B1 => n10, B2 => n1, A => n9, ZN => N11);
   U5 : OAI21_X1 port map( B1 => n5, B2 => n10, A => n9, ZN => N12);
   U3 : INV_X1 port map( A => reset, ZN => n2);

end SYN_bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity predictor_2_2 is

   port( clock, reset, enable, taken_i : in std_logic;  prediction_o : out 
         std_logic);

end predictor_2_2;

architecture SYN_bhe of predictor_2_2 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal prediction_o_port, next_STATE_1_port, next_STATE_0_port, N11, N12, n1
      , n2, n5, n7, n8, n9, n10, net246129 : std_logic;

begin
   prediction_o <= prediction_o_port;
   
   next_STATE_reg_0_inst : DLH_X1 port map( G => enable, D => N11, Q => 
                           next_STATE_0_port);
   STATE_reg_0_inst : DFFR_X1 port map( D => n7, CK => clock, RN => n2, Q => n1
                           , QN => n5);
   next_STATE_reg_1_inst : DLH_X1 port map( G => enable, D => N12, Q => 
                           next_STATE_1_port);
   STATE_reg_1_inst : DFFR_X1 port map( D => n8, CK => clock, RN => n2, Q => 
                           prediction_o_port, QN => net246129);
   U2 : MUX2_X1 port map( A => prediction_o_port, B => next_STATE_1_port, S => 
                           enable, Z => n8);
   U4 : MUX2_X1 port map( A => n1, B => next_STATE_0_port, S => enable, Z => n7
                           );
   U9 : NOR2_X1 port map( A1 => prediction_o_port, A2 => taken_i, ZN => n10);
   U7 : NAND2_X1 port map( A1 => prediction_o_port, A2 => taken_i, ZN => n9);
   U6 : OAI21_X1 port map( B1 => n10, B2 => n1, A => n9, ZN => N11);
   U5 : OAI21_X1 port map( B1 => n5, B2 => n10, A => n9, ZN => N12);
   U3 : INV_X1 port map( A => reset, ZN => n2);

end SYN_bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity predictor_2_1 is

   port( clock, reset, enable, taken_i : in std_logic;  prediction_o : out 
         std_logic);

end predictor_2_1;

architecture SYN_bhe of predictor_2_1 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal prediction_o_port, next_STATE_1_port, next_STATE_0_port, N11, N12, n1
      , n2, n5, n7, n8, n9, n10, net246128 : std_logic;

begin
   prediction_o <= prediction_o_port;
   
   next_STATE_reg_0_inst : DLH_X1 port map( G => enable, D => N11, Q => 
                           next_STATE_0_port);
   STATE_reg_0_inst : DFFR_X1 port map( D => n7, CK => clock, RN => n2, Q => n1
                           , QN => n5);
   next_STATE_reg_1_inst : DLH_X1 port map( G => enable, D => N12, Q => 
                           next_STATE_1_port);
   STATE_reg_1_inst : DFFR_X1 port map( D => n8, CK => clock, RN => n2, Q => 
                           prediction_o_port, QN => net246128);
   U2 : MUX2_X1 port map( A => prediction_o_port, B => next_STATE_1_port, S => 
                           enable, Z => n8);
   U4 : MUX2_X1 port map( A => n1, B => next_STATE_0_port, S => enable, Z => n7
                           );
   U9 : NOR2_X1 port map( A1 => prediction_o_port, A2 => taken_i, ZN => n10);
   U7 : NAND2_X1 port map( A1 => prediction_o_port, A2 => taken_i, ZN => n9);
   U6 : OAI21_X1 port map( B1 => n10, B2 => n1, A => n9, ZN => N11);
   U5 : OAI21_X1 port map( B1 => n5, B2 => n10, A => n9, ZN => N12);
   U3 : INV_X1 port map( A => reset, ZN => n2);

end SYN_bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity mux41_1 is

   port( IN0, IN1, IN2, IN3 : in std_logic_vector (31 downto 0);  CTRL : in 
         std_logic_vector (1 downto 0);  OUT1 : out std_logic_vector (31 downto
         0));

end mux41_1;

architecture SYN_bhe of mux41_1 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6, n7, n21, n22, n23, n24, n31, n32, n33, n34, n35, n36,
      n37, n38, n39, n40, n41, n42, n57, n58, n59, n60, n61, n62, n63, n64, n65
      , n66, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, 
      n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96
      , n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123 : std_logic;

begin
   
   U1 : AOI22_X1 port map( A1 => IN0(24), A2 => n110, B1 => IN1(24), B2 => n113
                           , ZN => n1);
   U2 : NAND2_X1 port map( A1 => n91, A2 => n1, ZN => OUT1(24));
   U3 : AOI22_X1 port map( A1 => IN0(25), A2 => n109, B1 => IN1(25), B2 => n113
                           , ZN => n2);
   U4 : NAND2_X1 port map( A1 => n107, A2 => n2, ZN => OUT1(25));
   U5 : AOI22_X1 port map( A1 => IN0(27), A2 => n110, B1 => IN1(27), B2 => n113
                           , ZN => n5);
   U6 : NAND2_X1 port map( A1 => n108, A2 => n5, ZN => OUT1(27));
   U7 : AOI22_X1 port map( A1 => IN0(30), A2 => n110, B1 => IN1(30), B2 => n112
                           , ZN => n6);
   U8 : NAND2_X1 port map( A1 => n89, A2 => n6, ZN => OUT1(30));
   U9 : AOI22_X1 port map( A1 => IN0(31), A2 => n109, B1 => IN1(31), B2 => n112
                           , ZN => n7);
   U10 : NAND2_X1 port map( A1 => n90, A2 => n7, ZN => OUT1(31));
   U11 : BUF_X2 port map( A => n21, Z => n119);
   U12 : BUF_X2 port map( A => n123, Z => n117);
   U13 : BUF_X2 port map( A => n123, Z => n115);
   U14 : BUF_X2 port map( A => n121, Z => n113);
   U15 : BUF_X2 port map( A => n123, Z => n116);
   U16 : BUF_X2 port map( A => n122, Z => n109);
   U17 : BUF_X2 port map( A => n121, Z => n112);
   U18 : INV_X1 port map( A => CTRL(0), ZN => n120);
   U19 : BUF_X2 port map( A => n122, Z => n111);
   U20 : BUF_X2 port map( A => n21, Z => n22);
   U21 : AND2_X1 port map( A1 => CTRL(1), A2 => CTRL(0), ZN => n123);
   U22 : BUF_X2 port map( A => n21, Z => n118);
   U23 : BUF_X2 port map( A => n122, Z => n110);
   U24 : AND2_X1 port map( A1 => CTRL(1), A2 => n120, ZN => n21);
   U25 : BUF_X1 port map( A => n121, Z => n114);
   U26 : AOI22_X1 port map( A1 => n116, A2 => IN3(16), B1 => n22, B2 => IN2(16)
                           , ZN => n72);
   U27 : AOI22_X1 port map( A1 => n115, A2 => IN3(6), B1 => n22, B2 => IN2(6), 
                           ZN => n74);
   U28 : AOI22_X1 port map( A1 => n115, A2 => IN3(10), B1 => n22, B2 => IN2(10)
                           , ZN => n76);
   U29 : AOI22_X1 port map( A1 => n115, A2 => IN3(2), B1 => n22, B2 => IN2(2), 
                           ZN => n78);
   U30 : AOI22_X1 port map( A1 => n115, A2 => IN3(8), B1 => n22, B2 => IN2(8), 
                           ZN => n79);
   U31 : AOI22_X1 port map( A1 => n115, A2 => IN3(21), B1 => n22, B2 => IN2(21)
                           , ZN => n82);
   U32 : AOI22_X1 port map( A1 => n116, A2 => IN3(1), B1 => n22, B2 => IN2(1), 
                           ZN => n84);
   U33 : AOI22_X1 port map( A1 => n115, A2 => IN3(18), B1 => n22, B2 => IN2(18)
                           , ZN => n86);
   U34 : AOI22_X1 port map( A1 => n116, A2 => IN3(19), B1 => n22, B2 => IN2(19)
                           , ZN => n88);
   U35 : AOI22_X1 port map( A1 => n22, A2 => IN2(30), B1 => n117, B2 => IN3(30)
                           , ZN => n89);
   U36 : AOI22_X1 port map( A1 => n22, A2 => IN2(31), B1 => n117, B2 => IN3(31)
                           , ZN => n90);
   U37 : NAND2_X1 port map( A1 => n77, A2 => n78, ZN => OUT1(2));
   U38 : NAND2_X1 port map( A1 => n73, A2 => n74, ZN => OUT1(6));
   U39 : NAND2_X1 port map( A1 => n83, A2 => n84, ZN => OUT1(1));
   U40 : AOI22_X1 port map( A1 => n116, A2 => IN3(4), B1 => n118, B2 => IN2(4),
                           ZN => n24);
   U41 : AOI22_X1 port map( A1 => n112, A2 => IN1(4), B1 => n111, B2 => IN0(4),
                           ZN => n23);
   U42 : NAND2_X1 port map( A1 => n23, A2 => n24, ZN => OUT1(4));
   U43 : AOI22_X1 port map( A1 => n115, A2 => IN3(13), B1 => n118, B2 => 
                           IN2(13), ZN => n32);
   U44 : AOI22_X1 port map( A1 => n114, A2 => IN1(13), B1 => n109, B2 => 
                           IN0(13), ZN => n31);
   U45 : NAND2_X1 port map( A1 => n31, A2 => n32, ZN => OUT1(13));
   U46 : AOI22_X1 port map( A1 => n116, A2 => IN3(0), B1 => n118, B2 => IN2(0),
                           ZN => n34);
   U47 : AOI22_X1 port map( A1 => n114, A2 => IN1(0), B1 => n109, B2 => IN0(0),
                           ZN => n33);
   U48 : NAND2_X1 port map( A1 => n33, A2 => n34, ZN => OUT1(0));
   U49 : AOI22_X1 port map( A1 => n115, A2 => IN3(9), B1 => n118, B2 => IN2(9),
                           ZN => n36);
   U50 : AOI22_X1 port map( A1 => n112, A2 => IN1(9), B1 => n110, B2 => IN0(9),
                           ZN => n35);
   U51 : NAND2_X1 port map( A1 => n35, A2 => n36, ZN => OUT1(9));
   U52 : AOI22_X1 port map( A1 => n116, A2 => IN3(14), B1 => n118, B2 => 
                           IN2(14), ZN => n38);
   U53 : AOI22_X1 port map( A1 => n114, A2 => IN1(14), B1 => n110, B2 => 
                           IN0(14), ZN => n37);
   U54 : NAND2_X1 port map( A1 => n37, A2 => n38, ZN => OUT1(14));
   U55 : AOI22_X1 port map( A1 => n115, A2 => IN3(3), B1 => n118, B2 => IN2(3),
                           ZN => n40);
   U56 : AOI22_X1 port map( A1 => n112, A2 => IN1(3), B1 => n111, B2 => IN0(3),
                           ZN => n39);
   U57 : NAND2_X1 port map( A1 => n39, A2 => n40, ZN => OUT1(3));
   U58 : AOI22_X1 port map( A1 => n116, A2 => IN3(7), B1 => n118, B2 => IN2(7),
                           ZN => n42);
   U59 : AOI22_X1 port map( A1 => n112, A2 => IN1(7), B1 => n110, B2 => IN0(7),
                           ZN => n41);
   U60 : NAND2_X1 port map( A1 => n41, A2 => n42, ZN => OUT1(7));
   U61 : AOI22_X1 port map( A1 => n115, A2 => IN3(12), B1 => n118, B2 => 
                           IN2(12), ZN => n58);
   U62 : AOI22_X1 port map( A1 => n114, A2 => IN1(12), B1 => n111, B2 => 
                           IN0(12), ZN => n57);
   U63 : NAND2_X1 port map( A1 => n57, A2 => n58, ZN => OUT1(12));
   U64 : AOI22_X1 port map( A1 => n116, A2 => IN3(28), B1 => n118, B2 => 
                           IN2(28), ZN => n60);
   U65 : AOI22_X1 port map( A1 => n112, A2 => IN1(28), B1 => n109, B2 => 
                           IN0(28), ZN => n59);
   U66 : NAND2_X1 port map( A1 => n59, A2 => n60, ZN => OUT1(28));
   U67 : AOI22_X1 port map( A1 => n116, A2 => IN3(5), B1 => n118, B2 => IN2(5),
                           ZN => n62);
   U68 : AOI22_X1 port map( A1 => n112, A2 => IN1(5), B1 => n109, B2 => IN0(5),
                           ZN => n61);
   U69 : NAND2_X1 port map( A1 => n61, A2 => n62, ZN => OUT1(5));
   U70 : AOI22_X1 port map( A1 => n115, A2 => IN3(29), B1 => n118, B2 => 
                           IN2(29), ZN => n64);
   U71 : AOI22_X1 port map( A1 => n112, A2 => IN1(29), B1 => n109, B2 => 
                           IN0(29), ZN => n63);
   U72 : NAND2_X1 port map( A1 => n63, A2 => n64, ZN => OUT1(29));
   U73 : AOI22_X1 port map( A1 => n116, A2 => IN3(20), B1 => n118, B2 => 
                           IN2(20), ZN => n66);
   U74 : AOI22_X1 port map( A1 => n113, A2 => IN1(20), B1 => n109, B2 => 
                           IN0(20), ZN => n65);
   U75 : NAND2_X1 port map( A1 => n65, A2 => n66, ZN => OUT1(20));
   U76 : AOI22_X1 port map( A1 => n116, A2 => IN3(17), B1 => n118, B2 => 
                           IN2(17), ZN => n70);
   U77 : AOI22_X1 port map( A1 => n113, A2 => IN1(17), B1 => n109, B2 => 
                           IN0(17), ZN => n69);
   U78 : NAND2_X1 port map( A1 => n69, A2 => n70, ZN => OUT1(17));
   U79 : AOI22_X1 port map( A1 => n114, A2 => IN1(16), B1 => n111, B2 => 
                           IN0(16), ZN => n71);
   U80 : NAND2_X1 port map( A1 => n71, A2 => n72, ZN => OUT1(16));
   U81 : AOI22_X1 port map( A1 => n112, A2 => IN1(6), B1 => n109, B2 => IN0(6),
                           ZN => n73);
   U82 : AOI22_X1 port map( A1 => n114, A2 => IN1(10), B1 => n110, B2 => 
                           IN0(10), ZN => n75);
   U83 : NAND2_X1 port map( A1 => n75, A2 => n76, ZN => OUT1(10));
   U84 : AOI22_X1 port map( A1 => n112, A2 => IN1(2), B1 => n110, B2 => IN0(2),
                           ZN => n77);
   U85 : AOI22_X1 port map( A1 => n112, A2 => IN1(8), B1 => n111, B2 => IN0(8),
                           ZN => n80);
   U86 : NAND2_X1 port map( A1 => n80, A2 => n79, ZN => OUT1(8));
   U87 : AOI22_X1 port map( A1 => n113, A2 => IN1(21), B1 => n109, B2 => 
                           IN0(21), ZN => n81);
   U88 : NAND2_X1 port map( A1 => n81, A2 => n82, ZN => OUT1(21));
   U89 : AOI22_X1 port map( A1 => n113, A2 => IN1(1), B1 => n110, B2 => IN0(1),
                           ZN => n83);
   U90 : AOI22_X1 port map( A1 => n113, A2 => IN1(18), B1 => n111, B2 => 
                           IN0(18), ZN => n85);
   U91 : NAND2_X1 port map( A1 => n85, A2 => n86, ZN => OUT1(18));
   U92 : AOI22_X1 port map( A1 => n113, A2 => IN1(19), B1 => n111, B2 => 
                           IN0(19), ZN => n87);
   U93 : NAND2_X1 port map( A1 => n87, A2 => n88, ZN => OUT1(19));
   U94 : AOI22_X1 port map( A1 => n117, A2 => IN3(24), B1 => n119, B2 => 
                           IN2(24), ZN => n91);
   U95 : NAND3_X1 port map( A1 => n92, A2 => n93, A3 => n94, ZN => OUT1(26));
   U96 : AOI22_X1 port map( A1 => n117, A2 => IN3(26), B1 => n119, B2 => 
                           IN2(26), ZN => n94);
   U97 : NAND2_X1 port map( A1 => n113, A2 => IN1(26), ZN => n93);
   U98 : NAND2_X1 port map( A1 => n111, A2 => IN0(26), ZN => n92);
   U99 : NAND3_X1 port map( A1 => n96, A2 => n95, A3 => n97, ZN => OUT1(11));
   U100 : AOI22_X1 port map( A1 => n116, A2 => IN3(11), B1 => n119, B2 => 
                           IN2(11), ZN => n96);
   U101 : NAND2_X1 port map( A1 => n114, A2 => IN1(11), ZN => n97);
   U102 : NAND2_X1 port map( A1 => n111, A2 => IN0(11), ZN => n95);
   U103 : NAND3_X1 port map( A1 => n99, A2 => n100, A3 => n98, ZN => OUT1(15));
   U104 : AOI22_X1 port map( A1 => n117, A2 => IN3(15), B1 => n119, B2 => 
                           IN2(15), ZN => n99);
   U105 : NAND2_X1 port map( A1 => n110, A2 => IN0(15), ZN => n98);
   U106 : NAND2_X1 port map( A1 => n114, A2 => IN1(15), ZN => n100);
   U107 : NAND3_X1 port map( A1 => n103, A2 => n102, A3 => n101, ZN => OUT1(22)
                           );
   U108 : AOI22_X1 port map( A1 => n117, A2 => IN3(22), B1 => n119, B2 => 
                           IN2(22), ZN => n103);
   U109 : NAND2_X1 port map( A1 => n110, A2 => IN0(22), ZN => n102);
   U110 : NAND2_X1 port map( A1 => n113, A2 => IN1(22), ZN => n101);
   U111 : NAND3_X1 port map( A1 => n106, A2 => n105, A3 => n104, ZN => OUT1(23)
                           );
   U112 : NAND2_X1 port map( A1 => n111, A2 => IN0(23), ZN => n104);
   U113 : NAND2_X1 port map( A1 => n113, A2 => IN1(23), ZN => n105);
   U114 : AOI22_X1 port map( A1 => n117, A2 => IN3(23), B1 => n119, B2 => 
                           IN2(23), ZN => n106);
   U115 : AOI22_X1 port map( A1 => n117, A2 => IN3(25), B1 => n119, B2 => 
                           IN2(25), ZN => n107);
   U116 : AOI22_X1 port map( A1 => n117, A2 => IN3(27), B1 => n119, B2 => 
                           IN2(27), ZN => n108);
   U117 : NOR2_X1 port map( A1 => CTRL(1), A2 => CTRL(0), ZN => n122);
   U118 : NOR2_X1 port map( A1 => CTRL(1), A2 => n120, ZN => n121);

end SYN_bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity ff32_en_1 is

   port( D : in std_logic_vector (31 downto 0);  en, clk, rst : in std_logic;  
         Q : out std_logic_vector (31 downto 0));

end ff32_en_1;

architecture SYN_behavioral of ff32_en_1 is

   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_ff32_en_1
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal net199618, n32, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44
      , n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, 
      n59, n60, n61, n62, n63, n64, n65 : std_logic;

begin
   
   Q_reg_31_inst : DFFR_X1 port map( D => D(31), CK => net199618, RN => n32, Q 
                           => Q(31), QN => n34);
   Q_reg_30_inst : DFFR_X1 port map( D => D(30), CK => net199618, RN => n32, Q 
                           => Q(30), QN => n35);
   Q_reg_29_inst : DFFR_X1 port map( D => D(29), CK => net199618, RN => n32, Q 
                           => Q(29), QN => n36);
   Q_reg_28_inst : DFFR_X1 port map( D => D(28), CK => net199618, RN => n32, Q 
                           => Q(28), QN => n37);
   Q_reg_27_inst : DFFR_X1 port map( D => D(27), CK => net199618, RN => n32, Q 
                           => Q(27), QN => n38);
   Q_reg_26_inst : DFFR_X1 port map( D => D(26), CK => net199618, RN => n32, Q 
                           => Q(26), QN => n39);
   Q_reg_25_inst : DFFR_X1 port map( D => D(25), CK => net199618, RN => n32, Q 
                           => Q(25), QN => n40);
   Q_reg_24_inst : DFFR_X1 port map( D => D(24), CK => net199618, RN => n32, Q 
                           => Q(24), QN => n41);
   Q_reg_23_inst : DFFR_X1 port map( D => D(23), CK => net199618, RN => n32, Q 
                           => Q(23), QN => n42);
   Q_reg_22_inst : DFFR_X1 port map( D => D(22), CK => net199618, RN => n32, Q 
                           => Q(22), QN => n43);
   Q_reg_21_inst : DFFR_X1 port map( D => D(21), CK => net199618, RN => n32, Q 
                           => Q(21), QN => n44);
   Q_reg_20_inst : DFFR_X1 port map( D => D(20), CK => net199618, RN => n32, Q 
                           => Q(20), QN => n45);
   Q_reg_19_inst : DFFR_X1 port map( D => D(19), CK => net199618, RN => n32, Q 
                           => Q(19), QN => n46);
   Q_reg_18_inst : DFFR_X1 port map( D => D(18), CK => net199618, RN => n32, Q 
                           => Q(18), QN => n47);
   Q_reg_17_inst : DFFR_X1 port map( D => D(17), CK => net199618, RN => n32, Q 
                           => Q(17), QN => n48);
   Q_reg_16_inst : DFFR_X1 port map( D => D(16), CK => net199618, RN => n32, Q 
                           => Q(16), QN => n49);
   Q_reg_15_inst : DFFR_X1 port map( D => D(15), CK => net199618, RN => n32, Q 
                           => Q(15), QN => n50);
   Q_reg_14_inst : DFFR_X1 port map( D => D(14), CK => net199618, RN => n32, Q 
                           => Q(14), QN => n51);
   Q_reg_13_inst : DFFR_X1 port map( D => D(13), CK => net199618, RN => n32, Q 
                           => Q(13), QN => n52);
   Q_reg_12_inst : DFFR_X1 port map( D => D(12), CK => net199618, RN => n32, Q 
                           => Q(12), QN => n53);
   Q_reg_11_inst : DFFR_X1 port map( D => D(11), CK => net199618, RN => n32, Q 
                           => Q(11), QN => n54);
   Q_reg_10_inst : DFFR_X1 port map( D => D(10), CK => net199618, RN => n32, Q 
                           => Q(10), QN => n55);
   Q_reg_9_inst : DFFR_X1 port map( D => D(9), CK => net199618, RN => n32, Q =>
                           Q(9), QN => n56);
   Q_reg_8_inst : DFFR_X1 port map( D => D(8), CK => net199618, RN => n32, Q =>
                           Q(8), QN => n57);
   Q_reg_7_inst : DFFR_X1 port map( D => D(7), CK => net199618, RN => n32, Q =>
                           Q(7), QN => n58);
   Q_reg_6_inst : DFFR_X1 port map( D => D(6), CK => net199618, RN => n32, Q =>
                           Q(6), QN => n59);
   Q_reg_5_inst : DFFR_X1 port map( D => D(5), CK => net199618, RN => n32, Q =>
                           Q(5), QN => n60);
   Q_reg_4_inst : DFFR_X1 port map( D => D(4), CK => net199618, RN => n32, Q =>
                           Q(4), QN => n61);
   Q_reg_3_inst : DFFR_X1 port map( D => D(3), CK => net199618, RN => n32, Q =>
                           Q(3), QN => n62);
   Q_reg_2_inst : DFFR_X1 port map( D => D(2), CK => net199618, RN => n32, Q =>
                           Q(2), QN => n63);
   Q_reg_1_inst : DFFR_X1 port map( D => D(1), CK => net199618, RN => n32, Q =>
                           Q(1), QN => n64);
   Q_reg_0_inst : DFFR_X1 port map( D => D(0), CK => net199618, RN => n32, Q =>
                           Q(0), QN => n65);
   clk_gate_Q_reg : SNPS_CLOCK_GATE_HIGH_ff32_en_1 port map( CLK => clk, EN => 
                           en, ENCLK => net199618);
   U2 : INV_X2 port map( A => rst, ZN => n32);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity FA_0 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_0;

architecture SYN_BEHAVIORAL of FA_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => S);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity mux21_SIZE4_0 is

   port( IN0, IN1 : in std_logic_vector (3 downto 0);  CTRL : in std_logic;  
         OUT1 : out std_logic_vector (3 downto 0));

end mux21_SIZE4_0;

architecture SYN_Bhe of mux21_SIZE4_0 is

begin
   OUT1 <= ( IN0(3), IN0(2), IN0(1), IN0(0) );

end SYN_Bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity RCA_N4_0 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_0;

architecture SYN_STRUCTURAL of RCA_N4_0 is

   component FA_125
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_126
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_127
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_0
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal n1, CTMP_3_port, CTMP_2_port, CTMP_1_port, net246127 : std_logic;

begin
   
   FAI_1 : FA_0 port map( A => A(0), B => B(0), Ci => n1, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_127 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_126 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_125 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => net246127);
   n1 <= '0';

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity shift_thirdLevel is

   port( sel : in std_logic_vector (2 downto 0);  A : in std_logic_vector (38 
         downto 0);  Y : out std_logic_vector (31 downto 0));

end shift_thirdLevel;

architecture SYN_behav of shift_thirdLevel is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, 
      n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32
      , n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, 
      n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61
      , n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, 
      n76, n77, n78 : std_logic;

begin
   
   U7 : MUX2_X1 port map( A => n7, B => n6, S => n72, Z => Y(30));
   U10 : MUX2_X1 port map( A => n6, B => n9, S => n72, Z => Y(29));
   U13 : MUX2_X1 port map( A => n9, B => n11, S => sel(0), Z => Y(28));
   U16 : MUX2_X1 port map( A => n11, B => n13, S => n71, Z => Y(27));
   U19 : MUX2_X1 port map( A => n13, B => n15, S => n72, Z => Y(26));
   U22 : MUX2_X1 port map( A => n15, B => n17, S => sel(0), Z => Y(25));
   U25 : MUX2_X1 port map( A => n17, B => n19, S => sel(0), Z => Y(24));
   U28 : MUX2_X1 port map( A => n19, B => n21, S => n71, Z => Y(23));
   U31 : MUX2_X1 port map( A => n21, B => n23, S => n71, Z => Y(22));
   U34 : MUX2_X1 port map( A => n23, B => n25, S => n72, Z => Y(21));
   U37 : MUX2_X1 port map( A => n25, B => n27, S => sel(0), Z => Y(20));
   U40 : MUX2_X1 port map( A => n27, B => n29, S => n72, Z => Y(19));
   U43 : MUX2_X1 port map( A => n29, B => n31, S => n71, Z => Y(18));
   U46 : MUX2_X1 port map( A => n31, B => n33, S => n71, Z => Y(17));
   U49 : MUX2_X1 port map( A => n33, B => n35, S => n71, Z => Y(16));
   U55 : MUX2_X1 port map( A => n37, B => n39, S => n71, Z => Y(14));
   U58 : MUX2_X1 port map( A => n39, B => n41, S => n71, Z => Y(13));
   U61 : MUX2_X1 port map( A => n41, B => n43, S => n71, Z => Y(12));
   U64 : MUX2_X1 port map( A => n43, B => n45, S => n71, Z => Y(11));
   U67 : MUX2_X1 port map( A => n45, B => n47, S => n71, Z => Y(10));
   U70 : MUX2_X1 port map( A => n47, B => n49, S => n71, Z => Y(9));
   U73 : MUX2_X1 port map( A => n49, B => n51, S => n71, Z => Y(8));
   U76 : MUX2_X1 port map( A => n51, B => n53, S => n71, Z => Y(7));
   U79 : MUX2_X1 port map( A => n53, B => n55, S => n72, Z => Y(6));
   U82 : MUX2_X1 port map( A => n55, B => n57, S => n72, Z => Y(5));
   U85 : MUX2_X1 port map( A => n57, B => n59, S => n72, Z => Y(4));
   U88 : MUX2_X1 port map( A => n59, B => n61, S => n72, Z => Y(3));
   U91 : MUX2_X1 port map( A => n61, B => n63, S => n72, Z => Y(2));
   U92 : MUX2_X1 port map( A => n63, B => n64, S => n72, Z => Y(1));
   U97 : MUX2_X1 port map( A => n64, B => n67, S => n72, Z => Y(0));
   U102 : MUX2_X1 port map( A => n70, B => n7, S => n72, Z => Y(31));
   U93 : AOI22_X1 port map( A1 => n78, A2 => A(1), B1 => A(5), B2 => n76, ZN =>
                           n65);
   U86 : AOI22_X1 port map( A1 => sel(2), A2 => A(3), B1 => A(7), B2 => n77, ZN
                           => n60);
   U94 : AOI22_X1 port map( A1 => n74, A2 => n65, B1 => n60, B2 => n73, ZN => 
                           n64);
   U95 : AOI22_X1 port map( A1 => n78, A2 => A(0), B1 => A(4), B2 => n77, ZN =>
                           n66);
   U89 : AOI22_X1 port map( A1 => sel(2), A2 => A(2), B1 => A(6), B2 => n76, ZN
                           => n62);
   U96 : AOI22_X1 port map( A1 => n74, A2 => n66, B1 => n62, B2 => n73, ZN => 
                           n67);
   U26 : AOI22_X1 port map( A1 => n78, A2 => A(23), B1 => A(27), B2 => n76, ZN 
                           => n20);
   U20 : AOI22_X1 port map( A1 => n78, A2 => A(25), B1 => A(29), B2 => n76, ZN 
                           => n16);
   U27 : AOI22_X1 port map( A1 => n75, A2 => n20, B1 => n16, B2 => n73, ZN => 
                           n21);
   U29 : AOI22_X1 port map( A1 => sel(2), A2 => A(22), B1 => A(26), B2 => n76, 
                           ZN => n22);
   U23 : AOI22_X1 port map( A1 => n78, A2 => A(24), B1 => A(28), B2 => n76, ZN 
                           => n18);
   U30 : AOI22_X1 port map( A1 => n74, A2 => n22, B1 => n18, B2 => n73, ZN => 
                           n23);
   U32 : AOI22_X1 port map( A1 => sel(2), A2 => A(21), B1 => A(25), B2 => n76, 
                           ZN => n24);
   U33 : AOI22_X1 port map( A1 => n74, A2 => n24, B1 => n20, B2 => n73, ZN => 
                           n25);
   U35 : AOI22_X1 port map( A1 => sel(2), A2 => A(20), B1 => A(24), B2 => n77, 
                           ZN => n26);
   U36 : AOI22_X1 port map( A1 => n74, A2 => n26, B1 => n22, B2 => n73, ZN => 
                           n27);
   U38 : AOI22_X1 port map( A1 => sel(2), A2 => A(19), B1 => A(23), B2 => n77, 
                           ZN => n28);
   U39 : AOI22_X1 port map( A1 => n74, A2 => n28, B1 => n24, B2 => n73, ZN => 
                           n29);
   U41 : AOI22_X1 port map( A1 => sel(2), A2 => A(18), B1 => A(22), B2 => n77, 
                           ZN => n30);
   U42 : AOI22_X1 port map( A1 => n74, A2 => n30, B1 => n26, B2 => n73, ZN => 
                           n31);
   U17 : AOI22_X1 port map( A1 => n78, A2 => A(26), B1 => A(30), B2 => n76, ZN 
                           => n14);
   U24 : AOI22_X1 port map( A1 => n75, A2 => n18, B1 => n14, B2 => n73, ZN => 
                           n19);
   U11 : AOI22_X1 port map( A1 => sel(2), A2 => A(28), B1 => A(32), B2 => n76, 
                           ZN => n10);
   U5 : AOI22_X1 port map( A1 => sel(2), A2 => A(30), B1 => A(34), B2 => n76, 
                           ZN => n5);
   U12 : AOI22_X1 port map( A1 => sel(1), A2 => n10, B1 => n5, B2 => n73, ZN =>
                           n11);
   U14 : AOI22_X1 port map( A1 => n78, A2 => A(27), B1 => A(31), B2 => n76, ZN 
                           => n12);
   U8 : AOI22_X1 port map( A1 => sel(2), A2 => A(29), B1 => A(33), B2 => n76, 
                           ZN => n8);
   U15 : AOI22_X1 port map( A1 => n75, A2 => n12, B1 => n8, B2 => n73, ZN => 
                           n13);
   U18 : AOI22_X1 port map( A1 => n75, A2 => n14, B1 => n10, B2 => n73, ZN => 
                           n15);
   U44 : AOI22_X1 port map( A1 => n78, A2 => A(17), B1 => A(21), B2 => n77, ZN 
                           => n32);
   U45 : AOI22_X1 port map( A1 => n75, A2 => n32, B1 => n28, B2 => n73, ZN => 
                           n33);
   U21 : AOI22_X1 port map( A1 => n74, A2 => n16, B1 => n12, B2 => n73, ZN => 
                           n17);
   U2 : AOI22_X1 port map( A1 => sel(2), A2 => A(32), B1 => A(36), B2 => n76, 
                           ZN => n2);
   U100 : AOI22_X1 port map( A1 => sel(2), A2 => A(34), B1 => A(38), B2 => n77,
                           ZN => n69);
   U101 : AOI22_X1 port map( A1 => n74, A2 => n2, B1 => n69, B2 => n73, ZN => 
                           n70);
   U4 : AOI22_X1 port map( A1 => sel(2), A2 => A(31), B1 => A(35), B2 => n76, 
                           ZN => n4);
   U98 : AOI22_X1 port map( A1 => sel(2), A2 => A(33), B1 => A(37), B2 => n76, 
                           ZN => n68);
   U99 : AOI22_X1 port map( A1 => n74, A2 => n4, B1 => n68, B2 => n73, ZN => n7
                           );
   U6 : AOI22_X1 port map( A1 => sel(1), A2 => n5, B1 => n2, B2 => n73, ZN => 
                           n6);
   U9 : AOI22_X1 port map( A1 => sel(1), A2 => n8, B1 => n4, B2 => n73, ZN => 
                           n9);
   U47 : AOI22_X1 port map( A1 => sel(2), A2 => A(16), B1 => A(20), B2 => n77, 
                           ZN => n34);
   U48 : AOI22_X1 port map( A1 => n75, A2 => n34, B1 => n30, B2 => n73, ZN => 
                           n35);
   U50 : AOI22_X1 port map( A1 => sel(2), A2 => A(15), B1 => A(19), B2 => n77, 
                           ZN => n36);
   U51 : AOI22_X1 port map( A1 => n75, A2 => n36, B1 => n32, B2 => n73, ZN => 
                           n37);
   U71 : AOI22_X1 port map( A1 => n78, A2 => A(8), B1 => A(12), B2 => n76, ZN 
                           => n50);
   U65 : AOI22_X1 port map( A1 => n78, A2 => A(10), B1 => A(14), B2 => n77, ZN 
                           => n46);
   U72 : AOI22_X1 port map( A1 => n75, A2 => n50, B1 => n46, B2 => n73, ZN => 
                           n51);
   U74 : AOI22_X1 port map( A1 => n78, A2 => A(7), B1 => A(11), B2 => n77, ZN 
                           => n52);
   U68 : AOI22_X1 port map( A1 => n78, A2 => A(9), B1 => A(13), B2 => n77, ZN 
                           => n48);
   U75 : AOI22_X1 port map( A1 => n75, A2 => n52, B1 => n48, B2 => n73, ZN => 
                           n53);
   U59 : AOI22_X1 port map( A1 => n78, A2 => A(12), B1 => A(16), B2 => n77, ZN 
                           => n42);
   U53 : AOI22_X1 port map( A1 => sel(2), A2 => A(14), B1 => A(18), B2 => n77, 
                           ZN => n38);
   U60 : AOI22_X1 port map( A1 => n75, A2 => n42, B1 => n38, B2 => n73, ZN => 
                           n43);
   U62 : AOI22_X1 port map( A1 => n78, A2 => A(11), B1 => A(15), B2 => n77, ZN 
                           => n44);
   U56 : AOI22_X1 port map( A1 => sel(2), A2 => A(13), B1 => A(17), B2 => n77, 
                           ZN => n40);
   U63 : AOI22_X1 port map( A1 => n75, A2 => n44, B1 => n40, B2 => n73, ZN => 
                           n45);
   U54 : AOI22_X1 port map( A1 => n75, A2 => n38, B1 => n34, B2 => n73, ZN => 
                           n39);
   U57 : AOI22_X1 port map( A1 => n75, A2 => n40, B1 => n36, B2 => n73, ZN => 
                           n41);
   U66 : AOI22_X1 port map( A1 => n74, A2 => n46, B1 => n42, B2 => n73, ZN => 
                           n47);
   U69 : AOI22_X1 port map( A1 => n74, A2 => n48, B1 => n44, B2 => n73, ZN => 
                           n49);
   U83 : AOI22_X1 port map( A1 => n78, A2 => A(4), B1 => A(8), B2 => n77, ZN =>
                           n58);
   U77 : AOI22_X1 port map( A1 => n78, A2 => A(6), B1 => A(10), B2 => n76, ZN 
                           => n54);
   U84 : AOI22_X1 port map( A1 => n74, A2 => n58, B1 => n54, B2 => n73, ZN => 
                           n59);
   U80 : AOI22_X1 port map( A1 => n78, A2 => A(5), B1 => A(9), B2 => n77, ZN =>
                           n56);
   U87 : AOI22_X1 port map( A1 => n75, A2 => n60, B1 => n56, B2 => n73, ZN => 
                           n61);
   U78 : AOI22_X1 port map( A1 => n75, A2 => n54, B1 => n50, B2 => n73, ZN => 
                           n55);
   U90 : AOI22_X1 port map( A1 => n74, A2 => n62, B1 => n58, B2 => n73, ZN => 
                           n63);
   U81 : AOI22_X1 port map( A1 => n74, A2 => n56, B1 => n52, B2 => n73, ZN => 
                           n57);
   U1 : MUX2_X1 port map( A => n35, B => n37, S => n71, Z => Y(15));
   U3 : INV_X1 port map( A => sel(2), ZN => n76);
   U52 : INV_X1 port map( A => sel(2), ZN => n77);
   U103 : BUF_X1 port map( A => sel(0), Z => n71);
   U104 : BUF_X1 port map( A => sel(1), Z => n75);
   U105 : BUF_X1 port map( A => sel(0), Z => n72);
   U106 : INV_X2 port map( A => sel(1), ZN => n73);
   U107 : BUF_X1 port map( A => sel(2), Z => n78);
   U108 : BUF_X1 port map( A => sel(1), Z => n74);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity shift_secondLevel is

   port( sel : in std_logic_vector (1 downto 0);  mask00, mask08, mask16 : in 
         std_logic_vector (38 downto 0);  Y : out std_logic_vector (38 downto 
         0));

end shift_secondLevel;

architecture SYN_behav of shift_secondLevel is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n42, n43, n44, n45, n46, n48, n49, n50, n51, n52, n53, n54, n55, n56,
      n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71
      , n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n1, n2
      , n3, n4 : std_logic;

begin
   
   U57 : AOI222_X1 port map( A1 => n3, A2 => mask00(1), B1 => n44, B2 => 
                           mask16(1), C1 => n2, C2 => mask08(1), ZN => n72);
   U11 : AOI222_X1 port map( A1 => n3, A2 => mask00(5), B1 => n44, B2 => 
                           mask16(5), C1 => n2, C2 => mask08(5), ZN => n49);
   U15 : AOI222_X1 port map( A1 => n3, A2 => mask00(3), B1 => n44, B2 => 
                           mask16(3), C1 => n2, C2 => mask08(3), ZN => n51);
   U79 : AOI222_X1 port map( A1 => n3, A2 => mask00(0), B1 => n44, B2 => 
                           mask16(0), C1 => n2, C2 => mask08(0), ZN => n83);
   U13 : AOI222_X1 port map( A1 => n3, A2 => mask00(4), B1 => n44, B2 => 
                           mask16(4), C1 => n2, C2 => mask08(4), ZN => n50);
   U35 : AOI222_X1 port map( A1 => n4, A2 => mask00(2), B1 => n44, B2 => 
                           mask16(2), C1 => n45, C2 => mask08(2), ZN => n61);
   U9 : AOI222_X1 port map( A1 => n3, A2 => mask00(6), B1 => n44, B2 => 
                           mask16(6), C1 => n2, C2 => mask08(6), ZN => n48);
   U49 : AOI222_X1 port map( A1 => n4, A2 => mask00(23), B1 => n44, B2 => 
                           mask16(23), C1 => n45, C2 => mask08(23), ZN => n68);
   U41 : AOI222_X1 port map( A1 => n4, A2 => mask00(27), B1 => n44, B2 => 
                           mask16(27), C1 => n45, C2 => mask08(27), ZN => n64);
   U45 : AOI222_X1 port map( A1 => n4, A2 => mask00(25), B1 => n44, B2 => 
                           mask16(25), C1 => n45, C2 => mask08(25), ZN => n66);
   U37 : AOI222_X1 port map( A1 => n4, A2 => mask00(29), B1 => n44, B2 => 
                           mask16(29), C1 => n45, C2 => mask08(29), ZN => n62);
   U51 : AOI222_X1 port map( A1 => n4, A2 => mask00(22), B1 => n44, B2 => 
                           mask16(22), C1 => n45, C2 => mask08(22), ZN => n69);
   U43 : AOI222_X1 port map( A1 => n4, A2 => mask00(26), B1 => n44, B2 => 
                           mask16(26), C1 => n45, C2 => mask08(26), ZN => n65);
   U47 : AOI222_X1 port map( A1 => n4, A2 => mask00(24), B1 => n44, B2 => 
                           mask16(24), C1 => n45, C2 => mask08(24), ZN => n67);
   U39 : AOI222_X1 port map( A1 => n4, A2 => mask00(28), B1 => n44, B2 => 
                           mask16(28), C1 => n45, C2 => mask08(28), ZN => n63);
   U53 : AOI222_X1 port map( A1 => n4, A2 => mask00(21), B1 => n44, B2 => 
                           mask16(21), C1 => n45, C2 => mask08(21), ZN => n70);
   U55 : AOI222_X1 port map( A1 => n4, A2 => mask00(20), B1 => n44, B2 => 
                           mask16(20), C1 => n45, C2 => mask08(20), ZN => n71);
   U59 : AOI222_X1 port map( A1 => n3, A2 => mask00(19), B1 => n44, B2 => 
                           mask16(19), C1 => n2, C2 => mask08(19), ZN => n73);
   U61 : AOI222_X1 port map( A1 => n3, A2 => mask00(18), B1 => n44, B2 => 
                           mask16(18), C1 => n2, C2 => mask08(18), ZN => n74);
   U33 : AOI222_X1 port map( A1 => n4, A2 => mask00(30), B1 => n44, B2 => 
                           mask16(30), C1 => n45, C2 => mask08(30), ZN => n60);
   U29 : AOI222_X1 port map( A1 => n3, A2 => mask00(32), B1 => n44, B2 => 
                           mask16(32), C1 => n2, C2 => mask08(32), ZN => n58);
   U25 : AOI222_X1 port map( A1 => n3, A2 => mask00(34), B1 => n44, B2 => 
                           mask16(34), C1 => n2, C2 => mask08(34), ZN => n56);
   U31 : AOI222_X1 port map( A1 => n3, A2 => mask00(31), B1 => n44, B2 => 
                           mask16(31), C1 => n2, C2 => mask08(31), ZN => n59);
   U27 : AOI222_X1 port map( A1 => n3, A2 => mask00(33), B1 => n44, B2 => 
                           mask16(33), C1 => n2, C2 => mask08(33), ZN => n57);
   U63 : AOI222_X1 port map( A1 => n3, A2 => mask00(17), B1 => n44, B2 => 
                           mask16(17), C1 => n2, C2 => mask08(17), ZN => n75);
   U21 : AOI222_X1 port map( A1 => n3, A2 => mask00(36), B1 => n44, B2 => 
                           mask16(36), C1 => n2, C2 => mask08(36), ZN => n54);
   U17 : AOI222_X1 port map( A1 => n3, A2 => mask00(38), B1 => n44, B2 => 
                           mask16(38), C1 => n2, C2 => mask08(38), ZN => n52);
   U23 : AOI222_X1 port map( A1 => n3, A2 => mask00(35), B1 => n44, B2 => 
                           mask16(35), C1 => n2, C2 => mask08(35), ZN => n55);
   U19 : AOI222_X1 port map( A1 => n3, A2 => mask00(37), B1 => n44, B2 => 
                           mask16(37), C1 => n2, C2 => mask08(37), ZN => n53);
   U65 : AOI222_X1 port map( A1 => n3, A2 => mask00(16), B1 => n44, B2 => 
                           mask16(16), C1 => n2, C2 => mask08(16), ZN => n76);
   U67 : AOI222_X1 port map( A1 => n3, A2 => mask00(15), B1 => n44, B2 => 
                           mask16(15), C1 => n2, C2 => mask08(15), ZN => n77);
   U5 : AOI222_X1 port map( A1 => n4, A2 => mask00(8), B1 => n44, B2 => 
                           mask16(8), C1 => n2, C2 => mask08(8), ZN => n46);
   U73 : AOI222_X1 port map( A1 => n3, A2 => mask00(12), B1 => n44, B2 => 
                           mask16(12), C1 => n2, C2 => mask08(12), ZN => n80);
   U77 : AOI222_X1 port map( A1 => n3, A2 => mask00(10), B1 => n44, B2 => 
                           mask16(10), C1 => n2, C2 => mask08(10), ZN => n82);
   U69 : AOI222_X1 port map( A1 => n3, A2 => mask00(14), B1 => n44, B2 => 
                           mask16(14), C1 => n2, C2 => mask08(14), ZN => n78);
   U75 : AOI222_X1 port map( A1 => n3, A2 => mask00(11), B1 => n44, B2 => 
                           mask16(11), C1 => n2, C2 => mask08(11), ZN => n81);
   U3 : AOI222_X1 port map( A1 => n3, A2 => mask00(9), B1 => n44, B2 => 
                           mask16(9), C1 => n45, C2 => mask08(9), ZN => n42);
   U71 : AOI222_X1 port map( A1 => n3, A2 => mask00(13), B1 => n44, B2 => 
                           mask16(13), C1 => n2, C2 => mask08(13), ZN => n79);
   U82 : INV_X1 port map( A => sel(0), ZN => n84);
   U60 : INV_X1 port map( A => n74, ZN => Y(18));
   U62 : INV_X1 port map( A => n75, ZN => Y(17));
   U4 : INV_X1 port map( A => n46, ZN => Y(8));
   U52 : INV_X1 port map( A => n70, ZN => Y(21));
   U14 : INV_X1 port map( A => n51, ZN => Y(3));
   U64 : INV_X1 port map( A => n76, ZN => Y(16));
   U58 : INV_X1 port map( A => n73, ZN => Y(19));
   U50 : INV_X1 port map( A => n69, ZN => Y(22));
   U10 : INV_X1 port map( A => n49, ZN => Y(5));
   U56 : INV_X1 port map( A => n72, ZN => Y(1));
   U54 : INV_X1 port map( A => n71, ZN => Y(20));
   U66 : INV_X1 port map( A => n77, ZN => Y(15));
   U72 : INV_X1 port map( A => n80, ZN => Y(12));
   U68 : INV_X1 port map( A => n78, ZN => Y(14));
   U8 : INV_X1 port map( A => n48, ZN => Y(6));
   U34 : INV_X1 port map( A => n61, ZN => Y(2));
   U12 : INV_X1 port map( A => n50, ZN => Y(4));
   U74 : INV_X1 port map( A => n81, ZN => Y(11));
   U76 : INV_X1 port map( A => n82, ZN => Y(10));
   U2 : INV_X1 port map( A => n42, ZN => Y(9));
   U70 : INV_X1 port map( A => n79, ZN => Y(13));
   U78 : INV_X1 port map( A => n83, ZN => Y(0));
   U24 : INV_X1 port map( A => n56, ZN => Y(34));
   U26 : INV_X1 port map( A => n57, ZN => Y(33));
   U18 : INV_X1 port map( A => n53, ZN => Y(37));
   U32 : INV_X1 port map( A => n60, ZN => Y(30));
   U22 : INV_X1 port map( A => n55, ZN => Y(35));
   U20 : INV_X1 port map( A => n54, ZN => Y(36));
   U46 : INV_X1 port map( A => n67, ZN => Y(24));
   U30 : INV_X1 port map( A => n59, ZN => Y(31));
   U38 : INV_X1 port map( A => n63, ZN => Y(28));
   U16 : INV_X1 port map( A => n52, ZN => Y(38));
   U40 : INV_X1 port map( A => n64, ZN => Y(27));
   U42 : INV_X1 port map( A => n65, ZN => Y(26));
   U48 : INV_X1 port map( A => n68, ZN => Y(23));
   U44 : INV_X1 port map( A => n66, ZN => Y(25));
   U36 : INV_X1 port map( A => n62, ZN => Y(29));
   U28 : INV_X1 port map( A => n58, ZN => Y(32));
   U6 : AOI222_X1 port map( A1 => mask00(7), A2 => n3, B1 => mask08(7), B2 => 
                           n2, C1 => mask16(7), C2 => n44, ZN => n1);
   U7 : INV_X1 port map( A => n1, ZN => Y(7));
   U80 : BUF_X1 port map( A => n45, Z => n2);
   U81 : NOR2_X2 port map( A1 => sel(1), A2 => n84, ZN => n45);
   U83 : BUF_X2 port map( A => n43, Z => n3);
   U84 : BUF_X1 port map( A => n43, Z => n4);
   U85 : AND2_X2 port map( A1 => n84, A2 => sel(1), ZN => n44);
   U86 : NOR2_X1 port map( A1 => sel(1), A2 => sel(0), ZN => n43);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity shift_firstLevel is

   port( A : in std_logic_vector (31 downto 0);  sel : in std_logic_vector (1 
         downto 0);  mask00, mask08, mask16 : out std_logic_vector (38 downto 
         0));

end shift_firstLevel;

architecture SYN_behav of shift_firstLevel is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal mask08_38_port, mask08_37_port, mask08_36_port, mask08_35_port, 
      mask08_34_port, mask08_33_port, mask08_32_port, mask08_31_port, 
      mask08_23_port, mask08_22_port, mask08_21_port, mask08_20_port, 
      mask08_19_port, mask08_18_port, mask08_17_port, mask08_16_port, 
      mask08_15_port, mask08_7_port, mask08_6_port, mask08_5_port, 
      mask08_4_port, mask08_3_port, mask08_2_port, mask08_1_port, mask08_0_port
      , mask16_38_port, mask16_37_port, mask16_36_port, mask16_35_port, 
      mask16_34_port, mask16_33_port, mask16_32_port, mask16_31_port, 
      mask16_30_port, mask16_29_port, mask16_28_port, mask16_27_port, 
      mask16_26_port, mask16_25_port, mask16_24_port, mask16_23_port, 
      mask16_15_port, mask16_14_port, mask16_13_port, mask16_12_port, 
      mask16_11_port, mask16_10_port, mask16_9_port, mask16_8_port, 
      mask16_7_port, mask16_6_port, mask16_5_port, mask16_4_port, mask16_3_port
      , mask16_2_port, mask16_1_port, mask16_0_port, n37, n38, n39, n40, n41, 
      n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56
      , n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, 
      n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85
      , n86, n89, n90, n91, n92, n93, n94, n95, n96, n1, n2, n3, mask16_16_port
      : std_logic;

begin
   mask08 <= ( mask08_38_port, mask08_37_port, mask08_36_port, mask08_35_port, 
      mask08_34_port, mask08_33_port, mask08_32_port, mask08_31_port, 
      mask16_38_port, mask16_37_port, mask16_36_port, mask16_35_port, 
      mask16_34_port, mask16_33_port, mask16_32_port, mask08_23_port, 
      mask08_22_port, mask08_21_port, mask08_20_port, mask08_19_port, 
      mask08_18_port, mask08_17_port, mask08_16_port, mask08_15_port, 
      mask16_6_port, mask16_5_port, mask16_4_port, mask16_3_port, mask16_2_port
      , mask16_1_port, mask16_0_port, mask08_7_port, mask08_6_port, 
      mask08_5_port, mask08_4_port, mask08_3_port, mask08_2_port, mask08_1_port
      , mask08_0_port );
   mask16 <= ( mask16_38_port, mask16_37_port, mask16_36_port, mask16_35_port, 
      mask16_34_port, mask16_33_port, mask16_32_port, mask16_31_port, 
      mask16_30_port, mask16_29_port, mask16_28_port, mask16_27_port, 
      mask16_26_port, mask16_25_port, mask16_24_port, mask16_23_port, 
      mask16_16_port, mask16_16_port, mask16_16_port, mask16_16_port, 
      mask16_16_port, mask16_16_port, mask16_16_port, mask16_15_port, 
      mask16_14_port, mask16_13_port, mask16_12_port, mask16_11_port, 
      mask16_10_port, mask16_9_port, mask16_8_port, mask16_7_port, 
      mask16_6_port, mask16_5_port, mask16_4_port, mask16_3_port, mask16_2_port
      , mask16_1_port, mask16_0_port );
   
   U134 : NAND2_X1 port map( A1 => sel(0), A2 => A(17), ZN => n55);
   U59 : NAND2_X1 port map( A1 => sel(0), A2 => A(9), ZN => n79);
   U122 : NAND2_X1 port map( A1 => sel(0), A2 => A(21), ZN => n81);
   U146 : NAND2_X1 port map( A1 => sel(0), A2 => A(13), ZN => n59);
   U129 : NAND2_X1 port map( A1 => sel(0), A2 => A(19), ZN => n83);
   U152 : NAND2_X1 port map( A1 => sel(0), A2 => A(11), ZN => n61);
   U157 : NOR2_X1 port map( A1 => sel(0), A2 => sel(1), ZN => n86);
   U67 : NAND2_X1 port map( A1 => n2, A2 => A(0), ZN => n49);
   U116 : NAND2_X1 port map( A1 => sel(0), A2 => A(23), ZN => n39);
   U140 : NAND2_X1 port map( A1 => sel(0), A2 => A(15), ZN => n57);
   U137 : NAND2_X1 port map( A1 => sel(0), A2 => A(16), ZN => n56);
   U62 : NAND2_X1 port map( A1 => sel(0), A2 => A(8), ZN => n85);
   U125 : NAND2_X1 port map( A1 => sel(0), A2 => A(20), ZN => n82);
   U149 : NAND2_X1 port map( A1 => sel(0), A2 => A(12), ZN => n60);
   U131 : NAND2_X1 port map( A1 => sel(0), A2 => A(18), ZN => n84);
   U155 : NAND2_X1 port map( A1 => sel(0), A2 => A(10), ZN => n71);
   U119 : NAND2_X1 port map( A1 => sel(0), A2 => A(22), ZN => n80);
   U143 : NAND2_X1 port map( A1 => sel(0), A2 => A(14), ZN => n58);
   U115 : NAND2_X1 port map( A1 => n2, A2 => A(16), ZN => n69);
   U114 : NAND2_X1 port map( A1 => n39, A2 => n69, ZN => mask00(23));
   U91 : NAND2_X1 port map( A1 => sel(0), A2 => A(31), ZN => n78);
   U13 : NAND2_X1 port map( A1 => n3, A2 => n49, ZN => mask16_23_port);
   U141 : NAND2_X1 port map( A1 => n86, A2 => A(8), ZN => n40);
   U42 : NAND2_X1 port map( A1 => n40, A2 => n78, ZN => mask08_23_port);
   U104 : NAND2_X1 port map( A1 => sel(0), A2 => A(27), ZN => n53);
   U103 : NAND2_X1 port map( A1 => n2, A2 => A(20), ZN => n65);
   U102 : NAND2_X1 port map( A1 => n53, A2 => n65, ZN => mask00(27));
   U153 : NAND2_X1 port map( A1 => n2, A2 => A(4), ZN => n45);
   U9 : NAND2_X1 port map( A1 => n45, A2 => n41, ZN => mask16_27_port);
   U128 : NAND2_X1 port map( A1 => n86, A2 => A(12), ZN => n74);
   U38 : NAND2_X1 port map( A1 => n74, A2 => n3, ZN => mask16_35_port);
   U110 : NAND2_X1 port map( A1 => sel(0), A2 => A(25), ZN => n37);
   U109 : NAND2_X1 port map( A1 => n2, A2 => A(18), ZN => n67);
   U108 : NAND2_X1 port map( A1 => n37, A2 => n67, ZN => mask00(25));
   U60 : NAND2_X1 port map( A1 => n2, A2 => A(2), ZN => n47);
   U11 : NAND2_X1 port map( A1 => n3, A2 => n47, ZN => mask16_25_port);
   U135 : NAND2_X1 port map( A1 => n2, A2 => A(10), ZN => n76);
   U40 : NAND2_X1 port map( A1 => n76, A2 => n3, ZN => mask16_33_port);
   U98 : NAND2_X1 port map( A1 => sel(0), A2 => A(29), ZN => n51);
   U97 : NAND2_X1 port map( A1 => n2, A2 => A(22), ZN => n63);
   U96 : NAND2_X1 port map( A1 => n51, A2 => n63, ZN => mask00(29));
   U147 : NAND2_X1 port map( A1 => n86, A2 => A(6), ZN => n43);
   U7 : NAND2_X1 port map( A1 => n43, A2 => n41, ZN => mask16_29_port);
   U121 : NAND2_X1 port map( A1 => n86, A2 => A(14), ZN => n72);
   U36 : NAND2_X1 port map( A1 => n72, A2 => n3, ZN => mask16_37_port);
   U118 : NAND2_X1 port map( A1 => n2, A2 => A(15), ZN => n70);
   U117 : NAND2_X1 port map( A1 => n80, A2 => n70, ZN => mask00(22));
   U144 : NAND2_X1 port map( A1 => n2, A2 => A(7), ZN => n42);
   U94 : NAND2_X1 port map( A1 => sel(0), A2 => A(30), ZN => n50);
   U43 : NAND2_X1 port map( A1 => n42, A2 => n50, ZN => mask08_22_port);
   U107 : NAND2_X1 port map( A1 => sel(0), A2 => A(26), ZN => n54);
   U106 : NAND2_X1 port map( A1 => n2, A2 => A(19), ZN => n66);
   U105 : NAND2_X1 port map( A1 => n54, A2 => n66, ZN => mask00(26));
   U156 : NAND2_X1 port map( A1 => n2, A2 => A(3), ZN => n46);
   U10 : NAND2_X1 port map( A1 => n46, A2 => n41, ZN => mask16_26_port);
   U132 : NAND2_X1 port map( A1 => n86, A2 => A(11), ZN => n75);
   U39 : NAND2_X1 port map( A1 => n75, A2 => n3, ZN => mask16_34_port);
   U113 : NAND2_X1 port map( A1 => sel(0), A2 => A(24), ZN => n38);
   U112 : NAND2_X1 port map( A1 => n2, A2 => A(17), ZN => n68);
   U111 : NAND2_X1 port map( A1 => n38, A2 => n68, ZN => mask00(24));
   U63 : NAND2_X1 port map( A1 => n2, A2 => A(1), ZN => n48);
   U12 : NAND2_X1 port map( A1 => n3, A2 => n48, ZN => mask16_24_port);
   U138 : NAND2_X1 port map( A1 => n2, A2 => A(9), ZN => n77);
   U41 : NAND2_X1 port map( A1 => n77, A2 => n3, ZN => mask16_32_port);
   U101 : NAND2_X1 port map( A1 => sel(0), A2 => A(28), ZN => n52);
   U100 : NAND2_X1 port map( A1 => n2, A2 => A(21), ZN => n64);
   U99 : NAND2_X1 port map( A1 => n52, A2 => n64, ZN => mask00(28));
   U150 : NAND2_X1 port map( A1 => n2, A2 => A(5), ZN => n44);
   U8 : NAND2_X1 port map( A1 => n44, A2 => n41, ZN => mask16_28_port);
   U124 : NAND2_X1 port map( A1 => n86, A2 => A(13), ZN => n73);
   U37 : NAND2_X1 port map( A1 => n73, A2 => n3, ZN => mask16_36_port);
   U120 : NAND2_X1 port map( A1 => n81, A2 => n72, ZN => mask00(21));
   U44 : NAND2_X1 port map( A1 => n43, A2 => n51, ZN => mask08_21_port);
   U123 : NAND2_X1 port map( A1 => n82, A2 => n73, ZN => mask00(20));
   U45 : NAND2_X1 port map( A1 => n44, A2 => n52, ZN => mask08_20_port);
   U127 : NAND2_X1 port map( A1 => n83, A2 => n74, ZN => mask00(19));
   U47 : NAND2_X1 port map( A1 => n45, A2 => n53, ZN => mask08_19_port);
   U130 : NAND2_X1 port map( A1 => n75, A2 => n84, ZN => mask00(18));
   U48 : NAND2_X1 port map( A1 => n46, A2 => n54, ZN => mask08_18_port);
   U93 : NAND2_X1 port map( A1 => n2, A2 => A(23), ZN => n62);
   U92 : NAND2_X1 port map( A1 => n50, A2 => n62, ZN => mask00(30));
   U6 : NAND2_X1 port map( A1 => n42, A2 => n41, ZN => mask16_30_port);
   U34 : NAND2_X1 port map( A1 => n70, A2 => n3, ZN => mask16_38_port);
   U85 : AOI21_X1 port map( B1 => A(25), B2 => n2, A => mask16_16_port, ZN => 
                           n95);
   U32 : NAND2_X1 port map( A1 => n68, A2 => n3, ZN => mask08_32_port);
   U81 : AOI21_X1 port map( B1 => A(27), B2 => n2, A => mask16_16_port, ZN => 
                           n93);
   U30 : NAND2_X1 port map( A1 => n66, A2 => n41, ZN => mask08_34_port);
   U89 : AOI21_X1 port map( B1 => A(24), B2 => n2, A => mask16_15_port, ZN => 
                           n96);
   U5 : NAND2_X1 port map( A1 => n40, A2 => n41, ZN => mask16_31_port);
   U33 : NAND2_X1 port map( A1 => n69, A2 => n3, ZN => mask08_31_port);
   U83 : AOI21_X1 port map( B1 => A(26), B2 => n2, A => mask16_16_port, ZN => 
                           n94);
   U31 : NAND2_X1 port map( A1 => n67, A2 => n3, ZN => mask08_33_port);
   U133 : NAND2_X1 port map( A1 => n76, A2 => n55, ZN => mask00(17));
   U49 : NAND2_X1 port map( A1 => n37, A2 => n47, ZN => mask08_17_port);
   U77 : AOI21_X1 port map( B1 => A(29), B2 => n2, A => mask16_16_port, ZN => 
                           n91);
   U28 : NAND2_X1 port map( A1 => n64, A2 => n41, ZN => mask08_36_port);
   U73 : AOI21_X1 port map( B1 => A(31), B2 => n2, A => mask16_16_port, ZN => 
                           n89);
   U26 : NAND2_X1 port map( A1 => n62, A2 => n41, ZN => mask08_38_port);
   U79 : AOI21_X1 port map( B1 => A(28), B2 => n2, A => mask16_16_port, ZN => 
                           n92);
   U29 : NAND2_X1 port map( A1 => n65, A2 => n41, ZN => mask08_35_port);
   U75 : AOI21_X1 port map( B1 => A(30), B2 => n2, A => mask16_16_port, ZN => 
                           n90);
   U27 : NAND2_X1 port map( A1 => n63, A2 => n41, ZN => mask08_37_port);
   U136 : NAND2_X1 port map( A1 => n77, A2 => n56, ZN => mask00(16));
   U50 : NAND2_X1 port map( A1 => n38, A2 => n48, ZN => mask08_16_port);
   U139 : NAND2_X1 port map( A1 => n40, A2 => n57, ZN => mask00(15));
   U51 : NAND2_X1 port map( A1 => n39, A2 => n49, ZN => mask08_15_port);
   U61 : NAND2_X1 port map( A1 => n48, A2 => n85, ZN => mask00(8));
   U148 : NAND2_X1 port map( A1 => n44, A2 => n60, ZN => mask00(12));
   U154 : NAND2_X1 port map( A1 => n46, A2 => n71, ZN => mask00(10));
   U142 : NAND2_X1 port map( A1 => n42, A2 => n58, ZN => mask00(14));
   U151 : NAND2_X1 port map( A1 => n45, A2 => n61, ZN => mask00(11));
   U58 : NAND2_X1 port map( A1 => n47, A2 => n79, ZN => mask00(9));
   U145 : NAND2_X1 port map( A1 => n43, A2 => n59, ZN => mask00(13));
   U70 : AND2_X1 port map( A1 => sel(0), A2 => A(4), ZN => mask00(4));
   U158 : AND2_X1 port map( A1 => sel(0), A2 => A(0), ZN => mask00(0));
   U95 : AND2_X1 port map( A1 => sel(0), A2 => A(2), ZN => mask00(2));
   U68 : AND2_X1 port map( A1 => sel(0), A2 => A(6), ZN => mask00(6));
   U69 : AND2_X1 port map( A1 => sel(0), A2 => A(5), ZN => mask00(5));
   U71 : AND2_X1 port map( A1 => sel(0), A2 => A(3), ZN => mask00(3));
   U126 : AND2_X1 port map( A1 => sel(0), A2 => A(1), ZN => mask00(1));
   U3 : INV_X1 port map( A => n38, ZN => mask16_8_port);
   U15 : INV_X1 port map( A => n51, ZN => mask16_13_port);
   U16 : INV_X1 port map( A => n52, ZN => mask16_12_port);
   U2 : INV_X1 port map( A => n37, ZN => mask16_9_port);
   U17 : INV_X1 port map( A => n53, ZN => mask16_11_port);
   U18 : INV_X1 port map( A => n54, ZN => mask16_10_port);
   U14 : INV_X1 port map( A => n50, ZN => mask16_14_port);
   U57 : INV_X1 port map( A => n85, ZN => mask08_0_port);
   U20 : INV_X1 port map( A => n56, ZN => mask16_0_port);
   U54 : INV_X1 port map( A => n82, ZN => mask16_4_port);
   U24 : INV_X1 port map( A => n60, ZN => mask08_4_port);
   U25 : INV_X1 port map( A => n61, ZN => mask08_3_port);
   U55 : INV_X1 port map( A => n83, ZN => mask16_3_port);
   U23 : INV_X1 port map( A => n59, ZN => mask08_5_port);
   U53 : INV_X1 port map( A => n81, ZN => mask16_5_port);
   U56 : INV_X1 port map( A => n84, ZN => mask16_2_port);
   U46 : INV_X1 port map( A => n79, ZN => mask08_1_port);
   U19 : INV_X1 port map( A => n55, ZN => mask16_1_port);
   U35 : INV_X1 port map( A => n71, ZN => mask08_2_port);
   U52 : INV_X1 port map( A => n80, ZN => mask16_6_port);
   U22 : INV_X1 port map( A => n58, ZN => mask08_6_port);
   U90 : INV_X1 port map( A => n78, ZN => mask16_15_port);
   U88 : INV_X1 port map( A => n96, ZN => mask00(31));
   U78 : INV_X1 port map( A => n92, ZN => mask00(35));
   U74 : INV_X1 port map( A => n90, ZN => mask00(37));
   U82 : INV_X1 port map( A => n94, ZN => mask00(33));
   U84 : INV_X1 port map( A => n95, ZN => mask00(32));
   U76 : INV_X1 port map( A => n91, ZN => mask00(36));
   U72 : INV_X1 port map( A => n89, ZN => mask00(38));
   U80 : INV_X1 port map( A => n93, ZN => mask00(34));
   U4 : INV_X1 port map( A => n57, ZN => mask08_7_port);
   U21 : INV_X1 port map( A => n39, ZN => mask16_7_port);
   U64 : NAND2_X1 port map( A1 => sel(0), A2 => A(7), ZN => n1);
   U65 : NAND2_X1 port map( A1 => n49, A2 => n1, ZN => mask00(7));
   U66 : INV_X1 port map( A => mask16_16_port, ZN => n3);
   U86 : INV_X1 port map( A => n41, ZN => mask16_16_port);
   U87 : NAND2_X1 port map( A1 => sel(1), A2 => mask16_15_port, ZN => n41);
   U159 : BUF_X1 port map( A => n86, Z => n2);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_simple_booth_add_ext_N16 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_simple_booth_add_ext_N16;

architecture SYN_USE_DEFA_ARCH_NAME of 
   SNPS_CLOCK_GATE_HIGH_simple_booth_add_ext_N16 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net199337 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net199337);
   main_gate : AND2_X1 port map( A1 => net199337, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity piso_r_2_N32 is

   port( Clock, ALOAD : in std_logic;  D : in std_logic_vector (31 downto 0);  
         SO : out std_logic_vector (31 downto 0));

end piso_r_2_N32;

architecture SYN_archi of piso_r_2_N32 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component SDFF_X1
      port( D, SI, SE, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal SO_31_port, SO_30_port, SO_29_port, SO_28_port, SO_27_port, 
      SO_26_port, SO_25_port, SO_24_port, SO_23_port, SO_22_port, SO_21_port, 
      SO_20_port, SO_19_port, SO_18_port, SO_17_port, SO_16_port, SO_15_port, 
      SO_14_port, SO_13_port, SO_12_port, SO_11_port, SO_10_port, SO_9_port, 
      SO_8_port, SO_7_port, SO_6_port, SO_5_port, SO_4_port, SO_3_port, 
      SO_2_port, SO_1_port, SO_0_port, N3, N4, n2, n3_port, n4_port, n5, n6, n7
      , n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22
      , n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33 : std_logic;

begin
   SO <= ( SO_31_port, SO_30_port, SO_29_port, SO_28_port, SO_27_port, 
      SO_26_port, SO_25_port, SO_24_port, SO_23_port, SO_22_port, SO_21_port, 
      SO_20_port, SO_19_port, SO_18_port, SO_17_port, SO_16_port, SO_15_port, 
      SO_14_port, SO_13_port, SO_12_port, SO_11_port, SO_10_port, SO_9_port, 
      SO_8_port, SO_7_port, SO_6_port, SO_5_port, SO_4_port, SO_3_port, 
      SO_2_port, SO_1_port, SO_0_port );
   
   tmp_reg_1_inst : DFF_X1 port map( D => N4, CK => Clock, Q => SO_1_port, QN 
                           => n33);
   tmp_reg_3_inst : SDFF_X1 port map( D => SO_1_port, SI => D(3), SE => ALOAD, 
                           CK => Clock, Q => SO_3_port, QN => n32);
   tmp_reg_5_inst : SDFF_X1 port map( D => SO_3_port, SI => D(5), SE => ALOAD, 
                           CK => Clock, Q => SO_5_port, QN => n31);
   tmp_reg_7_inst : SDFF_X1 port map( D => SO_5_port, SI => D(7), SE => ALOAD, 
                           CK => Clock, Q => SO_7_port, QN => n30);
   tmp_reg_9_inst : SDFF_X1 port map( D => SO_7_port, SI => D(9), SE => ALOAD, 
                           CK => Clock, Q => SO_9_port, QN => n29);
   tmp_reg_11_inst : SDFF_X1 port map( D => SO_9_port, SI => D(11), SE => ALOAD
                           , CK => Clock, Q => SO_11_port, QN => n28);
   tmp_reg_13_inst : SDFF_X1 port map( D => SO_11_port, SI => D(13), SE => 
                           ALOAD, CK => Clock, Q => SO_13_port, QN => n27);
   tmp_reg_15_inst : SDFF_X1 port map( D => SO_13_port, SI => D(15), SE => 
                           ALOAD, CK => Clock, Q => SO_15_port, QN => n26);
   tmp_reg_17_inst : SDFF_X1 port map( D => SO_15_port, SI => D(17), SE => 
                           ALOAD, CK => Clock, Q => SO_17_port, QN => n25);
   tmp_reg_19_inst : SDFF_X1 port map( D => SO_17_port, SI => D(19), SE => 
                           ALOAD, CK => Clock, Q => SO_19_port, QN => n24);
   tmp_reg_21_inst : SDFF_X1 port map( D => SO_19_port, SI => D(21), SE => 
                           ALOAD, CK => Clock, Q => SO_21_port, QN => n23);
   tmp_reg_23_inst : SDFF_X1 port map( D => SO_21_port, SI => D(23), SE => 
                           ALOAD, CK => Clock, Q => SO_23_port, QN => n22);
   tmp_reg_25_inst : SDFF_X1 port map( D => SO_23_port, SI => D(25), SE => 
                           ALOAD, CK => Clock, Q => SO_25_port, QN => n21);
   tmp_reg_27_inst : SDFF_X1 port map( D => SO_25_port, SI => D(27), SE => 
                           ALOAD, CK => Clock, Q => SO_27_port, QN => n20);
   tmp_reg_29_inst : SDFF_X1 port map( D => SO_27_port, SI => D(29), SE => 
                           ALOAD, CK => Clock, Q => SO_29_port, QN => n19);
   tmp_reg_31_inst : SDFF_X1 port map( D => SO_29_port, SI => D(31), SE => 
                           ALOAD, CK => Clock, Q => SO_31_port, QN => n18);
   tmp_reg_0_inst : DFF_X1 port map( D => N3, CK => Clock, Q => SO_0_port, QN 
                           => n17);
   tmp_reg_2_inst : SDFF_X1 port map( D => SO_0_port, SI => D(2), SE => ALOAD, 
                           CK => Clock, Q => SO_2_port, QN => n16);
   tmp_reg_4_inst : SDFF_X1 port map( D => SO_2_port, SI => D(4), SE => ALOAD, 
                           CK => Clock, Q => SO_4_port, QN => n15);
   tmp_reg_6_inst : SDFF_X1 port map( D => SO_4_port, SI => D(6), SE => ALOAD, 
                           CK => Clock, Q => SO_6_port, QN => n14);
   tmp_reg_8_inst : SDFF_X1 port map( D => SO_6_port, SI => D(8), SE => ALOAD, 
                           CK => Clock, Q => SO_8_port, QN => n13);
   tmp_reg_10_inst : SDFF_X1 port map( D => SO_8_port, SI => D(10), SE => ALOAD
                           , CK => Clock, Q => SO_10_port, QN => n12);
   tmp_reg_12_inst : SDFF_X1 port map( D => SO_10_port, SI => D(12), SE => 
                           ALOAD, CK => Clock, Q => SO_12_port, QN => n11);
   tmp_reg_14_inst : SDFF_X1 port map( D => SO_12_port, SI => D(14), SE => 
                           ALOAD, CK => Clock, Q => SO_14_port, QN => n10);
   tmp_reg_16_inst : SDFF_X1 port map( D => SO_14_port, SI => D(16), SE => 
                           ALOAD, CK => Clock, Q => SO_16_port, QN => n9);
   tmp_reg_18_inst : SDFF_X1 port map( D => SO_16_port, SI => D(18), SE => 
                           ALOAD, CK => Clock, Q => SO_18_port, QN => n8);
   tmp_reg_20_inst : SDFF_X1 port map( D => SO_18_port, SI => D(20), SE => 
                           ALOAD, CK => Clock, Q => SO_20_port, QN => n7);
   tmp_reg_22_inst : SDFF_X1 port map( D => SO_20_port, SI => D(22), SE => 
                           ALOAD, CK => Clock, Q => SO_22_port, QN => n6);
   tmp_reg_24_inst : SDFF_X1 port map( D => SO_22_port, SI => D(24), SE => 
                           ALOAD, CK => Clock, Q => SO_24_port, QN => n5);
   tmp_reg_26_inst : SDFF_X1 port map( D => SO_24_port, SI => D(26), SE => 
                           ALOAD, CK => Clock, Q => SO_26_port, QN => n4_port);
   tmp_reg_28_inst : SDFF_X1 port map( D => SO_26_port, SI => D(28), SE => 
                           ALOAD, CK => Clock, Q => SO_28_port, QN => n3_port);
   tmp_reg_30_inst : SDFF_X1 port map( D => SO_28_port, SI => D(30), SE => 
                           ALOAD, CK => Clock, Q => SO_30_port, QN => n2);
   U4 : AND2_X1 port map( A1 => ALOAD, A2 => D(0), ZN => N3);
   U3 : AND2_X1 port map( A1 => ALOAD, A2 => D(1), ZN => N4);

end SYN_archi;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity shift_N9_0 is

   port( Clock, ALOAD : in std_logic;  D : in std_logic_vector (8 downto 0);  
         SO : out std_logic);

end shift_N9_0;

architecture SYN_archi of shift_N9_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component SDFF_X2
      port( D, SI, SE, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component SDFF_X1
      port( D, SI, SE, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal tmp_8_port, tmp_7_port, tmp_6_port, tmp_5_port, tmp_4_port, 
      tmp_3_port, tmp_2_port, tmp_1_port, N11, n3, n4, n5, n6, n7, n8, n9, n10,
      n1 : std_logic;

begin
   
   tmp_reg_8_inst : DFF_X1 port map( D => N11, CK => Clock, Q => tmp_8_port, QN
                           => n10);
   tmp_reg_7_inst : SDFF_X1 port map( D => tmp_8_port, SI => D(7), SE => ALOAD,
                           CK => Clock, Q => tmp_7_port, QN => n9);
   tmp_reg_6_inst : SDFF_X1 port map( D => tmp_7_port, SI => D(6), SE => ALOAD,
                           CK => Clock, Q => tmp_6_port, QN => n8);
   tmp_reg_5_inst : SDFF_X1 port map( D => tmp_6_port, SI => D(5), SE => ALOAD,
                           CK => Clock, Q => tmp_5_port, QN => n7);
   tmp_reg_4_inst : SDFF_X1 port map( D => tmp_5_port, SI => D(4), SE => ALOAD,
                           CK => Clock, Q => tmp_4_port, QN => n6);
   tmp_reg_3_inst : SDFF_X1 port map( D => tmp_4_port, SI => D(3), SE => ALOAD,
                           CK => Clock, Q => tmp_3_port, QN => n5);
   tmp_reg_2_inst : SDFF_X1 port map( D => tmp_3_port, SI => D(2), SE => ALOAD,
                           CK => Clock, Q => tmp_2_port, QN => n4);
   tmp_reg_1_inst : SDFF_X1 port map( D => tmp_2_port, SI => D(1), SE => ALOAD,
                           CK => Clock, Q => tmp_1_port, QN => n3);
   tmp_reg_0_inst : SDFF_X2 port map( D => tmp_1_port, SI => D(0), SE => ALOAD,
                           CK => Clock, Q => SO, QN => n1);
   U3 : AND2_X1 port map( A1 => ALOAD, A2 => D(8), ZN => N11);

end SYN_archi;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity booth_encoder_0 is

   port( B_in : in std_logic_vector (2 downto 0);  A_out : out std_logic_vector
         (2 downto 0));

end booth_encoder_0;

architecture SYN_bhe of booth_encoder_0 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal N53, N57, n3, n4 : std_logic;

begin
   A_out <= ( N57, B_in(2), N53 );
   
   U3 : INV_X1 port map( A => B_in(1), ZN => n3);
   U4 : INV_X1 port map( A => B_in(2), ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n3, ZN => N57);
   U6 : NOR2_X1 port map( A1 => B_in(1), A2 => n4, ZN => N53);

end SYN_bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity carry_sel_gen_N4_0 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end carry_sel_gen_N4_0;

architecture SYN_STRUCTURAL of carry_sel_gen_N4_0 is

   component mux21_SIZE4_0
      port( IN0, IN1 : in std_logic_vector (3 downto 0);  CTRL : in std_logic; 
            OUT1 : out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_N4_0
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic0_port, n5, nocarry_sum_to_mux_3_port, 
      nocarry_sum_to_mux_2_port, nocarry_sum_to_mux_1_port, 
      nocarry_sum_to_mux_0_port, n1, n2, n3, n4, net246126 : std_logic;

begin
   
   X_Logic0_port <= '0';
   rca_nocarry : RCA_N4_0 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           nocarry_sum_to_mux_3_port, S(2) => 
                           nocarry_sum_to_mux_2_port, S(1) => 
                           nocarry_sum_to_mux_1_port, S(0) => 
                           nocarry_sum_to_mux_0_port, Co => net246126);
   outmux : mux21_SIZE4_0 port map( IN0(3) => nocarry_sum_to_mux_3_port, IN0(2)
                           => nocarry_sum_to_mux_2_port, IN0(1) => 
                           nocarry_sum_to_mux_1_port, IN0(0) => 
                           nocarry_sum_to_mux_0_port, IN1(3) => n1, IN1(2) => 
                           n2, IN1(1) => n3, IN1(0) => n4, CTRL => n5, OUT1(3) 
                           => S(3), OUT1(2) => S(2), OUT1(1) => S(1), OUT1(0) 
                           => S(0));
   n1 <= '0';
   n2 <= '0';
   n3 <= '0';
   n4 <= '0';
   n5 <= '0';

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_0 is

   port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic);

end pg_0;

architecture SYN_beh of pg_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U3 : AOI21_X1 port map( B1 => g_prec, B2 => p, A => g, ZN => n2);
   U1 : AND2_X1 port map( A1 => p, A2 => p_prec, ZN => p_out);
   U2 : INV_X1 port map( A => n2, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity g_0 is

   port( g, p, g_prec : in std_logic;  g_out : out std_logic);

end g_0;

architecture SYN_beh of g_0 is

begin
   g_out <= g;

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity pg_net_0 is

   port( a, b : in std_logic;  g_out, p_out : out std_logic);

end pg_net_0;

architecture SYN_beh of pg_net_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p_out);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g_out);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity logic_unit_SIZE32 is

   port( IN1, IN2 : in std_logic_vector (31 downto 0);  CTRL : in 
         std_logic_vector (1 downto 0);  OUT1 : out std_logic_vector (31 downto
         0));

end logic_unit_SIZE32;

architecture SYN_Bhe of logic_unit_SIZE32 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X4
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, 
      n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32
      , n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, 
      n47, n48, n49, n50, n51, n52, n53, n56, n57, n58, n59, n60, n61, n62, n63
      , n64, n65, n1, n2, n54, n55 : std_logic;

begin
   
   U55 : AOI21_X1 port map( B1 => IN2(22), B2 => IN1(22), A => CTRL(0), ZN => 
                           n38);
   U54 : OAI22_X1 port map( A1 => IN1(22), A2 => IN2(22), B1 => n3, B2 => n38, 
                           ZN => n39);
   U53 : AOI21_X1 port map( B1 => n3, B2 => n38, A => n39, ZN => OUT1(22));
   U58 : AOI21_X1 port map( B1 => IN2(21), B2 => IN1(21), A => CTRL(0), ZN => 
                           n40);
   U57 : OAI22_X1 port map( A1 => IN1(21), A2 => IN2(21), B1 => n3, B2 => n40, 
                           ZN => n41);
   U56 : AOI21_X1 port map( B1 => n3, B2 => n40, A => n41, ZN => OUT1(21));
   U67 : AOI21_X1 port map( B1 => IN2(19), B2 => IN1(19), A => CTRL(0), ZN => 
                           n46);
   U66 : OAI22_X1 port map( A1 => IN1(19), A2 => IN2(19), B1 => n3, B2 => n46, 
                           ZN => n47);
   U65 : AOI21_X1 port map( B1 => n3, B2 => n46, A => n47, ZN => OUT1(19));
   U70 : AOI21_X1 port map( B1 => IN2(18), B2 => IN1(18), A => CTRL(0), ZN => 
                           n48);
   U69 : OAI22_X1 port map( A1 => IN1(18), A2 => IN2(18), B1 => n3, B2 => n48, 
                           ZN => n49);
   U68 : AOI21_X1 port map( B1 => n3, B2 => n48, A => n49, ZN => OUT1(18));
   U50 : AOI21_X1 port map( B1 => n3, B2 => n36, A => n37, ZN => OUT1(23));
   U40 : AOI21_X1 port map( B1 => IN2(27), B2 => IN1(27), A => CTRL(0), ZN => 
                           n28);
   U39 : OAI22_X1 port map( A1 => IN1(27), A2 => IN2(27), B1 => n3, B2 => n28, 
                           ZN => n29);
   U38 : AOI21_X1 port map( B1 => n3, B2 => n28, A => n29, ZN => OUT1(27));
   U43 : AOI21_X1 port map( B1 => IN2(26), B2 => IN1(26), A => CTRL(0), ZN => 
                           n30);
   U42 : OAI22_X1 port map( A1 => IN1(26), A2 => IN2(26), B1 => n3, B2 => n30, 
                           ZN => n31);
   U41 : AOI21_X1 port map( B1 => n3, B2 => n30, A => n31, ZN => OUT1(26));
   U71 : AOI21_X1 port map( B1 => n3, B2 => n50, A => n51, ZN => OUT1(17));
   U49 : AOI21_X1 port map( B1 => IN2(24), B2 => IN1(24), A => CTRL(0), ZN => 
                           n34);
   U48 : OAI22_X1 port map( A1 => IN1(24), A2 => IN2(24), B1 => n3, B2 => n34, 
                           ZN => n35);
   U47 : AOI21_X1 port map( B1 => n3, B2 => n34, A => n35, ZN => OUT1(24));
   U61 : AOI21_X1 port map( B1 => IN2(20), B2 => IN1(20), A => CTRL(0), ZN => 
                           n42);
   U60 : OAI22_X1 port map( A1 => IN1(20), A2 => IN2(20), B1 => n3, B2 => n42, 
                           ZN => n43);
   U59 : AOI21_X1 port map( B1 => n3, B2 => n42, A => n43, ZN => OUT1(20));
   U46 : AOI21_X1 port map( B1 => IN2(25), B2 => IN1(25), A => CTRL(0), ZN => 
                           n32);
   U45 : OAI22_X1 port map( A1 => IN1(25), A2 => IN2(25), B1 => n3, B2 => n32, 
                           ZN => n33);
   U44 : AOI21_X1 port map( B1 => n3, B2 => n32, A => n33, ZN => OUT1(25));
   U25 : AOI21_X1 port map( B1 => IN2(31), B2 => IN1(31), A => CTRL(0), ZN => 
                           n18);
   U24 : OAI22_X1 port map( A1 => IN1(31), A2 => IN2(31), B1 => n3, B2 => n18, 
                           ZN => n19);
   U23 : AOI21_X1 port map( B1 => n3, B2 => n18, A => n19, ZN => OUT1(31));
   U28 : AOI21_X1 port map( B1 => IN2(30), B2 => IN1(30), A => CTRL(0), ZN => 
                           n20);
   U27 : OAI22_X1 port map( A1 => IN1(30), A2 => IN2(30), B1 => n3, B2 => n20, 
                           ZN => n21);
   U26 : AOI21_X1 port map( B1 => n3, B2 => n20, A => n21, ZN => OUT1(30));
   U34 : AOI21_X1 port map( B1 => IN2(29), B2 => IN1(29), A => CTRL(0), ZN => 
                           n24);
   U33 : OAI22_X1 port map( A1 => IN1(29), A2 => IN2(29), B1 => n3, B2 => n24, 
                           ZN => n25);
   U32 : AOI21_X1 port map( B1 => n3, B2 => n24, A => n25, ZN => OUT1(29));
   U37 : AOI21_X1 port map( B1 => IN2(28), B2 => IN1(28), A => CTRL(0), ZN => 
                           n26);
   U36 : OAI22_X1 port map( A1 => IN1(28), A2 => IN2(28), B1 => n3, B2 => n26, 
                           ZN => n27);
   U35 : AOI21_X1 port map( B1 => n3, B2 => n26, A => n27, ZN => OUT1(28));
   U76 : AOI21_X1 port map( B1 => IN2(16), B2 => IN1(16), A => CTRL(0), ZN => 
                           n52);
   U75 : OAI22_X1 port map( A1 => IN1(16), A2 => IN2(16), B1 => n3, B2 => n52, 
                           ZN => n53);
   U74 : AOI21_X1 port map( B1 => n3, B2 => n52, A => n53, ZN => OUT1(16));
   U8 : AOI21_X1 port map( B1 => n3, B2 => n8, A => n9, ZN => OUT1(7));
   U89 : AOI21_X1 port map( B1 => n3, B2 => n62, A => n63, ZN => OUT1(11));
   U83 : AOI21_X1 port map( B1 => n3, B2 => n58, A => n59, ZN => OUT1(13));
   U82 : AOI21_X1 port map( B1 => IN2(14), B2 => IN1(14), A => CTRL(0), ZN => 
                           n56);
   U81 : OAI22_X1 port map( A1 => IN1(14), A2 => IN2(14), B1 => n3, B2 => n56, 
                           ZN => n57);
   U80 : AOI21_X1 port map( B1 => n3, B2 => n56, A => n57, ZN => OUT1(14));
   U88 : AOI21_X1 port map( B1 => IN2(12), B2 => IN1(12), A => CTRL(0), ZN => 
                           n60);
   U87 : OAI22_X1 port map( A1 => IN1(12), A2 => IN2(12), B1 => n3, B2 => n60, 
                           ZN => n61);
   U86 : AOI21_X1 port map( B1 => n3, B2 => n60, A => n61, ZN => OUT1(12));
   U94 : AOI21_X1 port map( B1 => IN2(10), B2 => IN1(10), A => CTRL(0), ZN => 
                           n64);
   U93 : OAI22_X1 port map( A1 => IN1(10), A2 => IN2(10), B1 => n3, B2 => n64, 
                           ZN => n65);
   U92 : AOI21_X1 port map( B1 => n3, B2 => n64, A => n65, ZN => OUT1(10));
   U2 : AOI21_X1 port map( B1 => n3, B2 => n4, A => n5, ZN => OUT1(9));
   U22 : AOI21_X1 port map( B1 => IN2(3), B2 => IN1(3), A => CTRL(0), ZN => n16
                           );
   U21 : OAI22_X1 port map( A1 => IN1(3), A2 => IN2(3), B1 => n3, B2 => n16, ZN
                           => n17);
   U20 : AOI21_X1 port map( B1 => n3, B2 => n16, A => n17, ZN => OUT1(3));
   U11 : AOI21_X1 port map( B1 => n3, B2 => n10, A => n11, ZN => OUT1(6));
   U62 : AOI21_X1 port map( B1 => n3, B2 => n44, A => n45, ZN => OUT1(1));
   U29 : AOI21_X1 port map( B1 => n3, B2 => n22, A => n23, ZN => OUT1(2));
   U14 : AOI21_X1 port map( B1 => n3, B2 => n12, A => n13, ZN => OUT1(5));
   U17 : AOI21_X1 port map( B1 => n3, B2 => n14, A => n15, ZN => OUT1(4));
   U7 : AOI21_X1 port map( B1 => IN2(8), B2 => IN1(8), A => CTRL(0), ZN => n6);
   U6 : OAI22_X1 port map( A1 => IN1(8), A2 => IN2(8), B1 => n3, B2 => n6, ZN 
                           => n7);
   U5 : AOI21_X1 port map( B1 => n3, B2 => n6, A => n7, ZN => OUT1(8));
   U3 : AOI21_X1 port map( B1 => IN1(0), B2 => IN2(0), A => CTRL(0), ZN => n1);
   U4 : OAI22_X1 port map( A1 => IN2(0), A2 => IN1(0), B1 => n3, B2 => n1, ZN 
                           => n2);
   U9 : AOI21_X1 port map( B1 => n3, B2 => n1, A => n2, ZN => OUT1(0));
   U10 : AOI21_X1 port map( B1 => IN1(15), B2 => IN2(15), A => CTRL(0), ZN => 
                           n54);
   U12 : OAI22_X1 port map( A1 => IN2(15), A2 => IN1(15), B1 => n3, B2 => n54, 
                           ZN => n55);
   U13 : AOI21_X1 port map( B1 => n3, B2 => n54, A => n55, ZN => OUT1(15));
   U15 : INV_X4 port map( A => CTRL(1), ZN => n3);
   U16 : OAI22_X1 port map( A1 => IN1(13), A2 => IN2(13), B1 => n3, B2 => n58, 
                           ZN => n59);
   U18 : AOI21_X1 port map( B1 => IN2(13), B2 => IN1(13), A => CTRL(0), ZN => 
                           n58);
   U19 : OAI22_X1 port map( A1 => IN1(17), A2 => IN2(17), B1 => n3, B2 => n50, 
                           ZN => n51);
   U30 : AOI21_X1 port map( B1 => IN2(17), B2 => IN1(17), A => CTRL(0), ZN => 
                           n50);
   U31 : OAI22_X1 port map( A1 => IN1(9), A2 => IN2(9), B1 => n3, B2 => n4, ZN 
                           => n5);
   U51 : AOI21_X1 port map( B1 => IN2(9), B2 => IN1(9), A => CTRL(0), ZN => n4)
                           ;
   U52 : OAI22_X1 port map( A1 => IN1(23), A2 => IN2(23), B1 => n3, B2 => n36, 
                           ZN => n37);
   U63 : AOI21_X1 port map( B1 => IN2(23), B2 => IN1(23), A => CTRL(0), ZN => 
                           n36);
   U64 : OAI22_X1 port map( A1 => IN1(11), A2 => IN2(11), B1 => n3, B2 => n62, 
                           ZN => n63);
   U72 : AOI21_X1 port map( B1 => IN2(11), B2 => IN1(11), A => CTRL(0), ZN => 
                           n62);
   U73 : OAI22_X1 port map( A1 => IN1(7), A2 => IN2(7), B1 => n3, B2 => n8, ZN 
                           => n9);
   U77 : AOI21_X1 port map( B1 => IN2(7), B2 => IN1(7), A => CTRL(0), ZN => n8)
                           ;
   U78 : OAI22_X1 port map( A1 => IN1(4), A2 => IN2(4), B1 => n3, B2 => n14, ZN
                           => n15);
   U79 : AOI21_X1 port map( B1 => IN2(4), B2 => IN1(4), A => CTRL(0), ZN => n14
                           );
   U84 : OAI22_X1 port map( A1 => IN1(2), A2 => IN2(2), B1 => n3, B2 => n22, ZN
                           => n23);
   U85 : AOI21_X1 port map( B1 => IN2(2), B2 => IN1(2), A => CTRL(0), ZN => n22
                           );
   U90 : OAI22_X1 port map( A1 => IN1(6), A2 => IN2(6), B1 => n3, B2 => n10, ZN
                           => n11);
   U91 : AOI21_X1 port map( B1 => IN2(6), B2 => IN1(6), A => CTRL(0), ZN => n10
                           );
   U95 : OAI22_X1 port map( A1 => IN1(5), A2 => IN2(5), B1 => n3, B2 => n12, ZN
                           => n13);
   U96 : AOI21_X1 port map( B1 => IN2(5), B2 => IN1(5), A => CTRL(0), ZN => n12
                           );
   U97 : OAI22_X1 port map( A1 => IN1(1), A2 => IN2(1), B1 => n3, B2 => n44, ZN
                           => n45);
   U98 : AOI21_X1 port map( B1 => IN2(1), B2 => IN1(1), A => CTRL(0), ZN => n44
                           );

end SYN_Bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity shifter is

   port( A : in std_logic_vector (31 downto 0);  B : in std_logic_vector (4 
         downto 0);  LOGIC_ARITH, LEFT_RIGHT : in std_logic;  OUTPUT : out 
         std_logic_vector (31 downto 0));

end shifter;

architecture SYN_struct of shifter is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X2
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component shift_thirdLevel
      port( sel : in std_logic_vector (2 downto 0);  A : in std_logic_vector 
            (38 downto 0);  Y : out std_logic_vector (31 downto 0));
   end component;
   
   component shift_secondLevel
      port( sel : in std_logic_vector (1 downto 0);  mask00, mask08, mask16 : 
            in std_logic_vector (38 downto 0);  Y : out std_logic_vector (38 
            downto 0));
   end component;
   
   component shift_firstLevel
      port( A : in std_logic_vector (31 downto 0);  sel : in std_logic_vector 
            (1 downto 0);  mask00, mask08, mask16 : out std_logic_vector (38 
            downto 0));
   end component;
   
   signal s3_2_port, s3_1_port, s3_0_port, m0_38_port, m0_37_port, m0_36_port, 
      m0_35_port, m0_34_port, m0_33_port, m0_32_port, m0_31_port, m0_30_port, 
      m0_29_port, m0_28_port, m0_27_port, m0_26_port, m0_25_port, m0_24_port, 
      m0_23_port, m0_22_port, m0_21_port, m0_20_port, m0_19_port, m0_18_port, 
      m0_17_port, m0_16_port, m0_15_port, m0_14_port, m0_13_port, m0_12_port, 
      m0_11_port, m0_10_port, m0_9_port, m0_8_port, m0_7_port, m0_6_port, 
      m0_5_port, m0_4_port, m0_3_port, m0_2_port, m0_1_port, m0_0_port, 
      m8_38_port, m8_37_port, m8_36_port, m8_35_port, m8_34_port, m8_33_port, 
      m8_32_port, m8_31_port, m8_30_port, m8_29_port, m8_28_port, m8_27_port, 
      m8_26_port, m8_25_port, m8_24_port, m8_23_port, m8_22_port, m8_21_port, 
      m8_20_port, m8_19_port, m8_18_port, m8_17_port, m8_16_port, m8_15_port, 
      m8_14_port, m8_13_port, m8_12_port, m8_11_port, m8_10_port, m8_9_port, 
      m8_8_port, m8_7_port, m8_6_port, m8_5_port, m8_4_port, m8_3_port, 
      m8_2_port, m8_1_port, m8_0_port, m16_38_port, m16_37_port, m16_36_port, 
      m16_35_port, m16_34_port, m16_33_port, m16_32_port, m16_31_port, 
      m16_30_port, m16_29_port, m16_28_port, m16_27_port, m16_26_port, 
      m16_25_port, m16_24_port, m16_23_port, m16_22_port, m16_21_port, 
      m16_20_port, m16_19_port, m16_18_port, m16_17_port, m16_16_port, 
      m16_15_port, m16_14_port, m16_13_port, m16_12_port, m16_11_port, 
      m16_10_port, m16_9_port, m16_8_port, m16_7_port, m16_6_port, m16_5_port, 
      m16_4_port, m16_3_port, m16_2_port, m16_1_port, m16_0_port, y_38_port, 
      y_37_port, y_36_port, y_35_port, y_34_port, y_33_port, y_32_port, 
      y_31_port, y_30_port, y_29_port, y_28_port, y_27_port, y_26_port, 
      y_25_port, y_24_port, y_23_port, y_22_port, y_21_port, y_20_port, 
      y_19_port, y_18_port, y_17_port, y_16_port, y_15_port, y_14_port, 
      y_13_port, y_12_port, y_11_port, y_10_port, y_9_port, y_8_port, y_7_port,
      y_6_port, y_5_port, y_4_port, y_3_port, y_2_port, y_1_port, y_0_port, n6,
      n8, n9, n10, n1 : std_logic;

begin
   
   IL : shift_firstLevel port map( A(31) => A(31), A(30) => A(30), A(29) => 
                           A(29), A(28) => A(28), A(27) => A(27), A(26) => 
                           A(26), A(25) => A(25), A(24) => A(24), A(23) => 
                           A(23), A(22) => A(22), A(21) => A(21), A(20) => 
                           A(20), A(19) => A(19), A(18) => A(18), A(17) => 
                           A(17), A(16) => A(16), A(15) => A(15), A(14) => 
                           A(14), A(13) => A(13), A(12) => A(12), A(11) => 
                           A(11), A(10) => A(10), A(9) => A(9), A(8) => A(8), 
                           A(7) => A(7), A(6) => A(6), A(5) => A(5), A(4) => 
                           A(4), A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), sel(1) => LOGIC_ARITH, sel(0) => LEFT_RIGHT
                           , mask00(38) => m0_38_port, mask00(37) => m0_37_port
                           , mask00(36) => m0_36_port, mask00(35) => m0_35_port
                           , mask00(34) => m0_34_port, mask00(33) => m0_33_port
                           , mask00(32) => m0_32_port, mask00(31) => m0_31_port
                           , mask00(30) => m0_30_port, mask00(29) => m0_29_port
                           , mask00(28) => m0_28_port, mask00(27) => m0_27_port
                           , mask00(26) => m0_26_port, mask00(25) => m0_25_port
                           , mask00(24) => m0_24_port, mask00(23) => m0_23_port
                           , mask00(22) => m0_22_port, mask00(21) => m0_21_port
                           , mask00(20) => m0_20_port, mask00(19) => m0_19_port
                           , mask00(18) => m0_18_port, mask00(17) => m0_17_port
                           , mask00(16) => m0_16_port, mask00(15) => m0_15_port
                           , mask00(14) => m0_14_port, mask00(13) => m0_13_port
                           , mask00(12) => m0_12_port, mask00(11) => m0_11_port
                           , mask00(10) => m0_10_port, mask00(9) => m0_9_port, 
                           mask00(8) => m0_8_port, mask00(7) => m0_7_port, 
                           mask00(6) => m0_6_port, mask00(5) => m0_5_port, 
                           mask00(4) => m0_4_port, mask00(3) => m0_3_port, 
                           mask00(2) => m0_2_port, mask00(1) => m0_1_port, 
                           mask00(0) => m0_0_port, mask08(38) => m8_38_port, 
                           mask08(37) => m8_37_port, mask08(36) => m8_36_port, 
                           mask08(35) => m8_35_port, mask08(34) => m8_34_port, 
                           mask08(33) => m8_33_port, mask08(32) => m8_32_port, 
                           mask08(31) => m8_31_port, mask08(30) => m8_30_port, 
                           mask08(29) => m8_29_port, mask08(28) => m8_28_port, 
                           mask08(27) => m8_27_port, mask08(26) => m8_26_port, 
                           mask08(25) => m8_25_port, mask08(24) => m8_24_port, 
                           mask08(23) => m8_23_port, mask08(22) => m8_22_port, 
                           mask08(21) => m8_21_port, mask08(20) => m8_20_port, 
                           mask08(19) => m8_19_port, mask08(18) => m8_18_port, 
                           mask08(17) => m8_17_port, mask08(16) => m8_16_port, 
                           mask08(15) => m8_15_port, mask08(14) => m8_14_port, 
                           mask08(13) => m8_13_port, mask08(12) => m8_12_port, 
                           mask08(11) => m8_11_port, mask08(10) => m8_10_port, 
                           mask08(9) => m8_9_port, mask08(8) => m8_8_port, 
                           mask08(7) => m8_7_port, mask08(6) => m8_6_port, 
                           mask08(5) => m8_5_port, mask08(4) => m8_4_port, 
                           mask08(3) => m8_3_port, mask08(2) => m8_2_port, 
                           mask08(1) => m8_1_port, mask08(0) => m8_0_port, 
                           mask16(38) => m16_38_port, mask16(37) => m16_37_port
                           , mask16(36) => m16_36_port, mask16(35) => 
                           m16_35_port, mask16(34) => m16_34_port, mask16(33) 
                           => m16_33_port, mask16(32) => m16_32_port, 
                           mask16(31) => m16_31_port, mask16(30) => m16_30_port
                           , mask16(29) => m16_29_port, mask16(28) => 
                           m16_28_port, mask16(27) => m16_27_port, mask16(26) 
                           => m16_26_port, mask16(25) => m16_25_port, 
                           mask16(24) => m16_24_port, mask16(23) => m16_23_port
                           , mask16(22) => m16_22_port, mask16(21) => 
                           m16_21_port, mask16(20) => m16_20_port, mask16(19) 
                           => m16_19_port, mask16(18) => m16_18_port, 
                           mask16(17) => m16_17_port, mask16(16) => m16_16_port
                           , mask16(15) => m16_15_port, mask16(14) => 
                           m16_14_port, mask16(13) => m16_13_port, mask16(12) 
                           => m16_12_port, mask16(11) => m16_11_port, 
                           mask16(10) => m16_10_port, mask16(9) => m16_9_port, 
                           mask16(8) => m16_8_port, mask16(7) => m16_7_port, 
                           mask16(6) => m16_6_port, mask16(5) => m16_5_port, 
                           mask16(4) => m16_4_port, mask16(3) => m16_3_port, 
                           mask16(2) => m16_2_port, mask16(1) => m16_1_port, 
                           mask16(0) => m16_0_port);
   IIL : shift_secondLevel port map( sel(1) => B(4), sel(0) => B(3), mask00(38)
                           => m0_38_port, mask00(37) => m0_37_port, mask00(36) 
                           => m0_36_port, mask00(35) => m0_35_port, mask00(34) 
                           => m0_34_port, mask00(33) => m0_33_port, mask00(32) 
                           => m0_32_port, mask00(31) => m0_31_port, mask00(30) 
                           => m0_30_port, mask00(29) => m0_29_port, mask00(28) 
                           => m0_28_port, mask00(27) => m0_27_port, mask00(26) 
                           => m0_26_port, mask00(25) => m0_25_port, mask00(24) 
                           => m0_24_port, mask00(23) => m0_23_port, mask00(22) 
                           => m0_22_port, mask00(21) => m0_21_port, mask00(20) 
                           => m0_20_port, mask00(19) => m0_19_port, mask00(18) 
                           => m0_18_port, mask00(17) => m0_17_port, mask00(16) 
                           => m0_16_port, mask00(15) => m0_15_port, mask00(14) 
                           => m0_14_port, mask00(13) => m0_13_port, mask00(12) 
                           => m0_12_port, mask00(11) => m0_11_port, mask00(10) 
                           => m0_10_port, mask00(9) => m0_9_port, mask00(8) => 
                           m0_8_port, mask00(7) => m0_7_port, mask00(6) => 
                           m0_6_port, mask00(5) => m0_5_port, mask00(4) => 
                           m0_4_port, mask00(3) => m0_3_port, mask00(2) => 
                           m0_2_port, mask00(1) => m0_1_port, mask00(0) => 
                           m0_0_port, mask08(38) => m8_38_port, mask08(37) => 
                           m8_37_port, mask08(36) => m8_36_port, mask08(35) => 
                           m8_35_port, mask08(34) => m8_34_port, mask08(33) => 
                           m8_33_port, mask08(32) => m8_32_port, mask08(31) => 
                           m8_31_port, mask08(30) => m8_30_port, mask08(29) => 
                           m8_29_port, mask08(28) => m8_28_port, mask08(27) => 
                           m8_27_port, mask08(26) => m8_26_port, mask08(25) => 
                           m8_25_port, mask08(24) => m8_24_port, mask08(23) => 
                           m8_23_port, mask08(22) => m8_22_port, mask08(21) => 
                           m8_21_port, mask08(20) => m8_20_port, mask08(19) => 
                           m8_19_port, mask08(18) => m8_18_port, mask08(17) => 
                           m8_17_port, mask08(16) => m8_16_port, mask08(15) => 
                           m8_15_port, mask08(14) => m8_14_port, mask08(13) => 
                           m8_13_port, mask08(12) => m8_12_port, mask08(11) => 
                           m8_11_port, mask08(10) => m8_10_port, mask08(9) => 
                           m8_9_port, mask08(8) => m8_8_port, mask08(7) => 
                           m8_7_port, mask08(6) => m8_6_port, mask08(5) => 
                           m8_5_port, mask08(4) => m8_4_port, mask08(3) => 
                           m8_3_port, mask08(2) => m8_2_port, mask08(1) => 
                           m8_1_port, mask08(0) => m8_0_port, mask16(38) => 
                           m16_38_port, mask16(37) => m16_37_port, mask16(36) 
                           => m16_36_port, mask16(35) => m16_35_port, 
                           mask16(34) => m16_34_port, mask16(33) => m16_33_port
                           , mask16(32) => m16_32_port, mask16(31) => 
                           m16_31_port, mask16(30) => m16_30_port, mask16(29) 
                           => m16_29_port, mask16(28) => m16_28_port, 
                           mask16(27) => m16_27_port, mask16(26) => m16_26_port
                           , mask16(25) => m16_25_port, mask16(24) => 
                           m16_24_port, mask16(23) => m16_23_port, mask16(22) 
                           => m16_22_port, mask16(21) => m16_21_port, 
                           mask16(20) => m16_20_port, mask16(19) => m16_19_port
                           , mask16(18) => m16_18_port, mask16(17) => 
                           m16_17_port, mask16(16) => m16_16_port, mask16(15) 
                           => m16_15_port, mask16(14) => m16_14_port, 
                           mask16(13) => m16_13_port, mask16(12) => m16_12_port
                           , mask16(11) => m16_11_port, mask16(10) => 
                           m16_10_port, mask16(9) => m16_9_port, mask16(8) => 
                           m16_8_port, mask16(7) => m16_7_port, mask16(6) => 
                           m16_6_port, mask16(5) => m16_5_port, mask16(4) => 
                           m16_4_port, mask16(3) => m16_3_port, mask16(2) => 
                           m16_2_port, mask16(1) => m16_1_port, mask16(0) => 
                           m16_0_port, Y(38) => y_38_port, Y(37) => y_37_port, 
                           Y(36) => y_36_port, Y(35) => y_35_port, Y(34) => 
                           y_34_port, Y(33) => y_33_port, Y(32) => y_32_port, 
                           Y(31) => y_31_port, Y(30) => y_30_port, Y(29) => 
                           y_29_port, Y(28) => y_28_port, Y(27) => y_27_port, 
                           Y(26) => y_26_port, Y(25) => y_25_port, Y(24) => 
                           y_24_port, Y(23) => y_23_port, Y(22) => y_22_port, 
                           Y(21) => y_21_port, Y(20) => y_20_port, Y(19) => 
                           y_19_port, Y(18) => y_18_port, Y(17) => y_17_port, 
                           Y(16) => y_16_port, Y(15) => y_15_port, Y(14) => 
                           y_14_port, Y(13) => y_13_port, Y(12) => y_12_port, 
                           Y(11) => y_11_port, Y(10) => y_10_port, Y(9) => 
                           y_9_port, Y(8) => y_8_port, Y(7) => y_7_port, Y(6) 
                           => y_6_port, Y(5) => y_5_port, Y(4) => y_4_port, 
                           Y(3) => y_3_port, Y(2) => y_2_port, Y(1) => y_1_port
                           , Y(0) => y_0_port);
   IIIL : shift_thirdLevel port map( sel(2) => s3_2_port, sel(1) => s3_1_port, 
                           sel(0) => s3_0_port, A(38) => y_38_port, A(37) => 
                           y_37_port, A(36) => y_36_port, A(35) => y_35_port, 
                           A(34) => y_34_port, A(33) => y_33_port, A(32) => 
                           y_32_port, A(31) => y_31_port, A(30) => y_30_port, 
                           A(29) => y_29_port, A(28) => y_28_port, A(27) => 
                           y_27_port, A(26) => y_26_port, A(25) => y_25_port, 
                           A(24) => y_24_port, A(23) => y_23_port, A(22) => 
                           y_22_port, A(21) => y_21_port, A(20) => y_20_port, 
                           A(19) => y_19_port, A(18) => y_18_port, A(17) => 
                           y_17_port, A(16) => y_16_port, A(15) => y_15_port, 
                           A(14) => y_14_port, A(13) => y_13_port, A(12) => 
                           y_12_port, A(11) => y_11_port, A(10) => y_10_port, 
                           A(9) => y_9_port, A(8) => y_8_port, A(7) => y_7_port
                           , A(6) => y_6_port, A(5) => y_5_port, A(4) => 
                           y_4_port, A(3) => y_3_port, A(2) => y_2_port, A(1) 
                           => y_1_port, A(0) => y_0_port, Y(31) => OUTPUT(31), 
                           Y(30) => OUTPUT(30), Y(29) => OUTPUT(29), Y(28) => 
                           OUTPUT(28), Y(27) => OUTPUT(27), Y(26) => OUTPUT(26)
                           , Y(25) => OUTPUT(25), Y(24) => OUTPUT(24), Y(23) =>
                           OUTPUT(23), Y(22) => OUTPUT(22), Y(21) => OUTPUT(21)
                           , Y(20) => OUTPUT(20), Y(19) => OUTPUT(19), Y(18) =>
                           OUTPUT(18), Y(17) => OUTPUT(17), Y(16) => OUTPUT(16)
                           , Y(15) => OUTPUT(15), Y(14) => OUTPUT(14), Y(13) =>
                           OUTPUT(13), Y(12) => OUTPUT(12), Y(11) => OUTPUT(11)
                           , Y(10) => OUTPUT(10), Y(9) => OUTPUT(9), Y(8) => 
                           OUTPUT(8), Y(7) => OUTPUT(7), Y(6) => OUTPUT(6), 
                           Y(5) => OUTPUT(5), Y(4) => OUTPUT(4), Y(3) => 
                           OUTPUT(3), Y(2) => OUTPUT(2), Y(1) => OUTPUT(1), 
                           Y(0) => OUTPUT(0));
   U8 : OR2_X1 port map( A1 => LOGIC_ARITH, A2 => LEFT_RIGHT, ZN => n6);
   U1 : INV_X1 port map( A => B(0), ZN => n10);
   U2 : INV_X1 port map( A => B(1), ZN => n9);
   U3 : INV_X1 port map( A => B(2), ZN => n8);
   U4 : INV_X1 port map( A => LEFT_RIGHT, ZN => n1);
   U5 : AOI22_X2 port map( A1 => B(2), A2 => n6, B1 => n1, B2 => n8, ZN => 
                           s3_2_port);
   U6 : AOI22_X1 port map( A1 => B(1), A2 => n6, B1 => n1, B2 => n9, ZN => 
                           s3_1_port);
   U7 : AOI22_X1 port map( A1 => B(0), A2 => n6, B1 => n1, B2 => n10, ZN => 
                           s3_0_port);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity comparator_M32 is

   port( C, V : in std_logic;  SUM : in std_logic_vector (31 downto 0);  sel : 
         in std_logic_vector (2 downto 0);  sign : in std_logic;  S : out 
         std_logic);

end comparator_M32;

architecture SYN_BEHAVIORAL of comparator_M32 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n13, n12, n6, n1, n2, n3, n4, n5, n7, n8, n9, n10, n11, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37 : std_logic;

begin
   
   U1 : NOR4_X1 port map( A1 => SUM(14), A2 => SUM(13), A3 => SUM(15), A4 => 
                           SUM(16), ZN => n18);
   U2 : OR4_X1 port map( A1 => SUM(4), A2 => SUM(3), A3 => SUM(6), A4 => SUM(5)
                           , ZN => n15);
   U3 : OR2_X1 port map( A1 => C, A2 => sign, ZN => n7);
   U4 : OR2_X1 port map( A1 => SUM(7), A2 => SUM(8), ZN => n14);
   U5 : INV_X1 port map( A => n7, ZN => n1);
   U6 : NOR2_X1 port map( A1 => n31, A2 => n1, ZN => n5);
   U7 : OAI21_X1 port map( B1 => sel(2), B2 => sel(0), A => n31, ZN => n2);
   U8 : INV_X1 port map( A => n2, ZN => n3);
   U9 : INV_X1 port map( A => SUM(10), ZN => n25);
   U10 : INV_X1 port map( A => SUM(0), ZN => n26);
   U11 : INV_X1 port map( A => n36, ZN => n37);
   U12 : INV_X1 port map( A => sel(1), ZN => n35);
   U13 : INV_X1 port map( A => sel(2), ZN => n30);
   U14 : NAND2_X1 port map( A1 => n34, A2 => n3, ZN => n27);
   U15 : AND2_X1 port map( A1 => n12, A2 => n5, ZN => n32);
   U16 : OR2_X1 port map( A1 => n6, A2 => sel(0), ZN => n33);
   U17 : NAND2_X1 port map( A1 => n35, A2 => n30, ZN => n31);
   U18 : OAI21_X1 port map( B1 => sel(1), B2 => sel(0), A => sel(2), ZN => n36)
                           ;
   U19 : NOR4_X1 port map( A1 => SUM(31), A2 => SUM(9), A3 => n14, A4 => n15, 
                           ZN => n11);
   U20 : NOR2_X1 port map( A1 => SUM(19), A2 => SUM(1), ZN => n20);
   U21 : NOR2_X1 port map( A1 => SUM(18), A2 => SUM(17), ZN => n19);
   U22 : NOR3_X1 port map( A1 => SUM(11), A2 => SUM(12), A3 => n24, ZN => n22);
   U23 : NAND4_X1 port map( A1 => n8, A2 => n9, A3 => n10, A4 => n11, ZN => n6)
                           ;
   U24 : XNOR2_X1 port map( A => n6, B => n37, ZN => n34);
   U25 : NAND3_X1 port map( A1 => n4, A2 => n30, A3 => n31, ZN => n29);
   U26 : NAND2_X1 port map( A1 => n12, A2 => n7, ZN => n4);
   U27 : NAND3_X1 port map( A1 => n27, A2 => n28, A3 => n29, ZN => S);
   U28 : NAND2_X1 port map( A1 => SUM(31), A2 => V, ZN => n13);
   U29 : OAI211_X1 port map( C1 => V, C2 => SUM(31), A => n13, B => sign, ZN =>
                           n12);
   U30 : NAND3_X1 port map( A1 => n18, A2 => n19, A3 => n20, ZN => n17);
   U31 : NAND3_X1 port map( A1 => n21, A2 => n22, A3 => n23, ZN => n16);
   U32 : NOR2_X1 port map( A1 => SUM(23), A2 => SUM(22), ZN => n21);
   U33 : NAND2_X1 port map( A1 => n25, A2 => n26, ZN => n24);
   U34 : NOR2_X1 port map( A1 => SUM(21), A2 => SUM(20), ZN => n23);
   U35 : NOR2_X1 port map( A1 => n16, A2 => n17, ZN => n8);
   U36 : NOR4_X1 port map( A1 => SUM(27), A2 => SUM(26), A3 => SUM(25), A4 => 
                           SUM(24), ZN => n9);
   U37 : NOR4_X1 port map( A1 => SUM(29), A2 => SUM(30), A3 => SUM(28), A4 => 
                           SUM(2), ZN => n10);
   U38 : NAND2_X1 port map( A1 => n33, A2 => n32, ZN => n28);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity simple_booth_add_ext_N16 is

   port( Clock, Reset, sign, enable : in std_logic;  valid : out std_logic;  A,
         B : in std_logic_vector (15 downto 0);  A_to_add, B_to_add : out 
         std_logic_vector (31 downto 0);  sign_to_add : out std_logic;  
         final_out : out std_logic_vector (31 downto 0);  ACC_from_add : in 
         std_logic_vector (31 downto 0));

end simple_booth_add_ext_N16;

architecture SYN_struct of simple_booth_add_ext_N16 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X4
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_simple_booth_add_ext_N16
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component ff32_en_SIZE32_1
      port( D : in std_logic_vector (31 downto 0);  en, clk, rst : in std_logic
            ;  Q : out std_logic_vector (31 downto 0));
   end component;
   
   component mux21_1
      port( IN0, IN1 : in std_logic_vector (31 downto 0);  CTRL : in std_logic;
            OUT1 : out std_logic_vector (31 downto 0));
   end component;
   
   component piso_r_2_N32
      port( Clock, ALOAD : in std_logic;  D : in std_logic_vector (31 downto 0)
            ;  SO : out std_logic_vector (31 downto 0));
   end component;
   
   component shift_N9_1
      port( Clock, ALOAD : in std_logic;  D : in std_logic_vector (8 downto 0);
            SO : out std_logic);
   end component;
   
   component shift_N9_2
      port( Clock, ALOAD : in std_logic;  D : in std_logic_vector (8 downto 0);
            SO : out std_logic);
   end component;
   
   component shift_N9_0
      port( Clock, ALOAD : in std_logic;  D : in std_logic_vector (8 downto 0);
            SO : out std_logic);
   end component;
   
   component booth_encoder_1
      port( B_in : in std_logic_vector (2 downto 0);  A_out : out 
            std_logic_vector (2 downto 0));
   end component;
   
   component booth_encoder_2
      port( B_in : in std_logic_vector (2 downto 0);  A_out : out 
            std_logic_vector (2 downto 0));
   end component;
   
   component booth_encoder_3
      port( B_in : in std_logic_vector (2 downto 0);  A_out : out 
            std_logic_vector (2 downto 0));
   end component;
   
   component booth_encoder_4
      port( B_in : in std_logic_vector (2 downto 0);  A_out : out 
            std_logic_vector (2 downto 0));
   end component;
   
   component booth_encoder_5
      port( B_in : in std_logic_vector (2 downto 0);  A_out : out 
            std_logic_vector (2 downto 0));
   end component;
   
   component booth_encoder_6
      port( B_in : in std_logic_vector (2 downto 0);  A_out : out 
            std_logic_vector (2 downto 0));
   end component;
   
   component booth_encoder_7
      port( B_in : in std_logic_vector (2 downto 0);  A_out : out 
            std_logic_vector (2 downto 0));
   end component;
   
   component booth_encoder_8
      port( B_in : in std_logic_vector (2 downto 0);  A_out : out 
            std_logic_vector (2 downto 0));
   end component;
   
   component booth_encoder_0
      port( B_in : in std_logic_vector (2 downto 0);  A_out : out 
            std_logic_vector (2 downto 0));
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFS_X1
      port( D, CK, SN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal X_Logic0_port, valid_port, A_to_add_31_port, A_to_add_30_port, 
      A_to_add_29_port, A_to_add_28_port, A_to_add_27_port, A_to_add_26_port, 
      A_to_add_25_port, A_to_add_24_port, A_to_add_23_port, A_to_add_22_port, 
      A_to_add_21_port, A_to_add_20_port, A_to_add_19_port, A_to_add_18_port, 
      A_to_add_17_port, A_to_add_16_port, A_to_add_15_port, A_to_add_14_port, 
      A_to_add_13_port, A_to_add_12_port, A_to_add_11_port, A_to_add_10_port, 
      A_to_add_9_port, A_to_add_8_port, A_to_add_7_port, A_to_add_6_port, 
      A_to_add_5_port, A_to_add_4_port, A_to_add_3_port, A_to_add_2_port, 
      A_to_add_1_port, A_to_add_0_port, enc_N2_in_2_port, piso_0_in_8_port, 
      piso_0_in_7_port, piso_0_in_6_port, piso_0_in_5_port, piso_0_in_4_port, 
      piso_0_in_3_port, piso_0_in_2_port, piso_0_in_1_port, piso_0_in_0_port, 
      piso_1_in_8_port, piso_1_in_7_port, piso_1_in_6_port, piso_1_in_5_port, 
      piso_1_in_4_port, piso_1_in_3_port, piso_1_in_2_port, piso_1_in_1_port, 
      piso_1_in_0_port, piso_2_in_8_port, piso_2_in_7_port, piso_2_in_6_port, 
      piso_2_in_5_port, piso_2_in_4_port, piso_2_in_3_port, piso_2_in_2_port, 
      piso_2_in_1_port, piso_2_in_0_port, extend_vector_15_port, 
      A_to_mux_31_port, A_to_mux_30_port, A_to_mux_29_port, A_to_mux_28_port, 
      A_to_mux_27_port, A_to_mux_26_port, A_to_mux_25_port, A_to_mux_24_port, 
      A_to_mux_23_port, A_to_mux_22_port, A_to_mux_21_port, A_to_mux_20_port, 
      A_to_mux_19_port, A_to_mux_18_port, A_to_mux_17_port, A_to_mux_16_port, 
      A_to_mux_15_port, A_to_mux_14_port, A_to_mux_13_port, A_to_mux_12_port, 
      A_to_mux_11_port, A_to_mux_10_port, A_to_mux_9_port, A_to_mux_8_port, 
      A_to_mux_7_port, A_to_mux_6_port, A_to_mux_5_port, A_to_mux_4_port, 
      A_to_mux_3_port, A_to_mux_2_port, A_to_mux_1_port, A_to_mux_0_port, 
      input_mux_sel_2_port, input_mux_sel_0, next_accumulate_31_port, 
      next_accumulate_30_port, next_accumulate_29_port, next_accumulate_28_port
      , next_accumulate_27_port, next_accumulate_26_port, 
      next_accumulate_25_port, next_accumulate_24_port, next_accumulate_23_port
      , next_accumulate_22_port, next_accumulate_21_port, 
      next_accumulate_20_port, next_accumulate_19_port, next_accumulate_18_port
      , next_accumulate_17_port, next_accumulate_16_port, 
      next_accumulate_15_port, next_accumulate_14_port, next_accumulate_13_port
      , next_accumulate_12_port, next_accumulate_11_port, 
      next_accumulate_10_port, next_accumulate_9_port, next_accumulate_8_port, 
      next_accumulate_7_port, next_accumulate_6_port, next_accumulate_5_port, 
      next_accumulate_4_port, next_accumulate_3_port, next_accumulate_2_port, 
      next_accumulate_1_port, next_accumulate_0_port, reg_enable, count_4_port,
      count_3_port, count_2_port, count_1_port, count_0_port, N23, N37, N39, 
      N41, N43, N44, N45, net199343, n2, n3, n5, n8, n9, n10, n11, n1, n4, n6, 
      n7, n12, n13, n14, n15, n16, n17, n18 : std_logic;

begin
   valid <= valid_port;
   A_to_add <= ( A_to_add_31_port, A_to_add_30_port, A_to_add_29_port, 
      A_to_add_28_port, A_to_add_27_port, A_to_add_26_port, A_to_add_25_port, 
      A_to_add_24_port, A_to_add_23_port, A_to_add_22_port, A_to_add_21_port, 
      A_to_add_20_port, A_to_add_19_port, A_to_add_18_port, A_to_add_17_port, 
      A_to_add_16_port, A_to_add_15_port, A_to_add_14_port, A_to_add_13_port, 
      A_to_add_12_port, A_to_add_11_port, A_to_add_10_port, A_to_add_9_port, 
      A_to_add_8_port, A_to_add_7_port, A_to_add_6_port, A_to_add_5_port, 
      A_to_add_4_port, A_to_add_3_port, A_to_add_2_port, A_to_add_1_port, 
      A_to_add_0_port );
   
   X_Logic0_port <= '0';
   count_reg_0_inst : DFFS_X1 port map( D => N37, CK => net199343, SN => n18, Q
                           => count_0_port, QN => n13);
   count_reg_1_inst : DFFR_X1 port map( D => N39, CK => net199343, RN => n18, Q
                           => count_1_port, QN => n5);
   count_reg_2_inst : DFFR_X1 port map( D => N41, CK => net199343, RN => n18, Q
                           => count_2_port, QN => n14);
   count_reg_3_inst : DFFS_X1 port map( D => N43, CK => net199343, SN => n18, Q
                           => count_3_port, QN => n3);
   count_reg_4_inst : DFFR_X1 port map( D => N45, CK => net199343, RN => n18, Q
                           => count_4_port, QN => n2);
   U51 : MUX2_X1 port map( A => A_to_add_9_port, B => ACC_from_add(9), S => 
                           input_mux_sel_2_port, Z => final_out(9));
   U52 : MUX2_X1 port map( A => A_to_add_8_port, B => ACC_from_add(8), S => 
                           input_mux_sel_2_port, Z => final_out(8));
   U53 : MUX2_X1 port map( A => A_to_add_7_port, B => ACC_from_add(7), S => 
                           input_mux_sel_2_port, Z => final_out(7));
   U54 : MUX2_X1 port map( A => A_to_add_6_port, B => ACC_from_add(6), S => 
                           input_mux_sel_2_port, Z => final_out(6));
   U55 : MUX2_X1 port map( A => A_to_add_5_port, B => ACC_from_add(5), S => 
                           input_mux_sel_2_port, Z => final_out(5));
   U56 : MUX2_X1 port map( A => A_to_add_4_port, B => ACC_from_add(4), S => 
                           input_mux_sel_2_port, Z => final_out(4));
   U57 : MUX2_X1 port map( A => A_to_add_3_port, B => ACC_from_add(3), S => 
                           input_mux_sel_2_port, Z => final_out(3));
   U58 : MUX2_X1 port map( A => A_to_add_31_port, B => ACC_from_add(31), S => 
                           input_mux_sel_2_port, Z => final_out(31));
   U59 : MUX2_X1 port map( A => A_to_add_30_port, B => ACC_from_add(30), S => 
                           input_mux_sel_2_port, Z => final_out(30));
   U60 : MUX2_X1 port map( A => A_to_add_2_port, B => ACC_from_add(2), S => 
                           input_mux_sel_2_port, Z => final_out(2));
   U61 : MUX2_X1 port map( A => A_to_add_29_port, B => ACC_from_add(29), S => 
                           input_mux_sel_2_port, Z => final_out(29));
   U62 : MUX2_X1 port map( A => A_to_add_28_port, B => ACC_from_add(28), S => 
                           input_mux_sel_2_port, Z => final_out(28));
   U63 : MUX2_X1 port map( A => A_to_add_27_port, B => ACC_from_add(27), S => 
                           input_mux_sel_2_port, Z => final_out(27));
   U64 : MUX2_X1 port map( A => A_to_add_26_port, B => ACC_from_add(26), S => 
                           input_mux_sel_2_port, Z => final_out(26));
   U65 : MUX2_X1 port map( A => A_to_add_25_port, B => ACC_from_add(25), S => 
                           input_mux_sel_2_port, Z => final_out(25));
   U66 : MUX2_X1 port map( A => A_to_add_24_port, B => ACC_from_add(24), S => 
                           input_mux_sel_2_port, Z => final_out(24));
   U67 : MUX2_X1 port map( A => A_to_add_23_port, B => ACC_from_add(23), S => 
                           input_mux_sel_2_port, Z => final_out(23));
   U68 : MUX2_X1 port map( A => A_to_add_22_port, B => ACC_from_add(22), S => 
                           input_mux_sel_2_port, Z => final_out(22));
   U69 : MUX2_X1 port map( A => A_to_add_21_port, B => ACC_from_add(21), S => 
                           input_mux_sel_2_port, Z => final_out(21));
   U70 : MUX2_X1 port map( A => A_to_add_20_port, B => ACC_from_add(20), S => 
                           input_mux_sel_2_port, Z => final_out(20));
   U71 : MUX2_X1 port map( A => A_to_add_1_port, B => ACC_from_add(1), S => 
                           input_mux_sel_2_port, Z => final_out(1));
   U72 : MUX2_X1 port map( A => A_to_add_19_port, B => ACC_from_add(19), S => 
                           input_mux_sel_2_port, Z => final_out(19));
   U73 : MUX2_X1 port map( A => A_to_add_18_port, B => ACC_from_add(18), S => 
                           input_mux_sel_2_port, Z => final_out(18));
   U74 : MUX2_X1 port map( A => A_to_add_17_port, B => ACC_from_add(17), S => 
                           input_mux_sel_2_port, Z => final_out(17));
   U75 : MUX2_X1 port map( A => A_to_add_16_port, B => ACC_from_add(16), S => 
                           input_mux_sel_2_port, Z => final_out(16));
   U77 : MUX2_X1 port map( A => A_to_add_14_port, B => ACC_from_add(14), S => 
                           input_mux_sel_2_port, Z => final_out(14));
   U78 : MUX2_X1 port map( A => A_to_add_13_port, B => ACC_from_add(13), S => 
                           input_mux_sel_2_port, Z => final_out(13));
   U79 : MUX2_X1 port map( A => A_to_add_12_port, B => ACC_from_add(12), S => 
                           input_mux_sel_2_port, Z => final_out(12));
   U80 : MUX2_X1 port map( A => A_to_add_11_port, B => ACC_from_add(11), S => 
                           input_mux_sel_2_port, Z => final_out(11));
   U81 : MUX2_X1 port map( A => A_to_add_10_port, B => ACC_from_add(10), S => 
                           input_mux_sel_2_port, Z => final_out(10));
   encod_0_0 : booth_encoder_0 port map( B_in(2) => B(1), B_in(1) => B(0), 
                           B_in(0) => X_Logic0_port, A_out(2) => 
                           piso_2_in_0_port, A_out(1) => piso_1_in_0_port, 
                           A_out(0) => piso_0_in_0_port);
   encod_i_1 : booth_encoder_8 port map( B_in(2) => B(3), B_in(1) => B(2), 
                           B_in(0) => B(1), A_out(2) => piso_2_in_1_port, 
                           A_out(1) => piso_1_in_1_port, A_out(0) => 
                           piso_0_in_1_port);
   encod_i_2 : booth_encoder_7 port map( B_in(2) => B(5), B_in(1) => B(4), 
                           B_in(0) => B(3), A_out(2) => piso_2_in_2_port, 
                           A_out(1) => piso_1_in_2_port, A_out(0) => 
                           piso_0_in_2_port);
   encod_i_3 : booth_encoder_6 port map( B_in(2) => B(7), B_in(1) => B(6), 
                           B_in(0) => B(5), A_out(2) => piso_2_in_3_port, 
                           A_out(1) => piso_1_in_3_port, A_out(0) => 
                           piso_0_in_3_port);
   encod_i_4 : booth_encoder_5 port map( B_in(2) => B(9), B_in(1) => B(8), 
                           B_in(0) => B(7), A_out(2) => piso_2_in_4_port, 
                           A_out(1) => piso_1_in_4_port, A_out(0) => 
                           piso_0_in_4_port);
   encod_i_5 : booth_encoder_4 port map( B_in(2) => B(11), B_in(1) => B(10), 
                           B_in(0) => B(9), A_out(2) => piso_2_in_5_port, 
                           A_out(1) => piso_1_in_5_port, A_out(0) => 
                           piso_0_in_5_port);
   encod_i_6 : booth_encoder_3 port map( B_in(2) => B(13), B_in(1) => B(12), 
                           B_in(0) => B(11), A_out(2) => piso_2_in_6_port, 
                           A_out(1) => piso_1_in_6_port, A_out(0) => 
                           piso_0_in_6_port);
   encod_i_7 : booth_encoder_2 port map( B_in(2) => B(15), B_in(1) => B(14), 
                           B_in(0) => B(13), A_out(2) => piso_2_in_7_port, 
                           A_out(1) => piso_1_in_7_port, A_out(0) => 
                           piso_0_in_7_port);
   encod_i_8 : booth_encoder_1 port map( B_in(2) => enc_N2_in_2_port, B_in(1) 
                           => enc_N2_in_2_port, B_in(0) => B(15), A_out(2) => 
                           piso_2_in_8_port, A_out(1) => piso_1_in_8_port, 
                           A_out(0) => piso_0_in_8_port);
   piso_0 : shift_N9_0 port map( Clock => Clock, ALOAD => n17, D(8) => 
                           piso_0_in_8_port, D(7) => piso_0_in_7_port, D(6) => 
                           piso_0_in_6_port, D(5) => piso_0_in_5_port, D(4) => 
                           piso_0_in_4_port, D(3) => piso_0_in_3_port, D(2) => 
                           piso_0_in_2_port, D(1) => piso_0_in_1_port, D(0) => 
                           piso_0_in_0_port, SO => input_mux_sel_0);
   piso_1 : shift_N9_2 port map( Clock => Clock, ALOAD => n17, D(8) => 
                           piso_1_in_8_port, D(7) => piso_1_in_7_port, D(6) => 
                           piso_1_in_6_port, D(5) => piso_1_in_5_port, D(4) => 
                           piso_1_in_4_port, D(3) => piso_1_in_3_port, D(2) => 
                           piso_1_in_2_port, D(1) => piso_1_in_1_port, D(0) => 
                           piso_1_in_0_port, SO => sign_to_add);
   piso_2 : shift_N9_1 port map( Clock => Clock, ALOAD => n17, D(8) => 
                           piso_2_in_8_port, D(7) => piso_2_in_7_port, D(6) => 
                           piso_2_in_6_port, D(5) => piso_2_in_5_port, D(4) => 
                           piso_2_in_4_port, D(3) => piso_2_in_3_port, D(2) => 
                           piso_2_in_2_port, D(1) => piso_2_in_1_port, D(0) => 
                           piso_2_in_0_port, SO => input_mux_sel_2_port);
   A_reg : piso_r_2_N32 port map( Clock => Clock, ALOAD => n17, D(31) => 
                           extend_vector_15_port, D(30) => 
                           extend_vector_15_port, D(29) => 
                           extend_vector_15_port, D(28) => 
                           extend_vector_15_port, D(27) => 
                           extend_vector_15_port, D(26) => 
                           extend_vector_15_port, D(25) => 
                           extend_vector_15_port, D(24) => 
                           extend_vector_15_port, D(23) => 
                           extend_vector_15_port, D(22) => 
                           extend_vector_15_port, D(21) => 
                           extend_vector_15_port, D(20) => 
                           extend_vector_15_port, D(19) => 
                           extend_vector_15_port, D(18) => 
                           extend_vector_15_port, D(17) => 
                           extend_vector_15_port, D(16) => 
                           extend_vector_15_port, D(15) => A(15), D(14) => 
                           A(14), D(13) => A(13), D(12) => A(12), D(11) => 
                           A(11), D(10) => A(10), D(9) => A(9), D(8) => A(8), 
                           D(7) => A(7), D(6) => A(6), D(5) => A(5), D(4) => 
                           A(4), D(3) => A(3), D(2) => A(2), D(1) => A(1), D(0)
                           => A(0), SO(31) => A_to_mux_31_port, SO(30) => 
                           A_to_mux_30_port, SO(29) => A_to_mux_29_port, SO(28)
                           => A_to_mux_28_port, SO(27) => A_to_mux_27_port, 
                           SO(26) => A_to_mux_26_port, SO(25) => 
                           A_to_mux_25_port, SO(24) => A_to_mux_24_port, SO(23)
                           => A_to_mux_23_port, SO(22) => A_to_mux_22_port, 
                           SO(21) => A_to_mux_21_port, SO(20) => 
                           A_to_mux_20_port, SO(19) => A_to_mux_19_port, SO(18)
                           => A_to_mux_18_port, SO(17) => A_to_mux_17_port, 
                           SO(16) => A_to_mux_16_port, SO(15) => 
                           A_to_mux_15_port, SO(14) => A_to_mux_14_port, SO(13)
                           => A_to_mux_13_port, SO(12) => A_to_mux_12_port, 
                           SO(11) => A_to_mux_11_port, SO(10) => 
                           A_to_mux_10_port, SO(9) => A_to_mux_9_port, SO(8) =>
                           A_to_mux_8_port, SO(7) => A_to_mux_7_port, SO(6) => 
                           A_to_mux_6_port, SO(5) => A_to_mux_5_port, SO(4) => 
                           A_to_mux_4_port, SO(3) => A_to_mux_3_port, SO(2) => 
                           A_to_mux_2_port, SO(1) => A_to_mux_1_port, SO(0) => 
                           A_to_mux_0_port);
   INPUTMUX : mux21_1 port map( IN0(31) => A_to_mux_31_port, IN0(30) => 
                           A_to_mux_30_port, IN0(29) => A_to_mux_29_port, 
                           IN0(28) => A_to_mux_28_port, IN0(27) => 
                           A_to_mux_27_port, IN0(26) => A_to_mux_26_port, 
                           IN0(25) => A_to_mux_25_port, IN0(24) => 
                           A_to_mux_24_port, IN0(23) => A_to_mux_23_port, 
                           IN0(22) => A_to_mux_22_port, IN0(21) => 
                           A_to_mux_21_port, IN0(20) => A_to_mux_20_port, 
                           IN0(19) => A_to_mux_19_port, IN0(18) => 
                           A_to_mux_18_port, IN0(17) => A_to_mux_17_port, 
                           IN0(16) => A_to_mux_16_port, IN0(15) => 
                           A_to_mux_15_port, IN0(14) => A_to_mux_14_port, 
                           IN0(13) => A_to_mux_13_port, IN0(12) => 
                           A_to_mux_12_port, IN0(11) => A_to_mux_11_port, 
                           IN0(10) => A_to_mux_10_port, IN0(9) => 
                           A_to_mux_9_port, IN0(8) => A_to_mux_8_port, IN0(7) 
                           => A_to_mux_7_port, IN0(6) => A_to_mux_6_port, 
                           IN0(5) => A_to_mux_5_port, IN0(4) => A_to_mux_4_port
                           , IN0(3) => A_to_mux_3_port, IN0(2) => 
                           A_to_mux_2_port, IN0(1) => A_to_mux_1_port, IN0(0) 
                           => A_to_mux_0_port, IN1(31) => A_to_mux_30_port, 
                           IN1(30) => A_to_mux_29_port, IN1(29) => 
                           A_to_mux_28_port, IN1(28) => A_to_mux_27_port, 
                           IN1(27) => A_to_mux_26_port, IN1(26) => 
                           A_to_mux_25_port, IN1(25) => A_to_mux_24_port, 
                           IN1(24) => A_to_mux_23_port, IN1(23) => 
                           A_to_mux_22_port, IN1(22) => A_to_mux_21_port, 
                           IN1(21) => A_to_mux_20_port, IN1(20) => 
                           A_to_mux_19_port, IN1(19) => A_to_mux_18_port, 
                           IN1(18) => A_to_mux_17_port, IN1(17) => 
                           A_to_mux_16_port, IN1(16) => A_to_mux_15_port, 
                           IN1(15) => A_to_mux_14_port, IN1(14) => 
                           A_to_mux_13_port, IN1(13) => A_to_mux_12_port, 
                           IN1(12) => A_to_mux_11_port, IN1(11) => 
                           A_to_mux_10_port, IN1(10) => A_to_mux_9_port, IN1(9)
                           => A_to_mux_8_port, IN1(8) => A_to_mux_7_port, 
                           IN1(7) => A_to_mux_6_port, IN1(6) => A_to_mux_5_port
                           , IN1(5) => A_to_mux_4_port, IN1(4) => 
                           A_to_mux_3_port, IN1(3) => A_to_mux_2_port, IN1(2) 
                           => A_to_mux_1_port, IN1(1) => A_to_mux_0_port, 
                           IN1(0) => X_Logic0_port, CTRL => input_mux_sel_0, 
                           OUT1(31) => B_to_add(31), OUT1(30) => B_to_add(30), 
                           OUT1(29) => B_to_add(29), OUT1(28) => B_to_add(28), 
                           OUT1(27) => B_to_add(27), OUT1(26) => B_to_add(26), 
                           OUT1(25) => B_to_add(25), OUT1(24) => B_to_add(24), 
                           OUT1(23) => B_to_add(23), OUT1(22) => B_to_add(22), 
                           OUT1(21) => B_to_add(21), OUT1(20) => B_to_add(20), 
                           OUT1(19) => B_to_add(19), OUT1(18) => B_to_add(18), 
                           OUT1(17) => B_to_add(17), OUT1(16) => B_to_add(16), 
                           OUT1(15) => B_to_add(15), OUT1(14) => B_to_add(14), 
                           OUT1(13) => B_to_add(13), OUT1(12) => B_to_add(12), 
                           OUT1(11) => B_to_add(11), OUT1(10) => B_to_add(10), 
                           OUT1(9) => B_to_add(9), OUT1(8) => B_to_add(8), 
                           OUT1(7) => B_to_add(7), OUT1(6) => B_to_add(6), 
                           OUT1(5) => B_to_add(5), OUT1(4) => B_to_add(4), 
                           OUT1(3) => B_to_add(3), OUT1(2) => B_to_add(2), 
                           OUT1(1) => B_to_add(1), OUT1(0) => B_to_add(0));
   ACCUMULATOR : ff32_en_SIZE32_1 port map( D(31) => next_accumulate_31_port, 
                           D(30) => next_accumulate_30_port, D(29) => 
                           next_accumulate_29_port, D(28) => 
                           next_accumulate_28_port, D(27) => 
                           next_accumulate_27_port, D(26) => 
                           next_accumulate_26_port, D(25) => 
                           next_accumulate_25_port, D(24) => 
                           next_accumulate_24_port, D(23) => 
                           next_accumulate_23_port, D(22) => 
                           next_accumulate_22_port, D(21) => 
                           next_accumulate_21_port, D(20) => 
                           next_accumulate_20_port, D(19) => 
                           next_accumulate_19_port, D(18) => 
                           next_accumulate_18_port, D(17) => 
                           next_accumulate_17_port, D(16) => 
                           next_accumulate_16_port, D(15) => 
                           next_accumulate_15_port, D(14) => 
                           next_accumulate_14_port, D(13) => 
                           next_accumulate_13_port, D(12) => 
                           next_accumulate_12_port, D(11) => 
                           next_accumulate_11_port, D(10) => 
                           next_accumulate_10_port, D(9) => 
                           next_accumulate_9_port, D(8) => 
                           next_accumulate_8_port, D(7) => 
                           next_accumulate_7_port, D(6) => 
                           next_accumulate_6_port, D(5) => 
                           next_accumulate_5_port, D(4) => 
                           next_accumulate_4_port, D(3) => 
                           next_accumulate_3_port, D(2) => 
                           next_accumulate_2_port, D(1) => 
                           next_accumulate_1_port, D(0) => 
                           next_accumulate_0_port, en => reg_enable, clk => 
                           Clock, rst => Reset, Q(31) => A_to_add_31_port, 
                           Q(30) => A_to_add_30_port, Q(29) => A_to_add_29_port
                           , Q(28) => A_to_add_28_port, Q(27) => 
                           A_to_add_27_port, Q(26) => A_to_add_26_port, Q(25) 
                           => A_to_add_25_port, Q(24) => A_to_add_24_port, 
                           Q(23) => A_to_add_23_port, Q(22) => A_to_add_22_port
                           , Q(21) => A_to_add_21_port, Q(20) => 
                           A_to_add_20_port, Q(19) => A_to_add_19_port, Q(18) 
                           => A_to_add_18_port, Q(17) => A_to_add_17_port, 
                           Q(16) => A_to_add_16_port, Q(15) => A_to_add_15_port
                           , Q(14) => A_to_add_14_port, Q(13) => 
                           A_to_add_13_port, Q(12) => A_to_add_12_port, Q(11) 
                           => A_to_add_11_port, Q(10) => A_to_add_10_port, Q(9)
                           => A_to_add_9_port, Q(8) => A_to_add_8_port, Q(7) =>
                           A_to_add_7_port, Q(6) => A_to_add_6_port, Q(5) => 
                           A_to_add_5_port, Q(4) => A_to_add_4_port, Q(3) => 
                           A_to_add_3_port, Q(2) => A_to_add_2_port, Q(1) => 
                           A_to_add_1_port, Q(0) => A_to_add_0_port);
   clk_gate_count_reg : SNPS_CLOCK_GATE_HIGH_simple_booth_add_ext_N16 port map(
                           CLK => Clock, EN => N44, ENCLK => net199343);
   U41 : OR2_X1 port map( A1 => valid_port, A2 => enable, ZN => N44);
   U49 : NOR3_X1 port map( A1 => count_1_port, A2 => count_4_port, A3 => 
                           count_2_port, ZN => n9);
   U47 : NOR3_X1 port map( A1 => count_3_port, A2 => count_0_port, A3 => n11, 
                           ZN => valid_port);
   U48 : INV_X1 port map( A => n9, ZN => n11);
   U50 : NAND3_X2 port map( A1 => n9, A2 => count_3_port, A3 => count_0_port, 
                           ZN => n8);
   U46 : OR2_X1 port map( A1 => valid_port, A2 => n13, ZN => N37);
   U45 : INV_X1 port map( A => valid_port, ZN => n10);
   U4 : OR2_X1 port map( A1 => n17, A2 => input_mux_sel_2_port, ZN => 
                           reg_enable);
   U43 : AND2_X1 port map( A1 => N23, A2 => n10, ZN => N41);
   U38 : AND2_X1 port map( A1 => sign, A2 => A(15), ZN => extend_vector_15_port
                           );
   U36 : AND2_X1 port map( A1 => n8, A2 => ACC_from_add(0), ZN => 
                           next_accumulate_0_port);
   U35 : AND2_X1 port map( A1 => n8, A2 => ACC_from_add(10), ZN => 
                           next_accumulate_10_port);
   U34 : AND2_X1 port map( A1 => n8, A2 => ACC_from_add(11), ZN => 
                           next_accumulate_11_port);
   U33 : AND2_X1 port map( A1 => n8, A2 => ACC_from_add(12), ZN => 
                           next_accumulate_12_port);
   U3 : AND2_X1 port map( A1 => n8, A2 => ACC_from_add(21), ZN => 
                           next_accumulate_21_port);
   U5 : AND2_X1 port map( A1 => n8, A2 => ACC_from_add(28), ZN => 
                           next_accumulate_28_port);
   U6 : NOR2_X1 port map( A1 => count_3_port, A2 => n16, ZN => n1);
   U7 : OAI21_X1 port map( B1 => count_4_port, B2 => n1, A => n10, ZN => n4);
   U8 : AOI21_X1 port map( B1 => count_4_port, B2 => n1, A => n4, ZN => N45);
   U9 : AOI21_X1 port map( B1 => n16, B2 => count_3_port, A => valid_port, ZN 
                           => n6);
   U10 : OAI21_X1 port map( B1 => n16, B2 => count_3_port, A => n6, ZN => N43);
   U11 : MUX2_X1 port map( A => A_to_add_0_port, B => ACC_from_add(0), S => 
                           input_mux_sel_2_port, Z => final_out(0));
   U12 : MUX2_X1 port map( A => A_to_add_15_port, B => ACC_from_add(15), S => 
                           input_mux_sel_2_port, Z => final_out(15));
   U13 : INV_X1 port map( A => n10, ZN => n7);
   U14 : AOI21_X1 port map( B1 => count_1_port, B2 => count_0_port, A => n15, 
                           ZN => n12);
   U15 : NOR2_X1 port map( A1 => n12, A2 => n7, ZN => N39);
   U16 : INV_X1 port map( A => Reset, ZN => n18);
   U17 : AND2_X1 port map( A1 => n8, A2 => ACC_from_add(31), ZN => 
                           next_accumulate_31_port);
   U18 : AND2_X1 port map( A1 => n8, A2 => ACC_from_add(26), ZN => 
                           next_accumulate_26_port);
   U19 : AND2_X1 port map( A1 => n8, A2 => ACC_from_add(25), ZN => 
                           next_accumulate_25_port);
   U20 : AND2_X1 port map( A1 => n8, A2 => ACC_from_add(23), ZN => 
                           next_accumulate_23_port);
   U21 : AND2_X1 port map( A1 => n8, A2 => ACC_from_add(29), ZN => 
                           next_accumulate_29_port);
   U22 : AND2_X1 port map( A1 => n8, A2 => ACC_from_add(15), ZN => 
                           next_accumulate_15_port);
   U23 : AND2_X1 port map( A1 => n8, A2 => ACC_from_add(1), ZN => 
                           next_accumulate_1_port);
   U24 : AND2_X1 port map( A1 => n8, A2 => ACC_from_add(4), ZN => 
                           next_accumulate_4_port);
   U25 : AND2_X1 port map( A1 => n8, A2 => ACC_from_add(5), ZN => 
                           next_accumulate_5_port);
   U26 : AND2_X1 port map( A1 => n8, A2 => ACC_from_add(2), ZN => 
                           next_accumulate_2_port);
   U27 : AND2_X1 port map( A1 => n8, A2 => ACC_from_add(9), ZN => 
                           next_accumulate_9_port);
   U28 : AND2_X1 port map( A1 => n8, A2 => ACC_from_add(8), ZN => 
                           next_accumulate_8_port);
   U29 : AND2_X1 port map( A1 => n8, A2 => ACC_from_add(6), ZN => 
                           next_accumulate_6_port);
   U30 : AND2_X1 port map( A1 => n8, A2 => ACC_from_add(3), ZN => 
                           next_accumulate_3_port);
   U31 : AND2_X1 port map( A1 => n8, A2 => ACC_from_add(14), ZN => 
                           next_accumulate_14_port);
   U32 : AND2_X1 port map( A1 => n8, A2 => ACC_from_add(7), ZN => 
                           next_accumulate_7_port);
   U37 : AND2_X1 port map( A1 => n8, A2 => ACC_from_add(16), ZN => 
                           next_accumulate_16_port);
   U39 : AND2_X1 port map( A1 => n8, A2 => ACC_from_add(18), ZN => 
                           next_accumulate_18_port);
   U40 : AND2_X1 port map( A1 => n8, A2 => ACC_from_add(17), ZN => 
                           next_accumulate_17_port);
   U42 : AND2_X1 port map( A1 => n8, A2 => ACC_from_add(30), ZN => 
                           next_accumulate_30_port);
   U44 : AND2_X1 port map( A1 => n8, A2 => ACC_from_add(19), ZN => 
                           next_accumulate_19_port);
   U76 : AND2_X1 port map( A1 => n8, A2 => ACC_from_add(22), ZN => 
                           next_accumulate_22_port);
   U82 : AND2_X1 port map( A1 => n8, A2 => ACC_from_add(27), ZN => 
                           next_accumulate_27_port);
   U83 : INV_X4 port map( A => n8, ZN => n17);
   U84 : NOR2_X1 port map( A1 => count_0_port, A2 => count_1_port, ZN => n15);
   U85 : OR3_X1 port map( A1 => count_2_port, A2 => count_0_port, A3 => 
                           count_1_port, ZN => n16);
   U86 : OAI21_X1 port map( B1 => n15, B2 => n14, A => n16, ZN => N23);
   U87 : AND2_X1 port map( A1 => n8, A2 => ACC_from_add(13), ZN => 
                           next_accumulate_13_port);
   U88 : AND2_X1 port map( A1 => n8, A2 => ACC_from_add(24), ZN => 
                           next_accumulate_24_port);
   U89 : AND2_X1 port map( A1 => sign, A2 => B(15), ZN => enc_N2_in_2_port);
   U90 : AND2_X1 port map( A1 => n8, A2 => ACC_from_add(20), ZN => 
                           next_accumulate_20_port);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_ff32_en_SIZE13 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_ff32_en_SIZE13;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_ff32_en_SIZE13 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net199382 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net199382);
   main_gate : AND2_X1 port map( A1 => net199382, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_ff32_en_SIZE5_0 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_ff32_en_SIZE5_0;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_ff32_en_SIZE5_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net199367 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net199367);
   main_gate : AND2_X1 port map( A1 => net199367, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_ff32_en_SIZE32_0 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_ff32_en_SIZE32_0;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_ff32_en_SIZE32_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net199352 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net199352);
   main_gate : AND2_X1 port map( A1 => net199352, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity sum_gen_N32_0 is

   port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic_vector 
         (8 downto 0);  S : out std_logic_vector (31 downto 0));

end sum_gen_N32_0;

architecture SYN_STRUCTURAL of sum_gen_N32_0 is

   component carry_sel_gen_N4_9
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component carry_sel_gen_N4_10
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component carry_sel_gen_N4_11
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component carry_sel_gen_N4_12
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component carry_sel_gen_N4_13
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component carry_sel_gen_N4_14
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component carry_sel_gen_N4_15
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component carry_sel_gen_N4_0
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal n5, net199157, net199158, net199159, net199160, net199161, net199162,
      net199163, net199164 : std_logic;

begin
   
   csel_N_0 : carry_sel_gen_N4_0 port map( A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), Ci => n5, S(3) => S(3), S(2) 
                           => S(2), S(1) => S(1), S(0) => S(0), Co => net199164
                           );
   csel_N_1 : carry_sel_gen_N4_15 port map( A(3) => A(7), A(2) => A(6), A(1) =>
                           A(5), A(0) => A(4), B(3) => B(7), B(2) => B(6), B(1)
                           => B(5), B(0) => B(4), Ci => Cin(1), S(3) => S(7), 
                           S(2) => S(6), S(1) => S(5), S(0) => S(4), Co => 
                           net199163);
   csel_N_2 : carry_sel_gen_N4_14 port map( A(3) => A(11), A(2) => A(10), A(1) 
                           => A(9), A(0) => A(8), B(3) => B(11), B(2) => B(10),
                           B(1) => B(9), B(0) => B(8), Ci => Cin(2), S(3) => 
                           S(11), S(2) => S(10), S(1) => S(9), S(0) => S(8), Co
                           => net199162);
   csel_N_3 : carry_sel_gen_N4_13 port map( A(3) => A(15), A(2) => A(14), A(1) 
                           => A(13), A(0) => A(12), B(3) => B(15), B(2) => 
                           B(14), B(1) => B(13), B(0) => B(12), Ci => Cin(3), 
                           S(3) => S(15), S(2) => S(14), S(1) => S(13), S(0) =>
                           S(12), Co => net199161);
   csel_N_4 : carry_sel_gen_N4_12 port map( A(3) => A(19), A(2) => A(18), A(1) 
                           => A(17), A(0) => A(16), B(3) => B(19), B(2) => 
                           B(18), B(1) => B(17), B(0) => B(16), Ci => Cin(4), 
                           S(3) => S(19), S(2) => S(18), S(1) => S(17), S(0) =>
                           S(16), Co => net199160);
   csel_N_5 : carry_sel_gen_N4_11 port map( A(3) => A(23), A(2) => A(22), A(1) 
                           => A(21), A(0) => A(20), B(3) => B(23), B(2) => 
                           B(22), B(1) => B(21), B(0) => B(20), Ci => Cin(5), 
                           S(3) => S(23), S(2) => S(22), S(1) => S(21), S(0) =>
                           S(20), Co => net199159);
   csel_N_6 : carry_sel_gen_N4_10 port map( A(3) => A(27), A(2) => A(26), A(1) 
                           => A(25), A(0) => A(24), B(3) => B(27), B(2) => 
                           B(26), B(1) => B(25), B(0) => B(24), Ci => Cin(6), 
                           S(3) => S(27), S(2) => S(26), S(1) => S(25), S(0) =>
                           S(24), Co => net199158);
   csel_N_7 : carry_sel_gen_N4_9 port map( A(3) => A(31), A(2) => A(30), A(1) 
                           => A(29), A(0) => A(28), B(3) => B(31), B(2) => 
                           B(30), B(1) => B(29), B(0) => B(28), Ci => Cin(7), 
                           S(3) => S(31), S(2) => S(30), S(1) => S(29), S(0) =>
                           S(28), Co => net199157);
   n5 <= '0';

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity carry_tree_N32_logN5_0 is

   port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  Cout :
         out std_logic_vector (7 downto 0));

end carry_tree_N32_logN5_0;

architecture SYN_arch of carry_tree_N32_logN5_0 is

   component pg_29
      port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic
            );
   end component;
   
   component pg_31
      port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic
            );
   end component;
   
   component pg_32
      port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic
            );
   end component;
   
   component g_12
      port( g, p, g_prec : in std_logic;  g_out : out std_logic);
   end component;
   
   component g_13
      port( g, p, g_prec : in std_logic;  g_out : out std_logic);
   end component;
   
   component g_14
      port( g, p, g_prec : in std_logic;  g_out : out std_logic);
   end component;
   
   component g_15
      port( g, p, g_prec : in std_logic;  g_out : out std_logic);
   end component;
   
   component g_16
      port( g, p, g_prec : in std_logic;  g_out : out std_logic);
   end component;
   
   component g_17
      port( g, p, g_prec : in std_logic;  g_out : out std_logic);
   end component;
   
   component pg_34
      port( p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic;  
            g_BAR : in std_logic);
   end component;
   
   component pg_35
      port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic
            );
   end component;
   
   component pg_36
      port( p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic;  
            g_BAR : in std_logic);
   end component;
   
   component pg_37
      port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic
            );
   end component;
   
   component pg_38
      port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic
            );
   end component;
   
   component pg_39
      port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic
            );
   end component;
   
   component g_18
      port( g, p, g_prec : in std_logic;  g_out : out std_logic);
   end component;
   
   component pg_42
      port( g, p, g_prec, p_prec : in std_logic;  p_out, g_out_BAR : out 
            std_logic);
   end component;
   
   component pg_43
      port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic
            );
   end component;
   
   component pg_44
      port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic
            );
   end component;
   
   component pg_45
      port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic
            );
   end component;
   
   component pg_46
      port( g, p, g_prec, p_prec : in std_logic;  p_out, g_out_BAR : out 
            std_logic);
   end component;
   
   component pg_47
      port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic
            );
   end component;
   
   component pg_48
      port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic
            );
   end component;
   
   component pg_49
      port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic
            );
   end component;
   
   component pg_50
      port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic
            );
   end component;
   
   component pg_51
      port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic
            );
   end component;
   
   component pg_52
      port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic
            );
   end component;
   
   component pg_53
      port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic
            );
   end component;
   
   component pg_0
      port( g, p, g_prec, p_prec : in std_logic;  g_out, p_out : out std_logic
            );
   end component;
   
   component g_19
      port( g, p, g_prec : in std_logic;  g_out : out std_logic);
   end component;
   
   component g_0
      port( g, p, g_prec : in std_logic;  g_out : out std_logic);
   end component;
   
   component pg_net_33
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_38
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_39
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_40
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_41
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_42
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_43
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_44
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_45
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_46
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_47
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_48
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_49
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_50
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_51
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_52
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_53
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_54
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_55
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_56
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_57
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_58
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_59
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_60
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_61
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_62
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_63
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   component pg_net_0
      port( a, b : in std_logic;  g_out, p_out : out std_logic);
   end component;
   
   signal n3, Cout_6_port, Cout_5_port, Cout_4_port, Cout_3_port, Cout_2_port, 
      Cout_1_port, Cout_0_port, p_net_27_port, p_net_26_port, p_net_25_port, 
      p_net_24_port, p_net_23_port, p_net_22_port, p_net_21_port, p_net_20_port
      , p_net_19_port, p_net_18_port, p_net_17_port, p_net_16_port, 
      p_net_15_port, p_net_14_port, p_net_13_port, p_net_12_port, p_net_11_port
      , p_net_10_port, p_net_9_port, p_net_8_port, p_net_7_port, p_net_6_port, 
      p_net_5_port, p_net_4_port, p_net_3_port, p_net_2_port, p_net_1_port, 
      g_net_27_port, g_net_26_port, g_net_25_port, g_net_24_port, g_net_23_port
      , g_net_22_port, g_net_21_port, g_net_20_port, g_net_19_port, 
      g_net_18_port, g_net_17_port, g_net_16_port, g_net_15_port, g_net_14_port
      , g_net_13_port, g_net_12_port, g_net_11_port, g_net_10_port, 
      g_net_9_port, g_net_8_port, g_net_7_port, g_net_6_port, g_net_5_port, 
      g_net_4_port, g_net_3_port, g_net_2_port, g_net_1_port, g_net_0_port, 
      magic_pro_0_port, pg_1_13_1_port, pg_1_13_0_port, pg_1_12_1_port, 
      pg_1_12_0_port, pg_1_11_1_port, pg_1_11_0_port, pg_1_10_1_port, 
      pg_1_10_0_port, pg_1_9_1_port, pg_1_9_0_port, pg_1_8_1_port, 
      pg_1_8_0_port, pg_1_7_1_port, pg_1_7_0_port, pg_1_6_1_port, pg_1_6_0_port
      , pg_1_5_1_port, pg_1_5_0_port, pg_1_4_1_port, pg_1_4_0_port, 
      pg_1_3_1_port, pg_1_3_0_port, pg_1_2_1_port, pg_1_2_0_port, pg_1_1_1_port
      , pg_1_1_0_port, pg_1_0_0_port, pg_n_4_6_1_port, pg_n_4_6_0_port, 
      pg_n_3_5_1_port, pg_n_3_5_0_port, pg_n_3_3_1_port, pg_n_3_3_0_port, 
      pg_n_2_6_1_port, pg_n_2_6_0_port, pg_n_2_5_1_port, pg_n_2_5_0_port, 
      pg_n_2_4_1_port, pg_n_2_4_0_port, pg_n_2_3_1_port, pg_n_2_3_0_port, 
      pg_n_2_2_1_port, pg_n_2_2_0_port, pg_n_2_1_1_port, pg_n_2_1_0_port, n2, 
      net246125, n_1169 : std_logic;

begin
   Cout <= ( n_1169, Cout_6_port, Cout_5_port, Cout_4_port, Cout_3_port, 
      Cout_2_port, Cout_1_port, Cout_0_port );
   
   pg_net_x_1 : pg_net_0 port map( a => A(1), b => B(1), g_out => g_net_1_port,
                           p_out => p_net_1_port);
   pg_net_x_2 : pg_net_63 port map( a => A(2), b => B(2), g_out => g_net_2_port
                           , p_out => p_net_2_port);
   pg_net_x_3 : pg_net_62 port map( a => A(3), b => B(3), g_out => g_net_3_port
                           , p_out => p_net_3_port);
   pg_net_x_4 : pg_net_61 port map( a => A(4), b => B(4), g_out => g_net_4_port
                           , p_out => p_net_4_port);
   pg_net_x_5 : pg_net_60 port map( a => A(5), b => B(5), g_out => g_net_5_port
                           , p_out => p_net_5_port);
   pg_net_x_6 : pg_net_59 port map( a => A(6), b => B(6), g_out => g_net_6_port
                           , p_out => p_net_6_port);
   pg_net_x_7 : pg_net_58 port map( a => A(7), b => B(7), g_out => g_net_7_port
                           , p_out => p_net_7_port);
   pg_net_x_8 : pg_net_57 port map( a => A(8), b => B(8), g_out => g_net_8_port
                           , p_out => p_net_8_port);
   pg_net_x_9 : pg_net_56 port map( a => A(9), b => B(9), g_out => g_net_9_port
                           , p_out => p_net_9_port);
   pg_net_x_10 : pg_net_55 port map( a => A(10), b => B(10), g_out => 
                           g_net_10_port, p_out => p_net_10_port);
   pg_net_x_11 : pg_net_54 port map( a => A(11), b => B(11), g_out => 
                           g_net_11_port, p_out => p_net_11_port);
   pg_net_x_12 : pg_net_53 port map( a => A(12), b => B(12), g_out => 
                           g_net_12_port, p_out => p_net_12_port);
   pg_net_x_13 : pg_net_52 port map( a => A(13), b => B(13), g_out => 
                           g_net_13_port, p_out => p_net_13_port);
   pg_net_x_14 : pg_net_51 port map( a => A(14), b => B(14), g_out => 
                           g_net_14_port, p_out => p_net_14_port);
   pg_net_x_15 : pg_net_50 port map( a => A(15), b => B(15), g_out => 
                           g_net_15_port, p_out => p_net_15_port);
   pg_net_x_16 : pg_net_49 port map( a => A(16), b => B(16), g_out => 
                           g_net_16_port, p_out => p_net_16_port);
   pg_net_x_17 : pg_net_48 port map( a => A(17), b => B(17), g_out => 
                           g_net_17_port, p_out => p_net_17_port);
   pg_net_x_18 : pg_net_47 port map( a => A(18), b => B(18), g_out => 
                           g_net_18_port, p_out => p_net_18_port);
   pg_net_x_19 : pg_net_46 port map( a => A(19), b => B(19), g_out => 
                           g_net_19_port, p_out => p_net_19_port);
   pg_net_x_20 : pg_net_45 port map( a => A(20), b => B(20), g_out => 
                           g_net_20_port, p_out => p_net_20_port);
   pg_net_x_21 : pg_net_44 port map( a => A(21), b => B(21), g_out => 
                           g_net_21_port, p_out => p_net_21_port);
   pg_net_x_22 : pg_net_43 port map( a => A(22), b => B(22), g_out => 
                           g_net_22_port, p_out => p_net_22_port);
   pg_net_x_23 : pg_net_42 port map( a => A(23), b => B(23), g_out => 
                           g_net_23_port, p_out => p_net_23_port);
   pg_net_x_24 : pg_net_41 port map( a => A(24), b => B(24), g_out => 
                           g_net_24_port, p_out => p_net_24_port);
   pg_net_x_25 : pg_net_40 port map( a => A(25), b => B(25), g_out => 
                           g_net_25_port, p_out => p_net_25_port);
   pg_net_x_26 : pg_net_39 port map( a => A(26), b => B(26), g_out => 
                           g_net_26_port, p_out => p_net_26_port);
   pg_net_x_27 : pg_net_38 port map( a => A(27), b => B(27), g_out => 
                           g_net_27_port, p_out => p_net_27_port);
   pg_net_0_MAGIC : pg_net_33 port map( a => A(0), b => B(0), g_out => 
                           magic_pro_0_port, p_out => net246125);
   xG_0_0_MAGIC : g_0 port map( g => magic_pro_0_port, p => n2, g_prec => n3, 
                           g_out => g_net_0_port);
   xG_1_0 : g_19 port map( g => g_net_1_port, p => p_net_1_port, g_prec => 
                           g_net_0_port, g_out => pg_1_0_0_port);
   xPG_1_1 : pg_0 port map( g => g_net_3_port, p => p_net_3_port, g_prec => 
                           g_net_2_port, p_prec => p_net_2_port, g_out => 
                           pg_1_1_0_port, p_out => pg_1_1_1_port);
   xPG_1_2 : pg_53 port map( g => g_net_5_port, p => p_net_5_port, g_prec => 
                           g_net_4_port, p_prec => p_net_4_port, g_out => 
                           pg_1_2_0_port, p_out => pg_1_2_1_port);
   xPG_1_3 : pg_52 port map( g => g_net_7_port, p => p_net_7_port, g_prec => 
                           g_net_6_port, p_prec => p_net_6_port, g_out => 
                           pg_1_3_0_port, p_out => pg_1_3_1_port);
   xPG_1_4 : pg_51 port map( g => g_net_9_port, p => p_net_9_port, g_prec => 
                           g_net_8_port, p_prec => p_net_8_port, g_out => 
                           pg_1_4_0_port, p_out => pg_1_4_1_port);
   xPG_1_5 : pg_50 port map( g => g_net_11_port, p => p_net_11_port, g_prec => 
                           g_net_10_port, p_prec => p_net_10_port, g_out => 
                           pg_1_5_0_port, p_out => pg_1_5_1_port);
   xPG_1_6 : pg_49 port map( g => g_net_13_port, p => p_net_13_port, g_prec => 
                           g_net_12_port, p_prec => p_net_12_port, g_out => 
                           pg_1_6_0_port, p_out => pg_1_6_1_port);
   xPG_1_7 : pg_48 port map( g => g_net_15_port, p => p_net_15_port, g_prec => 
                           g_net_14_port, p_prec => p_net_14_port, g_out => 
                           pg_1_7_0_port, p_out => pg_1_7_1_port);
   xPG_1_8 : pg_47 port map( g => g_net_17_port, p => p_net_17_port, g_prec => 
                           g_net_16_port, p_prec => p_net_16_port, g_out => 
                           pg_1_8_0_port, p_out => pg_1_8_1_port);
   xPG_1_9 : pg_46 port map( g => g_net_19_port, p => p_net_19_port, g_prec => 
                           g_net_18_port, p_prec => p_net_18_port, p_out => 
                           pg_1_9_1_port, g_out_BAR => pg_1_9_0_port);
   xPG_1_10 : pg_45 port map( g => g_net_21_port, p => p_net_21_port, g_prec =>
                           g_net_20_port, p_prec => p_net_20_port, g_out => 
                           pg_1_10_0_port, p_out => pg_1_10_1_port);
   xPG_1_11 : pg_44 port map( g => g_net_23_port, p => p_net_23_port, g_prec =>
                           g_net_22_port, p_prec => p_net_22_port, g_out => 
                           pg_1_11_0_port, p_out => pg_1_11_1_port);
   xPG_1_12 : pg_43 port map( g => g_net_25_port, p => p_net_25_port, g_prec =>
                           g_net_24_port, p_prec => p_net_24_port, g_out => 
                           pg_1_12_0_port, p_out => pg_1_12_1_port);
   xPG_1_13 : pg_42 port map( g => g_net_27_port, p => p_net_27_port, g_prec =>
                           g_net_26_port, p_prec => p_net_26_port, p_out => 
                           pg_1_13_1_port, g_out_BAR => pg_1_13_0_port);
   xG_2_0 : g_18 port map( g => pg_1_1_0_port, p => pg_1_1_1_port, g_prec => 
                           pg_1_0_0_port, g_out => Cout_0_port);
   xPG_2_1 : pg_39 port map( g => pg_1_3_0_port, p => pg_1_3_1_port, g_prec => 
                           pg_1_2_0_port, p_prec => pg_1_2_1_port, g_out => 
                           pg_n_2_1_0_port, p_out => pg_n_2_1_1_port);
   xPG_2_2 : pg_38 port map( g => pg_1_5_0_port, p => pg_1_5_1_port, g_prec => 
                           pg_1_4_0_port, p_prec => pg_1_4_1_port, g_out => 
                           pg_n_2_2_0_port, p_out => pg_n_2_2_1_port);
   xPG_2_3 : pg_37 port map( g => pg_1_7_0_port, p => pg_1_7_1_port, g_prec => 
                           pg_1_6_0_port, p_prec => pg_1_6_1_port, g_out => 
                           pg_n_2_3_0_port, p_out => pg_n_2_3_1_port);
   xPG_2_4 : pg_36 port map( p => pg_1_9_1_port, g_prec => pg_1_8_0_port, 
                           p_prec => pg_1_8_1_port, g_out => pg_n_2_4_0_port, 
                           p_out => pg_n_2_4_1_port, g_BAR => pg_1_9_0_port);
   xPG_2_5 : pg_35 port map( g => pg_1_11_0_port, p => pg_1_11_1_port, g_prec 
                           => pg_1_10_0_port, p_prec => pg_1_10_1_port, g_out 
                           => pg_n_2_5_0_port, p_out => pg_n_2_5_1_port);
   xPG_2_6 : pg_34 port map( p => pg_1_13_1_port, g_prec => pg_1_12_0_port, 
                           p_prec => pg_1_12_1_port, g_out => pg_n_2_6_0_port, 
                           p_out => pg_n_2_6_1_port, g_BAR => pg_1_13_0_port);
   xG_3_1 : g_17 port map( g => pg_n_2_1_0_port, p => pg_n_2_1_1_port, g_prec 
                           => Cout_0_port, g_out => Cout_1_port);
   xG_4_2 : g_16 port map( g => pg_n_2_2_0_port, p => pg_n_2_2_1_port, g_prec 
                           => Cout_1_port, g_out => Cout_2_port);
   xG_4_3 : g_15 port map( g => pg_n_3_3_0_port, p => pg_n_3_3_1_port, g_prec 
                           => Cout_1_port, g_out => Cout_3_port);
   xG_5_4 : g_14 port map( g => pg_n_2_4_0_port, p => pg_n_2_4_1_port, g_prec 
                           => Cout_3_port, g_out => Cout_4_port);
   xG_5_5 : g_13 port map( g => pg_n_3_5_0_port, p => pg_n_3_5_1_port, g_prec 
                           => Cout_3_port, g_out => Cout_5_port);
   xG_5_6 : g_12 port map( g => pg_n_4_6_0_port, p => pg_n_4_6_1_port, g_prec 
                           => Cout_3_port, g_out => Cout_6_port);
   xPG_3_3 : pg_32 port map( g => pg_n_2_3_0_port, p => pg_n_2_3_1_port, g_prec
                           => pg_n_2_2_0_port, p_prec => pg_n_2_2_1_port, g_out
                           => pg_n_3_3_0_port, p_out => pg_n_3_3_1_port);
   xPG_3_5 : pg_31 port map( g => pg_n_2_5_0_port, p => pg_n_2_5_1_port, g_prec
                           => pg_n_2_4_0_port, p_prec => pg_n_2_4_1_port, g_out
                           => pg_n_3_5_0_port, p_out => pg_n_3_5_1_port);
   xPG_4_6 : pg_29 port map( g => pg_n_2_6_0_port, p => pg_n_2_6_1_port, g_prec
                           => pg_n_3_5_0_port, p_prec => pg_n_3_5_1_port, g_out
                           => pg_n_4_6_0_port, p_out => pg_n_4_6_1_port);
   n2 <= '0';
   n3 <= '0';

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity xor_gen_N32_0 is

   port( A : in std_logic_vector (31 downto 0);  B : in std_logic;  S : out 
         std_logic_vector (31 downto 0));

end xor_gen_N32_0;

architecture SYN_bhe of xor_gen_N32_0 is

begin
   S <= ( A(31), A(30), A(29), A(28), A(27), A(26), A(25), A(24), A(23), A(22),
      A(21), A(20), A(19), A(18), A(17), A(16), A(15), A(14), A(13), A(12), 
      A(11), A(10), A(9), A(8), A(7), A(6), A(5), A(4), A(3), A(2), A(1), A(0) 
      );

end SYN_bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_ff32_en_IR is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_ff32_en_IR;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_ff32_en_IR is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net199597 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net199597);
   main_gate : AND2_X1 port map( A1 => net199597, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_ff32_en_0 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_ff32_en_0;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_ff32_en_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net199612 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net199612);
   main_gate : AND2_X1 port map( A1 => net199612, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity ff32_SIZE5 is

   port( D : in std_logic_vector (4 downto 0);  clk, rst : in std_logic;  Q : 
         out std_logic_vector (4 downto 0));

end ff32_SIZE5;

architecture SYN_behavioral of ff32_SIZE5 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n6, n5 : std_logic;

begin
   
   Q_reg_4_inst : DFFR_X1 port map( D => D(4), CK => clk, RN => n5, Q => Q(4), 
                           QN => n6);
   Q_reg_3_inst : DFFR_X1 port map( D => D(3), CK => clk, RN => n5, Q => Q(3), 
                           QN => n4);
   Q_reg_2_inst : DFFR_X1 port map( D => D(2), CK => clk, RN => n5, Q => Q(2), 
                           QN => n3);
   Q_reg_1_inst : DFFR_X1 port map( D => D(1), CK => clk, RN => n5, Q => Q(1), 
                           QN => n2);
   Q_reg_0_inst : DFFR_X1 port map( D => D(0), CK => clk, RN => n5, Q => Q(0), 
                           QN => n1);
   U3 : INV_X1 port map( A => rst, ZN => n5);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity ff32_SIZE32 is

   port( D : in std_logic_vector (31 downto 0);  clk, rst : in std_logic;  Q : 
         out std_logic_vector (31 downto 0));

end ff32_SIZE32;

architecture SYN_behavioral of ff32_SIZE32 is

   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n33, n32 : std_logic;

begin
   
   Q_reg_31_inst : DFFR_X1 port map( D => D(31), CK => clk, RN => n32, Q => 
                           Q(31), QN => n33);
   Q_reg_30_inst : DFFR_X1 port map( D => D(30), CK => clk, RN => n32, Q => 
                           Q(30), QN => n31);
   Q_reg_29_inst : DFFR_X1 port map( D => D(29), CK => clk, RN => n32, Q => 
                           Q(29), QN => n30);
   Q_reg_28_inst : DFFR_X1 port map( D => D(28), CK => clk, RN => n32, Q => 
                           Q(28), QN => n29);
   Q_reg_27_inst : DFFR_X1 port map( D => D(27), CK => clk, RN => n32, Q => 
                           Q(27), QN => n28);
   Q_reg_26_inst : DFFR_X1 port map( D => D(26), CK => clk, RN => n32, Q => 
                           Q(26), QN => n27);
   Q_reg_25_inst : DFFR_X1 port map( D => D(25), CK => clk, RN => n32, Q => 
                           Q(25), QN => n26);
   Q_reg_24_inst : DFFR_X1 port map( D => D(24), CK => clk, RN => n32, Q => 
                           Q(24), QN => n25);
   Q_reg_23_inst : DFFR_X1 port map( D => D(23), CK => clk, RN => n32, Q => 
                           Q(23), QN => n24);
   Q_reg_22_inst : DFFR_X1 port map( D => D(22), CK => clk, RN => n32, Q => 
                           Q(22), QN => n23);
   Q_reg_21_inst : DFFR_X1 port map( D => D(21), CK => clk, RN => n32, Q => 
                           Q(21), QN => n22);
   Q_reg_20_inst : DFFR_X1 port map( D => D(20), CK => clk, RN => n32, Q => 
                           Q(20), QN => n21);
   Q_reg_19_inst : DFFR_X1 port map( D => D(19), CK => clk, RN => n32, Q => 
                           Q(19), QN => n20);
   Q_reg_18_inst : DFFR_X1 port map( D => D(18), CK => clk, RN => n32, Q => 
                           Q(18), QN => n19);
   Q_reg_17_inst : DFFR_X1 port map( D => D(17), CK => clk, RN => n32, Q => 
                           Q(17), QN => n18);
   Q_reg_16_inst : DFFR_X1 port map( D => D(16), CK => clk, RN => n32, Q => 
                           Q(16), QN => n17);
   Q_reg_15_inst : DFFR_X1 port map( D => D(15), CK => clk, RN => n32, Q => 
                           Q(15), QN => n16);
   Q_reg_14_inst : DFFR_X1 port map( D => D(14), CK => clk, RN => n32, Q => 
                           Q(14), QN => n15);
   Q_reg_13_inst : DFFR_X1 port map( D => D(13), CK => clk, RN => n32, Q => 
                           Q(13), QN => n14);
   Q_reg_12_inst : DFFR_X1 port map( D => D(12), CK => clk, RN => n32, Q => 
                           Q(12), QN => n13);
   Q_reg_11_inst : DFFR_X1 port map( D => D(11), CK => clk, RN => n32, Q => 
                           Q(11), QN => n12);
   Q_reg_10_inst : DFFR_X1 port map( D => D(10), CK => clk, RN => n32, Q => 
                           Q(10), QN => n11);
   Q_reg_9_inst : DFFR_X1 port map( D => D(9), CK => clk, RN => n32, Q => Q(9),
                           QN => n10);
   Q_reg_8_inst : DFFR_X1 port map( D => D(8), CK => clk, RN => n32, Q => Q(8),
                           QN => n9);
   Q_reg_7_inst : DFFR_X1 port map( D => D(7), CK => clk, RN => n32, Q => Q(7),
                           QN => n8);
   Q_reg_6_inst : DFFR_X1 port map( D => D(6), CK => clk, RN => n32, Q => Q(6),
                           QN => n7);
   Q_reg_5_inst : DFFR_X1 port map( D => D(5), CK => clk, RN => n32, Q => Q(5),
                           QN => n6);
   Q_reg_4_inst : DFFR_X1 port map( D => D(4), CK => clk, RN => n32, Q => Q(4),
                           QN => n5);
   Q_reg_3_inst : DFFR_X1 port map( D => D(3), CK => clk, RN => n32, Q => Q(3),
                           QN => n4);
   Q_reg_2_inst : DFFR_X1 port map( D => D(2), CK => clk, RN => n32, Q => Q(2),
                           QN => n3);
   Q_reg_1_inst : DFFR_X1 port map( D => D(1), CK => clk, RN => n32, Q => Q(1),
                           QN => n2);
   Q_reg_0_inst : DFFR_X1 port map( D => D(0), CK => clk, RN => n32, Q => Q(0),
                           QN => n1);
   U3 : INV_X2 port map( A => rst, ZN => n32);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity mux41_MUX_SIZE5 is

   port( IN0, IN1, IN2, IN3 : in std_logic_vector (4 downto 0);  CTRL : in 
         std_logic_vector (1 downto 0);  OUT1 : out std_logic_vector (4 downto 
         0));

end mux41_MUX_SIZE5;

architecture SYN_bhe of mux41_MUX_SIZE5 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7, n9, n10, n11, n12, n13, n14, n15, n16, n17 : 
      std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n3, A2 => n4, ZN => OUT1(4));
   U17 : AOI22_X1 port map( A1 => n6, A2 => IN2(0), B1 => n7, B2 => IN1(0), ZN 
                           => n15);
   U13 : NAND2_X1 port map( A1 => n15, A2 => n16, ZN => OUT1(0));
   U20 : INV_X1 port map( A => CTRL(1), ZN => n17);
   U16 : AND2_X1 port map( A1 => CTRL(0), A2 => CTRL(1), ZN => n5);
   U19 : NOR2_X1 port map( A1 => CTRL(0), A2 => n17, ZN => n6);
   U18 : AND2_X1 port map( A1 => n17, A2 => CTRL(0), ZN => n7);
   U2 : INV_X1 port map( A => n5, ZN => n16);
   U3 : NAND2_X1 port map( A1 => n13, A2 => n14, ZN => OUT1(1));
   U4 : AOI21_X1 port map( B1 => n6, B2 => IN2(1), A => n5, ZN => n14);
   U5 : NAND2_X1 port map( A1 => n7, A2 => IN1(1), ZN => n13);
   U6 : AOI21_X1 port map( B1 => n6, B2 => IN2(2), A => n5, ZN => n12);
   U7 : NAND2_X1 port map( A1 => n7, A2 => IN1(2), ZN => n11);
   U8 : AOI21_X1 port map( B1 => n6, B2 => IN2(3), A => n5, ZN => n10);
   U9 : NAND2_X1 port map( A1 => n7, A2 => IN1(3), ZN => n9);
   U10 : AOI21_X1 port map( B1 => n6, B2 => IN2(4), A => n5, ZN => n4);
   U11 : NAND2_X1 port map( A1 => n7, A2 => IN1(4), ZN => n3);
   U12 : NAND2_X1 port map( A1 => n9, A2 => n10, ZN => OUT1(3));
   U14 : NAND2_X1 port map( A1 => n11, A2 => n12, ZN => OUT1(2));

end SYN_bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity real_alu_DATA_SIZE32 is

   port( IN1, IN2 : in std_logic_vector (31 downto 0);  ALUW_i : in 
         std_logic_vector (12 downto 0);  DOUT : out std_logic_vector (31 
         downto 0);  stall_o : out std_logic;  Clock, Reset : in std_logic);

end real_alu_DATA_SIZE32;

architecture SYN_Bhe of real_alu_DATA_SIZE32 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X4
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X2
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component logic_unit_SIZE32
      port( IN1, IN2 : in std_logic_vector (31 downto 0);  CTRL : in 
            std_logic_vector (1 downto 0);  OUT1 : out std_logic_vector (31 
            downto 0));
   end component;
   
   component shifter
      port( A : in std_logic_vector (31 downto 0);  B : in std_logic_vector (4 
            downto 0);  LOGIC_ARITH, LEFT_RIGHT : in std_logic;  OUTPUT : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component comparator_M32
      port( C, V : in std_logic;  SUM : in std_logic_vector (31 downto 0);  sel
            : in std_logic_vector (2 downto 0);  sign : in std_logic;  S : out 
            std_logic);
   end component;
   
   component p4add_N32_logN5_1
      port( A, B : in std_logic_vector (31 downto 0);  Cin, sign : in std_logic
            ;  S : out std_logic_vector (31 downto 0);  Cout : out std_logic);
   end component;
   
   component simple_booth_add_ext_N16
      port( Clock, Reset, sign, enable : in std_logic;  valid : out std_logic; 
            A, B : in std_logic_vector (15 downto 0);  A_to_add, B_to_add : out
            std_logic_vector (31 downto 0);  sign_to_add : out std_logic;  
            final_out : out std_logic_vector (31 downto 0);  ACC_from_add : in 
            std_logic_vector (31 downto 0));
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal X_Logic0_port, mux_A_31_port, mux_A_30_port, mux_A_29_port, 
      mux_A_28_port, mux_A_27_port, mux_A_26_port, mux_A_25_port, mux_A_24_port
      , mux_A_23_port, mux_A_22_port, mux_A_21_port, mux_A_20_port, 
      mux_A_19_port, mux_A_18_port, mux_A_17_port, mux_A_16_port, mux_A_15_port
      , mux_A_14_port, mux_A_13_port, mux_A_12_port, mux_A_11_port, 
      mux_A_10_port, mux_A_9_port, mux_A_8_port, mux_A_7_port, mux_A_6_port, 
      mux_A_5_port, mux_A_4_port, mux_A_3_port, mux_A_2_port, mux_A_1_port, 
      mux_A_0_port, A_booth_to_add_31_port, A_booth_to_add_30_port, 
      A_booth_to_add_29_port, A_booth_to_add_28_port, A_booth_to_add_27_port, 
      A_booth_to_add_26_port, A_booth_to_add_25_port, A_booth_to_add_24_port, 
      A_booth_to_add_23_port, A_booth_to_add_22_port, A_booth_to_add_21_port, 
      A_booth_to_add_20_port, A_booth_to_add_19_port, A_booth_to_add_18_port, 
      A_booth_to_add_17_port, A_booth_to_add_16_port, A_booth_to_add_15_port, 
      A_booth_to_add_14_port, A_booth_to_add_13_port, A_booth_to_add_12_port, 
      A_booth_to_add_11_port, A_booth_to_add_10_port, A_booth_to_add_9_port, 
      A_booth_to_add_8_port, A_booth_to_add_7_port, A_booth_to_add_6_port, 
      A_booth_to_add_5_port, A_booth_to_add_4_port, A_booth_to_add_3_port, 
      A_booth_to_add_2_port, A_booth_to_add_1_port, A_booth_to_add_0_port, 
      mux_B_31_port, mux_B_30_port, mux_B_29_port, mux_B_28_port, mux_B_27_port
      , mux_B_26_port, mux_B_25_port, mux_B_24_port, mux_B_23_port, 
      mux_B_22_port, mux_B_21_port, mux_B_20_port, mux_B_19_port, mux_B_18_port
      , mux_B_17_port, mux_B_16_port, mux_B_15_port, mux_B_14_port, 
      mux_B_13_port, mux_B_12_port, mux_B_11_port, mux_B_10_port, mux_B_9_port,
      mux_B_8_port, mux_B_7_port, mux_B_6_port, mux_B_5_port, mux_B_4_port, 
      mux_B_3_port, mux_B_2_port, mux_B_1_port, mux_B_0_port, 
      B_booth_to_add_31_port, B_booth_to_add_30_port, B_booth_to_add_29_port, 
      B_booth_to_add_28_port, B_booth_to_add_27_port, B_booth_to_add_26_port, 
      B_booth_to_add_25_port, B_booth_to_add_24_port, B_booth_to_add_23_port, 
      B_booth_to_add_22_port, B_booth_to_add_21_port, B_booth_to_add_20_port, 
      B_booth_to_add_19_port, B_booth_to_add_18_port, B_booth_to_add_17_port, 
      B_booth_to_add_16_port, B_booth_to_add_15_port, B_booth_to_add_14_port, 
      B_booth_to_add_13_port, B_booth_to_add_12_port, B_booth_to_add_11_port, 
      B_booth_to_add_10_port, B_booth_to_add_9_port, B_booth_to_add_8_port, 
      B_booth_to_add_7_port, B_booth_to_add_6_port, B_booth_to_add_5_port, 
      B_booth_to_add_4_port, B_booth_to_add_3_port, B_booth_to_add_2_port, 
      B_booth_to_add_1_port, B_booth_to_add_0_port, mux_sign, sign_booth_to_add
      , valid_from_booth, mult_out_31_port, mult_out_30_port, mult_out_29_port,
      mult_out_28_port, mult_out_27_port, mult_out_26_port, mult_out_25_port, 
      mult_out_24_port, mult_out_23_port, mult_out_22_port, mult_out_21_port, 
      mult_out_20_port, mult_out_19_port, mult_out_18_port, mult_out_17_port, 
      mult_out_16_port, mult_out_15_port, mult_out_14_port, mult_out_13_port, 
      mult_out_12_port, mult_out_11_port, mult_out_10_port, mult_out_9_port, 
      mult_out_8_port, mult_out_7_port, mult_out_6_port, mult_out_5_port, 
      mult_out_4_port, mult_out_3_port, mult_out_2_port, mult_out_1_port, 
      mult_out_0_port, sum_out_31_port, sum_out_30_port, sum_out_29_port, 
      sum_out_28_port, sum_out_27_port, sum_out_26_port, sum_out_25_port, 
      sum_out_24_port, sum_out_23_port, sum_out_22_port, sum_out_21_port, 
      sum_out_20_port, sum_out_19_port, sum_out_18_port, sum_out_17_port, 
      sum_out_16_port, sum_out_15_port, sum_out_14_port, sum_out_13_port, 
      sum_out_12_port, sum_out_11_port, sum_out_10_port, sum_out_9_port, 
      sum_out_8_port, sum_out_7_port, sum_out_6_port, sum_out_5_port, 
      sum_out_4_port, sum_out_3_port, sum_out_2_port, sum_out_1_port, 
      sum_out_0_port, carry_from_adder, overflow, comp_out, shift_out_31_port, 
      shift_out_30_port, shift_out_29_port, shift_out_28_port, 
      shift_out_27_port, shift_out_26_port, shift_out_25_port, 
      shift_out_24_port, shift_out_23_port, shift_out_22_port, 
      shift_out_21_port, shift_out_20_port, shift_out_19_port, 
      shift_out_18_port, shift_out_17_port, shift_out_16_port, 
      shift_out_15_port, shift_out_14_port, shift_out_13_port, 
      shift_out_12_port, shift_out_11_port, shift_out_10_port, shift_out_9_port
      , shift_out_8_port, shift_out_7_port, shift_out_6_port, shift_out_5_port,
      shift_out_4_port, shift_out_3_port, shift_out_2_port, shift_out_1_port, 
      shift_out_0_port, lu_out_31_port, lu_out_30_port, lu_out_29_port, 
      lu_out_28_port, lu_out_27_port, lu_out_26_port, lu_out_25_port, 
      lu_out_24_port, lu_out_23_port, lu_out_22_port, lu_out_21_port, 
      lu_out_20_port, lu_out_19_port, lu_out_18_port, lu_out_17_port, 
      lu_out_16_port, lu_out_15_port, lu_out_14_port, lu_out_13_port, 
      lu_out_12_port, lu_out_11_port, lu_out_10_port, lu_out_9_port, 
      lu_out_8_port, lu_out_7_port, lu_out_6_port, lu_out_5_port, lu_out_4_port
      , lu_out_3_port, lu_out_2_port, lu_out_1_port, lu_out_0_port, n9, n13, 
      n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28
      , n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, 
      n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57
      , n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n71, n72, n73, 
      n74, n75, n76, n77, n78, n79, n80, n84, n85, n1, n2, n3, n4, n5, n6, n7, 
      n8, n10, n11, n12, n69, n70, n81, n82, n83, n86, n87, n88, n89, n90, n91,
      n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, 
      n105, n106 : std_logic;

begin
   
   X_Logic0_port <= '0';
   U113 : MUX2_X1 port map( A => B_booth_to_add_9_port, B => IN2(9), S => n9, Z
                           => mux_B_9_port);
   U116 : MUX2_X1 port map( A => B_booth_to_add_6_port, B => IN2(6), S => n9, Z
                           => mux_B_6_port);
   U120 : MUX2_X1 port map( A => B_booth_to_add_31_port, B => IN2(31), S => n9,
                           Z => mux_B_31_port);
   U121 : MUX2_X1 port map( A => B_booth_to_add_30_port, B => IN2(30), S => n9,
                           Z => mux_B_30_port);
   U123 : MUX2_X1 port map( A => B_booth_to_add_29_port, B => IN2(29), S => n9,
                           Z => mux_B_29_port);
   U124 : MUX2_X1 port map( A => B_booth_to_add_28_port, B => IN2(28), S => n9,
                           Z => mux_B_28_port);
   U125 : MUX2_X1 port map( A => B_booth_to_add_27_port, B => IN2(27), S => 
                           n106, Z => mux_B_27_port);
   U126 : MUX2_X1 port map( A => B_booth_to_add_26_port, B => IN2(26), S => 
                           n106, Z => mux_B_26_port);
   U127 : MUX2_X1 port map( A => B_booth_to_add_25_port, B => IN2(25), S => 
                           n106, Z => mux_B_25_port);
   U128 : MUX2_X1 port map( A => B_booth_to_add_24_port, B => IN2(24), S => 
                           n106, Z => mux_B_24_port);
   U129 : MUX2_X1 port map( A => B_booth_to_add_23_port, B => IN2(23), S => 
                           n106, Z => mux_B_23_port);
   U130 : MUX2_X1 port map( A => B_booth_to_add_22_port, B => IN2(22), S => 
                           n106, Z => mux_B_22_port);
   U132 : MUX2_X1 port map( A => B_booth_to_add_20_port, B => IN2(20), S => 
                           n106, Z => mux_B_20_port);
   U134 : MUX2_X1 port map( A => B_booth_to_add_19_port, B => IN2(19), S => 
                           n106, Z => mux_B_19_port);
   U135 : MUX2_X1 port map( A => B_booth_to_add_18_port, B => IN2(18), S => 
                           n106, Z => mux_B_18_port);
   U136 : MUX2_X1 port map( A => B_booth_to_add_17_port, B => IN2(17), S => 
                           n106, Z => mux_B_17_port);
   U137 : MUX2_X1 port map( A => B_booth_to_add_16_port, B => IN2(16), S => 
                           n106, Z => mux_B_16_port);
   U138 : MUX2_X1 port map( A => B_booth_to_add_15_port, B => IN2(15), S => 
                           n106, Z => mux_B_15_port);
   U139 : MUX2_X1 port map( A => B_booth_to_add_14_port, B => IN2(14), S => 
                           n106, Z => mux_B_14_port);
   U141 : MUX2_X1 port map( A => B_booth_to_add_12_port, B => IN2(12), S => 
                           n106, Z => mux_B_12_port);
   U142 : MUX2_X1 port map( A => B_booth_to_add_11_port, B => IN2(11), S => 
                           n106, Z => mux_B_11_port);
   U145 : MUX2_X1 port map( A => A_booth_to_add_9_port, B => IN1(9), S => n9, Z
                           => mux_A_9_port);
   U146 : MUX2_X1 port map( A => A_booth_to_add_8_port, B => IN1(8), S => n9, Z
                           => mux_A_8_port);
   U147 : MUX2_X1 port map( A => A_booth_to_add_7_port, B => IN1(7), S => n9, Z
                           => mux_A_7_port);
   U148 : MUX2_X1 port map( A => A_booth_to_add_6_port, B => IN1(6), S => n9, Z
                           => mux_A_6_port);
   U149 : MUX2_X1 port map( A => A_booth_to_add_5_port, B => IN1(5), S => n9, Z
                           => mux_A_5_port);
   U150 : MUX2_X1 port map( A => A_booth_to_add_4_port, B => IN1(4), S => n9, Z
                           => mux_A_4_port);
   U151 : MUX2_X1 port map( A => A_booth_to_add_3_port, B => IN1(3), S => n9, Z
                           => mux_A_3_port);
   U152 : MUX2_X1 port map( A => A_booth_to_add_31_port, B => IN1(31), S => n9,
                           Z => mux_A_31_port);
   U153 : MUX2_X1 port map( A => A_booth_to_add_30_port, B => IN1(30), S => n9,
                           Z => mux_A_30_port);
   U154 : MUX2_X1 port map( A => A_booth_to_add_2_port, B => IN1(2), S => n9, Z
                           => mux_A_2_port);
   U155 : MUX2_X1 port map( A => A_booth_to_add_29_port, B => IN1(29), S => n9,
                           Z => mux_A_29_port);
   U156 : MUX2_X1 port map( A => A_booth_to_add_28_port, B => IN1(28), S => n9,
                           Z => mux_A_28_port);
   U157 : MUX2_X1 port map( A => A_booth_to_add_27_port, B => IN1(27), S => n9,
                           Z => mux_A_27_port);
   U158 : MUX2_X1 port map( A => A_booth_to_add_26_port, B => IN1(26), S => n9,
                           Z => mux_A_26_port);
   U159 : MUX2_X1 port map( A => A_booth_to_add_25_port, B => IN1(25), S => n9,
                           Z => mux_A_25_port);
   U160 : MUX2_X1 port map( A => A_booth_to_add_24_port, B => IN1(24), S => n9,
                           Z => mux_A_24_port);
   U161 : MUX2_X1 port map( A => A_booth_to_add_23_port, B => IN1(23), S => n9,
                           Z => mux_A_23_port);
   U162 : MUX2_X1 port map( A => A_booth_to_add_22_port, B => IN1(22), S => n9,
                           Z => mux_A_22_port);
   U163 : MUX2_X1 port map( A => A_booth_to_add_21_port, B => IN1(21), S => n9,
                           Z => mux_A_21_port);
   U164 : MUX2_X1 port map( A => A_booth_to_add_20_port, B => IN1(20), S => n9,
                           Z => mux_A_20_port);
   U165 : MUX2_X1 port map( A => A_booth_to_add_1_port, B => IN1(1), S => n9, Z
                           => mux_A_1_port);
   U166 : MUX2_X1 port map( A => A_booth_to_add_19_port, B => IN1(19), S => n9,
                           Z => mux_A_19_port);
   U167 : MUX2_X1 port map( A => A_booth_to_add_18_port, B => IN1(18), S => n9,
                           Z => mux_A_18_port);
   U168 : MUX2_X1 port map( A => A_booth_to_add_17_port, B => IN1(17), S => n9,
                           Z => mux_A_17_port);
   U169 : MUX2_X1 port map( A => A_booth_to_add_16_port, B => IN1(16), S => n9,
                           Z => mux_A_16_port);
   U170 : MUX2_X1 port map( A => A_booth_to_add_15_port, B => IN1(15), S => n9,
                           Z => mux_A_15_port);
   U171 : MUX2_X1 port map( A => A_booth_to_add_14_port, B => IN1(14), S => n9,
                           Z => mux_A_14_port);
   U172 : MUX2_X1 port map( A => A_booth_to_add_13_port, B => IN1(13), S => n9,
                           Z => mux_A_13_port);
   U173 : MUX2_X1 port map( A => A_booth_to_add_12_port, B => IN1(12), S => n9,
                           Z => mux_A_12_port);
   U174 : MUX2_X1 port map( A => A_booth_to_add_11_port, B => IN1(11), S => n9,
                           Z => mux_A_11_port);
   U175 : MUX2_X1 port map( A => A_booth_to_add_10_port, B => IN1(10), S => n9,
                           Z => mux_A_10_port);
   U178 : NAND3_X1 port map( A1 => n84, A2 => n85, A3 => ALUW_i(12), ZN => n32)
                           ;
   MULT : simple_booth_add_ext_N16 port map( Clock => Clock, Reset => Reset, 
                           sign => ALUW_i(0), enable => ALUW_i(1), valid => 
                           valid_from_booth, A(15) => IN1(15), A(14) => IN1(14)
                           , A(13) => IN1(13), A(12) => IN1(12), A(11) => 
                           IN1(11), A(10) => IN1(10), A(9) => IN1(9), A(8) => 
                           IN1(8), A(7) => IN1(7), A(6) => IN1(6), A(5) => 
                           IN1(5), A(4) => IN1(4), A(3) => IN1(3), A(2) => 
                           IN1(2), A(1) => IN1(1), A(0) => IN1(0), B(15) => 
                           IN2(15), B(14) => IN2(14), B(13) => IN2(13), B(12) 
                           => IN2(12), B(11) => IN2(11), B(10) => IN2(10), B(9)
                           => IN2(9), B(8) => IN2(8), B(7) => n100, B(6) => 
                           IN2(6), B(5) => n98, B(4) => IN2(4), B(3) => n103, 
                           B(2) => IN2(2), B(1) => n101, B(0) => n102, 
                           A_to_add(31) => A_booth_to_add_31_port, A_to_add(30)
                           => A_booth_to_add_30_port, A_to_add(29) => 
                           A_booth_to_add_29_port, A_to_add(28) => 
                           A_booth_to_add_28_port, A_to_add(27) => 
                           A_booth_to_add_27_port, A_to_add(26) => 
                           A_booth_to_add_26_port, A_to_add(25) => 
                           A_booth_to_add_25_port, A_to_add(24) => 
                           A_booth_to_add_24_port, A_to_add(23) => 
                           A_booth_to_add_23_port, A_to_add(22) => 
                           A_booth_to_add_22_port, A_to_add(21) => 
                           A_booth_to_add_21_port, A_to_add(20) => 
                           A_booth_to_add_20_port, A_to_add(19) => 
                           A_booth_to_add_19_port, A_to_add(18) => 
                           A_booth_to_add_18_port, A_to_add(17) => 
                           A_booth_to_add_17_port, A_to_add(16) => 
                           A_booth_to_add_16_port, A_to_add(15) => 
                           A_booth_to_add_15_port, A_to_add(14) => 
                           A_booth_to_add_14_port, A_to_add(13) => 
                           A_booth_to_add_13_port, A_to_add(12) => 
                           A_booth_to_add_12_port, A_to_add(11) => 
                           A_booth_to_add_11_port, A_to_add(10) => 
                           A_booth_to_add_10_port, A_to_add(9) => 
                           A_booth_to_add_9_port, A_to_add(8) => 
                           A_booth_to_add_8_port, A_to_add(7) => 
                           A_booth_to_add_7_port, A_to_add(6) => 
                           A_booth_to_add_6_port, A_to_add(5) => 
                           A_booth_to_add_5_port, A_to_add(4) => 
                           A_booth_to_add_4_port, A_to_add(3) => 
                           A_booth_to_add_3_port, A_to_add(2) => 
                           A_booth_to_add_2_port, A_to_add(1) => 
                           A_booth_to_add_1_port, A_to_add(0) => 
                           A_booth_to_add_0_port, B_to_add(31) => 
                           B_booth_to_add_31_port, B_to_add(30) => 
                           B_booth_to_add_30_port, B_to_add(29) => 
                           B_booth_to_add_29_port, B_to_add(28) => 
                           B_booth_to_add_28_port, B_to_add(27) => 
                           B_booth_to_add_27_port, B_to_add(26) => 
                           B_booth_to_add_26_port, B_to_add(25) => 
                           B_booth_to_add_25_port, B_to_add(24) => 
                           B_booth_to_add_24_port, B_to_add(23) => 
                           B_booth_to_add_23_port, B_to_add(22) => 
                           B_booth_to_add_22_port, B_to_add(21) => 
                           B_booth_to_add_21_port, B_to_add(20) => 
                           B_booth_to_add_20_port, B_to_add(19) => 
                           B_booth_to_add_19_port, B_to_add(18) => 
                           B_booth_to_add_18_port, B_to_add(17) => 
                           B_booth_to_add_17_port, B_to_add(16) => 
                           B_booth_to_add_16_port, B_to_add(15) => 
                           B_booth_to_add_15_port, B_to_add(14) => 
                           B_booth_to_add_14_port, B_to_add(13) => 
                           B_booth_to_add_13_port, B_to_add(12) => 
                           B_booth_to_add_12_port, B_to_add(11) => 
                           B_booth_to_add_11_port, B_to_add(10) => 
                           B_booth_to_add_10_port, B_to_add(9) => 
                           B_booth_to_add_9_port, B_to_add(8) => 
                           B_booth_to_add_8_port, B_to_add(7) => 
                           B_booth_to_add_7_port, B_to_add(6) => 
                           B_booth_to_add_6_port, B_to_add(5) => 
                           B_booth_to_add_5_port, B_to_add(4) => 
                           B_booth_to_add_4_port, B_to_add(3) => 
                           B_booth_to_add_3_port, B_to_add(2) => 
                           B_booth_to_add_2_port, B_to_add(1) => 
                           B_booth_to_add_1_port, B_to_add(0) => 
                           B_booth_to_add_0_port, sign_to_add => 
                           sign_booth_to_add, final_out(31) => mult_out_31_port
                           , final_out(30) => mult_out_30_port, final_out(29) 
                           => mult_out_29_port, final_out(28) => 
                           mult_out_28_port, final_out(27) => mult_out_27_port,
                           final_out(26) => mult_out_26_port, final_out(25) => 
                           mult_out_25_port, final_out(24) => mult_out_24_port,
                           final_out(23) => mult_out_23_port, final_out(22) => 
                           mult_out_22_port, final_out(21) => mult_out_21_port,
                           final_out(20) => mult_out_20_port, final_out(19) => 
                           mult_out_19_port, final_out(18) => mult_out_18_port,
                           final_out(17) => mult_out_17_port, final_out(16) => 
                           mult_out_16_port, final_out(15) => mult_out_15_port,
                           final_out(14) => mult_out_14_port, final_out(13) => 
                           mult_out_13_port, final_out(12) => mult_out_12_port,
                           final_out(11) => mult_out_11_port, final_out(10) => 
                           mult_out_10_port, final_out(9) => mult_out_9_port, 
                           final_out(8) => mult_out_8_port, final_out(7) => 
                           mult_out_7_port, final_out(6) => mult_out_6_port, 
                           final_out(5) => mult_out_5_port, final_out(4) => 
                           mult_out_4_port, final_out(3) => mult_out_3_port, 
                           final_out(2) => mult_out_2_port, final_out(1) => 
                           mult_out_1_port, final_out(0) => mult_out_0_port, 
                           ACC_from_add(31) => n99, ACC_from_add(30) => 
                           sum_out_30_port, ACC_from_add(29) => sum_out_29_port
                           , ACC_from_add(28) => sum_out_28_port, 
                           ACC_from_add(27) => sum_out_27_port, 
                           ACC_from_add(26) => sum_out_26_port, 
                           ACC_from_add(25) => sum_out_25_port, 
                           ACC_from_add(24) => sum_out_24_port, 
                           ACC_from_add(23) => sum_out_23_port, 
                           ACC_from_add(22) => sum_out_22_port, 
                           ACC_from_add(21) => sum_out_21_port, 
                           ACC_from_add(20) => sum_out_20_port, 
                           ACC_from_add(19) => sum_out_19_port, 
                           ACC_from_add(18) => sum_out_18_port, 
                           ACC_from_add(17) => sum_out_17_port, 
                           ACC_from_add(16) => sum_out_16_port, 
                           ACC_from_add(15) => sum_out_15_port, 
                           ACC_from_add(14) => sum_out_14_port, 
                           ACC_from_add(13) => sum_out_13_port, 
                           ACC_from_add(12) => sum_out_12_port, 
                           ACC_from_add(11) => sum_out_11_port, 
                           ACC_from_add(10) => sum_out_10_port, ACC_from_add(9)
                           => sum_out_9_port, ACC_from_add(8) => sum_out_8_port
                           , ACC_from_add(7) => sum_out_7_port, ACC_from_add(6)
                           => sum_out_6_port, ACC_from_add(5) => sum_out_5_port
                           , ACC_from_add(4) => sum_out_4_port, ACC_from_add(3)
                           => sum_out_3_port, ACC_from_add(2) => sum_out_2_port
                           , ACC_from_add(1) => sum_out_1_port, ACC_from_add(0)
                           => sum_out_0_port);
   ADDER : p4add_N32_logN5_1 port map( A(31) => mux_A_31_port, A(30) => 
                           mux_A_30_port, A(29) => mux_A_29_port, A(28) => 
                           mux_A_28_port, A(27) => mux_A_27_port, A(26) => 
                           mux_A_26_port, A(25) => mux_A_25_port, A(24) => 
                           mux_A_24_port, A(23) => mux_A_23_port, A(22) => 
                           mux_A_22_port, A(21) => mux_A_21_port, A(20) => 
                           mux_A_20_port, A(19) => mux_A_19_port, A(18) => 
                           mux_A_18_port, A(17) => mux_A_17_port, A(16) => 
                           mux_A_16_port, A(15) => mux_A_15_port, A(14) => 
                           mux_A_14_port, A(13) => mux_A_13_port, A(12) => 
                           mux_A_12_port, A(11) => mux_A_11_port, A(10) => 
                           mux_A_10_port, A(9) => mux_A_9_port, A(8) => 
                           mux_A_8_port, A(7) => mux_A_7_port, A(6) => 
                           mux_A_6_port, A(5) => mux_A_5_port, A(4) => 
                           mux_A_4_port, A(3) => mux_A_3_port, A(2) => 
                           mux_A_2_port, A(1) => mux_A_1_port, A(0) => 
                           mux_A_0_port, B(31) => mux_B_31_port, B(30) => 
                           mux_B_30_port, B(29) => mux_B_29_port, B(28) => 
                           mux_B_28_port, B(27) => mux_B_27_port, B(26) => 
                           mux_B_26_port, B(25) => mux_B_25_port, B(24) => 
                           mux_B_24_port, B(23) => mux_B_23_port, B(22) => 
                           mux_B_22_port, B(21) => mux_B_21_port, B(20) => 
                           mux_B_20_port, B(19) => mux_B_19_port, B(18) => 
                           mux_B_18_port, B(17) => mux_B_17_port, B(16) => 
                           mux_B_16_port, B(15) => mux_B_15_port, B(14) => 
                           mux_B_14_port, B(13) => mux_B_13_port, B(12) => 
                           mux_B_12_port, B(11) => mux_B_11_port, B(10) => 
                           mux_B_10_port, B(9) => mux_B_9_port, B(8) => 
                           mux_B_8_port, B(7) => mux_B_7_port, B(6) => 
                           mux_B_6_port, B(5) => mux_B_5_port, B(4) => 
                           mux_B_4_port, B(3) => mux_B_3_port, B(2) => 
                           mux_B_2_port, B(1) => mux_B_1_port, B(0) => 
                           mux_B_0_port, Cin => X_Logic0_port, sign => mux_sign
                           , S(31) => sum_out_31_port, S(30) => sum_out_30_port
                           , S(29) => sum_out_29_port, S(28) => sum_out_28_port
                           , S(27) => sum_out_27_port, S(26) => sum_out_26_port
                           , S(25) => sum_out_25_port, S(24) => sum_out_24_port
                           , S(23) => sum_out_23_port, S(22) => sum_out_22_port
                           , S(21) => sum_out_21_port, S(20) => sum_out_20_port
                           , S(19) => sum_out_19_port, S(18) => sum_out_18_port
                           , S(17) => sum_out_17_port, S(16) => sum_out_16_port
                           , S(15) => sum_out_15_port, S(14) => sum_out_14_port
                           , S(13) => sum_out_13_port, S(12) => sum_out_12_port
                           , S(11) => sum_out_11_port, S(10) => sum_out_10_port
                           , S(9) => sum_out_9_port, S(8) => sum_out_8_port, 
                           S(7) => sum_out_7_port, S(6) => sum_out_6_port, S(5)
                           => sum_out_5_port, S(4) => sum_out_4_port, S(3) => 
                           sum_out_3_port, S(2) => sum_out_2_port, S(1) => 
                           sum_out_1_port, S(0) => sum_out_0_port, Cout => 
                           carry_from_adder);
   COMP : comparator_M32 port map( C => carry_from_adder, V => overflow, 
                           SUM(31) => sum_out_31_port, SUM(30) => 
                           sum_out_30_port, SUM(29) => sum_out_29_port, SUM(28)
                           => sum_out_28_port, SUM(27) => sum_out_27_port, 
                           SUM(26) => sum_out_26_port, SUM(25) => 
                           sum_out_25_port, SUM(24) => sum_out_24_port, SUM(23)
                           => sum_out_23_port, SUM(22) => sum_out_22_port, 
                           SUM(21) => sum_out_21_port, SUM(20) => 
                           sum_out_20_port, SUM(19) => sum_out_19_port, SUM(18)
                           => sum_out_18_port, SUM(17) => sum_out_17_port, 
                           SUM(16) => sum_out_16_port, SUM(15) => 
                           sum_out_15_port, SUM(14) => sum_out_14_port, SUM(13)
                           => sum_out_13_port, SUM(12) => sum_out_12_port, 
                           SUM(11) => sum_out_11_port, SUM(10) => 
                           sum_out_10_port, SUM(9) => sum_out_9_port, SUM(8) =>
                           sum_out_8_port, SUM(7) => sum_out_7_port, SUM(6) => 
                           sum_out_6_port, SUM(5) => sum_out_5_port, SUM(4) => 
                           sum_out_4_port, SUM(3) => sum_out_3_port, SUM(2) => 
                           sum_out_2_port, SUM(1) => sum_out_1_port, SUM(0) => 
                           sum_out_0_port, sel(2) => ALUW_i(4), sel(1) => 
                           ALUW_i(3), sel(0) => ALUW_i(2), sign => ALUW_i(0), S
                           => comp_out);
   SHIFT : shifter port map( A(31) => IN1(31), A(30) => IN1(30), A(29) => 
                           IN1(29), A(28) => IN1(28), A(27) => IN1(27), A(26) 
                           => IN1(26), A(25) => IN1(25), A(24) => IN1(24), 
                           A(23) => IN1(23), A(22) => IN1(22), A(21) => IN1(21)
                           , A(20) => IN1(20), A(19) => IN1(19), A(18) => 
                           IN1(18), A(17) => IN1(17), A(16) => IN1(16), A(15) 
                           => IN1(15), A(14) => IN1(14), A(13) => IN1(13), 
                           A(12) => IN1(12), A(11) => IN1(11), A(10) => IN1(10)
                           , A(9) => IN1(9), A(8) => IN1(8), A(7) => IN1(7), 
                           A(6) => IN1(6), A(5) => IN1(5), A(4) => IN1(4), A(3)
                           => IN1(3), A(2) => IN1(2), A(1) => IN1(1), A(0) => 
                           IN1(0), B(4) => IN2(4), B(3) => n103, B(2) => IN2(2)
                           , B(1) => n101, B(0) => n102, LOGIC_ARITH => 
                           ALUW_i(8), LEFT_RIGHT => ALUW_i(9), OUTPUT(31) => 
                           shift_out_31_port, OUTPUT(30) => shift_out_30_port, 
                           OUTPUT(29) => shift_out_29_port, OUTPUT(28) => 
                           shift_out_28_port, OUTPUT(27) => shift_out_27_port, 
                           OUTPUT(26) => shift_out_26_port, OUTPUT(25) => 
                           shift_out_25_port, OUTPUT(24) => shift_out_24_port, 
                           OUTPUT(23) => shift_out_23_port, OUTPUT(22) => 
                           shift_out_22_port, OUTPUT(21) => shift_out_21_port, 
                           OUTPUT(20) => shift_out_20_port, OUTPUT(19) => 
                           shift_out_19_port, OUTPUT(18) => shift_out_18_port, 
                           OUTPUT(17) => shift_out_17_port, OUTPUT(16) => 
                           shift_out_16_port, OUTPUT(15) => shift_out_15_port, 
                           OUTPUT(14) => shift_out_14_port, OUTPUT(13) => 
                           shift_out_13_port, OUTPUT(12) => shift_out_12_port, 
                           OUTPUT(11) => shift_out_11_port, OUTPUT(10) => 
                           shift_out_10_port, OUTPUT(9) => shift_out_9_port, 
                           OUTPUT(8) => shift_out_8_port, OUTPUT(7) => 
                           shift_out_7_port, OUTPUT(6) => shift_out_6_port, 
                           OUTPUT(5) => shift_out_5_port, OUTPUT(4) => 
                           shift_out_4_port, OUTPUT(3) => shift_out_3_port, 
                           OUTPUT(2) => shift_out_2_port, OUTPUT(1) => 
                           shift_out_1_port, OUTPUT(0) => shift_out_0_port);
   LU : logic_unit_SIZE32 port map( IN1(31) => IN1(31), IN1(30) => IN1(30), 
                           IN1(29) => IN1(29), IN1(28) => IN1(28), IN1(27) => 
                           IN1(27), IN1(26) => IN1(26), IN1(25) => IN1(25), 
                           IN1(24) => IN1(24), IN1(23) => IN1(23), IN1(22) => 
                           IN1(22), IN1(21) => IN1(21), IN1(20) => IN1(20), 
                           IN1(19) => IN1(19), IN1(18) => IN1(18), IN1(17) => 
                           IN1(17), IN1(16) => IN1(16), IN1(15) => IN1(15), 
                           IN1(14) => IN1(14), IN1(13) => IN1(13), IN1(12) => 
                           IN1(12), IN1(11) => IN1(11), IN1(10) => IN1(10), 
                           IN1(9) => IN1(9), IN1(8) => IN1(8), IN1(7) => IN1(7)
                           , IN1(6) => IN1(6), IN1(5) => IN1(5), IN1(4) => 
                           IN1(4), IN1(3) => IN1(3), IN1(2) => IN1(2), IN1(1) 
                           => IN1(1), IN1(0) => IN1(0), IN2(31) => IN2(31), 
                           IN2(30) => IN2(30), IN2(29) => IN2(29), IN2(28) => 
                           IN2(28), IN2(27) => IN2(27), IN2(26) => IN2(26), 
                           IN2(25) => IN2(25), IN2(24) => IN2(24), IN2(23) => 
                           IN2(23), IN2(22) => IN2(22), IN2(21) => IN2(21), 
                           IN2(20) => IN2(20), IN2(19) => IN2(19), IN2(18) => 
                           IN2(18), IN2(17) => IN2(17), IN2(16) => IN2(16), 
                           IN2(15) => IN2(15), IN2(14) => IN2(14), IN2(13) => 
                           IN2(13), IN2(12) => IN2(12), IN2(11) => IN2(11), 
                           IN2(10) => IN2(10), IN2(9) => IN2(9), IN2(8) => 
                           IN2(8), IN2(7) => n100, IN2(6) => IN2(6), IN2(5) => 
                           n98, IN2(4) => IN2(4), IN2(3) => n103, IN2(2) => 
                           IN2(2), IN2(1) => n101, IN2(0) => n102, CTRL(1) => 
                           ALUW_i(6), CTRL(0) => ALUW_i(5), OUT1(31) => 
                           lu_out_31_port, OUT1(30) => lu_out_30_port, OUT1(29)
                           => lu_out_29_port, OUT1(28) => lu_out_28_port, 
                           OUT1(27) => lu_out_27_port, OUT1(26) => 
                           lu_out_26_port, OUT1(25) => lu_out_25_port, OUT1(24)
                           => lu_out_24_port, OUT1(23) => lu_out_23_port, 
                           OUT1(22) => lu_out_22_port, OUT1(21) => 
                           lu_out_21_port, OUT1(20) => lu_out_20_port, OUT1(19)
                           => lu_out_19_port, OUT1(18) => lu_out_18_port, 
                           OUT1(17) => lu_out_17_port, OUT1(16) => 
                           lu_out_16_port, OUT1(15) => lu_out_15_port, OUT1(14)
                           => lu_out_14_port, OUT1(13) => lu_out_13_port, 
                           OUT1(12) => lu_out_12_port, OUT1(11) => 
                           lu_out_11_port, OUT1(10) => lu_out_10_port, OUT1(9) 
                           => lu_out_9_port, OUT1(8) => lu_out_8_port, OUT1(7) 
                           => lu_out_7_port, OUT1(6) => lu_out_6_port, OUT1(5) 
                           => lu_out_5_port, OUT1(4) => lu_out_4_port, OUT1(3) 
                           => lu_out_3_port, OUT1(2) => lu_out_2_port, OUT1(1) 
                           => lu_out_1_port, OUT1(0) => lu_out_0_port);
   U114 : MUX2_X1 port map( A => B_booth_to_add_8_port, B => IN2(8), S => n9, Z
                           => mux_B_8_port);
   U60 : AOI222_X1 port map( A1 => IN2(22), A2 => n17, B1 => n104, B2 => 
                           lu_out_22_port, C1 => n19, C2 => mult_out_22_port, 
                           ZN => n53);
   U59 : AOI22_X1 port map( A1 => n12, A2 => shift_out_22_port, B1 => n105, B2 
                           => sum_out_22_port, ZN => n54);
   U58 : NAND2_X1 port map( A1 => n53, A2 => n54, ZN => DOUT(22));
   U63 : AOI222_X1 port map( A1 => IN2(21), A2 => n17, B1 => n104, B2 => 
                           lu_out_21_port, C1 => n19, C2 => mult_out_21_port, 
                           ZN => n55);
   U62 : AOI22_X1 port map( A1 => n12, A2 => shift_out_21_port, B1 => n105, B2 
                           => sum_out_21_port, ZN => n56);
   U61 : NAND2_X1 port map( A1 => n55, A2 => n56, ZN => DOUT(21));
   U72 : AOI222_X1 port map( A1 => IN2(19), A2 => n17, B1 => n104, B2 => 
                           lu_out_19_port, C1 => n19, C2 => mult_out_19_port, 
                           ZN => n61);
   U71 : AOI22_X1 port map( A1 => n12, A2 => shift_out_19_port, B1 => n105, B2 
                           => sum_out_19_port, ZN => n62);
   U70 : NAND2_X1 port map( A1 => n61, A2 => n62, ZN => DOUT(19));
   U75 : AOI222_X1 port map( A1 => IN2(18), A2 => n17, B1 => n18, B2 => 
                           lu_out_18_port, C1 => n19, C2 => mult_out_18_port, 
                           ZN => n63);
   U74 : AOI22_X1 port map( A1 => n12, A2 => shift_out_18_port, B1 => n105, B2 
                           => sum_out_18_port, ZN => n64);
   U73 : NAND2_X1 port map( A1 => n63, A2 => n64, ZN => DOUT(18));
   U56 : AOI22_X1 port map( A1 => n12, A2 => shift_out_23_port, B1 => n105, B2 
                           => sum_out_23_port, ZN => n52);
   U55 : NAND2_X1 port map( A1 => n51, A2 => n52, ZN => DOUT(23));
   U45 : AOI222_X1 port map( A1 => IN2(27), A2 => n17, B1 => n104, B2 => 
                           lu_out_27_port, C1 => n19, C2 => mult_out_27_port, 
                           ZN => n43);
   U44 : AOI22_X1 port map( A1 => n12, A2 => shift_out_27_port, B1 => n105, B2 
                           => sum_out_27_port, ZN => n44);
   U43 : NAND2_X1 port map( A1 => n43, A2 => n44, ZN => DOUT(27));
   U48 : AOI222_X1 port map( A1 => IN2(26), A2 => n17, B1 => n104, B2 => 
                           lu_out_26_port, C1 => n19, C2 => mult_out_26_port, 
                           ZN => n45);
   U47 : AOI22_X1 port map( A1 => n12, A2 => shift_out_26_port, B1 => n105, B2 
                           => sum_out_26_port, ZN => n46);
   U46 : NAND2_X1 port map( A1 => n45, A2 => n46, ZN => DOUT(26));
   U77 : AOI22_X1 port map( A1 => n12, A2 => shift_out_17_port, B1 => n105, B2 
                           => sum_out_17_port, ZN => n66);
   U76 : NAND2_X1 port map( A1 => n65, A2 => n66, ZN => DOUT(17));
   U54 : AOI222_X1 port map( A1 => IN2(24), A2 => n17, B1 => n104, B2 => 
                           lu_out_24_port, C1 => n19, C2 => mult_out_24_port, 
                           ZN => n49);
   U52 : NAND2_X1 port map( A1 => n49, A2 => n50, ZN => DOUT(24));
   U66 : AOI222_X1 port map( A1 => IN2(20), A2 => n17, B1 => n104, B2 => 
                           lu_out_20_port, C1 => n19, C2 => mult_out_20_port, 
                           ZN => n57);
   U64 : NAND2_X1 port map( A1 => n57, A2 => n58, ZN => DOUT(20));
   U51 : AOI222_X1 port map( A1 => IN2(25), A2 => n17, B1 => n104, B2 => 
                           lu_out_25_port, C1 => n19, C2 => mult_out_25_port, 
                           ZN => n47);
   U49 : NAND2_X1 port map( A1 => n47, A2 => n48, ZN => DOUT(25));
   U28 : AOI22_X1 port map( A1 => n104, A2 => lu_out_31_port, B1 => n19, B2 => 
                           mult_out_31_port, ZN => n34);
   U27 : OAI211_X1 port map( C1 => n32, C2 => n94, A => n33, B => n34, ZN => 
                           DOUT(31));
   U33 : AOI222_X1 port map( A1 => IN2(30), A2 => n17, B1 => n104, B2 => 
                           lu_out_30_port, C1 => n19, C2 => mult_out_30_port, 
                           ZN => n35);
   U32 : AOI22_X1 port map( A1 => n12, A2 => shift_out_30_port, B1 => n105, B2 
                           => sum_out_30_port, ZN => n36);
   U31 : NAND2_X1 port map( A1 => n35, A2 => n36, ZN => DOUT(30));
   U39 : AOI222_X1 port map( A1 => IN2(29), A2 => n17, B1 => n104, B2 => 
                           lu_out_29_port, C1 => n19, C2 => mult_out_29_port, 
                           ZN => n39);
   U38 : AOI22_X1 port map( A1 => n12, A2 => shift_out_29_port, B1 => n105, B2 
                           => sum_out_29_port, ZN => n40);
   U37 : NAND2_X1 port map( A1 => n39, A2 => n40, ZN => DOUT(29));
   U42 : AOI222_X1 port map( A1 => IN2(28), A2 => n17, B1 => n104, B2 => 
                           lu_out_28_port, C1 => n19, C2 => mult_out_28_port, 
                           ZN => n41);
   U40 : NAND2_X1 port map( A1 => n41, A2 => n42, ZN => DOUT(28));
   U81 : AOI222_X1 port map( A1 => IN2(16), A2 => n17, B1 => n104, B2 => 
                           lu_out_16_port, C1 => n19, C2 => mult_out_16_port, 
                           ZN => n67);
   U80 : AOI22_X1 port map( A1 => n12, A2 => shift_out_16_port, B1 => n105, B2 
                           => sum_out_16_port, ZN => n68);
   U79 : NAND2_X1 port map( A1 => n67, A2 => n68, ZN => DOUT(16));
   U13 : AOI22_X1 port map( A1 => n15, A2 => shift_out_7_port, B1 => n105, B2 
                           => sum_out_7_port, ZN => n23);
   U12 : NAND2_X1 port map( A1 => n22, A2 => n23, ZN => DOUT(7));
   U95 : AOI22_X1 port map( A1 => n12, A2 => shift_out_11_port, B1 => n105, B2 
                           => sum_out_11_port, ZN => n78);
   U94 : NAND2_X1 port map( A1 => n77, A2 => n78, ZN => DOUT(11));
   U89 : AOI22_X1 port map( A1 => n12, A2 => shift_out_13_port, B1 => n105, B2 
                           => sum_out_13_port, ZN => n74);
   U88 : NAND2_X1 port map( A1 => n73, A2 => n74, ZN => DOUT(13));
   U87 : AOI222_X1 port map( A1 => IN2(14), A2 => n17, B1 => n104, B2 => 
                           lu_out_14_port, C1 => n19, C2 => mult_out_14_port, 
                           ZN => n71);
   U86 : AOI22_X1 port map( A1 => n12, A2 => shift_out_14_port, B1 => n105, B2 
                           => sum_out_14_port, ZN => n72);
   U85 : NAND2_X1 port map( A1 => n71, A2 => n72, ZN => DOUT(14));
   U93 : AOI222_X1 port map( A1 => IN2(12), A2 => n17, B1 => n104, B2 => 
                           lu_out_12_port, C1 => n19, C2 => mult_out_12_port, 
                           ZN => n75);
   U92 : AOI22_X1 port map( A1 => n12, A2 => shift_out_12_port, B1 => n105, B2 
                           => sum_out_12_port, ZN => n76);
   U91 : NAND2_X1 port map( A1 => n75, A2 => n76, ZN => DOUT(12));
   U98 : AOI22_X1 port map( A1 => n12, A2 => shift_out_10_port, B1 => n105, B2 
                           => sum_out_10_port, ZN => n80);
   U97 : NAND2_X1 port map( A1 => n79, A2 => n80, ZN => DOUT(10));
   U7 : AOI22_X1 port map( A1 => n12, A2 => shift_out_9_port, B1 => n105, B2 =>
                           sum_out_9_port, ZN => n14);
   U6 : NAND2_X1 port map( A1 => n13, A2 => n14, ZN => DOUT(9));
   U26 : AOI222_X1 port map( A1 => n103, A2 => n17, B1 => n104, B2 => 
                           lu_out_3_port, C1 => n19, C2 => mult_out_3_port, ZN 
                           => n30);
   U25 : AOI22_X1 port map( A1 => n12, A2 => shift_out_3_port, B1 => n105, B2 
                           => sum_out_3_port, ZN => n31);
   U24 : NAND2_X1 port map( A1 => n30, A2 => n31, ZN => DOUT(3));
   U16 : AOI22_X1 port map( A1 => n12, A2 => shift_out_6_port, B1 => n105, B2 
                           => sum_out_6_port, ZN => n25);
   U15 : NAND2_X1 port map( A1 => n24, A2 => n25, ZN => DOUT(6));
   U68 : AOI22_X1 port map( A1 => n12, A2 => shift_out_1_port, B1 => n105, B2 
                           => sum_out_1_port, ZN => n60);
   U67 : NAND2_X1 port map( A1 => n59, A2 => n60, ZN => DOUT(1));
   U35 : AOI22_X1 port map( A1 => n12, A2 => shift_out_2_port, B1 => n105, B2 
                           => sum_out_2_port, ZN => n38);
   U34 : NAND2_X1 port map( A1 => n37, A2 => n38, ZN => DOUT(2));
   U19 : AOI22_X1 port map( A1 => n12, A2 => shift_out_5_port, B1 => n105, B2 
                           => sum_out_5_port, ZN => n27);
   U18 : NAND2_X1 port map( A1 => n26, A2 => n27, ZN => DOUT(5));
   U22 : AOI22_X1 port map( A1 => n15, A2 => shift_out_4_port, B1 => n105, B2 
                           => sum_out_4_port, ZN => n29);
   U21 : NAND2_X1 port map( A1 => n28, A2 => n29, ZN => DOUT(4));
   U11 : AOI222_X1 port map( A1 => IN2(8), A2 => n17, B1 => n104, B2 => 
                           lu_out_8_port, C1 => n19, C2 => mult_out_8_port, ZN 
                           => n20);
   U10 : AOI22_X1 port map( A1 => n12, A2 => shift_out_8_port, B1 => n16, B2 =>
                           sum_out_8_port, ZN => n21);
   U9 : NAND2_X1 port map( A1 => n20, A2 => n21, ZN => DOUT(8));
   U101 : AND2_X2 port map( A1 => n32, A2 => ALUW_i(12), ZN => n19);
   U105 : INV_X2 port map( A => n32, ZN => n17);
   U2 : NOR2_X1 port map( A1 => valid_from_booth, A2 => n9, ZN => stall_o);
   U108 : INV_X1 port map( A => ALUW_i(11), ZN => n84);
   U3 : MUX2_X1 port map( A => B_booth_to_add_5_port, B => IN2(5), S => n9, Z 
                           => mux_B_5_port);
   U4 : MUX2_X1 port map( A => B_booth_to_add_4_port, B => IN2(4), S => n9, Z 
                           => mux_B_4_port);
   U5 : INV_X1 port map( A => ALUW_i(10), ZN => n1);
   U8 : NOR3_X1 port map( A1 => ALUW_i(12), A2 => n84, A3 => n1, ZN => n70);
   U14 : INV_X1 port map( A => IN2(2), ZN => n2);
   U17 : INV_X1 port map( A => n9, ZN => n3);
   U20 : AOI22_X1 port map( A1 => n9, A2 => n2, B1 => n86, B2 => n3, ZN => 
                           mux_B_2_port);
   U23 : INV_X1 port map( A => n9, ZN => n4);
   U29 : NAND2_X1 port map( A1 => B_booth_to_add_0_port, A2 => n4, ZN => n83);
   U30 : MUX2_X1 port map( A => B_booth_to_add_7_port, B => IN2(7), S => n9, Z 
                           => mux_B_7_port);
   U36 : MUX2_X1 port map( A => B_booth_to_add_21_port, B => IN2(21), S => n106
                           , Z => mux_B_21_port);
   U41 : AOI222_X1 port map( A1 => sum_out_0_port, A2 => n105, B1 => n102, B2 
                           => n17, C1 => n104, C2 => lu_out_0_port, ZN => n5);
   U50 : INV_X1 port map( A => n5, ZN => n6);
   U53 : AOI21_X1 port map( B1 => n19, B2 => mult_out_0_port, A => n6, ZN => 
                           n96);
   U57 : INV_X1 port map( A => IN2(15), ZN => n7);
   U65 : INV_X1 port map( A => n17, ZN => n8);
   U69 : AOI22_X1 port map( A1 => mult_out_15_port, A2 => n19, B1 => 
                           lu_out_15_port, B2 => n104, ZN => n10);
   U78 : AOI22_X1 port map( A1 => sum_out_15_port, A2 => n105, B1 => 
                           shift_out_15_port, B2 => n12, ZN => n11);
   U82 : OAI211_X1 port map( C1 => n7, C2 => n8, A => n10, B => n11, ZN => 
                           DOUT(15));
   U83 : MUX2_X2 port map( A => sign_booth_to_add, B => ALUW_i(7), S => n9, Z 
                           => mux_sign);
   U84 : BUF_X1 port map( A => IN2(5), Z => n98);
   U90 : BUF_X1 port map( A => IN2(3), Z => n103);
   U96 : OR2_X1 port map( A1 => n9, A2 => n90, ZN => n82);
   U99 : AOI222_X1 port map( A1 => IN2(10), A2 => n17, B1 => n104, B2 => 
                           lu_out_10_port, C1 => n19, C2 => mult_out_10_port, 
                           ZN => n79);
   U100 : AOI222_X1 port map( A1 => IN2(11), A2 => n17, B1 => n18, B2 => 
                           lu_out_11_port, C1 => n19, C2 => mult_out_11_port, 
                           ZN => n77);
   U102 : AND2_X1 port map( A1 => n97, A2 => n96, ZN => n69);
   U103 : INV_X1 port map( A => IN2(31), ZN => n94);
   U104 : BUF_X1 port map( A => IN2(1), Z => n101);
   U106 : OR2_X1 port map( A1 => n88, A2 => n9, ZN => n81);
   U107 : BUF_X2 port map( A => n15, Z => n12);
   U109 : BUF_X2 port map( A => n16, Z => n105);
   U110 : INV_X1 port map( A => ALUW_i(10), ZN => n85);
   U111 : INV_X1 port map( A => B_booth_to_add_10_port, ZN => n90);
   U112 : INV_X1 port map( A => B_booth_to_add_2_port, ZN => n86);
   U115 : INV_X1 port map( A => B_booth_to_add_3_port, ZN => n88);
   U117 : NAND2_X1 port map( A1 => n95, A2 => n69, ZN => DOUT(0));
   U118 : CLKBUF_X1 port map( A => IN2(0), Z => n102);
   U119 : AOI222_X1 port map( A1 => IN2(9), A2 => n17, B1 => n18, B2 => 
                           lu_out_9_port, C1 => n19, C2 => mult_out_9_port, ZN 
                           => n13);
   U122 : NAND2_X1 port map( A1 => comp_out, A2 => n70, ZN => n95);
   U131 : INV_X4 port map( A => ALUW_i(1), ZN => n9);
   U133 : BUF_X1 port map( A => n9, Z => n106);
   U140 : NOR3_X1 port map( A1 => ALUW_i(12), A2 => ALUW_i(10), A3 => n84, ZN 
                           => n15);
   U143 : BUF_X1 port map( A => n18, Z => n104);
   U144 : NOR3_X1 port map( A1 => ALUW_i(11), A2 => ALUW_i(12), A3 => n85, ZN 
                           => n18);
   U176 : NOR3_X1 port map( A1 => ALUW_i(11), A2 => ALUW_i(12), A3 => 
                           ALUW_i(10), ZN => n16);
   U177 : BUF_X1 port map( A => IN2(7), Z => n100);
   U179 : BUF_X1 port map( A => sum_out_31_port, Z => n99);
   U180 : AOI222_X1 port map( A1 => IN2(4), A2 => n17, B1 => n104, B2 => 
                           lu_out_4_port, C1 => n19, C2 => mult_out_4_port, ZN 
                           => n28);
   U181 : AOI222_X1 port map( A1 => n98, A2 => n17, B1 => n104, B2 => 
                           lu_out_5_port, C1 => n19, C2 => mult_out_5_port, ZN 
                           => n26);
   U182 : AOI222_X1 port map( A1 => IN2(2), A2 => n17, B1 => n104, B2 => 
                           lu_out_2_port, C1 => n19, C2 => mult_out_2_port, ZN 
                           => n37);
   U183 : AOI222_X1 port map( A1 => n101, A2 => n17, B1 => n18, B2 => 
                           lu_out_1_port, C1 => n19, C2 => mult_out_1_port, ZN 
                           => n59);
   U184 : AOI222_X1 port map( A1 => IN2(6), A2 => n17, B1 => n104, B2 => 
                           lu_out_6_port, C1 => n19, C2 => mult_out_6_port, ZN 
                           => n24);
   U185 : AOI222_X1 port map( A1 => n100, A2 => n17, B1 => n104, B2 => 
                           lu_out_7_port, C1 => n19, C2 => mult_out_7_port, ZN 
                           => n22);
   U186 : AOI222_X1 port map( A1 => IN2(17), A2 => n17, B1 => n104, B2 => 
                           lu_out_17_port, C1 => n19, C2 => mult_out_17_port, 
                           ZN => n65);
   U187 : AOI222_X1 port map( A1 => IN2(23), A2 => n17, B1 => n18, B2 => 
                           lu_out_23_port, C1 => n19, C2 => mult_out_23_port, 
                           ZN => n51);
   U188 : NAND2_X1 port map( A1 => shift_out_0_port, A2 => n12, ZN => n97);
   U189 : NAND2_X1 port map( A1 => n94, A2 => IN1(31), ZN => n92);
   U190 : MUX2_X1 port map( A => B_booth_to_add_1_port, B => IN2(1), S => n106,
                           Z => mux_B_1_port);
   U191 : MUX2_X1 port map( A => A_booth_to_add_0_port, B => IN1(0), S => n9, Z
                           => mux_A_0_port);
   U192 : MUX2_X1 port map( A => B_booth_to_add_13_port, B => IN2(13), S => 
                           n106, Z => mux_B_13_port);
   U193 : NAND2_X1 port map( A1 => n91, A2 => n83, ZN => mux_B_0_port);
   U194 : OAI22_X1 port map( A1 => sum_out_31_port, A2 => n92, B1 => n93, B2 =>
                           IN1(31), ZN => overflow);
   U195 : NAND2_X1 port map( A1 => IN2(3), A2 => n9, ZN => n87);
   U196 : NAND2_X1 port map( A1 => n87, A2 => n81, ZN => mux_B_3_port);
   U197 : NAND2_X1 port map( A1 => IN2(10), A2 => n9, ZN => n89);
   U198 : NAND2_X1 port map( A1 => n89, A2 => n82, ZN => mux_B_10_port);
   U199 : NAND2_X1 port map( A1 => IN2(0), A2 => n9, ZN => n91);
   U200 : NAND2_X1 port map( A1 => sum_out_31_port, A2 => IN2(31), ZN => n93);
   U201 : AOI222_X1 port map( A1 => IN2(13), A2 => n17, B1 => n18, B2 => 
                           lu_out_13_port, C1 => n19, C2 => mult_out_13_port, 
                           ZN => n73);
   U202 : AOI22_X1 port map( A1 => n12, A2 => shift_out_20_port, B1 => n16, B2 
                           => sum_out_20_port, ZN => n58);
   U203 : AOI22_X1 port map( A1 => n12, A2 => shift_out_25_port, B1 => n16, B2 
                           => sum_out_25_port, ZN => n48);
   U204 : AOI22_X1 port map( A1 => n12, A2 => shift_out_28_port, B1 => n16, B2 
                           => sum_out_28_port, ZN => n42);
   U205 : AOI22_X1 port map( A1 => n12, A2 => shift_out_24_port, B1 => n16, B2 
                           => sum_out_24_port, ZN => n50);
   U206 : AOI22_X1 port map( A1 => n12, A2 => shift_out_31_port, B1 => n99, B2 
                           => n105, ZN => n33);

end SYN_Bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity ff32_en_SIZE13 is

   port( D : in std_logic_vector (12 downto 0);  en, clk, rst : in std_logic;  
         Q : out std_logic_vector (12 downto 0));

end ff32_en_SIZE13;

architecture SYN_behavioral of ff32_en_SIZE13 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFR_X2
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_ff32_en_SIZE13
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   signal net199388, n1, n2, n3, n4, n5, n7, n8, n9, n12, n14, n6, n10, n11, 
      n13 : std_logic;

begin
   
   Q_reg_12_inst : DFFR_X1 port map( D => D(12), CK => net199388, RN => n13, Q 
                           => Q(12), QN => n14);
   Q_reg_11_inst : DFFR_X1 port map( D => D(11), CK => net199388, RN => n13, Q 
                           => Q(11), QN => n12);
   Q_reg_8_inst : DFFR_X1 port map( D => D(8), CK => net199388, RN => n13, Q =>
                           Q(8), QN => n9);
   Q_reg_7_inst : DFFR_X1 port map( D => D(7), CK => net199388, RN => n13, Q =>
                           Q(7), QN => n8);
   Q_reg_6_inst : DFFR_X1 port map( D => D(6), CK => net199388, RN => n13, Q =>
                           Q(6), QN => n7);
   Q_reg_4_inst : DFFR_X1 port map( D => D(4), CK => net199388, RN => n13, Q =>
                           Q(4), QN => n5);
   Q_reg_3_inst : DFFR_X1 port map( D => D(3), CK => net199388, RN => n13, Q =>
                           Q(3), QN => n4);
   Q_reg_2_inst : DFFR_X1 port map( D => D(2), CK => net199388, RN => n13, Q =>
                           Q(2), QN => n3);
   Q_reg_1_inst : DFFR_X1 port map( D => D(1), CK => net199388, RN => n13, Q =>
                           Q(1), QN => n2);
   Q_reg_0_inst : DFFR_X1 port map( D => D(0), CK => net199388, RN => n13, Q =>
                           Q(0), QN => n1);
   clk_gate_Q_reg : SNPS_CLOCK_GATE_HIGH_ff32_en_SIZE13 port map( CLK => clk, 
                           EN => en, ENCLK => net199388);
   Q_reg_5_inst : DFFR_X2 port map( D => D(5), CK => net199388, RN => n13, Q =>
                           Q(5), QN => n11);
   Q_reg_9_inst : DFFR_X2 port map( D => D(9), CK => net199388, RN => n13, Q =>
                           Q(9), QN => n10);
   Q_reg_10_inst : DFFR_X1 port map( D => D(10), CK => net199388, RN => n13, Q 
                           => Q(10), QN => n6);
   U2 : INV_X1 port map( A => rst, ZN => n13);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity ff32_en_SIZE5_0 is

   port( D : in std_logic_vector (4 downto 0);  en, clk, rst : in std_logic;  Q
         : out std_logic_vector (4 downto 0));

end ff32_en_SIZE5_0;

architecture SYN_behavioral of ff32_en_SIZE5_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_ff32_en_SIZE5_0
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal net199373, n1, n2, n3, n4, n6, n5 : std_logic;

begin
   
   Q_reg_4_inst : DFFR_X1 port map( D => D(4), CK => net199373, RN => n5, Q => 
                           Q(4), QN => n6);
   Q_reg_3_inst : DFFR_X1 port map( D => D(3), CK => net199373, RN => n5, Q => 
                           Q(3), QN => n4);
   Q_reg_2_inst : DFFR_X1 port map( D => D(2), CK => net199373, RN => n5, Q => 
                           Q(2), QN => n3);
   Q_reg_1_inst : DFFR_X1 port map( D => D(1), CK => net199373, RN => n5, Q => 
                           Q(1), QN => n2);
   Q_reg_0_inst : DFFR_X1 port map( D => D(0), CK => net199373, RN => n5, Q => 
                           Q(0), QN => n1);
   clk_gate_Q_reg : SNPS_CLOCK_GATE_HIGH_ff32_en_SIZE5_0 port map( CLK => clk, 
                           EN => en, ENCLK => net199373);
   U2 : INV_X1 port map( A => rst, ZN => n5);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity ff32_en_SIZE32_0 is

   port( D : in std_logic_vector (31 downto 0);  en, clk, rst : in std_logic;  
         Q : out std_logic_vector (31 downto 0));

end ff32_en_SIZE32_0;

architecture SYN_behavioral of ff32_en_SIZE32_0 is

   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_ff32_en_SIZE32_0
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal net199358, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, 
      n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28
      , n29, n30, n31, n33, n32 : std_logic;

begin
   
   Q_reg_31_inst : DFFR_X1 port map( D => D(31), CK => net199358, RN => n32, Q 
                           => Q(31), QN => n33);
   Q_reg_30_inst : DFFR_X1 port map( D => D(30), CK => net199358, RN => n32, Q 
                           => Q(30), QN => n31);
   Q_reg_29_inst : DFFR_X1 port map( D => D(29), CK => net199358, RN => n32, Q 
                           => Q(29), QN => n30);
   Q_reg_28_inst : DFFR_X1 port map( D => D(28), CK => net199358, RN => n32, Q 
                           => Q(28), QN => n29);
   Q_reg_27_inst : DFFR_X1 port map( D => D(27), CK => net199358, RN => n32, Q 
                           => Q(27), QN => n28);
   Q_reg_26_inst : DFFR_X1 port map( D => D(26), CK => net199358, RN => n32, Q 
                           => Q(26), QN => n27);
   Q_reg_25_inst : DFFR_X1 port map( D => D(25), CK => net199358, RN => n32, Q 
                           => Q(25), QN => n26);
   Q_reg_24_inst : DFFR_X1 port map( D => D(24), CK => net199358, RN => n32, Q 
                           => Q(24), QN => n25);
   Q_reg_23_inst : DFFR_X1 port map( D => D(23), CK => net199358, RN => n32, Q 
                           => Q(23), QN => n24);
   Q_reg_22_inst : DFFR_X1 port map( D => D(22), CK => net199358, RN => n32, Q 
                           => Q(22), QN => n23);
   Q_reg_21_inst : DFFR_X1 port map( D => D(21), CK => net199358, RN => n32, Q 
                           => Q(21), QN => n22);
   Q_reg_20_inst : DFFR_X1 port map( D => D(20), CK => net199358, RN => n32, Q 
                           => Q(20), QN => n21);
   Q_reg_19_inst : DFFR_X1 port map( D => D(19), CK => net199358, RN => n32, Q 
                           => Q(19), QN => n20);
   Q_reg_18_inst : DFFR_X1 port map( D => D(18), CK => net199358, RN => n32, Q 
                           => Q(18), QN => n19);
   Q_reg_17_inst : DFFR_X1 port map( D => D(17), CK => net199358, RN => n32, Q 
                           => Q(17), QN => n18);
   Q_reg_16_inst : DFFR_X1 port map( D => D(16), CK => net199358, RN => n32, Q 
                           => Q(16), QN => n17);
   Q_reg_15_inst : DFFR_X1 port map( D => D(15), CK => net199358, RN => n32, Q 
                           => Q(15), QN => n16);
   Q_reg_14_inst : DFFR_X1 port map( D => D(14), CK => net199358, RN => n32, Q 
                           => Q(14), QN => n15);
   Q_reg_13_inst : DFFR_X1 port map( D => D(13), CK => net199358, RN => n32, Q 
                           => Q(13), QN => n14);
   Q_reg_12_inst : DFFR_X1 port map( D => D(12), CK => net199358, RN => n32, Q 
                           => Q(12), QN => n13);
   Q_reg_11_inst : DFFR_X1 port map( D => D(11), CK => net199358, RN => n32, Q 
                           => Q(11), QN => n12);
   Q_reg_10_inst : DFFR_X1 port map( D => D(10), CK => net199358, RN => n32, Q 
                           => Q(10), QN => n11);
   Q_reg_9_inst : DFFR_X1 port map( D => D(9), CK => net199358, RN => n32, Q =>
                           Q(9), QN => n10);
   Q_reg_8_inst : DFFR_X1 port map( D => D(8), CK => net199358, RN => n32, Q =>
                           Q(8), QN => n9);
   Q_reg_7_inst : DFFR_X1 port map( D => D(7), CK => net199358, RN => n32, Q =>
                           Q(7), QN => n8);
   Q_reg_6_inst : DFFR_X1 port map( D => D(6), CK => net199358, RN => n32, Q =>
                           Q(6), QN => n7);
   Q_reg_5_inst : DFFR_X1 port map( D => D(5), CK => net199358, RN => n32, Q =>
                           Q(5), QN => n6);
   Q_reg_4_inst : DFFR_X1 port map( D => D(4), CK => net199358, RN => n32, Q =>
                           Q(4), QN => n5);
   Q_reg_3_inst : DFFR_X1 port map( D => D(3), CK => net199358, RN => n32, Q =>
                           Q(3), QN => n4);
   Q_reg_2_inst : DFFR_X1 port map( D => D(2), CK => net199358, RN => n32, Q =>
                           Q(2), QN => n3);
   Q_reg_1_inst : DFFR_X1 port map( D => D(1), CK => net199358, RN => n32, Q =>
                           Q(1), QN => n2);
   Q_reg_0_inst : DFFR_X1 port map( D => D(0), CK => net199358, RN => n32, Q =>
                           Q(0), QN => n1);
   clk_gate_Q_reg : SNPS_CLOCK_GATE_HIGH_ff32_en_SIZE32_0 port map( CLK => clk,
                           EN => en, ENCLK => net199358);
   U2 : INV_X2 port map( A => rst, ZN => n32);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_dlx_regfile_0 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_dlx_regfile_0;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_dlx_regfile_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net199397 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net199397);
   main_gate : AND2_X1 port map( A1 => net199397, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity 
   SNPS_CLOCK_GATE_HIGH_dlx_cu_MICROCODE_MEM_SIZE64_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE13_0 
   is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end 
   SNPS_CLOCK_GATE_HIGH_dlx_cu_MICROCODE_MEM_SIZE64_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE13_0;

architecture SYN_USE_DEFA_ARCH_NAME of 
   SNPS_CLOCK_GATE_HIGH_dlx_cu_MICROCODE_MEM_SIZE64_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE13_0 
   is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net199577 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net199577);
   main_gate : AND2_X1 port map( A1 => net199577, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity alu_ctrl is

   port( OP : in std_logic_vector (0 to 4);  ALU_WORD : out std_logic_vector 
         (12 downto 0));

end alu_ctrl;

architecture SYN_bhe of alu_ctrl is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal ALU_WORD_12_port, ALU_WORD_11_port, ALU_WORD_10_port, ALU_WORD_9_port
      , ALU_WORD_8_port, ALU_WORD_7_port, ALU_WORD_6_port, ALU_WORD_5_port, 
      ALU_WORD_4_port, ALU_WORD_3_port, ALU_WORD_2_port, ALU_WORD_1_port, 
      ALU_WORD_0_port, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, 
      N31, N32, N33, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, 
      n14, n15, n16, n17, n18, n19, n20_port, n21_port, n22_port, n23_port, 
      n24_port, n25_port, n26_port, n27_port, n28_port, n29_port, n30_port, 
      n31_port, n32_port, n33_port, n34, n35 : std_logic;

begin
   ALU_WORD <= ( ALU_WORD_12_port, ALU_WORD_11_port, ALU_WORD_10_port, 
      ALU_WORD_9_port, ALU_WORD_8_port, ALU_WORD_7_port, ALU_WORD_6_port, 
      ALU_WORD_5_port, ALU_WORD_4_port, ALU_WORD_3_port, ALU_WORD_2_port, 
      ALU_WORD_1_port, ALU_WORD_0_port );
   
   comp_sel_reg_2_inst : DLH_X1 port map( G => N32, D => N33, Q => 
                           ALU_WORD_4_port);
   comp_sel_reg_1_inst : DLH_X1 port map( G => N32, D => N31, Q => 
                           ALU_WORD_3_port);
   comp_sel_reg_0_inst : DLH_X1 port map( G => N32, D => N30, Q => 
                           ALU_WORD_2_port);
   sign_to_booth_reg : DLH_X1 port map( G => N20, D => N21, Q => 
                           ALU_WORD_0_port);
   left_right_reg : DLH_X1 port map( G => N23, D => N22, Q => ALU_WORD_9_port);
   logic_arith_reg : DLH_X1 port map( G => N23, D => N24, Q => ALU_WORD_8_port)
                           ;
   sign_to_adder_reg : DLH_X1 port map( G => N25, D => N26, Q => 
                           ALU_WORD_7_port);
   lu_ctrl_reg_1_inst : DLH_X1 port map( G => N28, D => N29, Q => 
                           ALU_WORD_6_port);
   lu_ctrl_reg_0_inst : DLH_X1 port map( G => N28, D => N27, Q => 
                           ALU_WORD_5_port);
   U53 : NAND3_X1 port map( A1 => n9, A2 => OP(3), A3 => n28_port, ZN => 
                           n30_port);
   U54 : NAND3_X1 port map( A1 => n15, A2 => n35, A3 => n22_port, ZN => n19);
   U48 : NOR3_X1 port map( A1 => OP(2), A2 => OP(4), A3 => n22_port, ZN => n10)
                           ;
   U45 : NOR3_X1 port map( A1 => OP(2), A2 => n35, A3 => n22_port, ZN => 
                           n33_port);
   U43 : NOR2_X1 port map( A1 => n3, A2 => n2, ZN => n32_port);
   U41 : NOR2_X1 port map( A1 => OP(4), A2 => n15, ZN => n28_port);
   U40 : NAND2_X1 port map( A1 => n28_port, A2 => n22_port, ZN => n1);
   U39 : NOR2_X1 port map( A1 => n19, A2 => OP(1), ZN => n34);
   U38 : NOR4_X1 port map( A1 => n15, A2 => n3, A3 => n35, A4 => n22_port, ZN 
                           => n8);
   U37 : AOI21_X1 port map( B1 => n34, B2 => OP(0), A => n8, ZN => n18);
   U36 : NAND2_X1 port map( A1 => n33_port, A2 => n26_port, ZN => n6);
   U35 : OAI211_X1 port map( C1 => n1, C2 => n16, A => n18, B => n6, ZN => N30)
                           ;
   U34 : AOI211_X1 port map( C1 => n26_port, C2 => n10, A => n32_port, B => N30
                           , ZN => n29_port);
   U33 : NAND2_X1 port map( A1 => OP(4), A2 => n22_port, ZN => n27_port);
   U32 : NOR2_X1 port map( A1 => n3, A2 => n27_port, ZN => n31_port);
   U31 : NAND2_X1 port map( A1 => OP(2), A2 => n31_port, ZN => n4);
   U29 : NOR2_X1 port map( A1 => OP(2), A2 => n27_port, ZN => n24_port);
   U28 : NAND2_X1 port map( A1 => n26_port, A2 => n24_port, ZN => n7);
   U27 : NAND4_X1 port map( A1 => n29_port, A2 => n4, A3 => n30_port, A4 => n7,
                           ZN => N32);
   U26 : AOI211_X1 port map( C1 => OP(4), C2 => OP(3), A => OP(2), B => n3, ZN 
                           => N28);
   U25 : NAND2_X1 port map( A1 => OP(3), A2 => n28_port, ZN => n17);
   U24 : OAI21_X1 port map( B1 => n27_port, B2 => n15, A => n17, ZN => n25_port
                           );
   U23 : NAND2_X1 port map( A1 => n25_port, A2 => n26_port, ZN => n20_port);
   U18 : NOR3_X1 port map( A1 => OP(2), A2 => n22_port, A3 => n13, ZN => N22);
   U16 : OAI21_X1 port map( B1 => n11, B2 => n13, A => n21_port, ZN => N23);
   U14 : OAI21_X1 port map( B1 => n19, B2 => n13, A => n20_port, ZN => 
                           ALU_WORD_12_port);
   U6 : NOR2_X1 port map( A1 => n3, A2 => n11, ZN => N27);
   U8 : NAND2_X1 port map( A1 => OP(2), A2 => OP(3), ZN => n12);
   U7 : OAI21_X1 port map( B1 => n12, B2 => n13, A => n14, ZN => N26);
   U11 : NOR2_X1 port map( A1 => n2, A2 => n13, ZN => N24);
   U12 : OAI211_X1 port map( C1 => n16, C2 => n17, A => n18, B => n4, ZN => N21
                           );
   U3 : NAND4_X1 port map( A1 => n4, A2 => n5, A3 => n6, A4 => n7, ZN => N31);
   U2 : AOI21_X1 port map( B1 => n1, B2 => n2, A => n3, ZN => N33);
   U9 : OAI21_X1 port map( B1 => n15, B2 => n13, A => n14, ZN => N25);
   U47 : NAND2_X1 port map( A1 => OP(1), A2 => n23_port, ZN => n3);
   U19 : NAND2_X1 port map( A1 => n23_port, A2 => n16, ZN => n13);
   U50 : NOR2_X1 port map( A1 => n23_port, A2 => n16, ZN => n26_port);
   U46 : INV_X1 port map( A => OP(4), ZN => n35);
   U42 : INV_X1 port map( A => OP(2), ZN => n15);
   U52 : INV_X1 port map( A => OP(0), ZN => n23_port);
   U51 : INV_X1 port map( A => OP(1), ZN => n16);
   U30 : INV_X1 port map( A => n3, ZN => n9);
   U49 : INV_X1 port map( A => OP(3), ZN => n22_port);
   U4 : INV_X1 port map( A => n8, ZN => n5);
   U44 : INV_X1 port map( A => n33_port, ZN => n2);
   U5 : AND2_X1 port map( A1 => n9, A2 => n10, ZN => N29);
   U17 : INV_X1 port map( A => N22, ZN => n21_port);
   U20 : INV_X1 port map( A => n24_port, ZN => n11);
   U22 : INV_X1 port map( A => n20_port, ZN => ALU_WORD_1_port);
   U15 : OR2_X1 port map( A1 => N32, A2 => N23, ZN => ALU_WORD_11_port);
   U21 : OR3_X1 port map( A1 => N32, A2 => N28, A3 => ALU_WORD_1_port, ZN => 
                           ALU_WORD_10_port);
   U10 : INV_X1 port map( A => N32, ZN => n14);
   U13 : OR2_X1 port map( A1 => N32, A2 => ALU_WORD_12_port, ZN => N20);

end SYN_bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity cw_mem_MICROCODE_MEM_SIZE64_OP_CODE_SIZE6_CW_SIZE13 is

   port( OPCODE_IN : in std_logic_vector (5 downto 0);  CW_OUT : out 
         std_logic_vector (12 downto 0));

end cw_mem_MICROCODE_MEM_SIZE64_OP_CODE_SIZE6_CW_SIZE13;

architecture SYN_bhe of cw_mem_MICROCODE_MEM_SIZE64_OP_CODE_SIZE6_CW_SIZE13 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal CW_OUT_12_port, CW_OUT_11_port, CW_OUT_10_port, CW_OUT_9_port, 
      CW_OUT_8_port, CW_OUT_7_port, CW_OUT_5_port, CW_OUT_4, CW_OUT_3, CW_OUT_2
      , CW_OUT_1, CW_OUT_0, n6, n7, n8, n9, n10, n11, n12, n13, n14, n17, n18, 
      n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n1, n2 : std_logic
      ;

begin
   CW_OUT <= ( CW_OUT_12_port, CW_OUT_11_port, CW_OUT_10_port, CW_OUT_9_port, 
      CW_OUT_8_port, CW_OUT_7_port, CW_OUT_5_port, CW_OUT_5_port, CW_OUT_4, 
      CW_OUT_3, CW_OUT_2, CW_OUT_1, CW_OUT_0 );
   
   U35 : NAND3_X1 port map( A1 => OPCODE_IN(3), A2 => n23, A3 => n24, ZN => n22
                           );
   U36 : NAND3_X1 port map( A1 => OPCODE_IN(4), A2 => n14, A3 => n25, ZN => n29
                           );
   U8 : NOR2_X1 port map( A1 => n10, A2 => n17, ZN => CW_OUT_8_port);
   U23 : OAI21_X1 port map( B1 => OPCODE_IN(3), B2 => n17, A => n29, ZN => 
                           CW_OUT_11_port);
   U5 : NAND2_X1 port map( A1 => n13, A2 => n14, ZN => n11);
   U4 : OAI22_X1 port map( A1 => OPCODE_IN(3), A2 => n11, B1 => n12, B2 => n10,
                           ZN => CW_OUT_4);
   U20 : NAND2_X1 port map( A1 => OPCODE_IN(5), A2 => n28, ZN => n8);
   U19 : NOR2_X1 port map( A1 => n7, A2 => n8, ZN => CW_OUT_3);
   U1 : NOR3_X1 port map( A1 => n6, A2 => n7, A3 => n8, ZN => CW_OUT_2);
   U16 : NAND2_X1 port map( A1 => OPCODE_IN(3), A2 => OPCODE_IN(4), ZN => n20);
   U15 : NAND2_X1 port map( A1 => n23, A2 => n7, ZN => n27);
   U3 : NOR2_X1 port map( A1 => n8, A2 => n10, ZN => CW_OUT_1);
   U22 : AOI21_X1 port map( B1 => n12, B2 => n17, A => OPCODE_IN(3), ZN => 
                           CW_OUT_12_port);
   U21 : INV_X1 port map( A => OPCODE_IN(0), ZN => n7);
   U25 : INV_X1 port map( A => OPCODE_IN(3), ZN => n6);
   U18 : NAND2_X1 port map( A1 => OPCODE_IN(0), A2 => n6, ZN => n10);
   U30 : INV_X1 port map( A => OPCODE_IN(5), ZN => n23);
   U29 : NAND2_X1 port map( A1 => n28, A2 => n23, ZN => n12);
   U10 : OR2_X1 port map( A1 => CW_OUT_7_port, A2 => n18, ZN => n9);
   U2 : OR3_X1 port map( A1 => n9, A2 => CW_OUT_4, A3 => CW_OUT_1, ZN => 
                           CW_OUT_0);
   U9 : OR2_X1 port map( A1 => CW_OUT_3, A2 => n9, ZN => CW_OUT_5_port);
   U6 : AND3_X1 port map( A1 => n23, A2 => n6, A3 => OPCODE_IN(1), ZN => n25);
   U7 : OR2_X1 port map( A1 => CW_OUT_12_port, A2 => n1, ZN => CW_OUT_9_port);
   U11 : NOR2_X1 port map( A1 => n19, A2 => OPCODE_IN(4), ZN => n28);
   U12 : INV_X1 port map( A => OPCODE_IN(2), ZN => n14);
   U13 : NAND2_X1 port map( A1 => OPCODE_IN(1), A2 => n14, ZN => n19);
   U14 : NOR3_X1 port map( A1 => OPCODE_IN(5), A2 => OPCODE_IN(1), A3 => 
                           OPCODE_IN(4), ZN => n13);
   U17 : NOR3_X1 port map( A1 => OPCODE_IN(5), A2 => n19, A3 => n10, ZN => 
                           CW_OUT_7_port);
   U24 : NOR2_X1 port map( A1 => n12, A2 => OPCODE_IN(3), ZN => CW_OUT_10_port)
                           ;
   U26 : NAND3_X1 port map( A1 => n13, A2 => OPCODE_IN(3), A3 => n14, ZN => n2)
                           ;
   U27 : AOI21_X1 port map( B1 => n12, B2 => n2, A => OPCODE_IN(0), ZN => n1);
   U28 : OAI211_X1 port map( C1 => n19, C2 => n20, A => n21, B => n22, ZN => 
                           n18);
   U31 : AOI21_X1 port map( B1 => n6, B2 => n27, A => OPCODE_IN(1), ZN => n26);
   U32 : OAI211_X1 port map( C1 => OPCODE_IN(4), C2 => OPCODE_IN(0), A => 
                           OPCODE_IN(1), B => OPCODE_IN(2), ZN => n24);
   U33 : OAI211_X1 port map( C1 => n25, C2 => n26, A => OPCODE_IN(2), B => 
                           OPCODE_IN(4), ZN => n21);
   U34 : NAND2_X1 port map( A1 => OPCODE_IN(2), A2 => n13, ZN => n17);

end SYN_bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity stall_logic_FUNC_SIZE11_OP_CODE_SIZE6 is

   port( OPCODE_i : in std_logic_vector (5 downto 0);  FUNC_i : in 
         std_logic_vector (10 downto 0);  rA_i, rB_i, D1_i, D2_i : in 
         std_logic_vector (4 downto 0);  S_mem_LOAD_i, S_exe_LOAD_i, 
         S_exe_WRITE_i : in std_logic;  S_MUX_PC_BUS_i : in std_logic_vector (1
         downto 0);  mispredict_i : in std_logic;  bubble_dec_o, bubble_exe_o, 
         stall_exe_o, stall_dec_o, stall_btb_o, stall_fetch_o : out std_logic);

end stall_logic_FUNC_SIZE11_OP_CODE_SIZE6;

architecture SYN_stall_logic_hw of stall_logic_FUNC_SIZE11_OP_CODE_SIZE6 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI33_X1
      port( A1, A2, A3, B1, B2, B3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal stall_fetch_o_port, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
      n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40
      , n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, 
      n55, n56, n57, n58 : std_logic;

begin
   stall_dec_o <= stall_fetch_o_port;
   stall_btb_o <= stall_fetch_o_port;
   stall_fetch_o <= stall_fetch_o_port;
   
   U46 : OAI33_X1 port map( A1 => OPCODE_i(2), A2 => n52, A3 => n53, B1 => n50,
                           B2 => OPCODE_i(4), B3 => OPCODE_i(1), ZN => n51);
   U43 : OAI22_X1 port map( A1 => n43, A2 => D2_i(3), B1 => n40, B2 => D2_i(1),
                           ZN => n58);
   U42 : AOI221_X1 port map( B1 => n43, B2 => D2_i(3), C1 => D2_i(1), C2 => n40
                           , A => n58, ZN => n54);
   U37 : XNOR2_X1 port map( A => rA_i(4), B => D2_i(4), ZN => n56);
   U36 : NAND4_X1 port map( A1 => S_mem_LOAD_i, A2 => n54, A3 => n55, A4 => n56
                           , ZN => n17);
   U35 : NOR2_X1 port map( A1 => OPCODE_i(5), A2 => OPCODE_i(3), ZN => n27);
   U31 : NAND2_X1 port map( A1 => n27, A2 => n51, ZN => n18);
   U30 : OAI21_X1 port map( B1 => OPCODE_i(0), B2 => n50, A => OPCODE_i(4), ZN 
                           => n48);
   U26 : AOI21_X1 port map( B1 => n27, B2 => n46, A => n47, ZN => n34);
   U23 : XNOR2_X1 port map( A => n31, B => rA_i(4), ZN => n37);
   U22 : AOI22_X1 port map( A1 => n43, A2 => D1_i(3), B1 => D1_i(2), B2 => n44,
                           ZN => n45);
   U21 : OAI221_X1 port map( B1 => n43, B2 => D1_i(3), C1 => n44, C2 => D1_i(2)
                           , A => n45, ZN => n38);
   U20 : AOI22_X1 port map( A1 => n40, A2 => D1_i(1), B1 => D1_i(0), B2 => n41,
                           ZN => n42);
   U19 : OAI221_X1 port map( B1 => n40, B2 => D1_i(1), C1 => n41, C2 => D1_i(0)
                           , A => n42, ZN => n39);
   U18 : NOR3_X1 port map( A1 => n37, A2 => n38, A3 => n39, ZN => n36);
   U17 : OAI221_X1 port map( B1 => n34, B2 => n35, C1 => n34, C2 => 
                           S_exe_WRITE_i, A => n36, ZN => n19);
   U15 : OAI22_X1 port map( A1 => n31, A2 => rB_i(4), B1 => n32, B2 => rB_i(2),
                           ZN => n33);
   U14 : AOI221_X1 port map( B1 => n31, B2 => rB_i(4), C1 => rB_i(2), C2 => n32
                           , A => n33, ZN => n21);
   U11 : OAI22_X1 port map( A1 => n28, A2 => rB_i(0), B1 => n29, B2 => rB_i(3),
                           ZN => n30);
   U10 : AOI221_X1 port map( B1 => n28, B2 => rB_i(0), C1 => rB_i(3), C2 => n29
                           , A => n30, ZN => n22);
   U7 : OAI211_X1 port map( C1 => n25, C2 => rB_i(1), A => S_exe_LOAD_i, B => 
                           n27, ZN => n26);
   U6 : AOI21_X1 port map( B1 => n25, B2 => rB_i(1), A => n26, ZN => n24);
   U5 : NAND4_X1 port map( A1 => n21, A2 => n22, A3 => n23, A4 => n24, ZN => 
                           n20);
   U2 : NOR2_X1 port map( A1 => stall_fetch_o_port, A2 => n16, ZN => 
                           bubble_dec_o);
   U40 : INV_X1 port map( A => rA_i(2), ZN => n44);
   U41 : INV_X1 port map( A => rA_i(0), ZN => n41);
   U34 : INV_X1 port map( A => OPCODE_i(4), ZN => n52);
   U45 : INV_X1 port map( A => rA_i(3), ZN => n43);
   U44 : INV_X1 port map( A => rA_i(1), ZN => n40);
   U27 : INV_X1 port map( A => S_exe_LOAD_i, ZN => n47);
   U25 : INV_X1 port map( A => n18, ZN => n35);
   U16 : INV_X1 port map( A => D1_i(2), ZN => n32);
   U13 : INV_X1 port map( A => D1_i(0), ZN => n28);
   U12 : INV_X1 port map( A => D1_i(3), ZN => n29);
   U8 : INV_X1 port map( A => D1_i(1), ZN => n25);
   U24 : INV_X1 port map( A => D1_i(4), ZN => n31);
   U4 : OAI211_X1 port map( C1 => n17, C2 => n18, A => n19, B => n20, ZN => 
                           stall_fetch_o_port);
   U3 : INV_X1 port map( A => mispredict_i, ZN => n16);
   U9 : INV_X1 port map( A => OPCODE_i(1), ZN => n53);
   U28 : AOI221_X1 port map( B1 => n41, B2 => D2_i(0), C1 => D2_i(2), C2 => n44
                           , A => n57, ZN => n55);
   U29 : OAI22_X1 port map( A1 => n41, A2 => D2_i(0), B1 => n44, B2 => D2_i(2),
                           ZN => n57);
   U32 : OAI22_X1 port map( A1 => OPCODE_i(1), A2 => n48, B1 => OPCODE_i(4), B2
                           => n49, ZN => n46);
   U33 : NAND2_X1 port map( A1 => OPCODE_i(1), A2 => n50, ZN => n49);
   U38 : NOR4_X1 port map( A1 => OPCODE_i(2), A2 => OPCODE_i(4), A3 => 
                           OPCODE_i(1), A4 => OPCODE_i(0), ZN => n23);
   U39 : INV_X1 port map( A => OPCODE_i(2), ZN => n50);

end SYN_stall_logic_hw;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity mux41_MUX_SIZE32_0 is

   port( IN0, IN1, IN2, IN3 : in std_logic_vector (31 downto 0);  CTRL : in 
         std_logic_vector (1 downto 0);  OUT1 : out std_logic_vector (31 downto
         0));

end mux41_MUX_SIZE32_0;

architecture SYN_bhe of mux41_MUX_SIZE32_0 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n6, n7, n8, n11, n12, n15, n16, n17, n18, n19, n20, n43, n44, n45, 
      n46, n59, n60, n63, n64, n67, n68, n71, n1, n2, n3, n4, n5, n9, n10, n13,
      n14, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34
      , n35, n36, n37, n38, n39, n40, n41, n42, n47, n48, n49, n50, n51, n52, 
      n53, n54, n55, n56, n57, n58, n61, n62, n65, n66, n69, n70, n72, n73, n74
      , n75, n76, n77, n78, n79 : std_logic;

begin
   
   U57 : AOI22_X1 port map( A1 => n76, A2 => IN1(21), B1 => n75, B2 => IN0(21),
                           ZN => n43);
   U55 : NAND2_X1 port map( A1 => n43, A2 => n44, ZN => OUT1(21));
   U60 : AOI22_X1 port map( A1 => n76, A2 => IN1(20), B1 => n75, B2 => IN0(20),
                           ZN => n45);
   U58 : NAND2_X1 port map( A1 => n45, A2 => n46, ZN => OUT1(20));
   U81 : AOI22_X1 port map( A1 => n7, A2 => IN1(14), B1 => n74, B2 => IN0(14), 
                           ZN => n59);
   U79 : NAND2_X1 port map( A1 => n59, A2 => n60, ZN => OUT1(14));
   U93 : AOI22_X1 port map( A1 => n7, A2 => IN1(10), B1 => n74, B2 => IN0(10), 
                           ZN => n67);
   U91 : NAND2_X1 port map( A1 => n67, A2 => n68, ZN => OUT1(10));
   U87 : AOI22_X1 port map( A1 => n7, A2 => IN1(12), B1 => n74, B2 => IN0(12), 
                           ZN => n63);
   U85 : NAND2_X1 port map( A1 => n63, A2 => n64, ZN => OUT1(12));
   U7 : NAND2_X1 port map( A1 => n11, A2 => n12, ZN => OUT1(7));
   U19 : NAND2_X1 port map( A1 => n19, A2 => n20, ZN => OUT1(3));
   U13 : NAND2_X1 port map( A1 => n15, A2 => n16, ZN => OUT1(5));
   U16 : NAND2_X1 port map( A1 => n17, A2 => n18, ZN => OUT1(4));
   U100 : AND2_X1 port map( A1 => n71, A2 => CTRL(0), ZN => n7);
   U1 : AOI222_X1 port map( A1 => n7, A2 => IN1(0), B1 => n74, B2 => IN0(0), C1
                           => IN2(0), C2 => n6, ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => OUT1(0));
   U3 : AOI22_X1 port map( A1 => IN1(2), A2 => n76, B1 => IN0(2), B2 => n75, ZN
                           => n2);
   U4 : NAND2_X1 port map( A1 => n56, A2 => n2, ZN => OUT1(2));
   U5 : AOI222_X1 port map( A1 => n77, A2 => IN1(6), B1 => n8, B2 => IN0(6), C1
                           => IN2(6), C2 => n6, ZN => n3);
   U6 : INV_X1 port map( A => n3, ZN => OUT1(6));
   U8 : AOI222_X1 port map( A1 => n77, A2 => IN1(13), B1 => n74, B2 => IN0(13),
                           C1 => IN2(13), C2 => n6, ZN => n4);
   U9 : INV_X1 port map( A => n4, ZN => OUT1(13));
   U10 : AOI22_X1 port map( A1 => IN1(27), A2 => n76, B1 => IN0(27), B2 => n75,
                           ZN => n5);
   U11 : NAND2_X1 port map( A1 => n62, A2 => n5, ZN => OUT1(27));
   U12 : BUF_X1 port map( A => n6, Z => n79);
   U14 : BUF_X1 port map( A => n8, Z => n75);
   U15 : BUF_X1 port map( A => n8, Z => n74);
   U17 : BUF_X2 port map( A => n7, Z => n77);
   U18 : BUF_X2 port map( A => n7, Z => n76);
   U20 : INV_X1 port map( A => CTRL(1), ZN => n71);
   U21 : BUF_X2 port map( A => n6, Z => n78);
   U22 : NOR2_X1 port map( A1 => n71, A2 => CTRL(0), ZN => n6);
   U23 : NOR2_X2 port map( A1 => CTRL(0), A2 => CTRL(1), ZN => n8);
   U24 : NAND2_X1 port map( A1 => n78, A2 => IN2(4), ZN => n18);
   U25 : NAND2_X1 port map( A1 => n78, A2 => IN2(5), ZN => n16);
   U26 : NAND2_X1 port map( A1 => n78, A2 => IN2(3), ZN => n20);
   U27 : NAND2_X1 port map( A1 => n75, A2 => IN0(28), ZN => n34);
   U28 : NAND2_X1 port map( A1 => n75, A2 => IN0(29), ZN => n27);
   U29 : NAND2_X1 port map( A1 => n78, A2 => IN2(7), ZN => n12);
   U30 : NAND2_X1 port map( A1 => n78, A2 => IN2(12), ZN => n64);
   U31 : NAND2_X1 port map( A1 => n78, A2 => IN2(10), ZN => n68);
   U32 : NAND2_X1 port map( A1 => n78, A2 => IN2(14), ZN => n60);
   U33 : NAND2_X1 port map( A1 => n74, A2 => IN0(19), ZN => n72);
   U34 : NAND2_X1 port map( A1 => n74, A2 => IN0(1), ZN => n58);
   U35 : NAND2_X1 port map( A1 => n78, A2 => IN2(20), ZN => n46);
   U36 : NAND2_X1 port map( A1 => n78, A2 => IN2(21), ZN => n44);
   U37 : AOI22_X1 port map( A1 => n77, A2 => IN1(31), B1 => n8, B2 => IN0(31), 
                           ZN => n10);
   U38 : NAND2_X1 port map( A1 => n9, A2 => n10, ZN => OUT1(31));
   U39 : NAND2_X1 port map( A1 => n78, A2 => IN2(31), ZN => n9);
   U40 : AOI22_X1 port map( A1 => n77, A2 => IN1(8), B1 => n8, B2 => IN0(8), ZN
                           => n14);
   U41 : NAND2_X1 port map( A1 => n13, A2 => n14, ZN => OUT1(8));
   U42 : NAND2_X1 port map( A1 => n78, A2 => IN2(8), ZN => n13);
   U43 : AOI22_X1 port map( A1 => n7, A2 => IN1(11), B1 => n74, B2 => IN0(11), 
                           ZN => n22);
   U44 : NAND2_X1 port map( A1 => n21, A2 => n22, ZN => OUT1(11));
   U45 : NAND2_X1 port map( A1 => n78, A2 => IN2(11), ZN => n21);
   U46 : AOI22_X1 port map( A1 => n7, A2 => IN1(18), B1 => n74, B2 => IN0(18), 
                           ZN => n24);
   U47 : NAND2_X1 port map( A1 => n23, A2 => n24, ZN => OUT1(18));
   U48 : NAND2_X1 port map( A1 => n78, A2 => IN2(18), ZN => n23);
   U49 : NAND3_X1 port map( A1 => n25, A2 => n26, A3 => n27, ZN => OUT1(29));
   U50 : NAND2_X1 port map( A1 => n79, A2 => IN2(29), ZN => n25);
   U51 : NAND2_X1 port map( A1 => n76, A2 => IN1(29), ZN => n26);
   U52 : AOI22_X1 port map( A1 => n77, A2 => IN1(16), B1 => n74, B2 => IN0(16),
                           ZN => n29);
   U53 : NAND2_X1 port map( A1 => n28, A2 => n29, ZN => OUT1(16));
   U54 : NAND2_X1 port map( A1 => n78, A2 => IN2(16), ZN => n28);
   U56 : NAND2_X1 port map( A1 => n78, A2 => IN2(9), ZN => n30);
   U59 : NAND2_X1 port map( A1 => n31, A2 => n30, ZN => OUT1(9));
   U61 : AOI22_X1 port map( A1 => n77, A2 => IN1(9), B1 => n75, B2 => IN0(9), 
                           ZN => n31);
   U62 : NAND3_X1 port map( A1 => n32, A2 => n33, A3 => n34, ZN => OUT1(28));
   U63 : NAND2_X1 port map( A1 => n79, A2 => IN2(28), ZN => n32);
   U64 : NAND2_X1 port map( A1 => n76, A2 => IN1(28), ZN => n33);
   U65 : AOI22_X1 port map( A1 => n7, A2 => IN1(17), B1 => n74, B2 => IN0(17), 
                           ZN => n36);
   U66 : NAND2_X1 port map( A1 => n35, A2 => n36, ZN => OUT1(17));
   U67 : NAND2_X1 port map( A1 => n79, A2 => IN2(17), ZN => n35);
   U68 : NAND3_X1 port map( A1 => n38, A2 => n37, A3 => n39, ZN => OUT1(25));
   U69 : NAND2_X1 port map( A1 => n76, A2 => IN1(25), ZN => n38);
   U70 : NAND2_X1 port map( A1 => n79, A2 => IN2(25), ZN => n37);
   U71 : NAND2_X1 port map( A1 => n75, A2 => IN0(25), ZN => n39);
   U72 : NAND2_X1 port map( A1 => n78, A2 => IN2(15), ZN => n40);
   U73 : NAND2_X1 port map( A1 => n41, A2 => n40, ZN => OUT1(15));
   U74 : AOI22_X1 port map( A1 => n77, A2 => IN1(15), B1 => n74, B2 => IN0(15),
                           ZN => n41);
   U75 : NAND3_X1 port map( A1 => n47, A2 => n42, A3 => n48, ZN => OUT1(24));
   U76 : NAND2_X1 port map( A1 => n76, A2 => IN1(24), ZN => n47);
   U77 : NAND2_X1 port map( A1 => n79, A2 => IN2(24), ZN => n42);
   U78 : NAND2_X1 port map( A1 => n75, A2 => IN0(24), ZN => n48);
   U80 : NAND2_X1 port map( A1 => n78, A2 => IN2(23), ZN => n49);
   U82 : NAND2_X1 port map( A1 => n49, A2 => n50, ZN => OUT1(23));
   U83 : AOI22_X1 port map( A1 => n76, A2 => IN1(23), B1 => n75, B2 => IN0(23),
                           ZN => n50);
   U84 : NAND3_X1 port map( A1 => n52, A2 => n51, A3 => n53, ZN => OUT1(30));
   U86 : NAND2_X1 port map( A1 => n79, A2 => IN2(30), ZN => n52);
   U88 : NAND2_X1 port map( A1 => n76, A2 => IN1(30), ZN => n51);
   U89 : NAND2_X1 port map( A1 => n75, A2 => IN0(30), ZN => n53);
   U90 : NAND2_X1 port map( A1 => n78, A2 => IN2(22), ZN => n54);
   U92 : NAND2_X1 port map( A1 => n54, A2 => n55, ZN => OUT1(22));
   U94 : AOI22_X1 port map( A1 => n76, A2 => IN1(22), B1 => n75, B2 => IN0(22),
                           ZN => n55);
   U95 : NAND2_X1 port map( A1 => n79, A2 => IN2(2), ZN => n56);
   U96 : NAND3_X1 port map( A1 => n57, A2 => n58, A3 => n61, ZN => OUT1(1));
   U97 : NAND2_X1 port map( A1 => n79, A2 => IN2(1), ZN => n57);
   U98 : NAND2_X1 port map( A1 => n76, A2 => IN1(1), ZN => n61);
   U99 : NAND2_X1 port map( A1 => n79, A2 => IN2(27), ZN => n62);
   U101 : NAND3_X1 port map( A1 => n66, A2 => n65, A3 => n69, ZN => OUT1(26));
   U102 : NAND2_X1 port map( A1 => n79, A2 => IN2(26), ZN => n66);
   U103 : NAND2_X1 port map( A1 => n76, A2 => IN1(26), ZN => n65);
   U104 : NAND2_X1 port map( A1 => n75, A2 => IN0(26), ZN => n69);
   U105 : NAND3_X1 port map( A1 => n70, A2 => n72, A3 => n73, ZN => OUT1(19));
   U106 : NAND2_X1 port map( A1 => n79, A2 => IN2(19), ZN => n70);
   U107 : NAND2_X1 port map( A1 => n77, A2 => IN1(19), ZN => n73);
   U108 : AOI22_X1 port map( A1 => n77, A2 => IN1(5), B1 => n8, B2 => IN0(5), 
                           ZN => n15);
   U109 : AOI22_X1 port map( A1 => n77, A2 => IN1(4), B1 => n74, B2 => IN0(4), 
                           ZN => n17);
   U110 : AOI22_X1 port map( A1 => n77, A2 => IN1(3), B1 => n8, B2 => IN0(3), 
                           ZN => n19);
   U111 : AOI22_X1 port map( A1 => n77, A2 => IN1(7), B1 => n8, B2 => IN0(7), 
                           ZN => n11);

end SYN_bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity zerocheck is

   port( IN0 : in std_logic_vector (31 downto 0);  CTRL : in std_logic;  OUT1 :
         out std_logic);

end zerocheck;

architecture SYN_Bhe of zerocheck is

   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25 : std_logic;

begin
   
   U1 : INV_X1 port map( A => IN0(28), ZN => n14);
   U2 : INV_X1 port map( A => IN0(29), ZN => n13);
   U3 : INV_X1 port map( A => IN0(21), ZN => n24);
   U4 : INV_X1 port map( A => IN0(20), ZN => n25);
   U5 : INV_X1 port map( A => IN0(24), ZN => n11);
   U6 : INV_X1 port map( A => IN0(18), ZN => n21);
   U7 : INV_X1 port map( A => IN0(17), ZN => n22);
   U8 : INV_X1 port map( A => IN0(25), ZN => n10);
   U9 : XNOR2_X1 port map( A => n1, B => CTRL, ZN => OUT1);
   U10 : NOR2_X1 port map( A1 => n2, A2 => n3, ZN => n1);
   U11 : NOR4_X1 port map( A1 => IN0(7), A2 => IN0(6), A3 => IN0(8), A4 => 
                           IN0(9), ZN => n4);
   U12 : NOR4_X1 port map( A1 => IN0(14), A2 => IN0(13), A3 => IN0(16), A4 => 
                           IN0(15), ZN => n16);
   U13 : NAND3_X1 port map( A1 => n4, A2 => n6, A3 => n5, ZN => n3);
   U14 : NAND3_X1 port map( A1 => n9, A2 => n10, A3 => n11, ZN => n8);
   U15 : NAND3_X1 port map( A1 => n12, A2 => n13, A3 => n14, ZN => n7);
   U16 : NAND3_X1 port map( A1 => n15, A2 => n16, A3 => n17, ZN => n2);
   U17 : NAND3_X1 port map( A1 => n20, A2 => n21, A3 => n22, ZN => n19);
   U18 : NAND3_X1 port map( A1 => n23, A2 => n24, A3 => n25, ZN => n18);
   U19 : NOR2_X1 port map( A1 => IN0(23), A2 => IN0(22), ZN => n23);
   U20 : NOR2_X1 port map( A1 => n18, A2 => n19, ZN => n15);
   U21 : NOR2_X1 port map( A1 => IN0(1), A2 => IN0(19), ZN => n20);
   U22 : NOR2_X1 port map( A1 => IN0(30), A2 => IN0(2), ZN => n12);
   U23 : NOR2_X1 port map( A1 => n7, A2 => n8, ZN => n6);
   U24 : NOR2_X1 port map( A1 => IN0(27), A2 => IN0(26), ZN => n9);
   U25 : NOR4_X1 port map( A1 => IN0(10), A2 => IN0(0), A3 => IN0(12), A4 => 
                           IN0(11), ZN => n17);
   U26 : NOR4_X1 port map( A1 => IN0(3), A2 => IN0(5), A3 => IN0(4), A4 => 
                           IN0(31), ZN => n5);

end SYN_Bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity mux21_0 is

   port( IN0, IN1 : in std_logic_vector (31 downto 0);  CTRL : in std_logic;  
         OUT1 : out std_logic_vector (31 downto 0));

end mux21_0;

architecture SYN_Bhe of mux21_0 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X4
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15 : 
      std_logic;

begin
   
   U14 : MUX2_X1 port map( A => IN0(26), B => IN1(26), S => n14, Z => OUT1(26))
                           ;
   U18 : MUX2_X1 port map( A => IN0(22), B => IN1(22), S => n14, Z => OUT1(22))
                           ;
   U20 : MUX2_X1 port map( A => IN0(20), B => IN1(20), S => n14, Z => OUT1(20))
                           ;
   U21 : MUX2_X1 port map( A => IN0(1), B => IN1(1), S => n14, Z => OUT1(1));
   U23 : MUX2_X1 port map( A => IN0(18), B => IN1(18), S => n14, Z => OUT1(18))
                           ;
   U24 : MUX2_X1 port map( A => IN0(17), B => IN1(17), S => n14, Z => OUT1(17))
                           ;
   U25 : MUX2_X1 port map( A => IN0(16), B => IN1(16), S => n15, Z => OUT1(16))
                           ;
   U27 : MUX2_X1 port map( A => IN0(14), B => IN1(14), S => n15, Z => OUT1(14))
                           ;
   U28 : MUX2_X1 port map( A => IN0(13), B => IN1(13), S => n15, Z => OUT1(13))
                           ;
   U29 : MUX2_X1 port map( A => IN0(12), B => IN1(12), S => n15, Z => OUT1(12))
                           ;
   U30 : MUX2_X1 port map( A => IN0(11), B => IN1(11), S => n15, Z => OUT1(11))
                           ;
   U31 : MUX2_X1 port map( A => IN0(10), B => IN1(10), S => n15, Z => OUT1(10))
                           ;
   U32 : MUX2_X1 port map( A => IN0(0), B => IN1(0), S => n15, Z => OUT1(0));
   U26 : MUX2_X1 port map( A => IN0(15), B => IN1(15), S => n15, Z => OUT1(15))
                           ;
   U22 : MUX2_X1 port map( A => IN0(19), B => IN1(19), S => n14, Z => OUT1(19))
                           ;
   U15 : MUX2_X1 port map( A => IN0(25), B => IN1(25), S => n14, Z => OUT1(25))
                           ;
   U1 : MUX2_X1 port map( A => IN0(9), B => IN1(9), S => n15, Z => OUT1(9));
   U3 : MUX2_X1 port map( A => IN0(7), B => IN1(7), S => n14, Z => OUT1(7));
   U5 : MUX2_X1 port map( A => IN0(5), B => IN1(5), S => n14, Z => OUT1(5));
   U7 : MUX2_X1 port map( A => IN0(3), B => IN1(3), S => n14, Z => OUT1(3));
   U10 : MUX2_X1 port map( A => IN0(2), B => IN1(2), S => n15, Z => OUT1(2));
   U12 : MUX2_X1 port map( A => IN0(28), B => IN1(28), S => n14, Z => OUT1(28))
                           ;
   U6 : MUX2_X1 port map( A => IN0(4), B => IN1(4), S => n14, Z => OUT1(4));
   U2 : MUX2_X1 port map( A => IN0(8), B => IN1(8), S => n15, Z => OUT1(8));
   U4 : MUX2_X1 port map( A => IN0(21), B => IN1(21), S => n14, Z => OUT1(21));
   U8 : INV_X1 port map( A => IN0(6), ZN => n6);
   U9 : BUF_X2 port map( A => CTRL, Z => n15);
   U11 : MUX2_X1 port map( A => IN0(29), B => IN1(29), S => n15, Z => OUT1(29))
                           ;
   U13 : INV_X1 port map( A => n14, ZN => n11);
   U16 : BUF_X4 port map( A => CTRL, Z => n14);
   U17 : NAND2_X1 port map( A1 => n14, A2 => IN1(30), ZN => n5);
   U19 : NAND2_X1 port map( A1 => n15, A2 => IN1(31), ZN => n8);
   U33 : NAND2_X1 port map( A1 => n14, A2 => IN1(27), ZN => n3);
   U34 : NAND2_X1 port map( A1 => n14, A2 => IN1(24), ZN => n10);
   U35 : OAI21_X1 port map( B1 => n14, B2 => n6, A => n1, ZN => OUT1(6));
   U36 : NAND2_X1 port map( A1 => n15, A2 => IN1(6), ZN => n1);
   U37 : NAND2_X1 port map( A1 => IN0(27), A2 => n11, ZN => n2);
   U38 : NAND2_X1 port map( A1 => n2, A2 => n3, ZN => OUT1(27));
   U39 : NAND2_X1 port map( A1 => IN0(30), A2 => n11, ZN => n4);
   U40 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => OUT1(30));
   U41 : NAND2_X1 port map( A1 => IN0(31), A2 => n11, ZN => n7);
   U42 : NAND2_X1 port map( A1 => n7, A2 => n8, ZN => OUT1(31));
   U43 : NAND2_X1 port map( A1 => IN0(24), A2 => n11, ZN => n9);
   U44 : NAND2_X1 port map( A1 => n9, A2 => n10, ZN => OUT1(24));
   U45 : NAND2_X1 port map( A1 => IN0(23), A2 => n11, ZN => n12);
   U46 : NAND2_X1 port map( A1 => n14, A2 => IN1(23), ZN => n13);
   U47 : NAND2_X1 port map( A1 => n12, A2 => n13, ZN => OUT1(23));

end SYN_Bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity p4add_N32_logN5_0 is

   port( A, B : in std_logic_vector (31 downto 0);  Cin, sign : in std_logic;  
         S : out std_logic_vector (31 downto 0);  Cout : out std_logic);

end p4add_N32_logN5_0;

architecture SYN_STRUCTURAL of p4add_N32_logN5_0 is

   component sum_gen_N32_0
      port( A, B : in std_logic_vector (31 downto 0);  Cin : in 
            std_logic_vector (8 downto 0);  S : out std_logic_vector (31 downto
            0));
   end component;
   
   component carry_tree_N32_logN5_0
      port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  
            Cout : out std_logic_vector (7 downto 0));
   end component;
   
   component xor_gen_N32_0
      port( A : in std_logic_vector (31 downto 0);  B : in std_logic;  S : out 
            std_logic_vector (31 downto 0));
   end component;
   
   signal n17, new_B_31_port, new_B_30_port, new_B_28_port, new_B_26_port, 
      new_B_24_port, new_B_23_port, new_B_22_port, new_B_21_port, new_B_20_port
      , new_B_19_port, new_B_18_port, new_B_17_port, new_B_16_port, 
      new_B_15_port, new_B_14_port, new_B_13_port, new_B_12_port, new_B_11_port
      , new_B_10_port, new_B_9_port, new_B_8_port, new_B_7_port, new_B_6_port, 
      new_B_5_port, new_B_4_port, new_B_3_port, new_B_2_port, new_B_1_port, 
      new_B_0_port, carry_pro_7_port, carry_pro_6_port, carry_pro_5_port, 
      carry_pro_4_port, carry_pro_3_port, carry_pro_2_port, carry_pro_1_port, 
      n1, n3, n5, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, net246124 : 
      std_logic;

begin
   
   xor32 : xor_gen_N32_0 port map( A(31) => B(31), A(30) => B(30), A(29) => 
                           B(29), A(28) => B(28), A(27) => B(27), A(26) => 
                           B(26), A(25) => B(25), A(24) => B(24), A(23) => 
                           B(23), A(22) => B(22), A(21) => B(21), A(20) => 
                           B(20), A(19) => B(19), A(18) => B(18), A(17) => 
                           B(17), A(16) => B(16), A(15) => B(15), A(14) => 
                           B(14), A(13) => B(13), A(12) => B(12), A(11) => 
                           B(11), A(10) => B(10), A(9) => B(9), A(8) => B(8), 
                           A(7) => B(7), A(6) => B(6), A(5) => B(5), A(4) => 
                           B(4), A(3) => B(3), A(2) => B(2), A(1) => B(1), A(0)
                           => B(0), B => n17, S(31) => new_B_31_port, S(30) => 
                           new_B_30_port, S(29) => n5, S(28) => new_B_28_port, 
                           S(27) => n3, S(26) => new_B_26_port, S(25) => n1, 
                           S(24) => new_B_24_port, S(23) => new_B_23_port, 
                           S(22) => new_B_22_port, S(21) => new_B_21_port, 
                           S(20) => new_B_20_port, S(19) => new_B_19_port, 
                           S(18) => new_B_18_port, S(17) => new_B_17_port, 
                           S(16) => new_B_16_port, S(15) => new_B_15_port, 
                           S(14) => new_B_14_port, S(13) => new_B_13_port, 
                           S(12) => new_B_12_port, S(11) => new_B_11_port, 
                           S(10) => new_B_10_port, S(9) => new_B_9_port, S(8) 
                           => new_B_8_port, S(7) => new_B_7_port, S(6) => 
                           new_B_6_port, S(5) => new_B_5_port, S(4) => 
                           new_B_4_port, S(3) => new_B_3_port, S(2) => 
                           new_B_2_port, S(1) => new_B_1_port, S(0) => 
                           new_B_0_port);
   ct : carry_tree_N32_logN5_0 port map( A(31) => n8, A(30) => n9, A(29) => n10
                           , A(28) => n11, A(27) => A(27), A(26) => A(26), 
                           A(25) => A(25), A(24) => A(24), A(23) => A(23), 
                           A(22) => A(22), A(21) => A(21), A(20) => A(20), 
                           A(19) => A(19), A(18) => A(18), A(17) => A(17), 
                           A(16) => A(16), A(15) => A(15), A(14) => A(14), 
                           A(13) => A(13), A(12) => A(12), A(11) => A(11), 
                           A(10) => A(10), A(9) => A(9), A(8) => A(8), A(7) => 
                           A(7), A(6) => A(6), A(5) => A(5), A(4) => A(4), A(3)
                           => A(3), A(2) => A(2), A(1) => A(1), A(0) => A(0), 
                           B(31) => n12, B(30) => n13, B(29) => n14, B(28) => 
                           n15, B(27) => new_B_31_port, B(26) => new_B_26_port,
                           B(25) => n1, B(24) => new_B_24_port, B(23) => 
                           new_B_23_port, B(22) => new_B_22_port, B(21) => 
                           new_B_21_port, B(20) => new_B_20_port, B(19) => 
                           new_B_19_port, B(18) => new_B_18_port, B(17) => 
                           new_B_17_port, B(16) => new_B_16_port, B(15) => 
                           new_B_15_port, B(14) => new_B_14_port, B(13) => 
                           new_B_13_port, B(12) => new_B_12_port, B(11) => 
                           new_B_11_port, B(10) => new_B_10_port, B(9) => 
                           new_B_9_port, B(8) => new_B_8_port, B(7) => 
                           new_B_7_port, B(6) => new_B_6_port, B(5) => 
                           new_B_5_port, B(4) => new_B_4_port, B(3) => 
                           new_B_3_port, B(2) => new_B_2_port, B(1) => 
                           new_B_1_port, B(0) => new_B_0_port, Cin => n7, 
                           Cout(7) => net246124, Cout(6) => carry_pro_7_port, 
                           Cout(5) => carry_pro_6_port, Cout(4) => 
                           carry_pro_5_port, Cout(3) => carry_pro_4_port, 
                           Cout(2) => carry_pro_3_port, Cout(1) => 
                           carry_pro_2_port, Cout(0) => carry_pro_1_port);
   add : sum_gen_N32_0 port map( A(31) => A(31), A(30) => A(30), A(29) => A(29)
                           , A(28) => A(28), A(27) => A(27), A(26) => A(26), 
                           A(25) => A(25), A(24) => A(24), A(23) => A(23), 
                           A(22) => A(22), A(21) => A(21), A(20) => A(20), 
                           A(19) => A(19), A(18) => A(18), A(17) => A(17), 
                           A(16) => A(16), A(15) => A(15), A(14) => A(14), 
                           A(13) => A(13), A(12) => A(12), A(11) => A(11), 
                           A(10) => A(10), A(9) => A(9), A(8) => A(8), A(7) => 
                           A(7), A(6) => A(6), A(5) => A(5), A(4) => A(4), A(3)
                           => A(3), A(2) => A(2), A(1) => A(1), A(0) => A(0), 
                           B(31) => new_B_31_port, B(30) => new_B_30_port, 
                           B(29) => n5, B(28) => new_B_28_port, B(27) => n3, 
                           B(26) => new_B_26_port, B(25) => n1, B(24) => 
                           new_B_24_port, B(23) => new_B_23_port, B(22) => 
                           new_B_22_port, B(21) => new_B_21_port, B(20) => 
                           new_B_20_port, B(19) => new_B_19_port, B(18) => 
                           new_B_18_port, B(17) => new_B_17_port, B(16) => 
                           new_B_16_port, B(15) => new_B_15_port, B(14) => 
                           new_B_14_port, B(13) => new_B_13_port, B(12) => 
                           new_B_12_port, B(11) => new_B_11_port, B(10) => 
                           new_B_10_port, B(9) => new_B_9_port, B(8) => 
                           new_B_8_port, B(7) => new_B_7_port, B(6) => 
                           new_B_6_port, B(5) => new_B_5_port, B(4) => 
                           new_B_4_port, B(3) => new_B_3_port, B(2) => 
                           new_B_2_port, B(1) => new_B_1_port, B(0) => 
                           new_B_0_port, Cin(8) => n16, Cin(7) => 
                           carry_pro_7_port, Cin(6) => carry_pro_6_port, Cin(5)
                           => carry_pro_5_port, Cin(4) => carry_pro_4_port, 
                           Cin(3) => carry_pro_3_port, Cin(2) => 
                           carry_pro_2_port, Cin(1) => carry_pro_1_port, Cin(0)
                           => n7, S(31) => S(31), S(30) => S(30), S(29) => 
                           S(29), S(28) => S(28), S(27) => S(27), S(26) => 
                           S(26), S(25) => S(25), S(24) => S(24), S(23) => 
                           S(23), S(22) => S(22), S(21) => S(21), S(20) => 
                           S(20), S(19) => S(19), S(18) => S(18), S(17) => 
                           S(17), S(16) => S(16), S(15) => S(15), S(14) => 
                           S(14), S(13) => S(13), S(12) => S(12), S(11) => 
                           S(11), S(10) => S(10), S(9) => S(9), S(8) => S(8), 
                           S(7) => S(7), S(6) => S(6), S(5) => S(5), S(4) => 
                           S(4), S(3) => S(3), S(2) => S(2), S(1) => S(1), S(0)
                           => S(0));
   n7 <= '0';
   n17 <= '0';
   n8 <= '0';
   n9 <= '0';
   n10 <= '0';
   n11 <= '0';
   n12 <= '0';
   n13 <= '0';
   n14 <= '0';
   n15 <= '0';
   n16 <= '0';

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity extender_32 is

   port( IN1 : in std_logic_vector (31 downto 0);  CTRL, SIGN : in std_logic;  
         OUT1 : out std_logic_vector (31 downto 0));

end extender_32;

architecture SYN_Bhe of extender_32 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X4
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n15, OUT1_24_port, OUT1_23_port, OUT1_22_port, OUT1_21_port, 
      OUT1_20_port, OUT1_19_port, OUT1_18_port, OUT1_17_port, OUT1_16_port, n3,
      n5, n6, n7, n9, n10, n11, n12, n13, n4, n14, n8, OUT1_29_port, 
      OUT1_31_port : std_logic;

begin
   OUT1 <= ( OUT1_31_port, OUT1_29_port, OUT1_29_port, OUT1_31_port, 
      OUT1_29_port, OUT1_31_port, OUT1_29_port, OUT1_24_port, OUT1_23_port, 
      OUT1_22_port, OUT1_21_port, OUT1_20_port, OUT1_19_port, OUT1_18_port, 
      OUT1_17_port, OUT1_16_port, IN1(15), IN1(14), IN1(13), IN1(12), IN1(11), 
      IN1(10), IN1(9), IN1(8), IN1(7), IN1(6), IN1(5), IN1(4), IN1(3), IN1(2), 
      IN1(1), IN1(0) );
   
   U2 : BUF_X4 port map( A => n15, Z => OUT1_29_port);
   U3 : NAND2_X2 port map( A1 => n3, A2 => n12, ZN => OUT1_17_port);
   U4 : NAND2_X1 port map( A1 => n3, A2 => n10, ZN => OUT1_19_port);
   U5 : INV_X1 port map( A => CTRL, ZN => n14);
   U6 : BUF_X2 port map( A => n15, Z => OUT1_31_port);
   U7 : NAND2_X1 port map( A1 => n3, A2 => n4, ZN => n15);
   U8 : NAND3_X2 port map( A1 => SIGN, A2 => IN1(15), A3 => n14, ZN => n3);
   U9 : NAND2_X1 port map( A1 => CTRL, A2 => IN1(21), ZN => n8);
   U10 : NAND2_X1 port map( A1 => n3, A2 => n8, ZN => OUT1_21_port);
   U11 : NAND2_X1 port map( A1 => CTRL, A2 => IN1(25), ZN => n4);
   U12 : NAND2_X1 port map( A1 => CTRL, A2 => IN1(20), ZN => n9);
   U13 : NAND2_X1 port map( A1 => CTRL, A2 => IN1(24), ZN => n5);
   U14 : NAND2_X1 port map( A1 => CTRL, A2 => IN1(16), ZN => n13);
   U15 : NAND2_X1 port map( A1 => CTRL, A2 => IN1(17), ZN => n12);
   U16 : NAND2_X1 port map( A1 => CTRL, A2 => IN1(22), ZN => n7);
   U17 : NAND2_X1 port map( A1 => CTRL, A2 => IN1(23), ZN => n6);
   U18 : NAND2_X1 port map( A1 => CTRL, A2 => IN1(18), ZN => n11);
   U19 : NAND2_X1 port map( A1 => CTRL, A2 => IN1(19), ZN => n10);
   U20 : NAND2_X1 port map( A1 => n3, A2 => n5, ZN => OUT1_24_port);
   U21 : NAND2_X1 port map( A1 => n3, A2 => n13, ZN => OUT1_16_port);
   U22 : NAND2_X1 port map( A1 => n3, A2 => n9, ZN => OUT1_20_port);
   U23 : NAND2_X1 port map( A1 => n3, A2 => n11, ZN => OUT1_18_port);
   U24 : NAND2_X1 port map( A1 => n3, A2 => n7, ZN => OUT1_22_port);
   U25 : NAND2_X1 port map( A1 => n3, A2 => n6, ZN => OUT1_23_port);

end SYN_Bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity ff32_en_IR is

   port( D : in std_logic_vector (31 downto 0);  en, clk, rst : in std_logic;  
         Q : out std_logic_vector (31 downto 0));

end ff32_en_IR;

architecture SYN_behavioral of ff32_en_IR is

   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFS_X2
      port( D, CK, SN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFR_X2
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFS_X1
      port( D, CK, SN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_ff32_en_IR
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal net199603, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, 
      n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n30
      , n33, n28, n29, n31, n32 : std_logic;

begin
   
   Q_reg_31_inst : DFFR_X1 port map( D => D(31), CK => net199603, RN => n32, Q 
                           => Q(31), QN => n33);
   Q_reg_29_inst : DFFR_X1 port map( D => D(29), CK => net199603, RN => n32, Q 
                           => Q(29), QN => n30);
   Q_reg_26_inst : DFFS_X1 port map( D => D(26), CK => net199603, SN => n32, Q 
                           => Q(26), QN => n27);
   Q_reg_25_inst : DFFR_X1 port map( D => D(25), CK => net199603, RN => n32, Q 
                           => Q(25), QN => n26);
   Q_reg_24_inst : DFFR_X1 port map( D => D(24), CK => net199603, RN => n32, Q 
                           => Q(24), QN => n25);
   Q_reg_23_inst : DFFR_X1 port map( D => D(23), CK => net199603, RN => n32, Q 
                           => Q(23), QN => n24);
   Q_reg_22_inst : DFFR_X1 port map( D => D(22), CK => net199603, RN => n32, Q 
                           => Q(22), QN => n23);
   Q_reg_21_inst : DFFR_X1 port map( D => D(21), CK => net199603, RN => n32, Q 
                           => Q(21), QN => n22);
   Q_reg_20_inst : DFFR_X1 port map( D => D(20), CK => net199603, RN => n32, Q 
                           => Q(20), QN => n21);
   Q_reg_19_inst : DFFR_X1 port map( D => D(19), CK => net199603, RN => n32, Q 
                           => Q(19), QN => n20);
   Q_reg_18_inst : DFFR_X1 port map( D => D(18), CK => net199603, RN => n32, Q 
                           => Q(18), QN => n19);
   Q_reg_17_inst : DFFR_X1 port map( D => D(17), CK => net199603, RN => n32, Q 
                           => Q(17), QN => n18);
   Q_reg_16_inst : DFFR_X1 port map( D => D(16), CK => net199603, RN => n32, Q 
                           => Q(16), QN => n17);
   Q_reg_15_inst : DFFR_X1 port map( D => D(15), CK => net199603, RN => n32, Q 
                           => Q(15), QN => n16);
   Q_reg_14_inst : DFFR_X1 port map( D => D(14), CK => net199603, RN => n32, Q 
                           => Q(14), QN => n15);
   Q_reg_13_inst : DFFR_X1 port map( D => D(13), CK => net199603, RN => n32, Q 
                           => Q(13), QN => n14);
   Q_reg_12_inst : DFFR_X1 port map( D => D(12), CK => net199603, RN => n32, Q 
                           => Q(12), QN => n13);
   Q_reg_11_inst : DFFR_X1 port map( D => D(11), CK => net199603, RN => n32, Q 
                           => Q(11), QN => n12);
   Q_reg_10_inst : DFFR_X1 port map( D => D(10), CK => net199603, RN => n32, Q 
                           => Q(10), QN => n11);
   Q_reg_9_inst : DFFR_X1 port map( D => D(9), CK => net199603, RN => n32, Q =>
                           Q(9), QN => n10);
   Q_reg_8_inst : DFFR_X1 port map( D => D(8), CK => net199603, RN => n32, Q =>
                           Q(8), QN => n9);
   Q_reg_7_inst : DFFR_X1 port map( D => D(7), CK => net199603, RN => n32, Q =>
                           Q(7), QN => n8);
   Q_reg_6_inst : DFFR_X1 port map( D => D(6), CK => net199603, RN => n32, Q =>
                           Q(6), QN => n7);
   Q_reg_5_inst : DFFR_X1 port map( D => D(5), CK => net199603, RN => n32, Q =>
                           Q(5), QN => n6);
   Q_reg_4_inst : DFFR_X1 port map( D => D(4), CK => net199603, RN => n32, Q =>
                           Q(4), QN => n5);
   Q_reg_3_inst : DFFR_X1 port map( D => D(3), CK => net199603, RN => n32, Q =>
                           Q(3), QN => n4);
   Q_reg_2_inst : DFFR_X1 port map( D => D(2), CK => net199603, RN => n32, Q =>
                           Q(2), QN => n3);
   Q_reg_1_inst : DFFR_X1 port map( D => D(1), CK => net199603, RN => n32, Q =>
                           Q(1), QN => n2);
   Q_reg_0_inst : DFFR_X1 port map( D => D(0), CK => net199603, RN => n32, Q =>
                           Q(0), QN => n1);
   clk_gate_Q_reg : SNPS_CLOCK_GATE_HIGH_ff32_en_IR port map( CLK => clk, EN =>
                           en, ENCLK => net199603);
   Q_reg_30_inst : DFFS_X1 port map( D => D(30), CK => net199603, SN => n32, Q 
                           => Q(30), QN => n31);
   Q_reg_27_inst : DFFR_X2 port map( D => D(27), CK => net199603, RN => n32, Q 
                           => Q(27), QN => n29);
   Q_reg_28_inst : DFFS_X2 port map( D => D(28), CK => net199603, SN => n32, Q 
                           => Q(28), QN => n28);
   U2 : INV_X2 port map( A => rst, ZN => n32);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_0 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_0;

architecture SYN_USE_DEFA_ARCH_NAME of 
   SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net199627 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net199627);
   main_gate : AND2_X1 port map( A1 => net199627, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity predictor_2_0 is

   port( clock, reset, enable, taken_i : in std_logic;  prediction_o : out 
         std_logic);

end predictor_2_0;

architecture SYN_bhe of predictor_2_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal prediction_o_port, next_STATE_1_port, next_STATE_0_port, N11, N12, n3
      , n4, n6, n8, n9, n1, n2, net246123 : std_logic;

begin
   prediction_o <= prediction_o_port;
   
   next_STATE_reg_0_inst : DLH_X1 port map( G => enable, D => N11, Q => 
                           next_STATE_0_port);
   STATE_reg_0_inst : DFFR_X1 port map( D => n8, CK => clock, RN => n2, Q => n1
                           , QN => n9);
   next_STATE_reg_1_inst : DLH_X1 port map( G => enable, D => N12, Q => 
                           next_STATE_1_port);
   STATE_reg_1_inst : DFFR_X1 port map( D => n6, CK => clock, RN => n2, Q => 
                           prediction_o_port, QN => net246123);
   U2 : MUX2_X1 port map( A => prediction_o_port, B => next_STATE_1_port, S => 
                           enable, Z => n6);
   U4 : MUX2_X1 port map( A => n1, B => next_STATE_0_port, S => enable, Z => n8
                           );
   U9 : NOR2_X1 port map( A1 => prediction_o_port, A2 => taken_i, ZN => n3);
   U7 : NAND2_X1 port map( A1 => prediction_o_port, A2 => taken_i, ZN => n4);
   U5 : OAI21_X1 port map( B1 => n9, B2 => n3, A => n4, ZN => N12);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n1, A => n4, ZN => N11);
   U3 : INV_X1 port map( A => reset, ZN => n2);

end SYN_bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity mux41_0 is

   port( IN0, IN1, IN2, IN3 : in std_logic_vector (31 downto 0);  CTRL : in 
         std_logic_vector (1 downto 0);  OUT1 : out std_logic_vector (31 downto
         0));

end mux41_0;

architecture SYN_bhe of mux41_0 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n6, n7, n8, n45, n46, n53, n54, n55, n56, n63, n64, n65, n66, n67
      , n68, n71, n38, n37, n1, n2, n3, n4, n9, n10, n11, n12, n13, n14, n15, 
      n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30
      , n31, n32, n34, n35, n36, n39, n40, n41, n43, n44, n47, n48, n49, n50, 
      n52, n57, n58, n60, n61, n62, n70, n72, n73, n74, n75, n76, n77, n78, n79
      , n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, 
      n94, n95, n96, n97, n98, n99, n100, n102, n103, n104, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125 : std_logic;

begin
   
   U87 : AOI22_X1 port map( A1 => n7, A2 => IN1(12), B1 => n124, B2 => IN0(12),
                           ZN => n63);
   U86 : AOI22_X1 port map( A1 => n9, A2 => IN3(12), B1 => n125, B2 => IN2(12),
                           ZN => n64);
   U72 : AOI22_X1 port map( A1 => n7, A2 => IN1(17), B1 => n124, B2 => IN0(17),
                           ZN => n53);
   U71 : AOI22_X1 port map( A1 => n9, A2 => IN3(17), B1 => n125, B2 => IN2(17),
                           ZN => n54);
   U75 : AOI22_X1 port map( A1 => n7, A2 => IN1(16), B1 => n124, B2 => IN0(16),
                           ZN => n55);
   U74 : AOI22_X1 port map( A1 => n9, A2 => IN3(16), B1 => n125, B2 => IN2(16),
                           ZN => n56);
   U93 : AOI22_X1 port map( A1 => n7, A2 => IN1(10), B1 => n124, B2 => IN0(10),
                           ZN => n67);
   U92 : AOI22_X1 port map( A1 => n9, A2 => IN3(10), B1 => n125, B2 => IN2(10),
                           ZN => n68);
   U90 : AOI22_X1 port map( A1 => n7, A2 => IN1(11), B1 => n124, B2 => IN0(11),
                           ZN => n65);
   U89 : AOI22_X1 port map( A1 => n9, A2 => IN3(11), B1 => n125, B2 => IN2(11),
                           ZN => n66);
   U48 : AOI22_X1 port map( A1 => n7, A2 => IN1(24), B1 => n124, B2 => IN0(24),
                           ZN => n37);
   U60 : AOI22_X1 port map( A1 => n7, A2 => IN1(20), B1 => n124, B2 => IN0(20),
                           ZN => n45);
   U59 : AOI22_X1 port map( A1 => n5, A2 => IN3(20), B1 => n6, B2 => IN2(20), 
                           ZN => n46);
   U85 : NAND2_X2 port map( A1 => n63, A2 => n64, ZN => OUT1(12));
   U70 : NAND2_X2 port map( A1 => n53, A2 => n54, ZN => OUT1(17));
   U73 : NAND2_X2 port map( A1 => n55, A2 => n56, ZN => OUT1(16));
   U91 : NAND2_X2 port map( A1 => n67, A2 => n68, ZN => OUT1(10));
   U88 : NAND2_X2 port map( A1 => n65, A2 => n66, ZN => OUT1(11));
   U58 : NAND2_X2 port map( A1 => n45, A2 => n46, ZN => OUT1(20));
   U101 : INV_X1 port map( A => CTRL(1), ZN => n71);
   U1 : AOI22_X1 port map( A1 => IN2(8), A2 => n6, B1 => IN3(8), B2 => n9, ZN 
                           => n1);
   U2 : AOI22_X1 port map( A1 => IN0(8), A2 => n8, B1 => IN1(8), B2 => n7, ZN 
                           => n2);
   U3 : NAND2_X1 port map( A1 => n1, A2 => n2, ZN => OUT1(8));
   U4 : AOI22_X1 port map( A1 => IN2(21), A2 => n6, B1 => IN3(21), B2 => n9, ZN
                           => n3);
   U5 : AOI22_X1 port map( A1 => IN0(21), A2 => n124, B1 => IN1(21), B2 => n7, 
                           ZN => n4);
   U6 : NAND2_X1 port map( A1 => n3, A2 => n4, ZN => OUT1(21));
   U7 : NAND3_X2 port map( A1 => n102, A2 => n103, A3 => n104, ZN => OUT1(7));
   U8 : NAND3_X2 port map( A1 => n43, A2 => n44, A3 => n47, ZN => OUT1(27));
   U9 : AND2_X2 port map( A1 => n71, A2 => CTRL(0), ZN => n7);
   U10 : BUF_X2 port map( A => n5, Z => n9);
   U11 : NAND3_X1 port map( A1 => n106, A2 => n107, A3 => n108, ZN => OUT1(19))
                           ;
   U12 : NAND3_X1 port map( A1 => n34, A2 => n35, A3 => n36, ZN => OUT1(18));
   U13 : AND2_X1 port map( A1 => n124, A2 => IN0(28), ZN => n24);
   U14 : AND2_X1 port map( A1 => n124, A2 => IN0(15), ZN => n29);
   U15 : AND2_X1 port map( A1 => n124, A2 => IN0(2), ZN => n21);
   U16 : AND2_X1 port map( A1 => n124, A2 => IN0(0), ZN => n27);
   U17 : AND2_X1 port map( A1 => n124, A2 => IN0(30), ZN => n23);
   U18 : AND2_X1 port map( A1 => n124, A2 => IN0(1), ZN => n26);
   U19 : AND2_X1 port map( A1 => n124, A2 => IN0(29), ZN => n25);
   U20 : AND2_X1 port map( A1 => n124, A2 => IN0(13), ZN => n12);
   U21 : AND2_X1 port map( A1 => n124, A2 => IN0(25), ZN => n18);
   U22 : AND2_X1 port map( A1 => n124, A2 => IN0(14), ZN => n14);
   U23 : AND2_X1 port map( A1 => n124, A2 => IN0(22), ZN => n17);
   U24 : AND2_X1 port map( A1 => n124, A2 => IN0(27), ZN => n19);
   U25 : AND2_X1 port map( A1 => n124, A2 => IN0(19), ZN => n28);
   U26 : AND2_X1 port map( A1 => n124, A2 => IN0(18), ZN => n16);
   U27 : AND2_X1 port map( A1 => n124, A2 => IN0(23), ZN => n22);
   U28 : AND2_X1 port map( A1 => n124, A2 => IN0(26), ZN => n20);
   U29 : AND2_X1 port map( A1 => n8, A2 => IN0(7), ZN => n30);
   U30 : AND2_X1 port map( A1 => n8, A2 => IN0(5), ZN => n13);
   U31 : AND2_X1 port map( A1 => n8, A2 => IN0(6), ZN => n10);
   U32 : AND2_X1 port map( A1 => n8, A2 => IN0(31), ZN => n31);
   U33 : AND2_X1 port map( A1 => n8, A2 => IN0(4), ZN => n15);
   U34 : AND2_X1 port map( A1 => n8, A2 => IN0(9), ZN => n11);
   U35 : AND2_X1 port map( A1 => n8, A2 => IN0(3), ZN => n32);
   U36 : AND2_X1 port map( A1 => CTRL(0), A2 => CTRL(1), ZN => n5);
   U37 : NOR2_X1 port map( A1 => CTRL(0), A2 => CTRL(1), ZN => n8);
   U38 : NAND3_X1 port map( A1 => n121, A2 => n122, A3 => n123, ZN => OUT1(29))
                           ;
   U39 : NAND3_X1 port map( A1 => n115, A2 => n116, A3 => n117, ZN => OUT1(28))
                           ;
   U40 : NAND3_X2 port map( A1 => n95, A2 => n96, A3 => n97, ZN => OUT1(6));
   U41 : NAND3_X2 port map( A1 => n112, A2 => n113, A3 => n114, ZN => OUT1(14))
                           ;
   U42 : NAND3_X2 port map( A1 => n118, A2 => n119, A3 => n120, ZN => OUT1(15))
                           ;
   U43 : BUF_X1 port map( A => n8, Z => n124);
   U44 : NOR2_X2 port map( A1 => CTRL(0), A2 => n71, ZN => n6);
   U45 : BUF_X1 port map( A => n6, Z => n125);
   U46 : NAND3_X2 port map( A1 => n109, A2 => n110, A3 => n111, ZN => OUT1(30))
                           ;
   U47 : NAND3_X2 port map( A1 => n98, A2 => n99, A3 => n100, ZN => OUT1(31));
   U49 : NAND3_X2 port map( A1 => n60, A2 => n61, A3 => n62, ZN => OUT1(26));
   U50 : NAND3_X2 port map( A1 => n39, A2 => n40, A3 => n41, ZN => OUT1(25));
   U51 : NAND2_X2 port map( A1 => n37, A2 => n38, ZN => OUT1(24));
   U52 : NAND3_X2 port map( A1 => n80, A2 => n81, A3 => n82, ZN => OUT1(0));
   U53 : NAND3_X2 port map( A1 => n77, A2 => n78, A3 => n79, ZN => OUT1(1));
   U54 : NAND3_X2 port map( A1 => n92, A2 => n93, A3 => n94, ZN => OUT1(5));
   U55 : NAND3_X2 port map( A1 => n83, A2 => n84, A3 => n85, ZN => OUT1(4));
   U56 : NAND3_X2 port map( A1 => n89, A2 => n90, A3 => n91, ZN => OUT1(22));
   U57 : NAND3_X2 port map( A1 => n86, A2 => n87, A3 => n88, ZN => OUT1(23));
   U61 : NAND3_X2 port map( A1 => n70, A2 => n72, A3 => n73, ZN => OUT1(13));
   U62 : NAND3_X2 port map( A1 => n74, A2 => n75, A3 => n76, ZN => OUT1(2));
   U63 : NAND3_X2 port map( A1 => n48, A2 => n49, A3 => n50, ZN => OUT1(3));
   U64 : NAND3_X2 port map( A1 => n52, A2 => n57, A3 => n58, ZN => OUT1(9));
   U65 : NAND2_X1 port map( A1 => IN2(30), A2 => n6, ZN => n111);
   U66 : AOI21_X1 port map( B1 => IN1(30), B2 => n7, A => n23, ZN => n110);
   U67 : AOI21_X1 port map( B1 => IN1(31), B2 => n7, A => n31, ZN => n99);
   U68 : AOI21_X1 port map( B1 => IN1(27), B2 => n7, A => n19, ZN => n44);
   U69 : AOI21_X1 port map( B1 => IN1(26), B2 => n7, A => n20, ZN => n61);
   U76 : NAND2_X1 port map( A1 => IN2(25), A2 => n125, ZN => n41);
   U77 : AOI21_X1 port map( B1 => IN1(25), B2 => n7, A => n18, ZN => n40);
   U78 : NAND2_X1 port map( A1 => n125, A2 => IN2(0), ZN => n82);
   U79 : AOI21_X1 port map( B1 => IN1(0), B2 => n7, A => n27, ZN => n81);
   U80 : NAND2_X1 port map( A1 => n125, A2 => IN2(1), ZN => n79);
   U81 : AOI21_X1 port map( B1 => IN1(1), B2 => n7, A => n26, ZN => n78);
   U82 : NAND2_X1 port map( A1 => IN2(7), A2 => n125, ZN => n104);
   U83 : AOI21_X1 port map( B1 => IN1(7), B2 => n7, A => n30, ZN => n103);
   U84 : NAND2_X1 port map( A1 => IN2(6), A2 => n6, ZN => n97);
   U94 : AOI21_X1 port map( B1 => IN1(6), B2 => n7, A => n10, ZN => n96);
   U95 : NAND2_X1 port map( A1 => n6, A2 => IN2(5), ZN => n94);
   U96 : AOI21_X1 port map( B1 => IN1(5), B2 => n7, A => n13, ZN => n93);
   U97 : NAND2_X1 port map( A1 => n6, A2 => IN2(4), ZN => n85);
   U98 : AOI21_X1 port map( B1 => IN1(4), B2 => n7, A => n15, ZN => n84);
   U99 : NAND2_X1 port map( A1 => IN2(22), A2 => n6, ZN => n91);
   U100 : AOI21_X1 port map( B1 => IN1(22), B2 => n7, A => n17, ZN => n90);
   U102 : NAND2_X1 port map( A1 => IN2(23), A2 => n6, ZN => n88);
   U103 : AOI21_X1 port map( B1 => IN1(23), B2 => n7, A => n22, ZN => n87);
   U104 : NAND2_X1 port map( A1 => IN2(18), A2 => n125, ZN => n36);
   U105 : AOI21_X1 port map( B1 => IN1(18), B2 => n7, A => n16, ZN => n35);
   U106 : NAND2_X1 port map( A1 => IN2(19), A2 => n125, ZN => n108);
   U107 : AOI21_X1 port map( B1 => IN1(19), B2 => n7, A => n28, ZN => n107);
   U108 : NAND2_X1 port map( A1 => IN2(29), A2 => n6, ZN => n123);
   U109 : AOI21_X1 port map( B1 => IN1(29), B2 => n7, A => n25, ZN => n122);
   U110 : NAND2_X1 port map( A1 => IN2(28), A2 => n6, ZN => n117);
   U111 : AOI21_X1 port map( B1 => IN1(28), B2 => n7, A => n24, ZN => n116);
   U112 : NAND2_X1 port map( A1 => IN2(13), A2 => n125, ZN => n73);
   U113 : AOI21_X1 port map( B1 => IN1(13), B2 => n7, A => n12, ZN => n72);
   U114 : NAND2_X1 port map( A1 => n6, A2 => IN2(2), ZN => n76);
   U115 : AOI21_X1 port map( B1 => IN1(2), B2 => n7, A => n21, ZN => n75);
   U116 : NAND2_X1 port map( A1 => n6, A2 => IN2(3), ZN => n50);
   U117 : AOI21_X1 port map( B1 => IN1(3), B2 => n7, A => n32, ZN => n49);
   U118 : NAND2_X1 port map( A1 => IN2(9), A2 => n6, ZN => n58);
   U119 : AOI21_X1 port map( B1 => IN1(9), B2 => n7, A => n11, ZN => n57);
   U120 : NAND2_X1 port map( A1 => IN2(15), A2 => n125, ZN => n120);
   U121 : AOI21_X1 port map( B1 => IN1(15), B2 => n7, A => n29, ZN => n119);
   U122 : NAND2_X1 port map( A1 => IN2(14), A2 => n125, ZN => n114);
   U123 : AOI21_X1 port map( B1 => IN1(14), B2 => n7, A => n14, ZN => n113);
   U124 : NAND2_X1 port map( A1 => IN3(18), A2 => n9, ZN => n34);
   U125 : NAND2_X1 port map( A1 => IN3(25), A2 => n9, ZN => n39);
   U126 : AOI22_X1 port map( A1 => n9, A2 => IN3(24), B1 => n6, B2 => IN2(24), 
                           ZN => n38);
   U127 : NAND2_X1 port map( A1 => IN3(27), A2 => n9, ZN => n43);
   U128 : NAND2_X1 port map( A1 => IN2(27), A2 => n6, ZN => n47);
   U129 : NAND2_X1 port map( A1 => IN3(3), A2 => n9, ZN => n48);
   U130 : NAND2_X1 port map( A1 => IN3(9), A2 => n9, ZN => n52);
   U131 : NAND2_X1 port map( A1 => IN3(26), A2 => n9, ZN => n60);
   U132 : NAND2_X1 port map( A1 => IN2(26), A2 => n6, ZN => n62);
   U133 : NAND2_X1 port map( A1 => IN3(13), A2 => n9, ZN => n70);
   U134 : NAND2_X1 port map( A1 => IN3(2), A2 => n9, ZN => n74);
   U135 : NAND2_X1 port map( A1 => IN3(1), A2 => n9, ZN => n77);
   U136 : NAND2_X1 port map( A1 => IN3(0), A2 => n9, ZN => n80);
   U137 : NAND2_X1 port map( A1 => IN3(4), A2 => n9, ZN => n83);
   U138 : NAND2_X1 port map( A1 => IN3(23), A2 => n9, ZN => n86);
   U139 : NAND2_X1 port map( A1 => IN3(22), A2 => n9, ZN => n89);
   U140 : NAND2_X1 port map( A1 => IN3(5), A2 => n9, ZN => n92);
   U141 : NAND2_X1 port map( A1 => IN3(6), A2 => n9, ZN => n95);
   U142 : NAND2_X1 port map( A1 => IN3(31), A2 => n9, ZN => n98);
   U143 : NAND2_X1 port map( A1 => IN2(31), A2 => n6, ZN => n100);
   U144 : NAND2_X1 port map( A1 => IN3(7), A2 => n9, ZN => n102);
   U145 : NAND2_X1 port map( A1 => IN3(19), A2 => n9, ZN => n106);
   U146 : NAND2_X1 port map( A1 => IN3(30), A2 => n5, ZN => n109);
   U147 : NAND2_X1 port map( A1 => IN3(14), A2 => n9, ZN => n112);
   U148 : NAND2_X1 port map( A1 => IN3(28), A2 => n5, ZN => n115);
   U149 : NAND2_X1 port map( A1 => IN3(15), A2 => n9, ZN => n118);
   U150 : NAND2_X1 port map( A1 => IN3(29), A2 => n5, ZN => n121);

end SYN_bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity add4 is

   port( IN1 : in std_logic_vector (31 downto 0);  OUT1 : out std_logic_vector 
         (31 downto 0));

end add4;

architecture SYN_bhe of add4 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal OUT1_31_port, OUT1_30_port, OUT1_29_port, OUT1_28_port, OUT1_27_port,
      OUT1_26_port, OUT1_25_port, OUT1_24_port, OUT1_23_port, OUT1_22_port, 
      OUT1_21_port, OUT1_20_port, OUT1_19_port, OUT1_18_port, OUT1_17_port, 
      OUT1_16_port, OUT1_15_port, OUT1_14_port, OUT1_13_port, OUT1_12_port, 
      OUT1_11_port, OUT1_10_port, OUT1_9_port, OUT1_8_port, OUT1_7_port, 
      OUT1_6_port, OUT1_5_port, OUT1_4_port, OUT1_3_port, OUT1_2_port, n1, n2, 
      n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, 
      n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33
      , n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47 : 
      std_logic;

begin
   OUT1 <= ( OUT1_31_port, OUT1_30_port, OUT1_29_port, OUT1_28_port, 
      OUT1_27_port, OUT1_26_port, OUT1_25_port, OUT1_24_port, OUT1_23_port, 
      OUT1_22_port, OUT1_21_port, OUT1_20_port, OUT1_19_port, OUT1_18_port, 
      OUT1_17_port, OUT1_16_port, OUT1_15_port, OUT1_14_port, OUT1_13_port, 
      OUT1_12_port, OUT1_11_port, OUT1_10_port, OUT1_9_port, OUT1_8_port, 
      OUT1_7_port, OUT1_6_port, OUT1_5_port, OUT1_4_port, OUT1_3_port, 
      OUT1_2_port, IN1(1), IN1(0) );
   
   U3 : NAND3_X1 port map( A1 => n16, A2 => n15, A3 => IN1(15), ZN => n1);
   U4 : NOR3_X1 port map( A1 => n17, A2 => n18, A3 => n1, ZN => n2);
   U5 : NAND3_X1 port map( A1 => IN1(13), A2 => IN1(14), A3 => n2, ZN => n20);
   U6 : INV_X1 port map( A => n40, ZN => n3);
   U7 : NAND2_X1 port map( A1 => IN1(30), A2 => n3, ZN => n4);
   U8 : XNOR2_X1 port map( A => IN1(31), B => n4, ZN => OUT1_31_port);
   U9 : XOR2_X1 port map( A => n27, B => IN1(21), Z => OUT1_21_port);
   U10 : NAND2_X1 port map( A1 => n44, A2 => IN1(6), ZN => n5);
   U11 : XNOR2_X1 port map( A => n5, B => IN1(7), ZN => OUT1_7_port);
   U12 : NOR2_X1 port map( A1 => n10, A2 => n9, ZN => n6);
   U13 : XOR2_X1 port map( A => IN1(11), B => n6, Z => OUT1_11_port);
   U14 : INV_X1 port map( A => n14, ZN => n7);
   U15 : NAND2_X1 port map( A1 => IN1(14), A2 => n7, ZN => n8);
   U16 : XNOR2_X1 port map( A => IN1(15), B => n8, ZN => OUT1_15_port);
   U17 : XOR2_X1 port map( A => n21, B => IN1(17), Z => OUT1_17_port);
   U18 : XOR2_X1 port map( A => n24, B => IN1(19), Z => OUT1_19_port);
   U19 : XOR2_X1 port map( A => n30, B => IN1(23), Z => OUT1_23_port);
   U20 : XOR2_X1 port map( A => n33, B => IN1(25), Z => OUT1_25_port);
   U21 : XOR2_X1 port map( A => n36, B => IN1(27), Z => OUT1_27_port);
   U22 : XOR2_X1 port map( A => n39, B => IN1(29), Z => OUT1_29_port);
   U23 : INV_X1 port map( A => n11, ZN => n12);
   U24 : INV_X1 port map( A => IN1(28), ZN => n37);
   U25 : INV_X1 port map( A => IN1(26), ZN => n34);
   U26 : INV_X1 port map( A => IN1(24), ZN => n31);
   U27 : INV_X1 port map( A => IN1(22), ZN => n28);
   U28 : INV_X1 port map( A => IN1(20), ZN => n25);
   U29 : INV_X1 port map( A => IN1(18), ZN => n22);
   U30 : INV_X1 port map( A => IN1(16), ZN => n19);
   U31 : INV_X1 port map( A => IN1(12), ZN => n18);
   U32 : INV_X1 port map( A => IN1(10), ZN => n9);
   U33 : INV_X1 port map( A => IN1(8), ZN => n46);
   U34 : XOR2_X1 port map( A => n9, B => n10, Z => OUT1_10_port);
   U35 : NAND4_X1 port map( A1 => IN1(8), A2 => IN1(9), A3 => IN1(10), A4 => 
                           IN1(11), ZN => n17);
   U36 : XNOR2_X1 port map( A => n11, B => n18, ZN => OUT1_12_port);
   U37 : XOR2_X1 port map( A => IN1(13), B => n13, Z => OUT1_13_port);
   U38 : XNOR2_X1 port map( A => n14, B => IN1(14), ZN => OUT1_14_port);
   U39 : XNOR2_X1 port map( A => n20, B => IN1(16), ZN => OUT1_16_port);
   U40 : XNOR2_X1 port map( A => n23, B => IN1(18), ZN => OUT1_18_port);
   U41 : XNOR2_X1 port map( A => n26, B => IN1(20), ZN => OUT1_20_port);
   U42 : XNOR2_X1 port map( A => n29, B => IN1(22), ZN => OUT1_22_port);
   U43 : XNOR2_X1 port map( A => n32, B => IN1(24), ZN => OUT1_24_port);
   U44 : XNOR2_X1 port map( A => n35, B => IN1(26), ZN => OUT1_26_port);
   U45 : XNOR2_X1 port map( A => n38, B => IN1(28), ZN => OUT1_28_port);
   U46 : XNOR2_X1 port map( A => n40, B => IN1(30), ZN => OUT1_30_port);
   U47 : XNOR2_X1 port map( A => IN1(2), B => n41, ZN => OUT1_3_port);
   U48 : XOR2_X1 port map( A => IN1(4), B => n15, Z => OUT1_4_port);
   U49 : XOR2_X1 port map( A => n42, B => n43, Z => OUT1_5_port);
   U50 : INV_X1 port map( A => IN1(5), ZN => n42);
   U51 : XOR2_X1 port map( A => IN1(6), B => n44, Z => OUT1_6_port);
   U52 : XOR2_X1 port map( A => n46, B => n45, Z => OUT1_8_port);
   U53 : XOR2_X1 port map( A => IN1(9), B => n47, Z => OUT1_9_port);
   U54 : NAND2_X1 port map( A1 => n13, A2 => IN1(13), ZN => n14);
   U55 : NAND2_X1 port map( A1 => n47, A2 => IN1(9), ZN => n10);
   U56 : NAND2_X1 port map( A1 => n15, A2 => IN1(4), ZN => n43);
   U57 : AND4_X1 port map( A1 => IN1(5), A2 => IN1(4), A3 => IN1(6), A4 => 
                           IN1(7), ZN => n16);
   U58 : NAND2_X1 port map( A1 => n39, A2 => IN1(29), ZN => n40);
   U59 : NAND2_X1 port map( A1 => n36, A2 => IN1(27), ZN => n38);
   U60 : INV_X1 port map( A => IN1(3), ZN => n41);
   U61 : NOR2_X1 port map( A1 => n43, A2 => n42, ZN => n44);
   U62 : INV_X1 port map( A => IN1(2), ZN => OUT1_2_port);
   U63 : NAND2_X1 port map( A1 => n15, A2 => n16, ZN => n45);
   U64 : NOR2_X1 port map( A1 => n45, A2 => n46, ZN => n47);
   U65 : NOR2_X1 port map( A1 => n45, A2 => n17, ZN => n11);
   U66 : NAND2_X1 port map( A1 => n33, A2 => IN1(25), ZN => n35);
   U67 : NAND2_X1 port map( A1 => n21, A2 => IN1(17), ZN => n23);
   U68 : NAND2_X1 port map( A1 => n24, A2 => IN1(19), ZN => n26);
   U69 : NOR2_X1 port map( A1 => n12, A2 => n18, ZN => n13);
   U70 : NAND2_X1 port map( A1 => n27, A2 => IN1(21), ZN => n29);
   U71 : NAND2_X1 port map( A1 => n30, A2 => IN1(23), ZN => n32);
   U72 : NOR2_X1 port map( A1 => n38, A2 => n37, ZN => n39);
   U73 : NOR2_X1 port map( A1 => n41, A2 => OUT1_2_port, ZN => n15);
   U74 : NOR2_X1 port map( A1 => n20, A2 => n19, ZN => n21);
   U75 : NOR2_X1 port map( A1 => n23, A2 => n22, ZN => n24);
   U76 : NOR2_X1 port map( A1 => n26, A2 => n25, ZN => n27);
   U77 : NOR2_X1 port map( A1 => n29, A2 => n28, ZN => n30);
   U78 : NOR2_X1 port map( A1 => n32, A2 => n31, ZN => n33);
   U79 : NOR2_X1 port map( A1 => n35, A2 => n34, ZN => n36);

end SYN_bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity ff32_en_0 is

   port( D : in std_logic_vector (31 downto 0);  en, clk, rst : in std_logic;  
         Q : out std_logic_vector (31 downto 0));

end ff32_en_0;

architecture SYN_behavioral of ff32_en_0 is

   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_ff32_en_0
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal net199618, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, 
      n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28
      , n29, n30, n31, n33, n32 : std_logic;

begin
   
   Q_reg_31_inst : DFFR_X1 port map( D => D(31), CK => net199618, RN => n32, Q 
                           => Q(31), QN => n33);
   Q_reg_30_inst : DFFR_X1 port map( D => D(30), CK => net199618, RN => n32, Q 
                           => Q(30), QN => n31);
   Q_reg_29_inst : DFFR_X1 port map( D => D(29), CK => net199618, RN => n32, Q 
                           => Q(29), QN => n30);
   Q_reg_28_inst : DFFR_X1 port map( D => D(28), CK => net199618, RN => n32, Q 
                           => Q(28), QN => n29);
   Q_reg_27_inst : DFFR_X1 port map( D => D(27), CK => net199618, RN => n32, Q 
                           => Q(27), QN => n28);
   Q_reg_26_inst : DFFR_X1 port map( D => D(26), CK => net199618, RN => n32, Q 
                           => Q(26), QN => n27);
   Q_reg_25_inst : DFFR_X1 port map( D => D(25), CK => net199618, RN => n32, Q 
                           => Q(25), QN => n26);
   Q_reg_24_inst : DFFR_X1 port map( D => D(24), CK => net199618, RN => n32, Q 
                           => Q(24), QN => n25);
   Q_reg_23_inst : DFFR_X1 port map( D => D(23), CK => net199618, RN => n32, Q 
                           => Q(23), QN => n24);
   Q_reg_22_inst : DFFR_X1 port map( D => D(22), CK => net199618, RN => n32, Q 
                           => Q(22), QN => n23);
   Q_reg_21_inst : DFFR_X1 port map( D => D(21), CK => net199618, RN => n32, Q 
                           => Q(21), QN => n22);
   Q_reg_20_inst : DFFR_X1 port map( D => D(20), CK => net199618, RN => n32, Q 
                           => Q(20), QN => n21);
   Q_reg_19_inst : DFFR_X1 port map( D => D(19), CK => net199618, RN => n32, Q 
                           => Q(19), QN => n20);
   Q_reg_18_inst : DFFR_X1 port map( D => D(18), CK => net199618, RN => n32, Q 
                           => Q(18), QN => n19);
   Q_reg_17_inst : DFFR_X1 port map( D => D(17), CK => net199618, RN => n32, Q 
                           => Q(17), QN => n18);
   Q_reg_16_inst : DFFR_X1 port map( D => D(16), CK => net199618, RN => n32, Q 
                           => Q(16), QN => n17);
   Q_reg_15_inst : DFFR_X1 port map( D => D(15), CK => net199618, RN => n32, Q 
                           => Q(15), QN => n16);
   Q_reg_14_inst : DFFR_X1 port map( D => D(14), CK => net199618, RN => n32, Q 
                           => Q(14), QN => n15);
   Q_reg_13_inst : DFFR_X1 port map( D => D(13), CK => net199618, RN => n32, Q 
                           => Q(13), QN => n14);
   Q_reg_12_inst : DFFR_X1 port map( D => D(12), CK => net199618, RN => n32, Q 
                           => Q(12), QN => n13);
   Q_reg_11_inst : DFFR_X1 port map( D => D(11), CK => net199618, RN => n32, Q 
                           => Q(11), QN => n12);
   Q_reg_10_inst : DFFR_X1 port map( D => D(10), CK => net199618, RN => n32, Q 
                           => Q(10), QN => n11);
   Q_reg_9_inst : DFFR_X1 port map( D => D(9), CK => net199618, RN => n32, Q =>
                           Q(9), QN => n10);
   Q_reg_8_inst : DFFR_X1 port map( D => D(8), CK => net199618, RN => n32, Q =>
                           Q(8), QN => n9);
   Q_reg_7_inst : DFFR_X1 port map( D => D(7), CK => net199618, RN => n32, Q =>
                           Q(7), QN => n8);
   Q_reg_6_inst : DFFR_X1 port map( D => D(6), CK => net199618, RN => n32, Q =>
                           Q(6), QN => n7);
   Q_reg_5_inst : DFFR_X1 port map( D => D(5), CK => net199618, RN => n32, Q =>
                           Q(5), QN => n6);
   Q_reg_4_inst : DFFR_X1 port map( D => D(4), CK => net199618, RN => n32, Q =>
                           Q(4), QN => n5);
   Q_reg_3_inst : DFFR_X1 port map( D => D(3), CK => net199618, RN => n32, Q =>
                           Q(3), QN => n4);
   Q_reg_2_inst : DFFR_X1 port map( D => D(2), CK => net199618, RN => n32, Q =>
                           Q(2), QN => n3);
   Q_reg_1_inst : DFFR_X1 port map( D => D(1), CK => net199618, RN => n32, Q =>
                           Q(1), QN => n2);
   Q_reg_0_inst : DFFR_X1 port map( D => D(0), CK => net199618, RN => n32, Q =>
                           Q(0), QN => n1);
   clk_gate_Q_reg : SNPS_CLOCK_GATE_HIGH_ff32_en_0 port map( CLK => clk, EN => 
                           en, ENCLK => net199618);
   U2 : INV_X2 port map( A => rst, ZN => n32);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity fw_logic is

   port( D1_i, rAdec_i, D2_i, D3_i, rA_i, rB_i : in std_logic_vector (4 downto 
         0);  S_mem_W, S_mem_LOAD, S_wb_W, S_exe_W : in std_logic;  S_FWAdec, 
         S_FWA, S_FWB : out std_logic_vector (1 downto 0));

end fw_logic;

architecture SYN_beh of fw_logic is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X2
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal S_FWAdec_1_port, S_FWAdec_0_port, S_FWA_1_port, S_FWA_0_port, n22, 
      n23, n25, n26, n29, n31, n34, n35, n55, n57, n58, n1, n2, n3, n4, n5, n6,
      n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, 
      n24, n27, n28, n30, n32, n33, n36, n37, n38, n39, n40, n41, n42, n43, n44
      , n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n56, n59, n60, n61, 
      n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76
      , n77, n78, n79, n80, n81, n82, n83 : std_logic;

begin
   S_FWAdec <= ( S_FWAdec_1_port, S_FWAdec_0_port );
   S_FWA <= ( S_FWA_1_port, S_FWA_0_port );
   
   U51 : NAND2_X1 port map( A1 => S_mem_W, A2 => n83, ZN => n31);
   U38 : INV_X1 port map( A => rA_i(3), ZN => n57);
   U33 : INV_X1 port map( A => rA_i(2), ZN => n55);
   U37 : INV_X1 port map( A => rA_i(1), ZN => n58);
   U2 : OR2_X1 port map( A1 => n34, A2 => rA_i(0), ZN => n30);
   U3 : OR2_X1 port map( A1 => n34, A2 => rB_i(0), ZN => n77);
   U4 : OR2_X1 port map( A1 => n34, A2 => rAdec_i(0), ZN => n60);
   U5 : NOR3_X1 port map( A1 => n73, A2 => n49, A3 => n72, ZN => S_FWB(0));
   U6 : OAI22_X1 port map( A1 => n29, A2 => rAdec_i(4), B1 => rAdec_i(0), B2 =>
                           n22, ZN => n1);
   U7 : AOI21_X1 port map( B1 => rAdec_i(0), B2 => n22, A => n1, ZN => n65);
   U8 : XNOR2_X1 port map( A => n23, B => rAdec_i(2), ZN => n70);
   U9 : INV_X1 port map( A => D3_i(0), ZN => n2);
   U10 : INV_X1 port map( A => rA_i(0), ZN => n3);
   U11 : OAI222_X1 port map( A1 => rA_i(0), A2 => n2, B1 => n3, B2 => D3_i(0), 
                           C1 => D3_i(1), C2 => n58, ZN => n4);
   U12 : AOI21_X1 port map( B1 => D3_i(3), B2 => n57, A => n4, ZN => n39);
   U13 : BUF_X1 port map( A => n50, Z => S_FWAdec_0_port);
   U14 : OR2_X1 port map( A1 => n80, A2 => rAdec_i(3), ZN => n62);
   U15 : NOR2_X1 port map( A1 => S_FWAdec_0_port, A2 => n63, ZN => 
                           S_FWAdec_1_port);
   U16 : INV_X1 port map( A => n42, ZN => n41);
   U17 : INV_X1 port map( A => n67, ZN => n66);
   U18 : OR2_X1 port map( A1 => n74, A2 => n31, ZN => n49);
   U19 : OR2_X1 port map( A1 => n80, A2 => rB_i(3), ZN => n79);
   U20 : INV_X1 port map( A => n31, ZN => n36);
   U21 : OR2_X1 port map( A1 => n80, A2 => rA_i(3), ZN => n33);
   U22 : INV_X1 port map( A => D2_i(3), ZN => n80);
   U23 : OR2_X1 port map( A1 => n35, A2 => rAdec_i(2), ZN => n56);
   U24 : OR2_X1 port map( A1 => n35, A2 => rA_i(2), ZN => n27);
   U25 : INV_X1 port map( A => D2_i(1), ZN => n81);
   U26 : OR2_X1 port map( A1 => n35, A2 => rB_i(2), ZN => n75);
   U27 : INV_X1 port map( A => rB_i(3), ZN => n19);
   U28 : INV_X1 port map( A => D3_i(1), ZN => n26);
   U29 : INV_X1 port map( A => D3_i(4), ZN => n29);
   U30 : INV_X1 port map( A => S_wb_W, ZN => n47);
   U31 : INV_X1 port map( A => D3_i(0), ZN => n22);
   U32 : INV_X1 port map( A => D2_i(0), ZN => n34);
   U34 : INV_X1 port map( A => D3_i(2), ZN => n23);
   U35 : INV_X1 port map( A => D3_i(3), ZN => n25);
   U36 : INV_X1 port map( A => D2_i(2), ZN => n35);
   U39 : INV_X1 port map( A => D2_i(1), ZN => n82);
   U40 : NOR2_X1 port map( A1 => S_FWA_0_port, A2 => n38, ZN => S_FWA_1_port);
   U41 : NOR4_X1 port map( A1 => n52, A2 => n51, A3 => n31, A4 => n53, ZN => 
                           n50);
   U42 : INV_X1 port map( A => rB_i(4), ZN => n15);
   U43 : INV_X1 port map( A => n72, ZN => n6);
   U44 : OAI211_X1 port map( C1 => n81, C2 => rB_i(1), A => n79, B => n78, ZN 
                           => n72);
   U45 : AOI21_X2 port map( B1 => n5, B2 => n6, A => n7, ZN => S_FWB(1));
   U46 : NOR3_X2 port map( A1 => n20, A2 => n21, A3 => n24, ZN => S_FWA_0_port)
                           ;
   U47 : OAI22_X1 port map( A1 => n29, A2 => rA_i(4), B1 => n57, B2 => D3_i(3),
                           ZN => n42);
   U48 : NOR2_X1 port map( A1 => n43, A2 => n44, ZN => n40);
   U49 : NAND2_X1 port map( A1 => n45, A2 => n46, ZN => n44);
   U50 : AOI21_X1 port map( B1 => n29, B2 => rA_i(4), A => n47, ZN => n46);
   U52 : NAND2_X1 port map( A1 => n55, A2 => D3_i(2), ZN => n45);
   U53 : OAI21_X1 port map( B1 => D3_i(2), B2 => n55, A => n48, ZN => n43);
   U54 : NAND2_X1 port map( A1 => n58, A2 => D3_i(1), ZN => n48);
   U55 : NAND2_X1 port map( A1 => n26, A2 => rAdec_i(1), ZN => n68);
   U56 : NOR2_X1 port map( A1 => n70, A2 => n71, ZN => n64);
   U57 : XNOR2_X1 port map( A => n25, B => rAdec_i(3), ZN => n71);
   U58 : OAI21_X1 port map( B1 => n15, B2 => D3_i(4), A => S_wb_W, ZN => n14);
   U59 : OAI222_X1 port map( A1 => n19, A2 => D3_i(3), B1 => rB_i(4), B2 => n29
                           , C1 => n22, C2 => rB_i(0), ZN => n16);
   U60 : AOI21_X1 port map( B1 => n26, B2 => rB_i(1), A => n14, ZN => n13);
   U61 : OAI21_X1 port map( B1 => n25, B2 => rB_i(3), A => n13, ZN => n10);
   U62 : NAND2_X1 port map( A1 => n22, A2 => rB_i(0), ZN => n18);
   U63 : OAI21_X1 port map( B1 => n23, B2 => rB_i(2), A => n18, ZN => n17);
   U64 : NOR2_X1 port map( A1 => n16, A2 => n17, ZN => n8);
   U65 : NAND2_X1 port map( A1 => n9, A2 => n8, ZN => n7);
   U66 : NAND2_X1 port map( A1 => n23, A2 => rB_i(2), ZN => n12);
   U67 : OAI21_X1 port map( B1 => n26, B2 => rB_i(1), A => n12, ZN => n11);
   U68 : NOR2_X1 port map( A1 => n10, A2 => n11, ZN => n9);
   U69 : NOR2_X1 port map( A1 => n73, A2 => n49, ZN => n5);
   U70 : NAND3_X1 port map( A1 => n27, A2 => n28, A3 => n30, ZN => n24);
   U71 : NAND2_X1 port map( A1 => n36, A2 => n37, ZN => n20);
   U72 : AOI22_X1 port map( A1 => n80, A2 => rA_i(3), B1 => n82, B2 => rA_i(1),
                           ZN => n32);
   U73 : OAI211_X1 port map( C1 => n82, C2 => rA_i(1), A => n32, B => n33, ZN 
                           => n21);
   U74 : AOI22_X1 port map( A1 => n35, A2 => rA_i(2), B1 => n34, B2 => rA_i(0),
                           ZN => n28);
   U75 : XNOR2_X1 port map( A => rA_i(4), B => D2_i(4), ZN => n37);
   U76 : NAND3_X1 port map( A1 => n39, A2 => n40, A3 => n41, ZN => n38);
   U77 : NAND3_X1 port map( A1 => n59, A2 => n56, A3 => n60, ZN => n52);
   U78 : AOI22_X1 port map( A1 => n80, A2 => rAdec_i(3), B1 => n82, B2 => 
                           rAdec_i(1), ZN => n61);
   U79 : OAI211_X1 port map( C1 => n82, C2 => rAdec_i(1), A => n62, B => n61, 
                           ZN => n51);
   U80 : AOI22_X1 port map( A1 => n35, A2 => rAdec_i(2), B1 => n34, B2 => 
                           rAdec_i(0), ZN => n59);
   U81 : INV_X1 port map( A => D2_i(4), ZN => n54);
   U82 : XNOR2_X1 port map( A => rAdec_i(4), B => n54, ZN => n53);
   U83 : NAND3_X1 port map( A1 => n64, A2 => n65, A3 => n66, ZN => n63);
   U84 : AOI21_X1 port map( B1 => rAdec_i(4), B2 => n29, A => n47, ZN => n69);
   U85 : OAI211_X1 port map( C1 => rAdec_i(1), C2 => n26, A => n68, B => n69, 
                           ZN => n67);
   U86 : XOR2_X1 port map( A => rB_i(4), B => D2_i(4), Z => n74);
   U87 : NAND3_X1 port map( A1 => n75, A2 => n76, A3 => n77, ZN => n73);
   U88 : AOI22_X1 port map( A1 => n80, A2 => rB_i(3), B1 => n81, B2 => rB_i(1),
                           ZN => n78);
   U89 : AOI22_X1 port map( A1 => n35, A2 => rB_i(2), B1 => n34, B2 => rB_i(0),
                           ZN => n76);
   U90 : INV_X1 port map( A => S_mem_LOAD, ZN => n83);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity mem_block is

   port( X_i, LOAD_i : in std_logic_vector (31 downto 0);  S_MUX_MEM_i : in 
         std_logic;  W_o : out std_logic_vector (31 downto 0));

end mem_block;

architecture SYN_struct of mem_block is

   component mux21_2
      port( IN0, IN1 : in std_logic_vector (31 downto 0);  CTRL : in std_logic;
            OUT1 : out std_logic_vector (31 downto 0));
   end component;

begin
   
   MUXMEM : mux21_2 port map( IN0(31) => X_i(31), IN0(30) => X_i(30), IN0(29) 
                           => X_i(29), IN0(28) => X_i(28), IN0(27) => X_i(27), 
                           IN0(26) => X_i(26), IN0(25) => X_i(25), IN0(24) => 
                           X_i(24), IN0(23) => X_i(23), IN0(22) => X_i(22), 
                           IN0(21) => X_i(21), IN0(20) => X_i(20), IN0(19) => 
                           X_i(19), IN0(18) => X_i(18), IN0(17) => X_i(17), 
                           IN0(16) => X_i(16), IN0(15) => X_i(15), IN0(14) => 
                           X_i(14), IN0(13) => X_i(13), IN0(12) => X_i(12), 
                           IN0(11) => X_i(11), IN0(10) => X_i(10), IN0(9) => 
                           X_i(9), IN0(8) => X_i(8), IN0(7) => X_i(7), IN0(6) 
                           => X_i(6), IN0(5) => X_i(5), IN0(4) => X_i(4), 
                           IN0(3) => X_i(3), IN0(2) => X_i(2), IN0(1) => X_i(1)
                           , IN0(0) => X_i(0), IN1(31) => LOAD_i(31), IN1(30) 
                           => LOAD_i(30), IN1(29) => LOAD_i(29), IN1(28) => 
                           LOAD_i(28), IN1(27) => LOAD_i(27), IN1(26) => 
                           LOAD_i(26), IN1(25) => LOAD_i(25), IN1(24) => 
                           LOAD_i(24), IN1(23) => LOAD_i(23), IN1(22) => 
                           LOAD_i(22), IN1(21) => LOAD_i(21), IN1(20) => 
                           LOAD_i(20), IN1(19) => LOAD_i(19), IN1(18) => 
                           LOAD_i(18), IN1(17) => LOAD_i(17), IN1(16) => 
                           LOAD_i(16), IN1(15) => LOAD_i(15), IN1(14) => 
                           LOAD_i(14), IN1(13) => LOAD_i(13), IN1(12) => 
                           LOAD_i(12), IN1(11) => LOAD_i(11), IN1(10) => 
                           LOAD_i(10), IN1(9) => LOAD_i(9), IN1(8) => LOAD_i(8)
                           , IN1(7) => LOAD_i(7), IN1(6) => LOAD_i(6), IN1(5) 
                           => LOAD_i(5), IN1(4) => LOAD_i(4), IN1(3) => 
                           LOAD_i(3), IN1(2) => LOAD_i(2), IN1(1) => LOAD_i(1),
                           IN1(0) => LOAD_i(0), CTRL => S_MUX_MEM_i, OUT1(31) 
                           => W_o(31), OUT1(30) => W_o(30), OUT1(29) => W_o(29)
                           , OUT1(28) => W_o(28), OUT1(27) => W_o(27), OUT1(26)
                           => W_o(26), OUT1(25) => W_o(25), OUT1(24) => W_o(24)
                           , OUT1(23) => W_o(23), OUT1(22) => W_o(22), OUT1(21)
                           => W_o(21), OUT1(20) => W_o(20), OUT1(19) => W_o(19)
                           , OUT1(18) => W_o(18), OUT1(17) => W_o(17), OUT1(16)
                           => W_o(16), OUT1(15) => W_o(15), OUT1(14) => W_o(14)
                           , OUT1(13) => W_o(13), OUT1(12) => W_o(12), OUT1(11)
                           => W_o(11), OUT1(10) => W_o(10), OUT1(9) => W_o(9), 
                           OUT1(8) => W_o(8), OUT1(7) => W_o(7), OUT1(6) => 
                           W_o(6), OUT1(5) => W_o(5), OUT1(4) => W_o(4), 
                           OUT1(3) => W_o(3), OUT1(2) => W_o(2), OUT1(1) => 
                           W_o(1), OUT1(0) => W_o(0));

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity mem_regs is

   port( W_i : in std_logic_vector (31 downto 0);  D3_i : in std_logic_vector 
         (4 downto 0);  W_o : out std_logic_vector (31 downto 0);  D3_o : out 
         std_logic_vector (4 downto 0);  clk, rst : in std_logic);

end mem_regs;

architecture SYN_Struct of mem_regs is

   component ff32_SIZE5
      port( D : in std_logic_vector (4 downto 0);  clk, rst : in std_logic;  Q 
            : out std_logic_vector (4 downto 0));
   end component;
   
   component ff32_SIZE32
      port( D : in std_logic_vector (31 downto 0);  clk, rst : in std_logic;  Q
            : out std_logic_vector (31 downto 0));
   end component;

begin
   
   W : ff32_SIZE32 port map( D(31) => W_i(31), D(30) => W_i(30), D(29) => 
                           W_i(29), D(28) => W_i(28), D(27) => W_i(27), D(26) 
                           => W_i(26), D(25) => W_i(25), D(24) => W_i(24), 
                           D(23) => W_i(23), D(22) => W_i(22), D(21) => W_i(21)
                           , D(20) => W_i(20), D(19) => W_i(19), D(18) => 
                           W_i(18), D(17) => W_i(17), D(16) => W_i(16), D(15) 
                           => W_i(15), D(14) => W_i(14), D(13) => W_i(13), 
                           D(12) => W_i(12), D(11) => W_i(11), D(10) => W_i(10)
                           , D(9) => W_i(9), D(8) => W_i(8), D(7) => W_i(7), 
                           D(6) => W_i(6), D(5) => W_i(5), D(4) => W_i(4), D(3)
                           => W_i(3), D(2) => W_i(2), D(1) => W_i(1), D(0) => 
                           W_i(0), clk => clk, rst => rst, Q(31) => W_o(31), 
                           Q(30) => W_o(30), Q(29) => W_o(29), Q(28) => W_o(28)
                           , Q(27) => W_o(27), Q(26) => W_o(26), Q(25) => 
                           W_o(25), Q(24) => W_o(24), Q(23) => W_o(23), Q(22) 
                           => W_o(22), Q(21) => W_o(21), Q(20) => W_o(20), 
                           Q(19) => W_o(19), Q(18) => W_o(18), Q(17) => W_o(17)
                           , Q(16) => W_o(16), Q(15) => W_o(15), Q(14) => 
                           W_o(14), Q(13) => W_o(13), Q(12) => W_o(12), Q(11) 
                           => W_o(11), Q(10) => W_o(10), Q(9) => W_o(9), Q(8) 
                           => W_o(8), Q(7) => W_o(7), Q(6) => W_o(6), Q(5) => 
                           W_o(5), Q(4) => W_o(4), Q(3) => W_o(3), Q(2) => 
                           W_o(2), Q(1) => W_o(1), Q(0) => W_o(0));
   D3 : ff32_SIZE5 port map( D(4) => D3_i(4), D(3) => D3_i(3), D(2) => D3_i(2),
                           D(1) => D3_i(1), D(0) => D3_i(0), clk => clk, rst =>
                           rst, Q(4) => D3_o(4), Q(3) => D3_o(3), Q(2) => 
                           D3_o(2), Q(1) => D3_o(1), Q(0) => D3_o(0));

end SYN_Struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity execute_block is

   port( IMM_i, A_i : in std_logic_vector (31 downto 0);  rB_i, rC_i : in 
         std_logic_vector (4 downto 0);  MUXED_B_i : in std_logic_vector (31 
         downto 0);  S_MUX_ALUIN_i : in std_logic;  FW_X_i, FW_W_i : in 
         std_logic_vector (31 downto 0);  S_FW_A_i, S_FW_B_i : in 
         std_logic_vector (1 downto 0);  muxed_dest : out std_logic_vector (4 
         downto 0);  muxed_B : out std_logic_vector (31 downto 0);  
         S_MUX_DEST_i : in std_logic_vector (1 downto 0);  OP : in 
         std_logic_vector (0 to 4);  ALUW_i : in std_logic_vector (12 downto 0)
         ;  DOUT : out std_logic_vector (31 downto 0);  stall_o : out std_logic
         ;  Clock, Reset : in std_logic);

end execute_block;

architecture SYN_struct of execute_block is

   component mux41_MUX_SIZE32_1
      port( IN0, IN1, IN2, IN3 : in std_logic_vector (31 downto 0);  CTRL : in 
            std_logic_vector (1 downto 0);  OUT1 : out std_logic_vector (31 
            downto 0));
   end component;
   
   component mux41_MUX_SIZE32_2
      port( IN0, IN1, IN2, IN3 : in std_logic_vector (31 downto 0);  CTRL : in 
            std_logic_vector (1 downto 0);  OUT1 : out std_logic_vector (31 
            downto 0));
   end component;
   
   component mux41_MUX_SIZE5
      port( IN0, IN1, IN2, IN3 : in std_logic_vector (4 downto 0);  CTRL : in 
            std_logic_vector (1 downto 0);  OUT1 : out std_logic_vector (4 
            downto 0));
   end component;
   
   component real_alu_DATA_SIZE32
      port( IN1, IN2 : in std_logic_vector (31 downto 0);  ALUW_i : in 
            std_logic_vector (12 downto 0);  DOUT : out std_logic_vector (31 
            downto 0);  stall_o : out std_logic;  Clock, Reset : in std_logic);
   end component;
   
   component mux21_3
      port( IN0, IN1 : in std_logic_vector (31 downto 0);  CTRL : in std_logic;
            OUT1 : out std_logic_vector (31 downto 0));
   end component;
   
   signal X_Logic1_port, X_Logic0_port, muxed_B_31_port, muxed_B_30_port, 
      muxed_B_29_port, muxed_B_28_port, muxed_B_27_port, muxed_B_26_port, 
      muxed_B_25_port, muxed_B_24_port, muxed_B_23_port, muxed_B_22_port, 
      muxed_B_21_port, muxed_B_20_port, muxed_B_19_port, muxed_B_18_port, 
      muxed_B_17_port, muxed_B_16_port, muxed_B_15_port, muxed_B_14_port, 
      muxed_B_13_port, muxed_B_12_port, muxed_B_11_port, muxed_B_10_port, 
      muxed_B_9_port, muxed_B_8_port, muxed_B_7_port, muxed_B_6_port, 
      muxed_B_5_port, muxed_B_4_port, muxed_B_2_port, muxed_B_1_port, 
      muxed_B_0_port, FWB2alu_31_port, FWB2alu_30_port, FWB2alu_29_port, 
      FWB2alu_28_port, FWB2alu_27_port, FWB2alu_26_port, FWB2alu_25_port, 
      FWB2alu_24_port, FWB2alu_23_port, FWB2alu_22_port, FWB2alu_21_port, 
      FWB2alu_20_port, FWB2alu_19_port, FWB2alu_18_port, FWB2alu_17_port, 
      FWB2alu_16_port, FWB2alu_15_port, FWB2alu_14_port, FWB2alu_13_port, 
      FWB2alu_12_port, FWB2alu_11_port, FWB2alu_10_port, FWB2alu_9_port, 
      FWB2alu_8_port, FWB2alu_7_port, FWB2alu_6_port, FWB2alu_5_port, 
      FWB2alu_4_port, FWB2alu_3_port, FWB2alu_2_port, FWB2alu_1_port, 
      FWB2alu_0_port, FWA2alu_31_port, FWA2alu_30_port, FWA2alu_29_port, 
      FWA2alu_28_port, FWA2alu_27_port, FWA2alu_26_port, FWA2alu_25_port, 
      FWA2alu_24_port, FWA2alu_23_port, FWA2alu_22_port, FWA2alu_21_port, 
      FWA2alu_20_port, FWA2alu_19_port, FWA2alu_18_port, FWA2alu_17_port, 
      FWA2alu_16_port, FWA2alu_15_port, FWA2alu_14_port, FWA2alu_13_port, 
      FWA2alu_12_port, FWA2alu_11_port, FWA2alu_10_port, FWA2alu_9_port, 
      FWA2alu_8_port, FWA2alu_7_port, FWA2alu_6_port, FWA2alu_5_port, 
      FWA2alu_4_port, FWA2alu_3_port, FWA2alu_2_port, FWA2alu_1_port, 
      FWA2alu_0_port, n1, muxed_B_3_port : std_logic;

begin
   muxed_B <= ( muxed_B_31_port, muxed_B_30_port, muxed_B_29_port, 
      muxed_B_28_port, muxed_B_27_port, muxed_B_26_port, muxed_B_25_port, 
      muxed_B_24_port, muxed_B_23_port, muxed_B_22_port, muxed_B_21_port, 
      muxed_B_20_port, muxed_B_19_port, muxed_B_18_port, muxed_B_17_port, 
      muxed_B_16_port, muxed_B_15_port, muxed_B_14_port, muxed_B_13_port, 
      muxed_B_12_port, muxed_B_11_port, muxed_B_10_port, muxed_B_9_port, 
      muxed_B_8_port, muxed_B_7_port, muxed_B_6_port, muxed_B_5_port, 
      muxed_B_4_port, muxed_B_3_port, muxed_B_2_port, muxed_B_1_port, 
      muxed_B_0_port );
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   n1 <= '0';
   ALUIN_MUX : mux21_3 port map( IN0(31) => muxed_B_31_port, IN0(30) => 
                           muxed_B_30_port, IN0(29) => muxed_B_29_port, IN0(28)
                           => muxed_B_28_port, IN0(27) => muxed_B_27_port, 
                           IN0(26) => muxed_B_26_port, IN0(25) => 
                           muxed_B_25_port, IN0(24) => muxed_B_24_port, IN0(23)
                           => muxed_B_23_port, IN0(22) => muxed_B_22_port, 
                           IN0(21) => muxed_B_21_port, IN0(20) => 
                           muxed_B_20_port, IN0(19) => muxed_B_19_port, IN0(18)
                           => muxed_B_18_port, IN0(17) => muxed_B_17_port, 
                           IN0(16) => muxed_B_16_port, IN0(15) => 
                           muxed_B_15_port, IN0(14) => muxed_B_14_port, IN0(13)
                           => muxed_B_13_port, IN0(12) => muxed_B_12_port, 
                           IN0(11) => muxed_B_11_port, IN0(10) => 
                           muxed_B_10_port, IN0(9) => muxed_B_9_port, IN0(8) =>
                           muxed_B_8_port, IN0(7) => muxed_B_7_port, IN0(6) => 
                           muxed_B_6_port, IN0(5) => muxed_B_5_port, IN0(4) => 
                           muxed_B_4_port, IN0(3) => muxed_B_3_port, IN0(2) => 
                           muxed_B_2_port, IN0(1) => muxed_B_1_port, IN0(0) => 
                           muxed_B_0_port, IN1(31) => IMM_i(31), IN1(30) => 
                           IMM_i(30), IN1(29) => IMM_i(29), IN1(28) => 
                           IMM_i(28), IN1(27) => IMM_i(27), IN1(26) => 
                           IMM_i(26), IN1(25) => IMM_i(25), IN1(24) => 
                           IMM_i(24), IN1(23) => IMM_i(23), IN1(22) => 
                           IMM_i(22), IN1(21) => IMM_i(21), IN1(20) => 
                           IMM_i(20), IN1(19) => IMM_i(19), IN1(18) => 
                           IMM_i(18), IN1(17) => IMM_i(17), IN1(16) => 
                           IMM_i(16), IN1(15) => IMM_i(15), IN1(14) => 
                           IMM_i(14), IN1(13) => IMM_i(13), IN1(12) => 
                           IMM_i(12), IN1(11) => IMM_i(11), IN1(10) => 
                           IMM_i(10), IN1(9) => IMM_i(9), IN1(8) => IMM_i(8), 
                           IN1(7) => IMM_i(7), IN1(6) => IMM_i(6), IN1(5) => 
                           IMM_i(5), IN1(4) => IMM_i(4), IN1(3) => IMM_i(3), 
                           IN1(2) => IMM_i(2), IN1(1) => IMM_i(1), IN1(0) => 
                           IMM_i(0), CTRL => S_MUX_ALUIN_i, OUT1(31) => 
                           FWB2alu_31_port, OUT1(30) => FWB2alu_30_port, 
                           OUT1(29) => FWB2alu_29_port, OUT1(28) => 
                           FWB2alu_28_port, OUT1(27) => FWB2alu_27_port, 
                           OUT1(26) => FWB2alu_26_port, OUT1(25) => 
                           FWB2alu_25_port, OUT1(24) => FWB2alu_24_port, 
                           OUT1(23) => FWB2alu_23_port, OUT1(22) => 
                           FWB2alu_22_port, OUT1(21) => FWB2alu_21_port, 
                           OUT1(20) => FWB2alu_20_port, OUT1(19) => 
                           FWB2alu_19_port, OUT1(18) => FWB2alu_18_port, 
                           OUT1(17) => FWB2alu_17_port, OUT1(16) => 
                           FWB2alu_16_port, OUT1(15) => FWB2alu_15_port, 
                           OUT1(14) => FWB2alu_14_port, OUT1(13) => 
                           FWB2alu_13_port, OUT1(12) => FWB2alu_12_port, 
                           OUT1(11) => FWB2alu_11_port, OUT1(10) => 
                           FWB2alu_10_port, OUT1(9) => FWB2alu_9_port, OUT1(8) 
                           => FWB2alu_8_port, OUT1(7) => FWB2alu_7_port, 
                           OUT1(6) => FWB2alu_6_port, OUT1(5) => FWB2alu_5_port
                           , OUT1(4) => FWB2alu_4_port, OUT1(3) => 
                           FWB2alu_3_port, OUT1(2) => FWB2alu_2_port, OUT1(1) 
                           => FWB2alu_1_port, OUT1(0) => FWB2alu_0_port);
   ALU : real_alu_DATA_SIZE32 port map( IN1(31) => FWA2alu_31_port, IN1(30) => 
                           FWA2alu_30_port, IN1(29) => FWA2alu_29_port, IN1(28)
                           => FWA2alu_28_port, IN1(27) => FWA2alu_27_port, 
                           IN1(26) => FWA2alu_26_port, IN1(25) => 
                           FWA2alu_25_port, IN1(24) => FWA2alu_24_port, IN1(23)
                           => FWA2alu_23_port, IN1(22) => FWA2alu_22_port, 
                           IN1(21) => FWA2alu_21_port, IN1(20) => 
                           FWA2alu_20_port, IN1(19) => FWA2alu_19_port, IN1(18)
                           => FWA2alu_18_port, IN1(17) => FWA2alu_17_port, 
                           IN1(16) => FWA2alu_16_port, IN1(15) => 
                           FWA2alu_15_port, IN1(14) => FWA2alu_14_port, IN1(13)
                           => FWA2alu_13_port, IN1(12) => FWA2alu_12_port, 
                           IN1(11) => FWA2alu_11_port, IN1(10) => 
                           FWA2alu_10_port, IN1(9) => FWA2alu_9_port, IN1(8) =>
                           FWA2alu_8_port, IN1(7) => FWA2alu_7_port, IN1(6) => 
                           FWA2alu_6_port, IN1(5) => FWA2alu_5_port, IN1(4) => 
                           FWA2alu_4_port, IN1(3) => FWA2alu_3_port, IN1(2) => 
                           FWA2alu_2_port, IN1(1) => FWA2alu_1_port, IN1(0) => 
                           FWA2alu_0_port, IN2(31) => FWB2alu_31_port, IN2(30) 
                           => FWB2alu_30_port, IN2(29) => FWB2alu_29_port, 
                           IN2(28) => FWB2alu_28_port, IN2(27) => 
                           FWB2alu_27_port, IN2(26) => FWB2alu_26_port, IN2(25)
                           => FWB2alu_25_port, IN2(24) => FWB2alu_24_port, 
                           IN2(23) => FWB2alu_23_port, IN2(22) => 
                           FWB2alu_22_port, IN2(21) => FWB2alu_21_port, IN2(20)
                           => FWB2alu_20_port, IN2(19) => FWB2alu_19_port, 
                           IN2(18) => FWB2alu_18_port, IN2(17) => 
                           FWB2alu_17_port, IN2(16) => FWB2alu_16_port, IN2(15)
                           => FWB2alu_15_port, IN2(14) => FWB2alu_14_port, 
                           IN2(13) => FWB2alu_13_port, IN2(12) => 
                           FWB2alu_12_port, IN2(11) => FWB2alu_11_port, IN2(10)
                           => FWB2alu_10_port, IN2(9) => FWB2alu_9_port, IN2(8)
                           => FWB2alu_8_port, IN2(7) => FWB2alu_7_port, IN2(6) 
                           => FWB2alu_6_port, IN2(5) => FWB2alu_5_port, IN2(4) 
                           => FWB2alu_4_port, IN2(3) => FWB2alu_3_port, IN2(2) 
                           => FWB2alu_2_port, IN2(1) => FWB2alu_1_port, IN2(0) 
                           => FWB2alu_0_port, ALUW_i(12) => ALUW_i(12), 
                           ALUW_i(11) => ALUW_i(11), ALUW_i(10) => ALUW_i(10), 
                           ALUW_i(9) => ALUW_i(9), ALUW_i(8) => ALUW_i(8), 
                           ALUW_i(7) => ALUW_i(7), ALUW_i(6) => ALUW_i(6), 
                           ALUW_i(5) => ALUW_i(5), ALUW_i(4) => ALUW_i(4), 
                           ALUW_i(3) => ALUW_i(3), ALUW_i(2) => ALUW_i(2), 
                           ALUW_i(1) => ALUW_i(1), ALUW_i(0) => ALUW_i(0), 
                           DOUT(31) => DOUT(31), DOUT(30) => DOUT(30), DOUT(29)
                           => DOUT(29), DOUT(28) => DOUT(28), DOUT(27) => 
                           DOUT(27), DOUT(26) => DOUT(26), DOUT(25) => DOUT(25)
                           , DOUT(24) => DOUT(24), DOUT(23) => DOUT(23), 
                           DOUT(22) => DOUT(22), DOUT(21) => DOUT(21), DOUT(20)
                           => DOUT(20), DOUT(19) => DOUT(19), DOUT(18) => 
                           DOUT(18), DOUT(17) => DOUT(17), DOUT(16) => DOUT(16)
                           , DOUT(15) => DOUT(15), DOUT(14) => DOUT(14), 
                           DOUT(13) => DOUT(13), DOUT(12) => DOUT(12), DOUT(11)
                           => DOUT(11), DOUT(10) => DOUT(10), DOUT(9) => 
                           DOUT(9), DOUT(8) => DOUT(8), DOUT(7) => DOUT(7), 
                           DOUT(6) => DOUT(6), DOUT(5) => DOUT(5), DOUT(4) => 
                           DOUT(4), DOUT(3) => DOUT(3), DOUT(2) => DOUT(2), 
                           DOUT(1) => DOUT(1), DOUT(0) => DOUT(0), stall_o => 
                           stall_o, Clock => Clock, Reset => Reset);
   MUXDEST : mux41_MUX_SIZE5 port map( IN0(4) => X_Logic0_port, IN0(3) => 
                           X_Logic0_port, IN0(2) => X_Logic0_port, IN0(1) => 
                           X_Logic0_port, IN0(0) => X_Logic0_port, IN1(4) => 
                           rC_i(4), IN1(3) => rC_i(3), IN1(2) => rC_i(2), 
                           IN1(1) => rC_i(1), IN1(0) => rC_i(0), IN2(4) => 
                           rB_i(4), IN2(3) => rB_i(3), IN2(2) => rB_i(2), 
                           IN2(1) => rB_i(1), IN2(0) => rB_i(0), IN3(4) => 
                           X_Logic1_port, IN3(3) => X_Logic1_port, IN3(2) => 
                           X_Logic1_port, IN3(1) => X_Logic1_port, IN3(0) => 
                           X_Logic1_port, CTRL(1) => S_MUX_DEST_i(1), CTRL(0) 
                           => S_MUX_DEST_i(0), OUT1(4) => muxed_dest(4), 
                           OUT1(3) => muxed_dest(3), OUT1(2) => muxed_dest(2), 
                           OUT1(1) => muxed_dest(1), OUT1(0) => muxed_dest(0));
   MUX_FWA : mux41_MUX_SIZE32_2 port map( IN0(31) => A_i(31), IN0(30) => 
                           A_i(30), IN0(29) => A_i(29), IN0(28) => A_i(28), 
                           IN0(27) => A_i(27), IN0(26) => A_i(26), IN0(25) => 
                           A_i(25), IN0(24) => A_i(24), IN0(23) => A_i(23), 
                           IN0(22) => A_i(22), IN0(21) => A_i(21), IN0(20) => 
                           A_i(20), IN0(19) => A_i(19), IN0(18) => A_i(18), 
                           IN0(17) => A_i(17), IN0(16) => A_i(16), IN0(15) => 
                           A_i(15), IN0(14) => A_i(14), IN0(13) => A_i(13), 
                           IN0(12) => A_i(12), IN0(11) => A_i(11), IN0(10) => 
                           A_i(10), IN0(9) => A_i(9), IN0(8) => A_i(8), IN0(7) 
                           => A_i(7), IN0(6) => A_i(6), IN0(5) => A_i(5), 
                           IN0(4) => A_i(4), IN0(3) => A_i(3), IN0(2) => A_i(2)
                           , IN0(1) => A_i(1), IN0(0) => A_i(0), IN1(31) => 
                           FW_X_i(31), IN1(30) => FW_X_i(30), IN1(29) => 
                           FW_X_i(29), IN1(28) => FW_X_i(28), IN1(27) => 
                           FW_X_i(27), IN1(26) => FW_X_i(26), IN1(25) => 
                           FW_X_i(25), IN1(24) => FW_X_i(24), IN1(23) => 
                           FW_X_i(23), IN1(22) => FW_X_i(22), IN1(21) => 
                           FW_X_i(21), IN1(20) => FW_X_i(20), IN1(19) => 
                           FW_X_i(19), IN1(18) => FW_X_i(18), IN1(17) => 
                           FW_X_i(17), IN1(16) => FW_X_i(16), IN1(15) => 
                           FW_X_i(15), IN1(14) => FW_X_i(14), IN1(13) => 
                           FW_X_i(13), IN1(12) => FW_X_i(12), IN1(11) => 
                           FW_X_i(11), IN1(10) => FW_X_i(10), IN1(9) => 
                           FW_X_i(9), IN1(8) => FW_X_i(8), IN1(7) => FW_X_i(7),
                           IN1(6) => FW_X_i(6), IN1(5) => FW_X_i(5), IN1(4) => 
                           FW_X_i(4), IN1(3) => FW_X_i(3), IN1(2) => FW_X_i(2),
                           IN1(1) => FW_X_i(1), IN1(0) => FW_X_i(0), IN2(31) =>
                           FW_W_i(31), IN2(30) => FW_W_i(30), IN2(29) => 
                           FW_W_i(29), IN2(28) => FW_W_i(28), IN2(27) => 
                           FW_W_i(27), IN2(26) => FW_W_i(26), IN2(25) => 
                           FW_W_i(25), IN2(24) => FW_W_i(24), IN2(23) => 
                           FW_W_i(23), IN2(22) => FW_W_i(22), IN2(21) => 
                           FW_W_i(21), IN2(20) => FW_W_i(20), IN2(19) => 
                           FW_W_i(19), IN2(18) => FW_W_i(18), IN2(17) => 
                           FW_W_i(17), IN2(16) => FW_W_i(16), IN2(15) => 
                           FW_W_i(15), IN2(14) => FW_W_i(14), IN2(13) => 
                           FW_W_i(13), IN2(12) => FW_W_i(12), IN2(11) => 
                           FW_W_i(11), IN2(10) => FW_W_i(10), IN2(9) => 
                           FW_W_i(9), IN2(8) => FW_W_i(8), IN2(7) => FW_W_i(7),
                           IN2(6) => FW_W_i(6), IN2(5) => FW_W_i(5), IN2(4) => 
                           FW_W_i(4), IN2(3) => FW_W_i(3), IN2(2) => FW_W_i(2),
                           IN2(1) => FW_W_i(1), IN2(0) => FW_W_i(0), IN3(31) =>
                           n1, IN3(30) => n1, IN3(29) => n1, IN3(28) => n1, 
                           IN3(27) => n1, IN3(26) => n1, IN3(25) => n1, IN3(24)
                           => n1, IN3(23) => n1, IN3(22) => n1, IN3(21) => n1, 
                           IN3(20) => n1, IN3(19) => n1, IN3(18) => n1, IN3(17)
                           => n1, IN3(16) => n1, IN3(15) => n1, IN3(14) => n1, 
                           IN3(13) => n1, IN3(12) => n1, IN3(11) => n1, IN3(10)
                           => n1, IN3(9) => n1, IN3(8) => n1, IN3(7) => n1, 
                           IN3(6) => n1, IN3(5) => n1, IN3(4) => n1, IN3(3) => 
                           n1, IN3(2) => n1, IN3(1) => n1, IN3(0) => n1, 
                           CTRL(1) => S_FW_A_i(1), CTRL(0) => S_FW_A_i(0), 
                           OUT1(31) => FWA2alu_31_port, OUT1(30) => 
                           FWA2alu_30_port, OUT1(29) => FWA2alu_29_port, 
                           OUT1(28) => FWA2alu_28_port, OUT1(27) => 
                           FWA2alu_27_port, OUT1(26) => FWA2alu_26_port, 
                           OUT1(25) => FWA2alu_25_port, OUT1(24) => 
                           FWA2alu_24_port, OUT1(23) => FWA2alu_23_port, 
                           OUT1(22) => FWA2alu_22_port, OUT1(21) => 
                           FWA2alu_21_port, OUT1(20) => FWA2alu_20_port, 
                           OUT1(19) => FWA2alu_19_port, OUT1(18) => 
                           FWA2alu_18_port, OUT1(17) => FWA2alu_17_port, 
                           OUT1(16) => FWA2alu_16_port, OUT1(15) => 
                           FWA2alu_15_port, OUT1(14) => FWA2alu_14_port, 
                           OUT1(13) => FWA2alu_13_port, OUT1(12) => 
                           FWA2alu_12_port, OUT1(11) => FWA2alu_11_port, 
                           OUT1(10) => FWA2alu_10_port, OUT1(9) => 
                           FWA2alu_9_port, OUT1(8) => FWA2alu_8_port, OUT1(7) 
                           => FWA2alu_7_port, OUT1(6) => FWA2alu_6_port, 
                           OUT1(5) => FWA2alu_5_port, OUT1(4) => FWA2alu_4_port
                           , OUT1(3) => FWA2alu_3_port, OUT1(2) => 
                           FWA2alu_2_port, OUT1(1) => FWA2alu_1_port, OUT1(0) 
                           => FWA2alu_0_port);
   MUX_FWB : mux41_MUX_SIZE32_1 port map( IN0(31) => MUXED_B_i(31), IN0(30) => 
                           MUXED_B_i(30), IN0(29) => MUXED_B_i(29), IN0(28) => 
                           MUXED_B_i(28), IN0(27) => MUXED_B_i(27), IN0(26) => 
                           MUXED_B_i(26), IN0(25) => MUXED_B_i(25), IN0(24) => 
                           MUXED_B_i(24), IN0(23) => MUXED_B_i(23), IN0(22) => 
                           MUXED_B_i(22), IN0(21) => MUXED_B_i(21), IN0(20) => 
                           MUXED_B_i(20), IN0(19) => MUXED_B_i(19), IN0(18) => 
                           MUXED_B_i(18), IN0(17) => MUXED_B_i(17), IN0(16) => 
                           MUXED_B_i(16), IN0(15) => MUXED_B_i(15), IN0(14) => 
                           MUXED_B_i(14), IN0(13) => MUXED_B_i(13), IN0(12) => 
                           MUXED_B_i(12), IN0(11) => MUXED_B_i(11), IN0(10) => 
                           MUXED_B_i(10), IN0(9) => MUXED_B_i(9), IN0(8) => 
                           MUXED_B_i(8), IN0(7) => MUXED_B_i(7), IN0(6) => 
                           MUXED_B_i(6), IN0(5) => MUXED_B_i(5), IN0(4) => 
                           MUXED_B_i(4), IN0(3) => MUXED_B_i(3), IN0(2) => 
                           MUXED_B_i(2), IN0(1) => MUXED_B_i(1), IN0(0) => 
                           MUXED_B_i(0), IN1(31) => FW_X_i(31), IN1(30) => 
                           FW_X_i(30), IN1(29) => FW_X_i(29), IN1(28) => 
                           FW_X_i(28), IN1(27) => FW_X_i(27), IN1(26) => 
                           FW_X_i(26), IN1(25) => FW_X_i(25), IN1(24) => 
                           FW_X_i(24), IN1(23) => FW_X_i(23), IN1(22) => 
                           FW_X_i(22), IN1(21) => FW_X_i(21), IN1(20) => 
                           FW_X_i(20), IN1(19) => FW_X_i(19), IN1(18) => 
                           FW_X_i(18), IN1(17) => FW_X_i(17), IN1(16) => 
                           FW_X_i(16), IN1(15) => FW_X_i(15), IN1(14) => 
                           FW_X_i(14), IN1(13) => FW_X_i(13), IN1(12) => 
                           FW_X_i(12), IN1(11) => FW_X_i(11), IN1(10) => 
                           FW_X_i(10), IN1(9) => FW_X_i(9), IN1(8) => FW_X_i(8)
                           , IN1(7) => FW_X_i(7), IN1(6) => FW_X_i(6), IN1(5) 
                           => FW_X_i(5), IN1(4) => FW_X_i(4), IN1(3) => 
                           FW_X_i(3), IN1(2) => FW_X_i(2), IN1(1) => FW_X_i(1),
                           IN1(0) => FW_X_i(0), IN2(31) => FW_W_i(31), IN2(30) 
                           => FW_W_i(30), IN2(29) => FW_W_i(29), IN2(28) => 
                           FW_W_i(28), IN2(27) => FW_W_i(27), IN2(26) => 
                           FW_W_i(26), IN2(25) => FW_W_i(25), IN2(24) => 
                           FW_W_i(24), IN2(23) => FW_W_i(23), IN2(22) => 
                           FW_W_i(22), IN2(21) => FW_W_i(21), IN2(20) => 
                           FW_W_i(20), IN2(19) => FW_W_i(19), IN2(18) => 
                           FW_W_i(18), IN2(17) => FW_W_i(17), IN2(16) => 
                           FW_W_i(16), IN2(15) => FW_W_i(15), IN2(14) => 
                           FW_W_i(14), IN2(13) => FW_W_i(13), IN2(12) => 
                           FW_W_i(12), IN2(11) => FW_W_i(11), IN2(10) => 
                           FW_W_i(10), IN2(9) => FW_W_i(9), IN2(8) => FW_W_i(8)
                           , IN2(7) => FW_W_i(7), IN2(6) => FW_W_i(6), IN2(5) 
                           => FW_W_i(5), IN2(4) => FW_W_i(4), IN2(3) => 
                           FW_W_i(3), IN2(2) => FW_W_i(2), IN2(1) => FW_W_i(1),
                           IN2(0) => FW_W_i(0), IN3(31) => n1, IN3(30) => n1, 
                           IN3(29) => n1, IN3(28) => n1, IN3(27) => n1, IN3(26)
                           => n1, IN3(25) => n1, IN3(24) => n1, IN3(23) => n1, 
                           IN3(22) => n1, IN3(21) => n1, IN3(20) => n1, IN3(19)
                           => n1, IN3(18) => n1, IN3(17) => n1, IN3(16) => n1, 
                           IN3(15) => n1, IN3(14) => n1, IN3(13) => n1, IN3(12)
                           => n1, IN3(11) => n1, IN3(10) => n1, IN3(9) => n1, 
                           IN3(8) => n1, IN3(7) => n1, IN3(6) => n1, IN3(5) => 
                           n1, IN3(4) => n1, IN3(3) => n1, IN3(2) => n1, IN3(1)
                           => n1, IN3(0) => n1, CTRL(1) => S_FW_B_i(1), CTRL(0)
                           => S_FW_B_i(0), OUT1(31) => muxed_B_31_port, 
                           OUT1(30) => muxed_B_30_port, OUT1(29) => 
                           muxed_B_29_port, OUT1(28) => muxed_B_28_port, 
                           OUT1(27) => muxed_B_27_port, OUT1(26) => 
                           muxed_B_26_port, OUT1(25) => muxed_B_25_port, 
                           OUT1(24) => muxed_B_24_port, OUT1(23) => 
                           muxed_B_23_port, OUT1(22) => muxed_B_22_port, 
                           OUT1(21) => muxed_B_21_port, OUT1(20) => 
                           muxed_B_20_port, OUT1(19) => muxed_B_19_port, 
                           OUT1(18) => muxed_B_18_port, OUT1(17) => 
                           muxed_B_17_port, OUT1(16) => muxed_B_16_port, 
                           OUT1(15) => muxed_B_15_port, OUT1(14) => 
                           muxed_B_14_port, OUT1(13) => muxed_B_13_port, 
                           OUT1(12) => muxed_B_12_port, OUT1(11) => 
                           muxed_B_11_port, OUT1(10) => muxed_B_10_port, 
                           OUT1(9) => muxed_B_9_port, OUT1(8) => muxed_B_8_port
                           , OUT1(7) => muxed_B_7_port, OUT1(6) => 
                           muxed_B_6_port, OUT1(5) => muxed_B_5_port, OUT1(4) 
                           => muxed_B_4_port, OUT1(3) => muxed_B_3_port, 
                           OUT1(2) => muxed_B_2_port, OUT1(1) => muxed_B_1_port
                           , OUT1(0) => muxed_B_0_port);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity execute_regs is

   port( X_i, S_i : in std_logic_vector (31 downto 0);  D2_i : in 
         std_logic_vector (4 downto 0);  X_o, S_o : out std_logic_vector (31 
         downto 0);  D2_o : out std_logic_vector (4 downto 0);  stall_i, clk, 
         rst : in std_logic);

end execute_regs;

architecture SYN_struct of execute_regs is

   component ff32_en_SIZE5_1
      port( D : in std_logic_vector (4 downto 0);  en, clk, rst : in std_logic;
            Q : out std_logic_vector (4 downto 0));
   end component;
   
   component ff32_en_SIZE32_2
      port( D : in std_logic_vector (31 downto 0);  en, clk, rst : in std_logic
            ;  Q : out std_logic_vector (31 downto 0));
   end component;
   
   component ff32_en_SIZE32_3
      port( D : in std_logic_vector (31 downto 0);  en, clk, rst : in std_logic
            ;  Q : out std_logic_vector (31 downto 0));
   end component;
   
   signal n2 : std_logic;

begin
   
   X : ff32_en_SIZE32_3 port map( D(31) => X_i(31), D(30) => X_i(30), D(29) => 
                           X_i(29), D(28) => X_i(28), D(27) => X_i(27), D(26) 
                           => X_i(26), D(25) => X_i(25), D(24) => X_i(24), 
                           D(23) => X_i(23), D(22) => X_i(22), D(21) => X_i(21)
                           , D(20) => X_i(20), D(19) => X_i(19), D(18) => 
                           X_i(18), D(17) => X_i(17), D(16) => X_i(16), D(15) 
                           => X_i(15), D(14) => X_i(14), D(13) => X_i(13), 
                           D(12) => X_i(12), D(11) => X_i(11), D(10) => X_i(10)
                           , D(9) => X_i(9), D(8) => X_i(8), D(7) => X_i(7), 
                           D(6) => X_i(6), D(5) => X_i(5), D(4) => X_i(4), D(3)
                           => X_i(3), D(2) => X_i(2), D(1) => X_i(1), D(0) => 
                           X_i(0), en => n2, clk => clk, rst => rst, Q(31) => 
                           X_o(31), Q(30) => X_o(30), Q(29) => X_o(29), Q(28) 
                           => X_o(28), Q(27) => X_o(27), Q(26) => X_o(26), 
                           Q(25) => X_o(25), Q(24) => X_o(24), Q(23) => X_o(23)
                           , Q(22) => X_o(22), Q(21) => X_o(21), Q(20) => 
                           X_o(20), Q(19) => X_o(19), Q(18) => X_o(18), Q(17) 
                           => X_o(17), Q(16) => X_o(16), Q(15) => X_o(15), 
                           Q(14) => X_o(14), Q(13) => X_o(13), Q(12) => X_o(12)
                           , Q(11) => X_o(11), Q(10) => X_o(10), Q(9) => X_o(9)
                           , Q(8) => X_o(8), Q(7) => X_o(7), Q(6) => X_o(6), 
                           Q(5) => X_o(5), Q(4) => X_o(4), Q(3) => X_o(3), Q(2)
                           => X_o(2), Q(1) => X_o(1), Q(0) => X_o(0));
   S : ff32_en_SIZE32_2 port map( D(31) => S_i(31), D(30) => S_i(30), D(29) => 
                           S_i(29), D(28) => S_i(28), D(27) => S_i(27), D(26) 
                           => S_i(26), D(25) => S_i(25), D(24) => S_i(24), 
                           D(23) => S_i(23), D(22) => S_i(22), D(21) => S_i(21)
                           , D(20) => S_i(20), D(19) => S_i(19), D(18) => 
                           S_i(18), D(17) => S_i(17), D(16) => S_i(16), D(15) 
                           => S_i(15), D(14) => S_i(14), D(13) => S_i(13), 
                           D(12) => S_i(12), D(11) => S_i(11), D(10) => S_i(10)
                           , D(9) => S_i(9), D(8) => S_i(8), D(7) => S_i(7), 
                           D(6) => S_i(6), D(5) => S_i(5), D(4) => S_i(4), D(3)
                           => S_i(3), D(2) => S_i(2), D(1) => S_i(1), D(0) => 
                           S_i(0), en => n2, clk => clk, rst => rst, Q(31) => 
                           S_o(31), Q(30) => S_o(30), Q(29) => S_o(29), Q(28) 
                           => S_o(28), Q(27) => S_o(27), Q(26) => S_o(26), 
                           Q(25) => S_o(25), Q(24) => S_o(24), Q(23) => S_o(23)
                           , Q(22) => S_o(22), Q(21) => S_o(21), Q(20) => 
                           S_o(20), Q(19) => S_o(19), Q(18) => S_o(18), Q(17) 
                           => S_o(17), Q(16) => S_o(16), Q(15) => S_o(15), 
                           Q(14) => S_o(14), Q(13) => S_o(13), Q(12) => S_o(12)
                           , Q(11) => S_o(11), Q(10) => S_o(10), Q(9) => S_o(9)
                           , Q(8) => S_o(8), Q(7) => S_o(7), Q(6) => S_o(6), 
                           Q(5) => S_o(5), Q(4) => S_o(4), Q(3) => S_o(3), Q(2)
                           => S_o(2), Q(1) => S_o(1), Q(0) => S_o(0));
   D2 : ff32_en_SIZE5_1 port map( D(4) => D2_i(4), D(3) => D2_i(3), D(2) => 
                           D2_i(2), D(1) => D2_i(1), D(0) => D2_i(0), en => n2,
                           clk => clk, rst => rst, Q(4) => D2_o(4), Q(3) => 
                           D2_o(3), Q(2) => D2_o(2), Q(1) => D2_o(1), Q(0) => 
                           D2_o(0));
   n2 <= '1';

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity decode_regs is

   port( A_i, B_i : in std_logic_vector (31 downto 0);  rA_i, rB_i, rC_i : in 
         std_logic_vector (4 downto 0);  IMM_i : in std_logic_vector (31 downto
         0);  ALUW_i : in std_logic_vector (12 downto 0);  A_o, B_o : out 
         std_logic_vector (31 downto 0);  rA_o, rB_o, rC_o : out 
         std_logic_vector (4 downto 0);  IMM_o : out std_logic_vector (31 
         downto 0);  ALUW_o : out std_logic_vector (12 downto 0);  stall_i, clk
         , rst : in std_logic);

end decode_regs;

architecture SYN_struct of decode_regs is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component ff32_en_SIZE13
      port( D : in std_logic_vector (12 downto 0);  en, clk, rst : in std_logic
            ;  Q : out std_logic_vector (12 downto 0));
   end component;
   
   component ff32_en_SIZE32_4
      port( D : in std_logic_vector (31 downto 0);  en, clk, rst : in std_logic
            ;  Q : out std_logic_vector (31 downto 0));
   end component;
   
   component ff32_en_SIZE5_2
      port( D : in std_logic_vector (4 downto 0);  en, clk, rst : in std_logic;
            Q : out std_logic_vector (4 downto 0));
   end component;
   
   component ff32_en_SIZE5_3
      port( D : in std_logic_vector (4 downto 0);  en, clk, rst : in std_logic;
            Q : out std_logic_vector (4 downto 0));
   end component;
   
   component ff32_en_SIZE5_0
      port( D : in std_logic_vector (4 downto 0);  en, clk, rst : in std_logic;
            Q : out std_logic_vector (4 downto 0));
   end component;
   
   component ff32_en_SIZE32_5
      port( D : in std_logic_vector (31 downto 0);  en, clk, rst : in std_logic
            ;  Q : out std_logic_vector (31 downto 0));
   end component;
   
   component ff32_en_SIZE32_0
      port( D : in std_logic_vector (31 downto 0);  en, clk, rst : in std_logic
            ;  Q : out std_logic_vector (31 downto 0));
   end component;
   
   signal enable : std_logic;

begin
   
   A : ff32_en_SIZE32_0 port map( D(31) => A_i(31), D(30) => A_i(30), D(29) => 
                           A_i(29), D(28) => A_i(28), D(27) => A_i(27), D(26) 
                           => A_i(26), D(25) => A_i(25), D(24) => A_i(24), 
                           D(23) => A_i(23), D(22) => A_i(22), D(21) => A_i(21)
                           , D(20) => A_i(20), D(19) => A_i(19), D(18) => 
                           A_i(18), D(17) => A_i(17), D(16) => A_i(16), D(15) 
                           => A_i(15), D(14) => A_i(14), D(13) => A_i(13), 
                           D(12) => A_i(12), D(11) => A_i(11), D(10) => A_i(10)
                           , D(9) => A_i(9), D(8) => A_i(8), D(7) => A_i(7), 
                           D(6) => A_i(6), D(5) => A_i(5), D(4) => A_i(4), D(3)
                           => A_i(3), D(2) => A_i(2), D(1) => A_i(1), D(0) => 
                           A_i(0), en => enable, clk => clk, rst => rst, Q(31) 
                           => A_o(31), Q(30) => A_o(30), Q(29) => A_o(29), 
                           Q(28) => A_o(28), Q(27) => A_o(27), Q(26) => A_o(26)
                           , Q(25) => A_o(25), Q(24) => A_o(24), Q(23) => 
                           A_o(23), Q(22) => A_o(22), Q(21) => A_o(21), Q(20) 
                           => A_o(20), Q(19) => A_o(19), Q(18) => A_o(18), 
                           Q(17) => A_o(17), Q(16) => A_o(16), Q(15) => A_o(15)
                           , Q(14) => A_o(14), Q(13) => A_o(13), Q(12) => 
                           A_o(12), Q(11) => A_o(11), Q(10) => A_o(10), Q(9) =>
                           A_o(9), Q(8) => A_o(8), Q(7) => A_o(7), Q(6) => 
                           A_o(6), Q(5) => A_o(5), Q(4) => A_o(4), Q(3) => 
                           A_o(3), Q(2) => A_o(2), Q(1) => A_o(1), Q(0) => 
                           A_o(0));
   B : ff32_en_SIZE32_5 port map( D(31) => B_i(31), D(30) => B_i(30), D(29) => 
                           B_i(29), D(28) => B_i(28), D(27) => B_i(27), D(26) 
                           => B_i(26), D(25) => B_i(25), D(24) => B_i(24), 
                           D(23) => B_i(23), D(22) => B_i(22), D(21) => B_i(21)
                           , D(20) => B_i(20), D(19) => B_i(19), D(18) => 
                           B_i(18), D(17) => B_i(17), D(16) => B_i(16), D(15) 
                           => B_i(15), D(14) => B_i(14), D(13) => B_i(13), 
                           D(12) => B_i(12), D(11) => B_i(11), D(10) => B_i(10)
                           , D(9) => B_i(9), D(8) => B_i(8), D(7) => B_i(7), 
                           D(6) => B_i(6), D(5) => B_i(5), D(4) => B_i(4), D(3)
                           => B_i(3), D(2) => B_i(2), D(1) => B_i(1), D(0) => 
                           B_i(0), en => enable, clk => clk, rst => rst, Q(31) 
                           => B_o(31), Q(30) => B_o(30), Q(29) => B_o(29), 
                           Q(28) => B_o(28), Q(27) => B_o(27), Q(26) => B_o(26)
                           , Q(25) => B_o(25), Q(24) => B_o(24), Q(23) => 
                           B_o(23), Q(22) => B_o(22), Q(21) => B_o(21), Q(20) 
                           => B_o(20), Q(19) => B_o(19), Q(18) => B_o(18), 
                           Q(17) => B_o(17), Q(16) => B_o(16), Q(15) => B_o(15)
                           , Q(14) => B_o(14), Q(13) => B_o(13), Q(12) => 
                           B_o(12), Q(11) => B_o(11), Q(10) => B_o(10), Q(9) =>
                           B_o(9), Q(8) => B_o(8), Q(7) => B_o(7), Q(6) => 
                           B_o(6), Q(5) => B_o(5), Q(4) => B_o(4), Q(3) => 
                           B_o(3), Q(2) => B_o(2), Q(1) => B_o(1), Q(0) => 
                           B_o(0));
   rA : ff32_en_SIZE5_0 port map( D(4) => rA_i(4), D(3) => rA_i(3), D(2) => 
                           rA_i(2), D(1) => rA_i(1), D(0) => rA_i(0), en => 
                           enable, clk => clk, rst => rst, Q(4) => rA_o(4), 
                           Q(3) => rA_o(3), Q(2) => rA_o(2), Q(1) => rA_o(1), 
                           Q(0) => rA_o(0));
   rB : ff32_en_SIZE5_3 port map( D(4) => rB_i(4), D(3) => rB_i(3), D(2) => 
                           rB_i(2), D(1) => rB_i(1), D(0) => rB_i(0), en => 
                           enable, clk => clk, rst => rst, Q(4) => rB_o(4), 
                           Q(3) => rB_o(3), Q(2) => rB_o(2), Q(1) => rB_o(1), 
                           Q(0) => rB_o(0));
   rC : ff32_en_SIZE5_2 port map( D(4) => rC_i(4), D(3) => rC_i(3), D(2) => 
                           rC_i(2), D(1) => rC_i(1), D(0) => rC_i(0), en => 
                           enable, clk => clk, rst => rst, Q(4) => rC_o(4), 
                           Q(3) => rC_o(3), Q(2) => rC_o(2), Q(1) => rC_o(1), 
                           Q(0) => rC_o(0));
   IMM : ff32_en_SIZE32_4 port map( D(31) => IMM_i(31), D(30) => IMM_i(30), 
                           D(29) => IMM_i(29), D(28) => IMM_i(28), D(27) => 
                           IMM_i(27), D(26) => IMM_i(26), D(25) => IMM_i(25), 
                           D(24) => IMM_i(24), D(23) => IMM_i(23), D(22) => 
                           IMM_i(22), D(21) => IMM_i(21), D(20) => IMM_i(20), 
                           D(19) => IMM_i(19), D(18) => IMM_i(18), D(17) => 
                           IMM_i(17), D(16) => IMM_i(16), D(15) => IMM_i(15), 
                           D(14) => IMM_i(14), D(13) => IMM_i(13), D(12) => 
                           IMM_i(12), D(11) => IMM_i(11), D(10) => IMM_i(10), 
                           D(9) => IMM_i(9), D(8) => IMM_i(8), D(7) => IMM_i(7)
                           , D(6) => IMM_i(6), D(5) => IMM_i(5), D(4) => 
                           IMM_i(4), D(3) => IMM_i(3), D(2) => IMM_i(2), D(1) 
                           => IMM_i(1), D(0) => IMM_i(0), en => enable, clk => 
                           clk, rst => rst, Q(31) => IMM_o(31), Q(30) => 
                           IMM_o(30), Q(29) => IMM_o(29), Q(28) => IMM_o(28), 
                           Q(27) => IMM_o(27), Q(26) => IMM_o(26), Q(25) => 
                           IMM_o(25), Q(24) => IMM_o(24), Q(23) => IMM_o(23), 
                           Q(22) => IMM_o(22), Q(21) => IMM_o(21), Q(20) => 
                           IMM_o(20), Q(19) => IMM_o(19), Q(18) => IMM_o(18), 
                           Q(17) => IMM_o(17), Q(16) => IMM_o(16), Q(15) => 
                           IMM_o(15), Q(14) => IMM_o(14), Q(13) => IMM_o(13), 
                           Q(12) => IMM_o(12), Q(11) => IMM_o(11), Q(10) => 
                           IMM_o(10), Q(9) => IMM_o(9), Q(8) => IMM_o(8), Q(7) 
                           => IMM_o(7), Q(6) => IMM_o(6), Q(5) => IMM_o(5), 
                           Q(4) => IMM_o(4), Q(3) => IMM_o(3), Q(2) => IMM_o(2)
                           , Q(1) => IMM_o(1), Q(0) => IMM_o(0));
   ALUW : ff32_en_SIZE13 port map( D(12) => ALUW_i(12), D(11) => ALUW_i(11), 
                           D(10) => ALUW_i(10), D(9) => ALUW_i(9), D(8) => 
                           ALUW_i(8), D(7) => ALUW_i(7), D(6) => ALUW_i(6), 
                           D(5) => ALUW_i(5), D(4) => ALUW_i(4), D(3) => 
                           ALUW_i(3), D(2) => ALUW_i(2), D(1) => ALUW_i(1), 
                           D(0) => ALUW_i(0), en => enable, clk => clk, rst => 
                           rst, Q(12) => ALUW_o(12), Q(11) => ALUW_o(11), Q(10)
                           => ALUW_o(10), Q(9) => ALUW_o(9), Q(8) => ALUW_o(8),
                           Q(7) => ALUW_o(7), Q(6) => ALUW_o(6), Q(5) => 
                           ALUW_o(5), Q(4) => ALUW_o(4), Q(3) => ALUW_o(3), 
                           Q(2) => ALUW_o(2), Q(1) => ALUW_o(1), Q(0) => 
                           ALUW_o(0));
   U1 : INV_X1 port map( A => stall_i, ZN => enable);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity dlx_regfile is

   port( Clk, Rst, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, 
         ADD_RD2 : in std_logic_vector (4 downto 0);  DATAIN : in 
         std_logic_vector (31 downto 0);  OUT1, OUT2 : out std_logic_vector (31
         downto 0));

end dlx_regfile;

architecture SYN_A of dlx_regfile is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_dlx_regfile_1
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_dlx_regfile_2
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_dlx_regfile_3
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_dlx_regfile_4
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_dlx_regfile_5
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_dlx_regfile_6
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_dlx_regfile_7
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_dlx_regfile_8
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_dlx_regfile_9
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_dlx_regfile_10
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_dlx_regfile_11
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_dlx_regfile_12
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_dlx_regfile_13
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_dlx_regfile_14
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_dlx_regfile_15
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_dlx_regfile_16
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_dlx_regfile_17
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_dlx_regfile_18
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_dlx_regfile_19
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_dlx_regfile_20
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_dlx_regfile_21
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_dlx_regfile_22
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_dlx_regfile_23
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_dlx_regfile_24
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_dlx_regfile_25
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_dlx_regfile_26
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_dlx_regfile_27
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_dlx_regfile_28
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_dlx_regfile_29
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_dlx_regfile_30
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_dlx_regfile_31
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_dlx_regfile_32
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_dlx_regfile_33
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_dlx_regfile_0
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal N2503, N2567, N2631, N2695, N2759, N2823, N2887, N2951, N3015, N3079,
      N3143, N3207, N3271, N3335, N3399, N3463, N3527, N3591, N3655, N3719, 
      N3783, N3847, N3911, N3975, N4039, N4103, N4167, N4231, N4295, N4359, 
      N4423, N4490, N4492, N4494, N4496, N4498, N4500, N4502, N4504, N4506, 
      N4508, N4510, N4512, N4514, N4516, N4518, N4520, N4522, N4524, N4526, 
      N4528, N4530, N4532, N4534, N4536, N4538, N4540, N4542, N4544, N4546, 
      N4548, N4550, N4552, N4554, N4556, N4558, N4560, N4562, N4564, N4566, 
      N4568, N4570, N4572, N4574, N4576, N4578, N4580, N4582, N4584, N4586, 
      N4588, N4590, N4592, N4594, N4596, N4598, N4600, N4602, N4604, N4606, 
      N4608, N4610, N4612, N4614, N4615, N4616, net199403, net199408, net199413
      , net199418, net199423, net199428, net199433, net199438, net199443, 
      net199448, net199453, net199458, net199463, net199468, net199473, 
      net199478, net199483, net199488, net199493, net199498, net199503, 
      net199508, net199513, net199518, net199523, net199528, net199533, 
      net199538, net199543, net199548, net199553, net199558, net199563, 
      net199568, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17
      , n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, 
      n32, n33, n34, n35, n36, n38, n40, n42, n44, n46, n48, n50, n52, n54, n56
      , n58, n60, n62, n64, n66, n68, n70, n72, n74, n76, n78, n80, n82, n84, 
      n86, n88, n90, n92, n94, n96, n98, n1094, n1150, n1172, n1194, n1216, 
      n1238, n1260, n1282, n1304, n1326, n1348, n1370, n1392, n1414, n1436, 
      n1458, n1480, n1502, n1524, n1546, n1568, n1590, n1612, n1634, n1656, 
      n1678, n1700, n1722, n1744, n1766, n1788, n1810, n1, n2, n3, n37, n39, 
      n41, n43, n45, n47, n49, n51, n53, n55, n57, n59, n61, n63, n65, n67, n69
      , n71, n73, n75, n77, n79, n81, n83, n85, n87, n89, n91, n93, n95, n97, 
      n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, 
      n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, 
      n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, 
      n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, 
      n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, 
      n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, 
      n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, 
      n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, 
      n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, 
      n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, 
      n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, 
      n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, 
      n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, 
      n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, 
      n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, 
      n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, 
      n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, 
      n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, 
      n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, 
      n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, 
      n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, 
      n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, 
      n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, 
      n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, 
      n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, 
      n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, 
      n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, 
      n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, 
      n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, 
      n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, 
      n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, 
      n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, 
      n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, 
      n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, 
      n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, 
      n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, 
      n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, 
      n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, 
      n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, 
      n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, 
      n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, 
      n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, 
      n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, 
      n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, 
      n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, 
      n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, 
      n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, 
      n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, 
      n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, 
      n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, 
      n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, 
      n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, 
      n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, 
      n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, 
      n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, 
      n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, 
      n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, 
      n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, 
      n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, 
      n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, 
      n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, 
      n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, 
      n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, 
      n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, 
      n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, 
      n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, 
      n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, 
      n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, 
      n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, 
      n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, 
      n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, 
      n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, 
      n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, 
      n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, 
      n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, 
      n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, 
      n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, 
      n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, 
      n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, 
      n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, 
      n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, 
      n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, 
      n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, 
      n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, 
      n1089, n1090, n1091, n1092, n1093, n1095, n1096, n1097, n1098, n1099, 
      n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, 
      n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, 
      n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, 
      n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, 
      n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, 
      n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, 
      n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, 
      n1171, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, 
      n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, 
      n1192, n1193, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, 
      n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, 
      n1213, n1214, n1215, n1217, n1218, n1219, n1220, n1221, n1222, n1223, 
      n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, 
      n1234, n1235, n1236, n1237, n1239, n1240, n1241, n1242, n1243, n1244, 
      n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, 
      n1255, n1256, n1257, n1258, n1259, n1261, n1262, n1263, n1264, n1265, 
      n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, 
      n1276, n1277, n1278, n1279, n1280, n1281, n1283, n1284, n1285, n1286, 
      n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, 
      n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1305, n1306, n1307, 
      n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, 
      n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1327, n1328, 
      n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, 
      n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1349, 
      n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, 
      n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, 
      n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, 
      n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, 
      n1391, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, 
      n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, 
      n1412, n1413, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, 
      n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, 
      n1433, n1434, n1435, n1437, n1438, n1439, n1440, n1441, n1442, n1443, 
      n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, 
      n1454, n1455, n1456, n1457, n1459, n1460, n1461, n1462, n1463, n1464, 
      n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, 
      n1475, n1476, n1477, n1478, n1479, n1481, n1482, n1483, n1484, n1485, 
      n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, 
      n1496, n1497, n1498, n1499, n1500, n1501, n1503, n1504, n1505, n1506, 
      n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, 
      n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1525, n1526, n1527, 
      n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, 
      n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1547, n1548, 
      n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, 
      n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1569, 
      n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, 
      n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, 
      n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, 
      n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, 
      n1611, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, 
      n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, 
      n1632, n1633, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, 
      n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, 
      n1653, n1654, n1655, n1657, n1658, n1659, n1660, n1661, n1662, n1663, 
      n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, 
      n1674, n1675, n1676, n1677, n1679, n1680, n1681, n1682, n1683, n1684, 
      n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, 
      n1695, n1696, n1697, n1698, n1699, n1701, n1702, n1703, n1704, n1705, 
      n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, 
      n1716, n1717, n1718, n1719, n1720, n1721, n1723, n1724, n1725, n1726, 
      n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, 
      n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1745, n1746, n1747, 
      n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, 
      n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1767, n1768, 
      n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, 
      n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1789, 
      n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, 
      n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, 
      n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, 
      n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, 
      n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, 
      n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, 
      n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, 
      n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, 
      n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, 
      n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, 
      n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, 
      n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, 
      n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, 
      n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, 
      n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, 
      n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, 
      n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, 
      n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, 
      n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, 
      n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, 
      n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, 
      n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, 
      n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, 
      n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, 
      n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, 
      n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, 
      n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, 
      n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, 
      n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, 
      n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, 
      n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, 
      n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, 
      n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, 
      n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, 
      n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, 
      n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, 
      n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, 
      n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, 
      n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, 
      n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, 
      n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, 
      n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, 
      n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, 
      n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, 
      n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, 
      n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, 
      n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, 
      n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, 
      n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, 
      n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, 
      n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, 
      n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, 
      n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, 
      n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, 
      n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, 
      n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, 
      n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, 
      n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, 
      n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, 
      n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, 
      n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, 
      n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, 
      n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, 
      n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, 
      n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, 
      n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, 
      n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, 
      n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, 
      n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, 
      n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, 
      n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, 
      n2501, n2502, n2503_port, n2504, n2505, n2506, n2507, n2508, n2509, n2510
      , n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, 
      n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, 
      n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, 
      n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, 
      n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, 
      n2561, n2562, n2563, n2564, n2565, n2566, n2567_port, n2568, n2569, n2570
      , n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, 
      n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, 
      n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, 
      n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, 
      net245099, net245100, net245101, net245102, net245103, net245104, 
      net245105, net245106, net245107, net245108, net245109, net245110, 
      net245111, net245112, net245113, net245114, net245115, net245116, 
      net245117, net245118, net245119, net245120, net245121, net245122, 
      net245123, net245124, net245125, net245126, net245127, net245128, 
      net245129, net245130, net245131, net245132, net245133, net245134, 
      net245135, net245136, net245137, net245138, net245139, net245140, 
      net245141, net245142, net245143, net245144, net245145, net245146, 
      net245147, net245148, net245149, net245150, net245151, net245152, 
      net245153, net245154, net245155, net245156, net245157, net245158, 
      net245159, net245160, net245161, net245162, net245163, net245164, 
      net245165, net245166, net245167, net245168, net245169, net245170, 
      net245171, net245172, net245173, net245174, net245175, net245176, 
      net245177, net245178, net245179, net245180, net245181, net245182, 
      net245183, net245184, net245185, net245186, net245187, net245188, 
      net245189, net245190, net245191, net245192, net245193, net245194, 
      net245195, net245196, net245197, net245198, net245199, net245200, 
      net245201, net245202, net245203, net245204, net245205, net245206, 
      net245207, net245208, net245209, net245210, net245211, net245212, 
      net245213, net245214, net245215, net245216, net245217, net245218, 
      net245219, net245220, net245221, net245222, net245223, net245224, 
      net245225, net245226, net245227, net245228, net245229, net245230, 
      net245231, net245232, net245233, net245234, net245235, net245236, 
      net245237, net245238, net245239, net245240, net245241, net245242, 
      net245243, net245244, net245245, net245246, net245247, net245248, 
      net245249, net245250, net245251, net245252, net245253, net245254, 
      net245255, net245256, net245257, net245258, net245259, net245260, 
      net245261, net245262, net245263, net245264, net245265, net245266, 
      net245267, net245268, net245269, net245270, net245271, net245272, 
      net245273, net245274, net245275, net245276, net245277, net245278, 
      net245279, net245280, net245281, net245282, net245283, net245284, 
      net245285, net245286, net245287, net245288, net245289, net245290, 
      net245291, net245292, net245293, net245294, net245295, net245296, 
      net245297, net245298, net245299, net245300, net245301, net245302, 
      net245303, net245304, net245305, net245306, net245307, net245308, 
      net245309, net245310, net245311, net245312, net245313, net245314, 
      net245315, net245316, net245317, net245318, net245319, net245320, 
      net245321, net245322, net245323, net245324, net245325, net245326, 
      net245327, net245328, net245329, net245330, net245331, net245332, 
      net245333, net245334, net245335, net245336, net245337, net245338, 
      net245339, net245340, net245341, net245342, net245343, net245344, 
      net245345, net245346, net245347, net245348, net245349, net245350, 
      net245351, net245352, net245353, net245354, net245355, net245356, 
      net245357, net245358, net245359, net245360, net245361, net245362, 
      net245363, net245364, net245365, net245366, net245367, net245368, 
      net245369, net245370, net245371, net245372, net245373, net245374, 
      net245375, net245376, net245377, net245378, net245379, net245380, 
      net245381, net245382, net245383, net245384, net245385, net245386, 
      net245387, net245388, net245389, net245390, net245391, net245392, 
      net245393, net245394, net245395, net245396, net245397, net245398, 
      net245399, net245400, net245401, net245402, net245403, net245404, 
      net245405, net245406, net245407, net245408, net245409, net245410, 
      net245411, net245412, net245413, net245414, net245415, net245416, 
      net245417, net245418, net245419, net245420, net245421, net245422, 
      net245423, net245424, net245425, net245426, net245427, net245428, 
      net245429, net245430, net245431, net245432, net245433, net245434, 
      net245435, net245436, net245437, net245438, net245439, net245440, 
      net245441, net245442, net245443, net245444, net245445, net245446, 
      net245447, net245448, net245449, net245450, net245451, net245452, 
      net245453, net245454, net245455, net245456, net245457, net245458, 
      net245459, net245460, net245461, net245462, net245463, net245464, 
      net245465, net245466, net245467, net245468, net245469, net245470, 
      net245471, net245472, net245473, net245474, net245475, net245476, 
      net245477, net245478, net245479, net245480, net245481, net245482, 
      net245483, net245484, net245485, net245486, net245487, net245488, 
      net245489, net245490, net245491, net245492, net245493, net245494, 
      net245495, net245496, net245497, net245498, net245499, net245500, 
      net245501, net245502, net245503, net245504, net245505, net245506, 
      net245507, net245508, net245509, net245510, net245511, net245512, 
      net245513, net245514, net245515, net245516, net245517, net245518, 
      net245519, net245520, net245521, net245522, net245523, net245524, 
      net245525, net245526, net245527, net245528, net245529, net245530, 
      net245531, net245532, net245533, net245534, net245535, net245536, 
      net245537, net245538, net245539, net245540, net245541, net245542, 
      net245543, net245544, net245545, net245546, net245547, net245548, 
      net245549, net245550, net245551, net245552, net245553, net245554, 
      net245555, net245556, net245557, net245558, net245559, net245560, 
      net245561, net245562, net245563, net245564, net245565, net245566, 
      net245567, net245568, net245569, net245570, net245571, net245572, 
      net245573, net245574, net245575, net245576, net245577, net245578, 
      net245579, net245580, net245581, net245582, net245583, net245584, 
      net245585, net245586, net245587, net245588, net245589, net245590, 
      net245591, net245592, net245593, net245594, net245595, net245596, 
      net245597, net245598, net245599, net245600, net245601, net245602, 
      net245603, net245604, net245605, net245606, net245607, net245608, 
      net245609, net245610, net245611, net245612, net245613, net245614, 
      net245615, net245616, net245617, net245618, net245619, net245620, 
      net245621, net245622, net245623, net245624, net245625, net245626, 
      net245627, net245628, net245629, net245630, net245631, net245632, 
      net245633, net245634, net245635, net245636, net245637, net245638, 
      net245639, net245640, net245641, net245642, net245643, net245644, 
      net245645, net245646, net245647, net245648, net245649, net245650, 
      net245651, net245652, net245653, net245654, net245655, net245656, 
      net245657, net245658, net245659, net245660, net245661, net245662, 
      net245663, net245664, net245665, net245666, net245667, net245668, 
      net245669, net245670, net245671, net245672, net245673, net245674, 
      net245675, net245676, net245677, net245678, net245679, net245680, 
      net245681, net245682, net245683, net245684, net245685, net245686, 
      net245687, net245688, net245689, net245690, net245691, net245692, 
      net245693, net245694, net245695, net245696, net245697, net245698, 
      net245699, net245700, net245701, net245702, net245703, net245704, 
      net245705, net245706, net245707, net245708, net245709, net245710, 
      net245711, net245712, net245713, net245714, net245715, net245716, 
      net245717, net245718, net245719, net245720, net245721, net245722, 
      net245723, net245724, net245725, net245726, net245727, net245728, 
      net245729, net245730, net245731, net245732, net245733, net245734, 
      net245735, net245736, net245737, net245738, net245739, net245740, 
      net245741, net245742, net245743, net245744, net245745, net245746, 
      net245747, net245748, net245749, net245750, net245751, net245752, 
      net245753, net245754, net245755, net245756, net245757, net245758, 
      net245759, net245760, net245761, net245762, net245763, net245764, 
      net245765, net245766, net245767, net245768, net245769, net245770, 
      net245771, net245772, net245773, net245774, net245775, net245776, 
      net245777, net245778, net245779, net245780, net245781, net245782, 
      net245783, net245784, net245785, net245786, net245787, net245788, 
      net245789, net245790, net245791, net245792, net245793, net245794, 
      net245795, net245796, net245797, net245798, net245799, net245800, 
      net245801, net245802, net245803, net245804, net245805, net245806, 
      net245807, net245808, net245809, net245810, net245811, net245812, 
      net245813, net245814, net245815, net245816, net245817, net245818, 
      net245819, net245820, net245821, net245822, net245823, net245824, 
      net245825, net245826, net245827, net245828, net245829, net245830, 
      net245831, net245832, net245833, net245834, net245835, net245836, 
      net245837, net245838, net245839, net245840, net245841, net245842, 
      net245843, net245844, net245845, net245846, net245847, net245848, 
      net245849, net245850, net245851, net245852, net245853, net245854, 
      net245855, net245856, net245857, net245858, net245859, net245860, 
      net245861, net245862, net245863, net245864, net245865, net245866, 
      net245867, net245868, net245869, net245870, net245871, net245872, 
      net245873, net245874, net245875, net245876, net245877, net245878, 
      net245879, net245880, net245881, net245882, net245883, net245884, 
      net245885, net245886, net245887, net245888, net245889, net245890, 
      net245891, net245892, net245893, net245894, net245895, net245896, 
      net245897, net245898, net245899, net245900, net245901, net245902, 
      net245903, net245904, net245905, net245906, net245907, net245908, 
      net245909, net245910, net245911, net245912, net245913, net245914, 
      net245915, net245916, net245917, net245918, net245919, net245920, 
      net245921, net245922, net245923, net245924, net245925, net245926, 
      net245927, net245928, net245929, net245930, net245931, net245932, 
      net245933, net245934, net245935, net245936, net245937, net245938, 
      net245939, net245940, net245941, net245942, net245943, net245944, 
      net245945, net245946, net245947, net245948, net245949, net245950, 
      net245951, net245952, net245953, net245954, net245955, net245956, 
      net245957, net245958, net245959, net245960, net245961, net245962, 
      net245963, net245964, net245965, net245966, net245967, net245968, 
      net245969, net245970, net245971, net245972, net245973, net245974, 
      net245975, net245976, net245977, net245978, net245979, net245980, 
      net245981, net245982, net245983, net245984, net245985, net245986, 
      net245987, net245988, net245989, net245990, net245991, net245992, 
      net245993, net245994, net245995, net245996, net245997, net245998, 
      net245999, net246000, net246001, net246002, net246003, net246004, 
      net246005, net246006, net246007, net246008, net246009, net246010, 
      net246011, net246012, net246013, net246014, net246015, net246016, 
      net246017, net246018, net246019, net246020, net246021, net246022, 
      net246023, net246024, net246025, net246026, net246027, net246028, 
      net246029, net246030, net246031, net246032, net246033, net246034, 
      net246035, net246036, net246037, net246038, net246039, net246040, 
      net246041, net246042, net246043, net246044, net246045, net246046, 
      net246047, net246048, net246049, net246050, net246051, net246052, 
      net246053, net246054, net246055, net246056, net246057, net246058, 
      net246059, net246060, net246061, net246062, net246063, net246064, 
      net246065, net246066, net246067, net246068, net246069, net246070, 
      net246071, net246072, net246073, net246074, net246075, net246076, 
      net246077, net246078, net246079, net246080, net246081, net246082, 
      net246083, net246084, net246085, net246086, net246087, net246088, 
      net246089, net246090, net246091, net246092, net246093, net246094, 
      net246095, net246096, net246097, net246098, net246099, net246100, 
      net246101, net246102, net246103, net246104, net246105, net246106, 
      net246107, net246108, net246109, net246110, net246111, net246112, 
      net246113, net246114, net246115, net246116, net246117, net246118, 
      net246119, net246120, net246121, net246122 : std_logic;

begin
   
   REGISTERS_reg_0_31_inst : DFF_X1 port map( D => n1094, CK => net199408, Q =>
                           n178, QN => net246122);
   REGISTERS_reg_0_30_inst : DFF_X1 port map( D => n1150, CK => net199408, Q =>
                           n177, QN => net246121);
   REGISTERS_reg_0_29_inst : DFF_X1 port map( D => n1172, CK => net199408, Q =>
                           n175, QN => net246120);
   REGISTERS_reg_0_28_inst : DFF_X1 port map( D => n1194, CK => net199408, Q =>
                           n174, QN => net246119);
   REGISTERS_reg_0_27_inst : DFF_X1 port map( D => n1216, CK => net199408, Q =>
                           n173, QN => net246118);
   REGISTERS_reg_0_26_inst : DFF_X1 port map( D => n1238, CK => net199408, Q =>
                           n172, QN => net246117);
   REGISTERS_reg_0_25_inst : DFF_X1 port map( D => n1260, CK => net199408, Q =>
                           n171, QN => net246116);
   REGISTERS_reg_0_24_inst : DFF_X1 port map( D => n1282, CK => net199408, Q =>
                           n170, QN => net246115);
   REGISTERS_reg_0_23_inst : DFF_X1 port map( D => n1304, CK => net199408, Q =>
                           n169, QN => net246114);
   REGISTERS_reg_0_22_inst : DFF_X1 port map( D => n1326, CK => net199408, Q =>
                           n168, QN => net246113);
   REGISTERS_reg_0_21_inst : DFF_X1 port map( D => n1348, CK => net199408, Q =>
                           n167, QN => net246112);
   REGISTERS_reg_0_20_inst : DFF_X1 port map( D => n1370, CK => net199408, Q =>
                           n166, QN => net246111);
   REGISTERS_reg_0_19_inst : DFF_X1 port map( D => n1392, CK => net199408, Q =>
                           n164, QN => net246110);
   REGISTERS_reg_0_18_inst : DFF_X1 port map( D => n1414, CK => net199408, Q =>
                           n163, QN => net246109);
   REGISTERS_reg_0_17_inst : DFF_X1 port map( D => n1436, CK => net199408, Q =>
                           n162, QN => net246108);
   REGISTERS_reg_0_16_inst : DFF_X1 port map( D => n1458, CK => net199408, Q =>
                           n161, QN => net246107);
   REGISTERS_reg_0_15_inst : DFF_X1 port map( D => n1480, CK => net199408, Q =>
                           n160, QN => net246106);
   REGISTERS_reg_0_14_inst : DFF_X1 port map( D => n1502, CK => net199408, Q =>
                           n159, QN => net246105);
   REGISTERS_reg_0_13_inst : DFF_X1 port map( D => n1524, CK => net199408, Q =>
                           n158, QN => net246104);
   REGISTERS_reg_0_12_inst : DFF_X1 port map( D => n1546, CK => net199408, Q =>
                           n157, QN => net246103);
   REGISTERS_reg_0_11_inst : DFF_X1 port map( D => n1568, CK => net199408, Q =>
                           n156, QN => net246102);
   REGISTERS_reg_0_10_inst : DFF_X1 port map( D => n1590, CK => net199408, Q =>
                           n155, QN => net246101);
   REGISTERS_reg_0_9_inst : DFF_X1 port map( D => n1612, CK => net199408, Q => 
                           n153, QN => net246100);
   REGISTERS_reg_0_8_inst : DFF_X1 port map( D => n1634, CK => net199408, Q => 
                           n152, QN => net246099);
   REGISTERS_reg_0_7_inst : DFF_X1 port map( D => n1656, CK => net199408, Q => 
                           n151, QN => net246098);
   REGISTERS_reg_0_6_inst : DFF_X1 port map( D => n1678, CK => net199408, Q => 
                           n150, QN => net246097);
   REGISTERS_reg_0_5_inst : DFF_X1 port map( D => n1700, CK => net199408, Q => 
                           n149, QN => net246096);
   REGISTERS_reg_0_4_inst : DFF_X1 port map( D => n1722, CK => net199408, Q => 
                           n148, QN => net246095);
   REGISTERS_reg_0_3_inst : DFF_X1 port map( D => n1744, CK => net199408, Q => 
                           n147, QN => net246094);
   REGISTERS_reg_0_2_inst : DFF_X1 port map( D => n1766, CK => net199408, Q => 
                           n146, QN => net246093);
   REGISTERS_reg_0_1_inst : DFF_X1 port map( D => n1788, CK => net199408, Q => 
                           n145, QN => net246092);
   REGISTERS_reg_0_0_inst : DFF_X1 port map( D => n1810, CK => net199408, Q => 
                           n144, QN => net246091);
   REGISTERS_reg_1_31_inst : DFF_X1 port map( D => n1094, CK => net199413, Q =>
                           n142, QN => net246090);
   REGISTERS_reg_1_30_inst : DFF_X1 port map( D => n1150, CK => net199413, Q =>
                           n141, QN => net246089);
   REGISTERS_reg_1_29_inst : DFF_X1 port map( D => n1172, CK => net199413, Q =>
                           n140, QN => net246088);
   REGISTERS_reg_1_28_inst : DFF_X1 port map( D => n1194, CK => net199413, Q =>
                           n139, QN => net246087);
   REGISTERS_reg_1_27_inst : DFF_X1 port map( D => n1216, CK => net199413, Q =>
                           n138, QN => net246086);
   REGISTERS_reg_1_26_inst : DFF_X1 port map( D => n1238, CK => net199413, Q =>
                           n137, QN => net246085);
   REGISTERS_reg_1_25_inst : DFF_X1 port map( D => n1260, CK => net199413, Q =>
                           n136, QN => net246084);
   REGISTERS_reg_1_24_inst : DFF_X1 port map( D => n1282, CK => net199413, Q =>
                           n135, QN => net246083);
   REGISTERS_reg_1_23_inst : DFF_X1 port map( D => n1304, CK => net199413, Q =>
                           n134, QN => net246082);
   REGISTERS_reg_1_22_inst : DFF_X1 port map( D => n1326, CK => net199413, Q =>
                           n133, QN => net246081);
   REGISTERS_reg_1_21_inst : DFF_X1 port map( D => n1348, CK => net199413, Q =>
                           n131, QN => net246080);
   REGISTERS_reg_1_20_inst : DFF_X1 port map( D => n1370, CK => net199413, Q =>
                           n130, QN => net246079);
   REGISTERS_reg_1_19_inst : DFF_X1 port map( D => n1392, CK => net199413, Q =>
                           n129, QN => net246078);
   REGISTERS_reg_1_18_inst : DFF_X1 port map( D => n1414, CK => net199413, Q =>
                           n128, QN => net246077);
   REGISTERS_reg_1_17_inst : DFF_X1 port map( D => n1436, CK => net199413, Q =>
                           n127, QN => net246076);
   REGISTERS_reg_1_16_inst : DFF_X1 port map( D => n1458, CK => net199413, Q =>
                           n126, QN => net246075);
   REGISTERS_reg_1_15_inst : DFF_X1 port map( D => n1480, CK => net199413, Q =>
                           n125, QN => net246074);
   REGISTERS_reg_1_14_inst : DFF_X1 port map( D => n1502, CK => net199413, Q =>
                           n124, QN => net246073);
   REGISTERS_reg_1_13_inst : DFF_X1 port map( D => n1524, CK => net199413, Q =>
                           n123, QN => net246072);
   REGISTERS_reg_1_12_inst : DFF_X1 port map( D => n1546, CK => net199413, Q =>
                           n122, QN => net246071);
   REGISTERS_reg_1_11_inst : DFF_X1 port map( D => n1568, CK => net199413, Q =>
                           n120, QN => net246070);
   REGISTERS_reg_1_10_inst : DFF_X1 port map( D => n1590, CK => net199413, Q =>
                           n119, QN => net246069);
   REGISTERS_reg_1_9_inst : DFF_X1 port map( D => n1612, CK => net199413, Q => 
                           n118, QN => net246068);
   REGISTERS_reg_1_8_inst : DFF_X1 port map( D => n1634, CK => net199413, Q => 
                           n117, QN => net246067);
   REGISTERS_reg_1_7_inst : DFF_X1 port map( D => n1656, CK => net199413, Q => 
                           n116, QN => net246066);
   REGISTERS_reg_1_6_inst : DFF_X1 port map( D => n1678, CK => net199413, Q => 
                           n115, QN => net246065);
   REGISTERS_reg_1_5_inst : DFF_X1 port map( D => n1700, CK => net199413, Q => 
                           n114, QN => net246064);
   REGISTERS_reg_1_4_inst : DFF_X1 port map( D => n1722, CK => net199413, Q => 
                           n113, QN => net246063);
   REGISTERS_reg_1_3_inst : DFF_X1 port map( D => n1744, CK => net199413, Q => 
                           n112, QN => net246062);
   REGISTERS_reg_1_2_inst : DFF_X1 port map( D => n1766, CK => net199413, Q => 
                           n111, QN => net246061);
   REGISTERS_reg_1_1_inst : DFF_X1 port map( D => n1788, CK => net199413, Q => 
                           n109, QN => net246060);
   REGISTERS_reg_1_0_inst : DFF_X1 port map( D => n1810, CK => net199413, Q => 
                           n108, QN => net246059);
   REGISTERS_reg_2_31_inst : DFF_X1 port map( D => n1094, CK => net199418, Q =>
                           n107, QN => net246058);
   REGISTERS_reg_2_30_inst : DFF_X1 port map( D => n1150, CK => net199418, Q =>
                           n106, QN => net246057);
   REGISTERS_reg_2_29_inst : DFF_X1 port map( D => n1172, CK => net199418, Q =>
                           n105, QN => net246056);
   REGISTERS_reg_2_28_inst : DFF_X1 port map( D => n1194, CK => net199418, Q =>
                           n104, QN => net246055);
   REGISTERS_reg_2_27_inst : DFF_X1 port map( D => n1216, CK => net199418, Q =>
                           n103, QN => net246054);
   REGISTERS_reg_2_26_inst : DFF_X1 port map( D => n1238, CK => net199418, Q =>
                           n102, QN => net246053);
   REGISTERS_reg_2_25_inst : DFF_X1 port map( D => n1260, CK => net199418, Q =>
                           n101, QN => net246052);
   REGISTERS_reg_2_24_inst : DFF_X1 port map( D => n1282, CK => net199418, Q =>
                           n100, QN => net246051);
   REGISTERS_reg_2_23_inst : DFF_X1 port map( D => n1304, CK => net199418, Q =>
                           n97, QN => net246050);
   REGISTERS_reg_2_22_inst : DFF_X1 port map( D => n1326, CK => net199418, Q =>
                           n95, QN => net246049);
   REGISTERS_reg_2_21_inst : DFF_X1 port map( D => n1348, CK => net199418, Q =>
                           n93, QN => net246048);
   REGISTERS_reg_2_20_inst : DFF_X1 port map( D => n1370, CK => net199418, Q =>
                           n91, QN => net246047);
   REGISTERS_reg_2_19_inst : DFF_X1 port map( D => n1392, CK => net199418, Q =>
                           n89, QN => net246046);
   REGISTERS_reg_2_18_inst : DFF_X1 port map( D => n1414, CK => net199418, Q =>
                           n87, QN => net246045);
   REGISTERS_reg_2_17_inst : DFF_X1 port map( D => n1436, CK => net199418, Q =>
                           n85, QN => net246044);
   REGISTERS_reg_2_16_inst : DFF_X1 port map( D => n1458, CK => net199418, Q =>
                           n83, QN => net246043);
   REGISTERS_reg_2_15_inst : DFF_X1 port map( D => n1480, CK => net199418, Q =>
                           n81, QN => net246042);
   REGISTERS_reg_2_14_inst : DFF_X1 port map( D => n1502, CK => net199418, Q =>
                           n79, QN => net246041);
   REGISTERS_reg_2_13_inst : DFF_X1 port map( D => n1524, CK => net199418, Q =>
                           n75, QN => net246040);
   REGISTERS_reg_2_12_inst : DFF_X1 port map( D => n1546, CK => net199418, Q =>
                           n73, QN => net246039);
   REGISTERS_reg_2_11_inst : DFF_X1 port map( D => n1568, CK => net199418, Q =>
                           n71, QN => net246038);
   REGISTERS_reg_2_10_inst : DFF_X1 port map( D => n1590, CK => net199418, Q =>
                           n69, QN => net246037);
   REGISTERS_reg_2_9_inst : DFF_X1 port map( D => n1612, CK => net199418, Q => 
                           n67, QN => net246036);
   REGISTERS_reg_2_8_inst : DFF_X1 port map( D => n1634, CK => net199418, Q => 
                           n65, QN => net246035);
   REGISTERS_reg_2_7_inst : DFF_X1 port map( D => n1656, CK => net199418, Q => 
                           n63, QN => net246034);
   REGISTERS_reg_2_6_inst : DFF_X1 port map( D => n1678, CK => net199418, Q => 
                           n61, QN => net246033);
   REGISTERS_reg_2_5_inst : DFF_X1 port map( D => n1700, CK => net199418, Q => 
                           n59, QN => net246032);
   REGISTERS_reg_2_4_inst : DFF_X1 port map( D => n1722, CK => net199418, Q => 
                           n57, QN => net246031);
   REGISTERS_reg_2_3_inst : DFF_X1 port map( D => n1744, CK => net199418, Q => 
                           n1101, QN => net246030);
   REGISTERS_reg_2_2_inst : DFF_X1 port map( D => n1766, CK => net199418, Q => 
                           n1100, QN => net246029);
   REGISTERS_reg_2_1_inst : DFF_X1 port map( D => n1788, CK => net199418, Q => 
                           n1099, QN => net246028);
   REGISTERS_reg_2_0_inst : DFF_X1 port map( D => n1810, CK => net199418, Q => 
                           n1098, QN => net246027);
   REGISTERS_reg_3_31_inst : DFF_X1 port map( D => n1094, CK => net199423, Q =>
                           n1097, QN => net246026);
   REGISTERS_reg_3_30_inst : DFF_X1 port map( D => n1150, CK => net199423, Q =>
                           n1096, QN => net246025);
   REGISTERS_reg_3_29_inst : DFF_X1 port map( D => n1172, CK => net199423, Q =>
                           n1095, QN => net246024);
   REGISTERS_reg_3_28_inst : DFF_X1 port map( D => n1194, CK => net199423, Q =>
                           n1093, QN => net246023);
   REGISTERS_reg_3_27_inst : DFF_X1 port map( D => n1216, CK => net199423, Q =>
                           n1092, QN => net246022);
   REGISTERS_reg_3_26_inst : DFF_X1 port map( D => n1238, CK => net199423, Q =>
                           n1091, QN => net246021);
   REGISTERS_reg_3_25_inst : DFF_X1 port map( D => n1260, CK => net199423, Q =>
                           n1089, QN => net246020);
   REGISTERS_reg_3_24_inst : DFF_X1 port map( D => n1282, CK => net199423, Q =>
                           n1088, QN => net246019);
   REGISTERS_reg_3_23_inst : DFF_X1 port map( D => n1304, CK => net199423, Q =>
                           n1087, QN => net246018);
   REGISTERS_reg_3_22_inst : DFF_X1 port map( D => n1326, CK => net199423, Q =>
                           n1086, QN => net246017);
   REGISTERS_reg_3_21_inst : DFF_X1 port map( D => n1348, CK => net199423, Q =>
                           n1085, QN => net246016);
   REGISTERS_reg_3_20_inst : DFF_X1 port map( D => n1370, CK => net199423, Q =>
                           n1084, QN => net246015);
   REGISTERS_reg_3_19_inst : DFF_X1 port map( D => n1392, CK => net199423, Q =>
                           n1083, QN => net246014);
   REGISTERS_reg_3_18_inst : DFF_X1 port map( D => n1414, CK => net199423, Q =>
                           n1082, QN => net246013);
   REGISTERS_reg_3_17_inst : DFF_X1 port map( D => n1436, CK => net199423, Q =>
                           n1081, QN => net246012);
   REGISTERS_reg_3_16_inst : DFF_X1 port map( D => n1458, CK => net199423, Q =>
                           n1080, QN => net246011);
   REGISTERS_reg_3_15_inst : DFF_X1 port map( D => n1480, CK => net199423, Q =>
                           n1079, QN => net246010);
   REGISTERS_reg_3_14_inst : DFF_X1 port map( D => n1502, CK => net199423, Q =>
                           n1078, QN => net246009);
   REGISTERS_reg_3_13_inst : DFF_X1 port map( D => n1524, CK => net199423, Q =>
                           n1077, QN => net246008);
   REGISTERS_reg_3_12_inst : DFF_X1 port map( D => n1546, CK => net199423, Q =>
                           n1076, QN => net246007);
   REGISTERS_reg_3_11_inst : DFF_X1 port map( D => n1568, CK => net199423, Q =>
                           n1075, QN => net246006);
   REGISTERS_reg_3_10_inst : DFF_X1 port map( D => n1590, CK => net199423, Q =>
                           n1074, QN => net246005);
   REGISTERS_reg_3_9_inst : DFF_X1 port map( D => n1612, CK => net199423, Q => 
                           n1073, QN => net246004);
   REGISTERS_reg_3_8_inst : DFF_X1 port map( D => n1634, CK => net199423, Q => 
                           n1072, QN => net246003);
   REGISTERS_reg_3_7_inst : DFF_X1 port map( D => n1656, CK => net199423, Q => 
                           n1071, QN => net246002);
   REGISTERS_reg_3_6_inst : DFF_X1 port map( D => n1678, CK => net199423, Q => 
                           n1070, QN => net246001);
   REGISTERS_reg_3_5_inst : DFF_X1 port map( D => n1700, CK => net199423, Q => 
                           n1068, QN => net246000);
   REGISTERS_reg_3_4_inst : DFF_X1 port map( D => n1722, CK => net199423, Q => 
                           n1067, QN => net245999);
   REGISTERS_reg_3_3_inst : DFF_X1 port map( D => n1744, CK => net199423, Q => 
                           n1066, QN => net245998);
   REGISTERS_reg_3_2_inst : DFF_X1 port map( D => n1766, CK => net199423, Q => 
                           n1065, QN => net245997);
   REGISTERS_reg_3_1_inst : DFF_X1 port map( D => n1788, CK => net199423, Q => 
                           n1064, QN => net245996);
   REGISTERS_reg_3_0_inst : DFF_X1 port map( D => n1810, CK => net199423, Q => 
                           n1063, QN => net245995);
   REGISTERS_reg_4_31_inst : DFF_X1 port map( D => n1094, CK => net199428, Q =>
                           n1062, QN => net245994);
   REGISTERS_reg_4_30_inst : DFF_X1 port map( D => n1150, CK => net199428, Q =>
                           n1061, QN => net245993);
   REGISTERS_reg_4_29_inst : DFF_X1 port map( D => n1172, CK => net199428, Q =>
                           n1060, QN => net245992);
   REGISTERS_reg_4_28_inst : DFF_X1 port map( D => n1194, CK => net199428, Q =>
                           n1059, QN => net245991);
   REGISTERS_reg_4_27_inst : DFF_X1 port map( D => n1216, CK => net199428, Q =>
                           n1058, QN => net245990);
   REGISTERS_reg_4_26_inst : DFF_X1 port map( D => n1238, CK => net199428, Q =>
                           n1057, QN => net245989);
   REGISTERS_reg_4_25_inst : DFF_X1 port map( D => n1260, CK => net199428, Q =>
                           n1056, QN => net245988);
   REGISTERS_reg_4_24_inst : DFF_X1 port map( D => n1282, CK => net199428, Q =>
                           n1055, QN => net245987);
   REGISTERS_reg_4_23_inst : DFF_X1 port map( D => n1304, CK => net199428, Q =>
                           n1054, QN => net245986);
   REGISTERS_reg_4_22_inst : DFF_X1 port map( D => n1326, CK => net199428, Q =>
                           n1053, QN => net245985);
   REGISTERS_reg_4_21_inst : DFF_X1 port map( D => n1348, CK => net199428, Q =>
                           n1052, QN => net245984);
   REGISTERS_reg_4_20_inst : DFF_X1 port map( D => n1370, CK => net199428, Q =>
                           n1051, QN => net245983);
   REGISTERS_reg_4_19_inst : DFF_X1 port map( D => n1392, CK => net199428, Q =>
                           n1050, QN => net245982);
   REGISTERS_reg_4_18_inst : DFF_X1 port map( D => n1414, CK => net199428, Q =>
                           n1049, QN => net245981);
   REGISTERS_reg_4_17_inst : DFF_X1 port map( D => n1436, CK => net199428, Q =>
                           n1047, QN => net245980);
   REGISTERS_reg_4_16_inst : DFF_X1 port map( D => n1458, CK => net199428, Q =>
                           n1046, QN => net245979);
   REGISTERS_reg_4_15_inst : DFF_X1 port map( D => n1480, CK => net199428, Q =>
                           n1045, QN => net245978);
   REGISTERS_reg_4_14_inst : DFF_X1 port map( D => n1502, CK => net199428, Q =>
                           n1044, QN => net245977);
   REGISTERS_reg_4_13_inst : DFF_X1 port map( D => n1524, CK => net199428, Q =>
                           n1043, QN => net245976);
   REGISTERS_reg_4_12_inst : DFF_X1 port map( D => n1546, CK => net199428, Q =>
                           n1042, QN => net245975);
   REGISTERS_reg_4_11_inst : DFF_X1 port map( D => n1568, CK => net199428, Q =>
                           n1041, QN => net245974);
   REGISTERS_reg_4_10_inst : DFF_X1 port map( D => n1590, CK => net199428, Q =>
                           n1040, QN => net245973);
   REGISTERS_reg_4_9_inst : DFF_X1 port map( D => n1612, CK => net199428, Q => 
                           n1039, QN => net245972);
   REGISTERS_reg_4_8_inst : DFF_X1 port map( D => n1634, CK => net199428, Q => 
                           n1038, QN => net245971);
   REGISTERS_reg_4_7_inst : DFF_X1 port map( D => n1656, CK => net199428, Q => 
                           n1037, QN => net245970);
   REGISTERS_reg_4_6_inst : DFF_X1 port map( D => n1678, CK => net199428, Q => 
                           n1036, QN => net245969);
   REGISTERS_reg_4_5_inst : DFF_X1 port map( D => n1700, CK => net199428, Q => 
                           n1035, QN => net245968);
   REGISTERS_reg_4_4_inst : DFF_X1 port map( D => n1722, CK => net199428, Q => 
                           n1034, QN => net245967);
   REGISTERS_reg_4_3_inst : DFF_X1 port map( D => n1744, CK => net199428, Q => 
                           n1033, QN => net245966);
   REGISTERS_reg_4_2_inst : DFF_X1 port map( D => n1766, CK => net199428, Q => 
                           n1032, QN => net245965);
   REGISTERS_reg_4_1_inst : DFF_X1 port map( D => n1788, CK => net199428, Q => 
                           n1031, QN => net245964);
   REGISTERS_reg_4_0_inst : DFF_X1 port map( D => n1810, CK => net199428, Q => 
                           n1030, QN => net245963);
   REGISTERS_reg_5_31_inst : DFF_X1 port map( D => n1094, CK => net199433, Q =>
                           n1029, QN => net245962);
   REGISTERS_reg_5_30_inst : DFF_X1 port map( D => n1150, CK => net199433, Q =>
                           n1028, QN => net245961);
   REGISTERS_reg_5_29_inst : DFF_X1 port map( D => n1172, CK => net199433, Q =>
                           n1026, QN => net245960);
   REGISTERS_reg_5_28_inst : DFF_X1 port map( D => n1194, CK => net199433, Q =>
                           n1025, QN => net245959);
   REGISTERS_reg_5_27_inst : DFF_X1 port map( D => n1216, CK => net199433, Q =>
                           n1024, QN => net245958);
   REGISTERS_reg_5_26_inst : DFF_X1 port map( D => n1238, CK => net199433, Q =>
                           n1023, QN => net245957);
   REGISTERS_reg_5_25_inst : DFF_X1 port map( D => n1260, CK => net199433, Q =>
                           n1022, QN => net245956);
   REGISTERS_reg_5_24_inst : DFF_X1 port map( D => n1282, CK => net199433, Q =>
                           n1021, QN => net245955);
   REGISTERS_reg_5_23_inst : DFF_X1 port map( D => n1304, CK => net199433, Q =>
                           n1020, QN => net245954);
   REGISTERS_reg_5_22_inst : DFF_X1 port map( D => n1326, CK => net199433, Q =>
                           n1019, QN => net245953);
   REGISTERS_reg_5_21_inst : DFF_X1 port map( D => n1348, CK => net199433, Q =>
                           n1018, QN => net245952);
   REGISTERS_reg_5_20_inst : DFF_X1 port map( D => n1370, CK => net199433, Q =>
                           n1017, QN => net245951);
   REGISTERS_reg_5_19_inst : DFF_X1 port map( D => n1392, CK => net199433, Q =>
                           n1016, QN => net245950);
   REGISTERS_reg_5_18_inst : DFF_X1 port map( D => n1414, CK => net199433, Q =>
                           n1015, QN => net245949);
   REGISTERS_reg_5_17_inst : DFF_X1 port map( D => n1436, CK => net199433, Q =>
                           n1014, QN => net245948);
   REGISTERS_reg_5_16_inst : DFF_X1 port map( D => n1458, CK => net199433, Q =>
                           n1013, QN => net245947);
   REGISTERS_reg_5_15_inst : DFF_X1 port map( D => n1480, CK => net199433, Q =>
                           n1012, QN => net245946);
   REGISTERS_reg_5_14_inst : DFF_X1 port map( D => n1502, CK => net199433, Q =>
                           n1011, QN => net245945);
   REGISTERS_reg_5_13_inst : DFF_X1 port map( D => n1524, CK => net199433, Q =>
                           n1010, QN => net245944);
   REGISTERS_reg_5_12_inst : DFF_X1 port map( D => n1546, CK => net199433, Q =>
                           n1009, QN => net245943);
   REGISTERS_reg_5_11_inst : DFF_X1 port map( D => n1568, CK => net199433, Q =>
                           n1008, QN => net245942);
   REGISTERS_reg_5_10_inst : DFF_X1 port map( D => n1590, CK => net199433, Q =>
                           n1007, QN => net245941);
   REGISTERS_reg_5_9_inst : DFF_X1 port map( D => n1612, CK => net199433, Q => 
                           n1005, QN => net245940);
   REGISTERS_reg_5_8_inst : DFF_X1 port map( D => n1634, CK => net199433, Q => 
                           n1004, QN => net245939);
   REGISTERS_reg_5_7_inst : DFF_X1 port map( D => n1656, CK => net199433, Q => 
                           n1003, QN => net245938);
   REGISTERS_reg_5_6_inst : DFF_X1 port map( D => n1678, CK => net199433, Q => 
                           n1002, QN => net245937);
   REGISTERS_reg_5_5_inst : DFF_X1 port map( D => n1700, CK => net199433, Q => 
                           n1001, QN => net245936);
   REGISTERS_reg_5_4_inst : DFF_X1 port map( D => n1722, CK => net199433, Q => 
                           n1000, QN => net245935);
   REGISTERS_reg_5_3_inst : DFF_X1 port map( D => n1744, CK => net199433, Q => 
                           n999, QN => net245934);
   REGISTERS_reg_5_2_inst : DFF_X1 port map( D => n1766, CK => net199433, Q => 
                           n998, QN => net245933);
   REGISTERS_reg_5_1_inst : DFF_X1 port map( D => n1788, CK => net199433, Q => 
                           n997, QN => net245932);
   REGISTERS_reg_5_0_inst : DFF_X1 port map( D => n1810, CK => net199433, Q => 
                           n996, QN => net245931);
   REGISTERS_reg_6_31_inst : DFF_X1 port map( D => n1094, CK => net199438, Q =>
                           n995, QN => net245930);
   REGISTERS_reg_6_30_inst : DFF_X1 port map( D => n1150, CK => net199438, Q =>
                           n994, QN => net245929);
   REGISTERS_reg_6_29_inst : DFF_X1 port map( D => n1172, CK => net199438, Q =>
                           n993, QN => net245928);
   REGISTERS_reg_6_28_inst : DFF_X1 port map( D => n1194, CK => net199438, Q =>
                           n992, QN => net245927);
   REGISTERS_reg_6_27_inst : DFF_X1 port map( D => n1216, CK => net199438, Q =>
                           n991, QN => net245926);
   REGISTERS_reg_6_26_inst : DFF_X1 port map( D => n1238, CK => net199438, Q =>
                           n990, QN => net245925);
   REGISTERS_reg_6_25_inst : DFF_X1 port map( D => n1260, CK => net199438, Q =>
                           n989, QN => net245924);
   REGISTERS_reg_6_24_inst : DFF_X1 port map( D => n1282, CK => net199438, Q =>
                           n988, QN => net245923);
   REGISTERS_reg_6_23_inst : DFF_X1 port map( D => n1304, CK => net199438, Q =>
                           n987, QN => net245922);
   REGISTERS_reg_6_22_inst : DFF_X1 port map( D => n1326, CK => net199438, Q =>
                           n986, QN => net245921);
   REGISTERS_reg_6_21_inst : DFF_X1 port map( D => n1348, CK => net199438, Q =>
                           n984, QN => net245920);
   REGISTERS_reg_6_20_inst : DFF_X1 port map( D => n1370, CK => net199438, Q =>
                           n983, QN => net245919);
   REGISTERS_reg_6_19_inst : DFF_X1 port map( D => n1392, CK => net199438, Q =>
                           n982, QN => net245918);
   REGISTERS_reg_6_18_inst : DFF_X1 port map( D => n1414, CK => net199438, Q =>
                           n981, QN => net245917);
   REGISTERS_reg_6_17_inst : DFF_X1 port map( D => n1436, CK => net199438, Q =>
                           n980, QN => net245916);
   REGISTERS_reg_6_16_inst : DFF_X1 port map( D => n1458, CK => net199438, Q =>
                           n979, QN => net245915);
   REGISTERS_reg_6_15_inst : DFF_X1 port map( D => n1480, CK => net199438, Q =>
                           n978, QN => net245914);
   REGISTERS_reg_6_14_inst : DFF_X1 port map( D => n1502, CK => net199438, Q =>
                           n977, QN => net245913);
   REGISTERS_reg_6_13_inst : DFF_X1 port map( D => n1524, CK => net199438, Q =>
                           n976, QN => net245912);
   REGISTERS_reg_6_12_inst : DFF_X1 port map( D => n1546, CK => net199438, Q =>
                           n975, QN => net245911);
   REGISTERS_reg_6_11_inst : DFF_X1 port map( D => n1568, CK => net199438, Q =>
                           n974, QN => net245910);
   REGISTERS_reg_6_10_inst : DFF_X1 port map( D => n1590, CK => net199438, Q =>
                           n973, QN => net245909);
   REGISTERS_reg_6_9_inst : DFF_X1 port map( D => n1612, CK => net199438, Q => 
                           n972, QN => net245908);
   REGISTERS_reg_6_8_inst : DFF_X1 port map( D => n1634, CK => net199438, Q => 
                           n971, QN => net245907);
   REGISTERS_reg_6_7_inst : DFF_X1 port map( D => n1656, CK => net199438, Q => 
                           n970, QN => net245906);
   REGISTERS_reg_6_6_inst : DFF_X1 port map( D => n1678, CK => net199438, Q => 
                           n969, QN => net245905);
   REGISTERS_reg_6_5_inst : DFF_X1 port map( D => n1700, CK => net199438, Q => 
                           n968, QN => net245904);
   REGISTERS_reg_6_4_inst : DFF_X1 port map( D => n1722, CK => net199438, Q => 
                           n967, QN => net245903);
   REGISTERS_reg_6_3_inst : DFF_X1 port map( D => n1744, CK => net199438, Q => 
                           n966, QN => net245902);
   REGISTERS_reg_6_2_inst : DFF_X1 port map( D => n1766, CK => net199438, Q => 
                           n965, QN => net245901);
   REGISTERS_reg_6_1_inst : DFF_X1 port map( D => n1788, CK => net199438, Q => 
                           n963, QN => net245900);
   REGISTERS_reg_6_0_inst : DFF_X1 port map( D => n1810, CK => net199438, Q => 
                           n962, QN => net245899);
   REGISTERS_reg_7_31_inst : DFF_X1 port map( D => n1094, CK => net199443, Q =>
                           n961, QN => net245898);
   REGISTERS_reg_7_30_inst : DFF_X1 port map( D => n1150, CK => net199443, Q =>
                           n960, QN => net245897);
   REGISTERS_reg_7_29_inst : DFF_X1 port map( D => n1172, CK => net199443, Q =>
                           n959, QN => net245896);
   REGISTERS_reg_7_28_inst : DFF_X1 port map( D => n1194, CK => net199443, Q =>
                           n958, QN => net245895);
   REGISTERS_reg_7_27_inst : DFF_X1 port map( D => n1216, CK => net199443, Q =>
                           n957, QN => net245894);
   REGISTERS_reg_7_26_inst : DFF_X1 port map( D => n1238, CK => net199443, Q =>
                           n956, QN => net245893);
   REGISTERS_reg_7_25_inst : DFF_X1 port map( D => n1260, CK => net199443, Q =>
                           n955, QN => net245892);
   REGISTERS_reg_7_24_inst : DFF_X1 port map( D => n1282, CK => net199443, Q =>
                           n954, QN => net245891);
   REGISTERS_reg_7_23_inst : DFF_X1 port map( D => n1304, CK => net199443, Q =>
                           n953, QN => net245890);
   REGISTERS_reg_7_22_inst : DFF_X1 port map( D => n1326, CK => net199443, Q =>
                           n952, QN => net245889);
   REGISTERS_reg_7_21_inst : DFF_X1 port map( D => n1348, CK => net199443, Q =>
                           n951, QN => net245888);
   REGISTERS_reg_7_20_inst : DFF_X1 port map( D => n1370, CK => net199443, Q =>
                           n950, QN => net245887);
   REGISTERS_reg_7_19_inst : DFF_X1 port map( D => n1392, CK => net199443, Q =>
                           n949, QN => net245886);
   REGISTERS_reg_7_18_inst : DFF_X1 port map( D => n1414, CK => net199443, Q =>
                           n948, QN => net245885);
   REGISTERS_reg_7_17_inst : DFF_X1 port map( D => n1436, CK => net199443, Q =>
                           n947, QN => net245884);
   REGISTERS_reg_7_16_inst : DFF_X1 port map( D => n1458, CK => net199443, Q =>
                           n946, QN => net245883);
   REGISTERS_reg_7_15_inst : DFF_X1 port map( D => n1480, CK => net199443, Q =>
                           n945, QN => net245882);
   REGISTERS_reg_7_14_inst : DFF_X1 port map( D => n1502, CK => net199443, Q =>
                           n944, QN => net245881);
   REGISTERS_reg_7_13_inst : DFF_X1 port map( D => n1524, CK => net199443, Q =>
                           n942, QN => net245880);
   REGISTERS_reg_7_12_inst : DFF_X1 port map( D => n1546, CK => net199443, Q =>
                           n941, QN => net245879);
   REGISTERS_reg_7_11_inst : DFF_X1 port map( D => n1568, CK => net199443, Q =>
                           n940, QN => net245878);
   REGISTERS_reg_7_10_inst : DFF_X1 port map( D => n1590, CK => net199443, Q =>
                           n939, QN => net245877);
   REGISTERS_reg_7_9_inst : DFF_X1 port map( D => n1612, CK => net199443, Q => 
                           n938, QN => net245876);
   REGISTERS_reg_7_8_inst : DFF_X1 port map( D => n1634, CK => net199443, Q => 
                           n937, QN => net245875);
   REGISTERS_reg_7_7_inst : DFF_X1 port map( D => n1656, CK => net199443, Q => 
                           n936, QN => net245874);
   REGISTERS_reg_7_6_inst : DFF_X1 port map( D => n1678, CK => net199443, Q => 
                           n935, QN => net245873);
   REGISTERS_reg_7_5_inst : DFF_X1 port map( D => n1700, CK => net199443, Q => 
                           n934, QN => net245872);
   REGISTERS_reg_7_4_inst : DFF_X1 port map( D => n1722, CK => net199443, Q => 
                           n933, QN => net245871);
   REGISTERS_reg_7_3_inst : DFF_X1 port map( D => n1744, CK => net199443, Q => 
                           n932, QN => net245870);
   REGISTERS_reg_7_2_inst : DFF_X1 port map( D => n1766, CK => net199443, Q => 
                           n931, QN => net245869);
   REGISTERS_reg_7_1_inst : DFF_X1 port map( D => n1788, CK => net199443, Q => 
                           n930, QN => net245868);
   REGISTERS_reg_7_0_inst : DFF_X1 port map( D => n1810, CK => net199443, Q => 
                           n929, QN => net245867);
   REGISTERS_reg_8_31_inst : DFF_X1 port map( D => n1094, CK => net199448, Q =>
                           n928, QN => net245866);
   REGISTERS_reg_8_30_inst : DFF_X1 port map( D => n1150, CK => net199448, Q =>
                           n927, QN => net245865);
   REGISTERS_reg_8_29_inst : DFF_X1 port map( D => n1172, CK => net199448, Q =>
                           n926, QN => net245864);
   REGISTERS_reg_8_28_inst : DFF_X1 port map( D => n1194, CK => net199448, Q =>
                           n925, QN => net245863);
   REGISTERS_reg_8_27_inst : DFF_X1 port map( D => n1216, CK => net199448, Q =>
                           n924, QN => net245862);
   REGISTERS_reg_8_26_inst : DFF_X1 port map( D => n1238, CK => net199448, Q =>
                           n923, QN => net245861);
   REGISTERS_reg_8_25_inst : DFF_X1 port map( D => n1260, CK => net199448, Q =>
                           n921, QN => net245860);
   REGISTERS_reg_8_24_inst : DFF_X1 port map( D => n1282, CK => net199448, Q =>
                           n920, QN => net245859);
   REGISTERS_reg_8_23_inst : DFF_X1 port map( D => n1304, CK => net199448, Q =>
                           n919, QN => net245858);
   REGISTERS_reg_8_22_inst : DFF_X1 port map( D => n1326, CK => net199448, Q =>
                           n918, QN => net245857);
   REGISTERS_reg_8_21_inst : DFF_X1 port map( D => n1348, CK => net199448, Q =>
                           n917, QN => net245856);
   REGISTERS_reg_8_20_inst : DFF_X1 port map( D => n1370, CK => net199448, Q =>
                           n916, QN => net245855);
   REGISTERS_reg_8_19_inst : DFF_X1 port map( D => n1392, CK => net199448, Q =>
                           n915, QN => net245854);
   REGISTERS_reg_8_18_inst : DFF_X1 port map( D => n1414, CK => net199448, Q =>
                           n914, QN => net245853);
   REGISTERS_reg_8_17_inst : DFF_X1 port map( D => n1436, CK => net199448, Q =>
                           n913, QN => net245852);
   REGISTERS_reg_8_16_inst : DFF_X1 port map( D => n1458, CK => net199448, Q =>
                           n912, QN => net245851);
   REGISTERS_reg_8_15_inst : DFF_X1 port map( D => n1480, CK => net199448, Q =>
                           n911, QN => net245850);
   REGISTERS_reg_8_14_inst : DFF_X1 port map( D => n1502, CK => net199448, Q =>
                           n910, QN => net245849);
   REGISTERS_reg_8_13_inst : DFF_X1 port map( D => n1524, CK => net199448, Q =>
                           n909, QN => net245848);
   REGISTERS_reg_8_12_inst : DFF_X1 port map( D => n1546, CK => net199448, Q =>
                           n908, QN => net245847);
   REGISTERS_reg_8_11_inst : DFF_X1 port map( D => n1568, CK => net199448, Q =>
                           n907, QN => net245846);
   REGISTERS_reg_8_10_inst : DFF_X1 port map( D => n1590, CK => net199448, Q =>
                           n906, QN => net245845);
   REGISTERS_reg_8_9_inst : DFF_X1 port map( D => n1612, CK => net199448, Q => 
                           n905, QN => net245844);
   REGISTERS_reg_8_8_inst : DFF_X1 port map( D => n1634, CK => net199448, Q => 
                           n904, QN => net245843);
   REGISTERS_reg_8_7_inst : DFF_X1 port map( D => n1656, CK => net199448, Q => 
                           n903, QN => net245842);
   REGISTERS_reg_8_6_inst : DFF_X1 port map( D => n1678, CK => net199448, Q => 
                           n902, QN => net245841);
   REGISTERS_reg_8_5_inst : DFF_X1 port map( D => n1700, CK => net199448, Q => 
                           n900, QN => net245840);
   REGISTERS_reg_8_4_inst : DFF_X1 port map( D => n1722, CK => net199448, Q => 
                           n899, QN => net245839);
   REGISTERS_reg_8_3_inst : DFF_X1 port map( D => n1744, CK => net199448, Q => 
                           n898, QN => net245838);
   REGISTERS_reg_8_2_inst : DFF_X1 port map( D => n1766, CK => net199448, Q => 
                           n897, QN => net245837);
   REGISTERS_reg_8_1_inst : DFF_X1 port map( D => n1788, CK => net199448, Q => 
                           n896, QN => net245836);
   REGISTERS_reg_8_0_inst : DFF_X1 port map( D => n1810, CK => net199448, Q => 
                           n895, QN => net245835);
   REGISTERS_reg_9_31_inst : DFF_X1 port map( D => n1094, CK => net199453, Q =>
                           n894, QN => net245834);
   REGISTERS_reg_9_30_inst : DFF_X1 port map( D => n1150, CK => net199453, Q =>
                           n893, QN => net245833);
   REGISTERS_reg_9_29_inst : DFF_X1 port map( D => n1172, CK => net199453, Q =>
                           n892, QN => net245832);
   REGISTERS_reg_9_28_inst : DFF_X1 port map( D => n1194, CK => net199453, Q =>
                           n891, QN => net245831);
   REGISTERS_reg_9_27_inst : DFF_X1 port map( D => n1216, CK => net199453, Q =>
                           n890, QN => net245830);
   REGISTERS_reg_9_26_inst : DFF_X1 port map( D => n1238, CK => net199453, Q =>
                           n889, QN => net245829);
   REGISTERS_reg_9_25_inst : DFF_X1 port map( D => n1260, CK => net199453, Q =>
                           n888, QN => net245828);
   REGISTERS_reg_9_24_inst : DFF_X1 port map( D => n1282, CK => net199453, Q =>
                           n887, QN => net245827);
   REGISTERS_reg_9_23_inst : DFF_X1 port map( D => n1304, CK => net199453, Q =>
                           n886, QN => net245826);
   REGISTERS_reg_9_22_inst : DFF_X1 port map( D => n1326, CK => net199453, Q =>
                           n885, QN => net245825);
   REGISTERS_reg_9_21_inst : DFF_X1 port map( D => n1348, CK => net199453, Q =>
                           n884, QN => net245824);
   REGISTERS_reg_9_20_inst : DFF_X1 port map( D => n1370, CK => net199453, Q =>
                           n883, QN => net245823);
   REGISTERS_reg_9_19_inst : DFF_X1 port map( D => n1392, CK => net199453, Q =>
                           n882, QN => net245822);
   REGISTERS_reg_9_18_inst : DFF_X1 port map( D => n1414, CK => net199453, Q =>
                           n881, QN => net245821);
   REGISTERS_reg_9_17_inst : DFF_X1 port map( D => n1436, CK => net199453, Q =>
                           n879, QN => net245820);
   REGISTERS_reg_9_16_inst : DFF_X1 port map( D => n1458, CK => net199453, Q =>
                           n878, QN => net245819);
   REGISTERS_reg_9_15_inst : DFF_X1 port map( D => n1480, CK => net199453, Q =>
                           n877, QN => net245818);
   REGISTERS_reg_9_14_inst : DFF_X1 port map( D => n1502, CK => net199453, Q =>
                           n876, QN => net245817);
   REGISTERS_reg_9_13_inst : DFF_X1 port map( D => n1524, CK => net199453, Q =>
                           n875, QN => net245816);
   REGISTERS_reg_9_12_inst : DFF_X1 port map( D => n1546, CK => net199453, Q =>
                           n874, QN => net245815);
   REGISTERS_reg_9_11_inst : DFF_X1 port map( D => n1568, CK => net199453, Q =>
                           n873, QN => net245814);
   REGISTERS_reg_9_10_inst : DFF_X1 port map( D => n1590, CK => net199453, Q =>
                           n872, QN => net245813);
   REGISTERS_reg_9_9_inst : DFF_X1 port map( D => n1612, CK => net199453, Q => 
                           n871, QN => net245812);
   REGISTERS_reg_9_8_inst : DFF_X1 port map( D => n1634, CK => net199453, Q => 
                           n870, QN => net245811);
   REGISTERS_reg_9_7_inst : DFF_X1 port map( D => n1656, CK => net199453, Q => 
                           n869, QN => net245810);
   REGISTERS_reg_9_6_inst : DFF_X1 port map( D => n1678, CK => net199453, Q => 
                           n868, QN => net245809);
   REGISTERS_reg_9_5_inst : DFF_X1 port map( D => n1700, CK => net199453, Q => 
                           n867, QN => net245808);
   REGISTERS_reg_9_4_inst : DFF_X1 port map( D => n1722, CK => net199453, Q => 
                           n866, QN => net245807);
   REGISTERS_reg_9_3_inst : DFF_X1 port map( D => n1744, CK => net199453, Q => 
                           n865, QN => net245806);
   REGISTERS_reg_9_2_inst : DFF_X1 port map( D => n1766, CK => net199453, Q => 
                           n864, QN => net245805);
   REGISTERS_reg_9_1_inst : DFF_X1 port map( D => n1788, CK => net199453, Q => 
                           n863, QN => net245804);
   REGISTERS_reg_9_0_inst : DFF_X1 port map( D => n1810, CK => net199453, Q => 
                           n862, QN => net245803);
   REGISTERS_reg_10_31_inst : DFF_X1 port map( D => n1094, CK => net199458, Q 
                           => n861, QN => net245802);
   REGISTERS_reg_10_30_inst : DFF_X1 port map( D => n1150, CK => net199458, Q 
                           => n860, QN => net245801);
   REGISTERS_reg_10_29_inst : DFF_X1 port map( D => n1172, CK => net199458, Q 
                           => n858, QN => net245800);
   REGISTERS_reg_10_28_inst : DFF_X1 port map( D => n1194, CK => net199458, Q 
                           => n857, QN => net245799);
   REGISTERS_reg_10_27_inst : DFF_X1 port map( D => n1216, CK => net199458, Q 
                           => n856, QN => net245798);
   REGISTERS_reg_10_26_inst : DFF_X1 port map( D => n1238, CK => net199458, Q 
                           => n855, QN => net245797);
   REGISTERS_reg_10_25_inst : DFF_X1 port map( D => n1260, CK => net199458, Q 
                           => n854, QN => net245796);
   REGISTERS_reg_10_24_inst : DFF_X1 port map( D => n1282, CK => net199458, Q 
                           => n853, QN => net245795);
   REGISTERS_reg_10_23_inst : DFF_X1 port map( D => n1304, CK => net199458, Q 
                           => n852, QN => net245794);
   REGISTERS_reg_10_22_inst : DFF_X1 port map( D => n1326, CK => net199458, Q 
                           => n851, QN => net245793);
   REGISTERS_reg_10_21_inst : DFF_X1 port map( D => n1348, CK => net199458, Q 
                           => n850, QN => net245792);
   REGISTERS_reg_10_20_inst : DFF_X1 port map( D => n1370, CK => net199458, Q 
                           => n849, QN => net245791);
   REGISTERS_reg_10_19_inst : DFF_X1 port map( D => n1392, CK => net199458, Q 
                           => n848, QN => net245790);
   REGISTERS_reg_10_18_inst : DFF_X1 port map( D => n1414, CK => net199458, Q 
                           => n847, QN => net245789);
   REGISTERS_reg_10_17_inst : DFF_X1 port map( D => n1436, CK => net199458, Q 
                           => n846, QN => net245788);
   REGISTERS_reg_10_16_inst : DFF_X1 port map( D => n1458, CK => net199458, Q 
                           => n845, QN => net245787);
   REGISTERS_reg_10_15_inst : DFF_X1 port map( D => n1480, CK => net199458, Q 
                           => n844, QN => net245786);
   REGISTERS_reg_10_14_inst : DFF_X1 port map( D => n1502, CK => net199458, Q 
                           => n843, QN => net245785);
   REGISTERS_reg_10_13_inst : DFF_X1 port map( D => n1524, CK => net199458, Q 
                           => n842, QN => net245784);
   REGISTERS_reg_10_12_inst : DFF_X1 port map( D => n1546, CK => net199458, Q 
                           => n841, QN => net245783);
   REGISTERS_reg_10_11_inst : DFF_X1 port map( D => n1568, CK => net199458, Q 
                           => n840, QN => net245782);
   REGISTERS_reg_10_10_inst : DFF_X1 port map( D => n1590, CK => net199458, Q 
                           => n839, QN => net245781);
   REGISTERS_reg_10_9_inst : DFF_X1 port map( D => n1612, CK => net199458, Q =>
                           n837, QN => net245780);
   REGISTERS_reg_10_8_inst : DFF_X1 port map( D => n1634, CK => net199458, Q =>
                           n836, QN => net245779);
   REGISTERS_reg_10_7_inst : DFF_X1 port map( D => n1656, CK => net199458, Q =>
                           n835, QN => net245778);
   REGISTERS_reg_10_6_inst : DFF_X1 port map( D => n1678, CK => net199458, Q =>
                           n834, QN => net245777);
   REGISTERS_reg_10_5_inst : DFF_X1 port map( D => n1700, CK => net199458, Q =>
                           n833, QN => net245776);
   REGISTERS_reg_10_4_inst : DFF_X1 port map( D => n1722, CK => net199458, Q =>
                           n832, QN => net245775);
   REGISTERS_reg_10_3_inst : DFF_X1 port map( D => n1744, CK => net199458, Q =>
                           n831, QN => net245774);
   REGISTERS_reg_10_2_inst : DFF_X1 port map( D => n1766, CK => net199458, Q =>
                           n830, QN => net245773);
   REGISTERS_reg_10_1_inst : DFF_X1 port map( D => n1788, CK => net199458, Q =>
                           n829, QN => net245772);
   REGISTERS_reg_10_0_inst : DFF_X1 port map( D => n1810, CK => net199458, Q =>
                           n828, QN => net245771);
   REGISTERS_reg_11_31_inst : DFF_X1 port map( D => n1094, CK => net199463, Q 
                           => n827, QN => net245770);
   REGISTERS_reg_11_30_inst : DFF_X1 port map( D => n1150, CK => net199463, Q 
                           => n826, QN => net245769);
   REGISTERS_reg_11_29_inst : DFF_X1 port map( D => n1172, CK => net199463, Q 
                           => n825, QN => net245768);
   REGISTERS_reg_11_28_inst : DFF_X1 port map( D => n1194, CK => net199463, Q 
                           => n824, QN => net245767);
   REGISTERS_reg_11_27_inst : DFF_X1 port map( D => n1216, CK => net199463, Q 
                           => n823, QN => net245766);
   REGISTERS_reg_11_26_inst : DFF_X1 port map( D => n1238, CK => net199463, Q 
                           => n822, QN => net245765);
   REGISTERS_reg_11_25_inst : DFF_X1 port map( D => n1260, CK => net199463, Q 
                           => n821, QN => net245764);
   REGISTERS_reg_11_24_inst : DFF_X1 port map( D => n1282, CK => net199463, Q 
                           => n820, QN => net245763);
   REGISTERS_reg_11_23_inst : DFF_X1 port map( D => n1304, CK => net199463, Q 
                           => n819, QN => net245762);
   REGISTERS_reg_11_22_inst : DFF_X1 port map( D => n1326, CK => net199463, Q 
                           => n818, QN => net245761);
   REGISTERS_reg_11_21_inst : DFF_X1 port map( D => n1348, CK => net199463, Q 
                           => n816, QN => net245760);
   REGISTERS_reg_11_20_inst : DFF_X1 port map( D => n1370, CK => net199463, Q 
                           => n815, QN => net245759);
   REGISTERS_reg_11_19_inst : DFF_X1 port map( D => n1392, CK => net199463, Q 
                           => n814, QN => net245758);
   REGISTERS_reg_11_18_inst : DFF_X1 port map( D => n1414, CK => net199463, Q 
                           => n813, QN => net245757);
   REGISTERS_reg_11_17_inst : DFF_X1 port map( D => n1436, CK => net199463, Q 
                           => n812, QN => net245756);
   REGISTERS_reg_11_16_inst : DFF_X1 port map( D => n1458, CK => net199463, Q 
                           => n811, QN => net245755);
   REGISTERS_reg_11_15_inst : DFF_X1 port map( D => n1480, CK => net199463, Q 
                           => n810, QN => net245754);
   REGISTERS_reg_11_14_inst : DFF_X1 port map( D => n1502, CK => net199463, Q 
                           => n809, QN => net245753);
   REGISTERS_reg_11_13_inst : DFF_X1 port map( D => n1524, CK => net199463, Q 
                           => n808, QN => net245752);
   REGISTERS_reg_11_12_inst : DFF_X1 port map( D => n1546, CK => net199463, Q 
                           => n807, QN => net245751);
   REGISTERS_reg_11_11_inst : DFF_X1 port map( D => n1568, CK => net199463, Q 
                           => n806, QN => net245750);
   REGISTERS_reg_11_10_inst : DFF_X1 port map( D => n1590, CK => net199463, Q 
                           => n805, QN => net245749);
   REGISTERS_reg_11_9_inst : DFF_X1 port map( D => n1612, CK => net199463, Q =>
                           n804, QN => net245748);
   REGISTERS_reg_11_8_inst : DFF_X1 port map( D => n1634, CK => net199463, Q =>
                           n803, QN => net245747);
   REGISTERS_reg_11_7_inst : DFF_X1 port map( D => n1656, CK => net199463, Q =>
                           n802, QN => net245746);
   REGISTERS_reg_11_6_inst : DFF_X1 port map( D => n1678, CK => net199463, Q =>
                           n801, QN => net245745);
   REGISTERS_reg_11_5_inst : DFF_X1 port map( D => n1700, CK => net199463, Q =>
                           n800, QN => net245744);
   REGISTERS_reg_11_4_inst : DFF_X1 port map( D => n1722, CK => net199463, Q =>
                           n799, QN => net245743);
   REGISTERS_reg_11_3_inst : DFF_X1 port map( D => n1744, CK => net199463, Q =>
                           n798, QN => net245742);
   REGISTERS_reg_11_2_inst : DFF_X1 port map( D => n1766, CK => net199463, Q =>
                           n797, QN => net245741);
   REGISTERS_reg_11_1_inst : DFF_X1 port map( D => n1788, CK => net199463, Q =>
                           n795, QN => net245740);
   REGISTERS_reg_11_0_inst : DFF_X1 port map( D => n1810, CK => net199463, Q =>
                           n794, QN => net245739);
   REGISTERS_reg_12_31_inst : DFF_X1 port map( D => n1094, CK => net199468, Q 
                           => n793, QN => net245738);
   REGISTERS_reg_12_30_inst : DFF_X1 port map( D => n1150, CK => net199468, Q 
                           => n792, QN => net245737);
   REGISTERS_reg_12_29_inst : DFF_X1 port map( D => n1172, CK => net199468, Q 
                           => n791, QN => net245736);
   REGISTERS_reg_12_28_inst : DFF_X1 port map( D => n1194, CK => net199468, Q 
                           => n790, QN => net245735);
   REGISTERS_reg_12_27_inst : DFF_X1 port map( D => n1216, CK => net199468, Q 
                           => n789, QN => net245734);
   REGISTERS_reg_12_26_inst : DFF_X1 port map( D => n1238, CK => net199468, Q 
                           => n788, QN => net245733);
   REGISTERS_reg_12_25_inst : DFF_X1 port map( D => n1260, CK => net199468, Q 
                           => n787, QN => net245732);
   REGISTERS_reg_12_24_inst : DFF_X1 port map( D => n1282, CK => net199468, Q 
                           => n786, QN => net245731);
   REGISTERS_reg_12_23_inst : DFF_X1 port map( D => n1304, CK => net199468, Q 
                           => n785, QN => net245730);
   REGISTERS_reg_12_22_inst : DFF_X1 port map( D => n1326, CK => net199468, Q 
                           => n784, QN => net245729);
   REGISTERS_reg_12_21_inst : DFF_X1 port map( D => n1348, CK => net199468, Q 
                           => n783, QN => net245728);
   REGISTERS_reg_12_20_inst : DFF_X1 port map( D => n1370, CK => net199468, Q 
                           => n782, QN => net245727);
   REGISTERS_reg_12_19_inst : DFF_X1 port map( D => n1392, CK => net199468, Q 
                           => n781, QN => net245726);
   REGISTERS_reg_12_18_inst : DFF_X1 port map( D => n1414, CK => net199468, Q 
                           => n780, QN => net245725);
   REGISTERS_reg_12_17_inst : DFF_X1 port map( D => n1436, CK => net199468, Q 
                           => n779, QN => net245724);
   REGISTERS_reg_12_16_inst : DFF_X1 port map( D => n1458, CK => net199468, Q 
                           => n778, QN => net245723);
   REGISTERS_reg_12_15_inst : DFF_X1 port map( D => n1480, CK => net199468, Q 
                           => n777, QN => net245722);
   REGISTERS_reg_12_14_inst : DFF_X1 port map( D => n1502, CK => net199468, Q 
                           => n776, QN => net245721);
   REGISTERS_reg_12_13_inst : DFF_X1 port map( D => n1524, CK => net199468, Q 
                           => n774, QN => net245720);
   REGISTERS_reg_12_12_inst : DFF_X1 port map( D => n1546, CK => net199468, Q 
                           => n773, QN => net245719);
   REGISTERS_reg_12_11_inst : DFF_X1 port map( D => n1568, CK => net199468, Q 
                           => n772, QN => net245718);
   REGISTERS_reg_12_10_inst : DFF_X1 port map( D => n1590, CK => net199468, Q 
                           => n771, QN => net245717);
   REGISTERS_reg_12_9_inst : DFF_X1 port map( D => n1612, CK => net199468, Q =>
                           n770, QN => net245716);
   REGISTERS_reg_12_8_inst : DFF_X1 port map( D => n1634, CK => net199468, Q =>
                           n769, QN => net245715);
   REGISTERS_reg_12_7_inst : DFF_X1 port map( D => n1656, CK => net199468, Q =>
                           n768, QN => net245714);
   REGISTERS_reg_12_6_inst : DFF_X1 port map( D => n1678, CK => net199468, Q =>
                           n767, QN => net245713);
   REGISTERS_reg_12_5_inst : DFF_X1 port map( D => n1700, CK => net199468, Q =>
                           n766, QN => net245712);
   REGISTERS_reg_12_4_inst : DFF_X1 port map( D => n1722, CK => net199468, Q =>
                           n765, QN => net245711);
   REGISTERS_reg_12_3_inst : DFF_X1 port map( D => n1744, CK => net199468, Q =>
                           n764, QN => net245710);
   REGISTERS_reg_12_2_inst : DFF_X1 port map( D => n1766, CK => net199468, Q =>
                           n763, QN => net245709);
   REGISTERS_reg_12_1_inst : DFF_X1 port map( D => n1788, CK => net199468, Q =>
                           n762, QN => net245708);
   REGISTERS_reg_12_0_inst : DFF_X1 port map( D => n1810, CK => net199468, Q =>
                           n761, QN => net245707);
   REGISTERS_reg_13_31_inst : DFF_X1 port map( D => n1094, CK => net199473, Q 
                           => n760, QN => net245706);
   REGISTERS_reg_13_30_inst : DFF_X1 port map( D => n1150, CK => net199473, Q 
                           => n759, QN => net245705);
   REGISTERS_reg_13_29_inst : DFF_X1 port map( D => n1172, CK => net199473, Q 
                           => n758, QN => net245704);
   REGISTERS_reg_13_28_inst : DFF_X1 port map( D => n1194, CK => net199473, Q 
                           => n757, QN => net245703);
   REGISTERS_reg_13_27_inst : DFF_X1 port map( D => n1216, CK => net199473, Q 
                           => n756, QN => net245702);
   REGISTERS_reg_13_26_inst : DFF_X1 port map( D => n1238, CK => net199473, Q 
                           => n755, QN => net245701);
   REGISTERS_reg_13_25_inst : DFF_X1 port map( D => n1260, CK => net199473, Q 
                           => n753, QN => net245700);
   REGISTERS_reg_13_24_inst : DFF_X1 port map( D => n1282, CK => net199473, Q 
                           => n752, QN => net245699);
   REGISTERS_reg_13_23_inst : DFF_X1 port map( D => n1304, CK => net199473, Q 
                           => n751, QN => net245698);
   REGISTERS_reg_13_22_inst : DFF_X1 port map( D => n1326, CK => net199473, Q 
                           => n750, QN => net245697);
   REGISTERS_reg_13_21_inst : DFF_X1 port map( D => n1348, CK => net199473, Q 
                           => n749, QN => net245696);
   REGISTERS_reg_13_20_inst : DFF_X1 port map( D => n1370, CK => net199473, Q 
                           => n748, QN => net245695);
   REGISTERS_reg_13_19_inst : DFF_X1 port map( D => n1392, CK => net199473, Q 
                           => n747, QN => net245694);
   REGISTERS_reg_13_18_inst : DFF_X1 port map( D => n1414, CK => net199473, Q 
                           => n746, QN => net245693);
   REGISTERS_reg_13_17_inst : DFF_X1 port map( D => n1436, CK => net199473, Q 
                           => n745, QN => net245692);
   REGISTERS_reg_13_16_inst : DFF_X1 port map( D => n1458, CK => net199473, Q 
                           => n744, QN => net245691);
   REGISTERS_reg_13_15_inst : DFF_X1 port map( D => n1480, CK => net199473, Q 
                           => n743, QN => net245690);
   REGISTERS_reg_13_14_inst : DFF_X1 port map( D => n1502, CK => net199473, Q 
                           => n742, QN => net245689);
   REGISTERS_reg_13_13_inst : DFF_X1 port map( D => n1524, CK => net199473, Q 
                           => n741, QN => net245688);
   REGISTERS_reg_13_12_inst : DFF_X1 port map( D => n1546, CK => net199473, Q 
                           => n740, QN => net245687);
   REGISTERS_reg_13_11_inst : DFF_X1 port map( D => n1568, CK => net199473, Q 
                           => n739, QN => net245686);
   REGISTERS_reg_13_10_inst : DFF_X1 port map( D => n1590, CK => net199473, Q 
                           => n738, QN => net245685);
   REGISTERS_reg_13_9_inst : DFF_X1 port map( D => n1612, CK => net199473, Q =>
                           n737, QN => net245684);
   REGISTERS_reg_13_8_inst : DFF_X1 port map( D => n1634, CK => net199473, Q =>
                           n736, QN => net245683);
   REGISTERS_reg_13_7_inst : DFF_X1 port map( D => n1656, CK => net199473, Q =>
                           n735, QN => net245682);
   REGISTERS_reg_13_6_inst : DFF_X1 port map( D => n1678, CK => net199473, Q =>
                           n734, QN => net245681);
   REGISTERS_reg_13_5_inst : DFF_X1 port map( D => n1700, CK => net199473, Q =>
                           n732, QN => net245680);
   REGISTERS_reg_13_4_inst : DFF_X1 port map( D => n1722, CK => net199473, Q =>
                           n731, QN => net245679);
   REGISTERS_reg_13_3_inst : DFF_X1 port map( D => n1744, CK => net199473, Q =>
                           n730, QN => net245678);
   REGISTERS_reg_13_2_inst : DFF_X1 port map( D => n1766, CK => net199473, Q =>
                           n729, QN => net245677);
   REGISTERS_reg_13_1_inst : DFF_X1 port map( D => n1788, CK => net199473, Q =>
                           n728, QN => net245676);
   REGISTERS_reg_13_0_inst : DFF_X1 port map( D => n1810, CK => net199473, Q =>
                           n727, QN => net245675);
   REGISTERS_reg_14_31_inst : DFF_X1 port map( D => n1094, CK => net199478, Q 
                           => n726, QN => net245674);
   REGISTERS_reg_14_30_inst : DFF_X1 port map( D => n1150, CK => net199478, Q 
                           => n725, QN => net245673);
   REGISTERS_reg_14_29_inst : DFF_X1 port map( D => n1172, CK => net199478, Q 
                           => n724, QN => net245672);
   REGISTERS_reg_14_28_inst : DFF_X1 port map( D => n1194, CK => net199478, Q 
                           => n723, QN => net245671);
   REGISTERS_reg_14_27_inst : DFF_X1 port map( D => n1216, CK => net199478, Q 
                           => n722, QN => net245670);
   REGISTERS_reg_14_26_inst : DFF_X1 port map( D => n1238, CK => net199478, Q 
                           => n721, QN => net245669);
   REGISTERS_reg_14_25_inst : DFF_X1 port map( D => n1260, CK => net199478, Q 
                           => n720, QN => net245668);
   REGISTERS_reg_14_24_inst : DFF_X1 port map( D => n1282, CK => net199478, Q 
                           => n719, QN => net245667);
   REGISTERS_reg_14_23_inst : DFF_X1 port map( D => n1304, CK => net199478, Q 
                           => n718, QN => net245666);
   REGISTERS_reg_14_22_inst : DFF_X1 port map( D => n1326, CK => net199478, Q 
                           => n717, QN => net245665);
   REGISTERS_reg_14_21_inst : DFF_X1 port map( D => n1348, CK => net199478, Q 
                           => n716, QN => net245664);
   REGISTERS_reg_14_20_inst : DFF_X1 port map( D => n1370, CK => net199478, Q 
                           => n715, QN => net245663);
   REGISTERS_reg_14_19_inst : DFF_X1 port map( D => n1392, CK => net199478, Q 
                           => n714, QN => net245662);
   REGISTERS_reg_14_18_inst : DFF_X1 port map( D => n1414, CK => net199478, Q 
                           => n713, QN => net245661);
   REGISTERS_reg_14_17_inst : DFF_X1 port map( D => n1436, CK => net199478, Q 
                           => n711, QN => net245660);
   REGISTERS_reg_14_16_inst : DFF_X1 port map( D => n1458, CK => net199478, Q 
                           => n710, QN => net245659);
   REGISTERS_reg_14_15_inst : DFF_X1 port map( D => n1480, CK => net199478, Q 
                           => n709, QN => net245658);
   REGISTERS_reg_14_14_inst : DFF_X1 port map( D => n1502, CK => net199478, Q 
                           => n708, QN => net245657);
   REGISTERS_reg_14_13_inst : DFF_X1 port map( D => n1524, CK => net199478, Q 
                           => n707, QN => net245656);
   REGISTERS_reg_14_12_inst : DFF_X1 port map( D => n1546, CK => net199478, Q 
                           => n706, QN => net245655);
   REGISTERS_reg_14_11_inst : DFF_X1 port map( D => n1568, CK => net199478, Q 
                           => n705, QN => net245654);
   REGISTERS_reg_14_10_inst : DFF_X1 port map( D => n1590, CK => net199478, Q 
                           => n704, QN => net245653);
   REGISTERS_reg_14_9_inst : DFF_X1 port map( D => n1612, CK => net199478, Q =>
                           n703, QN => net245652);
   REGISTERS_reg_14_8_inst : DFF_X1 port map( D => n1634, CK => net199478, Q =>
                           n702, QN => net245651);
   REGISTERS_reg_14_7_inst : DFF_X1 port map( D => n1656, CK => net199478, Q =>
                           n701, QN => net245650);
   REGISTERS_reg_14_6_inst : DFF_X1 port map( D => n1678, CK => net199478, Q =>
                           n700, QN => net245649);
   REGISTERS_reg_14_5_inst : DFF_X1 port map( D => n1700, CK => net199478, Q =>
                           n699, QN => net245648);
   REGISTERS_reg_14_4_inst : DFF_X1 port map( D => n1722, CK => net199478, Q =>
                           n698, QN => net245647);
   REGISTERS_reg_14_3_inst : DFF_X1 port map( D => n1744, CK => net199478, Q =>
                           n697, QN => net245646);
   REGISTERS_reg_14_2_inst : DFF_X1 port map( D => n1766, CK => net199478, Q =>
                           n696, QN => net245645);
   REGISTERS_reg_14_1_inst : DFF_X1 port map( D => n1788, CK => net199478, Q =>
                           n695, QN => net245644);
   REGISTERS_reg_14_0_inst : DFF_X1 port map( D => n1810, CK => net199478, Q =>
                           n694, QN => net245643);
   REGISTERS_reg_15_31_inst : DFF_X1 port map( D => n1094, CK => net199483, Q 
                           => n693, QN => net245642);
   REGISTERS_reg_15_30_inst : DFF_X1 port map( D => n1150, CK => net199483, Q 
                           => n692, QN => net245641);
   REGISTERS_reg_15_29_inst : DFF_X1 port map( D => n1172, CK => net199483, Q 
                           => n690, QN => net245640);
   REGISTERS_reg_15_28_inst : DFF_X1 port map( D => n1194, CK => net199483, Q 
                           => n689, QN => net245639);
   REGISTERS_reg_15_27_inst : DFF_X1 port map( D => n1216, CK => net199483, Q 
                           => n688, QN => net245638);
   REGISTERS_reg_15_26_inst : DFF_X1 port map( D => n1238, CK => net199483, Q 
                           => n687, QN => net245637);
   REGISTERS_reg_15_25_inst : DFF_X1 port map( D => n1260, CK => net199483, Q 
                           => n686, QN => net245636);
   REGISTERS_reg_15_24_inst : DFF_X1 port map( D => n1282, CK => net199483, Q 
                           => n685, QN => net245635);
   REGISTERS_reg_15_23_inst : DFF_X1 port map( D => n1304, CK => net199483, Q 
                           => n684, QN => net245634);
   REGISTERS_reg_15_22_inst : DFF_X1 port map( D => n1326, CK => net199483, Q 
                           => n683, QN => net245633);
   REGISTERS_reg_15_21_inst : DFF_X1 port map( D => n1348, CK => net199483, Q 
                           => n682, QN => net245632);
   REGISTERS_reg_15_20_inst : DFF_X1 port map( D => n1370, CK => net199483, Q 
                           => n681, QN => net245631);
   REGISTERS_reg_15_19_inst : DFF_X1 port map( D => n1392, CK => net199483, Q 
                           => n680, QN => net245630);
   REGISTERS_reg_15_18_inst : DFF_X1 port map( D => n1414, CK => net199483, Q 
                           => n679, QN => net245629);
   REGISTERS_reg_15_17_inst : DFF_X1 port map( D => n1436, CK => net199483, Q 
                           => n678, QN => net245628);
   REGISTERS_reg_15_16_inst : DFF_X1 port map( D => n1458, CK => net199483, Q 
                           => n677, QN => net245627);
   REGISTERS_reg_15_15_inst : DFF_X1 port map( D => n1480, CK => net199483, Q 
                           => n676, QN => net245626);
   REGISTERS_reg_15_14_inst : DFF_X1 port map( D => n1502, CK => net199483, Q 
                           => n675, QN => net245625);
   REGISTERS_reg_15_13_inst : DFF_X1 port map( D => n1524, CK => net199483, Q 
                           => n674, QN => net245624);
   REGISTERS_reg_15_12_inst : DFF_X1 port map( D => n1546, CK => net199483, Q 
                           => n673, QN => net245623);
   REGISTERS_reg_15_11_inst : DFF_X1 port map( D => n1568, CK => net199483, Q 
                           => n672, QN => net245622);
   REGISTERS_reg_15_10_inst : DFF_X1 port map( D => n1590, CK => net199483, Q 
                           => n671, QN => net245621);
   REGISTERS_reg_15_9_inst : DFF_X1 port map( D => n1612, CK => net199483, Q =>
                           n669, QN => net245620);
   REGISTERS_reg_15_8_inst : DFF_X1 port map( D => n1634, CK => net199483, Q =>
                           n668, QN => net245619);
   REGISTERS_reg_15_7_inst : DFF_X1 port map( D => n1656, CK => net199483, Q =>
                           n667, QN => net245618);
   REGISTERS_reg_15_6_inst : DFF_X1 port map( D => n1678, CK => net199483, Q =>
                           n666, QN => net245617);
   REGISTERS_reg_15_5_inst : DFF_X1 port map( D => n1700, CK => net199483, Q =>
                           n665, QN => net245616);
   REGISTERS_reg_15_4_inst : DFF_X1 port map( D => n1722, CK => net199483, Q =>
                           n664, QN => net245615);
   REGISTERS_reg_15_3_inst : DFF_X1 port map( D => n1744, CK => net199483, Q =>
                           n663, QN => net245614);
   REGISTERS_reg_15_2_inst : DFF_X1 port map( D => n1766, CK => net199483, Q =>
                           n662, QN => net245613);
   REGISTERS_reg_15_1_inst : DFF_X1 port map( D => n1788, CK => net199483, Q =>
                           n661, QN => net245612);
   REGISTERS_reg_15_0_inst : DFF_X1 port map( D => n1810, CK => net199483, Q =>
                           n660, QN => net245611);
   REGISTERS_reg_16_31_inst : DFF_X1 port map( D => n1094, CK => net199488, Q 
                           => n659, QN => net245610);
   REGISTERS_reg_16_30_inst : DFF_X1 port map( D => n1150, CK => net199488, Q 
                           => n658, QN => net245609);
   REGISTERS_reg_16_29_inst : DFF_X1 port map( D => n1172, CK => net199488, Q 
                           => n657, QN => net245608);
   REGISTERS_reg_16_28_inst : DFF_X1 port map( D => n1194, CK => net199488, Q 
                           => n656, QN => net245607);
   REGISTERS_reg_16_27_inst : DFF_X1 port map( D => n1216, CK => net199488, Q 
                           => n655, QN => net245606);
   REGISTERS_reg_16_26_inst : DFF_X1 port map( D => n1238, CK => net199488, Q 
                           => n654, QN => net245605);
   REGISTERS_reg_16_25_inst : DFF_X1 port map( D => n1260, CK => net199488, Q 
                           => n653, QN => net245604);
   REGISTERS_reg_16_24_inst : DFF_X1 port map( D => n1282, CK => net199488, Q 
                           => n652, QN => net245603);
   REGISTERS_reg_16_23_inst : DFF_X1 port map( D => n1304, CK => net199488, Q 
                           => n651, QN => net245602);
   REGISTERS_reg_16_22_inst : DFF_X1 port map( D => n1326, CK => net199488, Q 
                           => n650, QN => net245601);
   REGISTERS_reg_16_21_inst : DFF_X1 port map( D => n1348, CK => net199488, Q 
                           => n648, QN => net245600);
   REGISTERS_reg_16_20_inst : DFF_X1 port map( D => n1370, CK => net199488, Q 
                           => n647, QN => net245599);
   REGISTERS_reg_16_19_inst : DFF_X1 port map( D => n1392, CK => net199488, Q 
                           => n646, QN => net245598);
   REGISTERS_reg_16_18_inst : DFF_X1 port map( D => n1414, CK => net199488, Q 
                           => n645, QN => net245597);
   REGISTERS_reg_16_17_inst : DFF_X1 port map( D => n1436, CK => net199488, Q 
                           => n644, QN => net245596);
   REGISTERS_reg_16_16_inst : DFF_X1 port map( D => n1458, CK => net199488, Q 
                           => n643, QN => net245595);
   REGISTERS_reg_16_15_inst : DFF_X1 port map( D => n1480, CK => net199488, Q 
                           => n642, QN => net245594);
   REGISTERS_reg_16_14_inst : DFF_X1 port map( D => n1502, CK => net199488, Q 
                           => n641, QN => net245593);
   REGISTERS_reg_16_13_inst : DFF_X1 port map( D => n1524, CK => net199488, Q 
                           => n640, QN => net245592);
   REGISTERS_reg_16_12_inst : DFF_X1 port map( D => n1546, CK => net199488, Q 
                           => n639, QN => net245591);
   REGISTERS_reg_16_11_inst : DFF_X1 port map( D => n1568, CK => net199488, Q 
                           => n638, QN => net245590);
   REGISTERS_reg_16_10_inst : DFF_X1 port map( D => n1590, CK => net199488, Q 
                           => n637, QN => net245589);
   REGISTERS_reg_16_9_inst : DFF_X1 port map( D => n1612, CK => net199488, Q =>
                           n636, QN => net245588);
   REGISTERS_reg_16_8_inst : DFF_X1 port map( D => n1634, CK => net199488, Q =>
                           n635, QN => net245587);
   REGISTERS_reg_16_7_inst : DFF_X1 port map( D => n1656, CK => net199488, Q =>
                           n634, QN => net245586);
   REGISTERS_reg_16_6_inst : DFF_X1 port map( D => n1678, CK => net199488, Q =>
                           n633, QN => net245585);
   REGISTERS_reg_16_5_inst : DFF_X1 port map( D => n1700, CK => net199488, Q =>
                           n632, QN => net245584);
   REGISTERS_reg_16_4_inst : DFF_X1 port map( D => n1722, CK => net199488, Q =>
                           n631, QN => net245583);
   REGISTERS_reg_16_3_inst : DFF_X1 port map( D => n1744, CK => net199488, Q =>
                           n630, QN => net245582);
   REGISTERS_reg_16_2_inst : DFF_X1 port map( D => n1766, CK => net199488, Q =>
                           n629, QN => net245581);
   REGISTERS_reg_16_1_inst : DFF_X1 port map( D => n1788, CK => net199488, Q =>
                           n627, QN => net245580);
   REGISTERS_reg_16_0_inst : DFF_X1 port map( D => n1810, CK => net199488, Q =>
                           n626, QN => net245579);
   REGISTERS_reg_17_31_inst : DFF_X1 port map( D => n1094, CK => net199493, Q 
                           => n625, QN => net245578);
   REGISTERS_reg_17_30_inst : DFF_X1 port map( D => n1150, CK => net199493, Q 
                           => n624, QN => net245577);
   REGISTERS_reg_17_29_inst : DFF_X1 port map( D => n1172, CK => net199493, Q 
                           => n623, QN => net245576);
   REGISTERS_reg_17_28_inst : DFF_X1 port map( D => n1194, CK => net199493, Q 
                           => n622, QN => net245575);
   REGISTERS_reg_17_27_inst : DFF_X1 port map( D => n1216, CK => net199493, Q 
                           => n621, QN => net245574);
   REGISTERS_reg_17_26_inst : DFF_X1 port map( D => n1238, CK => net199493, Q 
                           => n620, QN => net245573);
   REGISTERS_reg_17_25_inst : DFF_X1 port map( D => n1260, CK => net199493, Q 
                           => n619, QN => net245572);
   REGISTERS_reg_17_24_inst : DFF_X1 port map( D => n1282, CK => net199493, Q 
                           => n618, QN => net245571);
   REGISTERS_reg_17_23_inst : DFF_X1 port map( D => n1304, CK => net199493, Q 
                           => n617, QN => net245570);
   REGISTERS_reg_17_22_inst : DFF_X1 port map( D => n1326, CK => net199493, Q 
                           => n616, QN => net245569);
   REGISTERS_reg_17_21_inst : DFF_X1 port map( D => n1348, CK => net199493, Q 
                           => n615, QN => net245568);
   REGISTERS_reg_17_20_inst : DFF_X1 port map( D => n1370, CK => net199493, Q 
                           => n614, QN => net245567);
   REGISTERS_reg_17_19_inst : DFF_X1 port map( D => n1392, CK => net199493, Q 
                           => n613, QN => net245566);
   REGISTERS_reg_17_18_inst : DFF_X1 port map( D => n1414, CK => net199493, Q 
                           => n612, QN => net245565);
   REGISTERS_reg_17_17_inst : DFF_X1 port map( D => n1436, CK => net199493, Q 
                           => n611, QN => net245564);
   REGISTERS_reg_17_16_inst : DFF_X1 port map( D => n1458, CK => net199493, Q 
                           => n610, QN => net245563);
   REGISTERS_reg_17_15_inst : DFF_X1 port map( D => n1480, CK => net199493, Q 
                           => n609, QN => net245562);
   REGISTERS_reg_17_14_inst : DFF_X1 port map( D => n1502, CK => net199493, Q 
                           => n608, QN => net245561);
   REGISTERS_reg_17_13_inst : DFF_X1 port map( D => n1524, CK => net199493, Q 
                           => n606, QN => net245560);
   REGISTERS_reg_17_12_inst : DFF_X1 port map( D => n1546, CK => net199493, Q 
                           => n605, QN => net245559);
   REGISTERS_reg_17_11_inst : DFF_X1 port map( D => n1568, CK => net199493, Q 
                           => n604, QN => net245558);
   REGISTERS_reg_17_10_inst : DFF_X1 port map( D => n1590, CK => net199493, Q 
                           => n603, QN => net245557);
   REGISTERS_reg_17_9_inst : DFF_X1 port map( D => n1612, CK => net199493, Q =>
                           n602, QN => net245556);
   REGISTERS_reg_17_8_inst : DFF_X1 port map( D => n1634, CK => net199493, Q =>
                           n601, QN => net245555);
   REGISTERS_reg_17_7_inst : DFF_X1 port map( D => n1656, CK => net199493, Q =>
                           n600, QN => net245554);
   REGISTERS_reg_17_6_inst : DFF_X1 port map( D => n1678, CK => net199493, Q =>
                           n599, QN => net245553);
   REGISTERS_reg_17_5_inst : DFF_X1 port map( D => n1700, CK => net199493, Q =>
                           n598, QN => net245552);
   REGISTERS_reg_17_4_inst : DFF_X1 port map( D => n1722, CK => net199493, Q =>
                           n597, QN => net245551);
   REGISTERS_reg_17_3_inst : DFF_X1 port map( D => n1744, CK => net199493, Q =>
                           n596, QN => net245550);
   REGISTERS_reg_17_2_inst : DFF_X1 port map( D => n1766, CK => net199493, Q =>
                           n595, QN => net245549);
   REGISTERS_reg_17_1_inst : DFF_X1 port map( D => n1788, CK => net199493, Q =>
                           n594, QN => net245548);
   REGISTERS_reg_17_0_inst : DFF_X1 port map( D => n1810, CK => net199493, Q =>
                           n593, QN => net245547);
   REGISTERS_reg_18_31_inst : DFF_X1 port map( D => n1094, CK => net199498, Q 
                           => n592, QN => net245546);
   REGISTERS_reg_18_30_inst : DFF_X1 port map( D => n1150, CK => net199498, Q 
                           => n591, QN => net245545);
   REGISTERS_reg_18_29_inst : DFF_X1 port map( D => n1172, CK => net199498, Q 
                           => n590, QN => net245544);
   REGISTERS_reg_18_28_inst : DFF_X1 port map( D => n1194, CK => net199498, Q 
                           => n589, QN => net245543);
   REGISTERS_reg_18_27_inst : DFF_X1 port map( D => n1216, CK => net199498, Q 
                           => n588, QN => net245542);
   REGISTERS_reg_18_26_inst : DFF_X1 port map( D => n1238, CK => net199498, Q 
                           => n587, QN => net245541);
   REGISTERS_reg_18_25_inst : DFF_X1 port map( D => n1260, CK => net199498, Q 
                           => n585, QN => net245540);
   REGISTERS_reg_18_24_inst : DFF_X1 port map( D => n1282, CK => net199498, Q 
                           => n584, QN => net245539);
   REGISTERS_reg_18_23_inst : DFF_X1 port map( D => n1304, CK => net199498, Q 
                           => n583, QN => net245538);
   REGISTERS_reg_18_22_inst : DFF_X1 port map( D => n1326, CK => net199498, Q 
                           => n582, QN => net245537);
   REGISTERS_reg_18_21_inst : DFF_X1 port map( D => n1348, CK => net199498, Q 
                           => n581, QN => net245536);
   REGISTERS_reg_18_20_inst : DFF_X1 port map( D => n1370, CK => net199498, Q 
                           => n580, QN => net245535);
   REGISTERS_reg_18_19_inst : DFF_X1 port map( D => n1392, CK => net199498, Q 
                           => n579, QN => net245534);
   REGISTERS_reg_18_18_inst : DFF_X1 port map( D => n1414, CK => net199498, Q 
                           => n578, QN => net245533);
   REGISTERS_reg_18_17_inst : DFF_X1 port map( D => n1436, CK => net199498, Q 
                           => n577, QN => net245532);
   REGISTERS_reg_18_16_inst : DFF_X1 port map( D => n1458, CK => net199498, Q 
                           => n576, QN => net245531);
   REGISTERS_reg_18_15_inst : DFF_X1 port map( D => n1480, CK => net199498, Q 
                           => n575, QN => net245530);
   REGISTERS_reg_18_14_inst : DFF_X1 port map( D => n1502, CK => net199498, Q 
                           => n574, QN => net245529);
   REGISTERS_reg_18_13_inst : DFF_X1 port map( D => n1524, CK => net199498, Q 
                           => n573, QN => net245528);
   REGISTERS_reg_18_12_inst : DFF_X1 port map( D => n1546, CK => net199498, Q 
                           => n572, QN => net245527);
   REGISTERS_reg_18_11_inst : DFF_X1 port map( D => n1568, CK => net199498, Q 
                           => n571, QN => net245526);
   REGISTERS_reg_18_10_inst : DFF_X1 port map( D => n1590, CK => net199498, Q 
                           => n570, QN => net245525);
   REGISTERS_reg_18_9_inst : DFF_X1 port map( D => n1612, CK => net199498, Q =>
                           n569, QN => net245524);
   REGISTERS_reg_18_8_inst : DFF_X1 port map( D => n1634, CK => net199498, Q =>
                           n568, QN => net245523);
   REGISTERS_reg_18_7_inst : DFF_X1 port map( D => n1656, CK => net199498, Q =>
                           n567, QN => net245522);
   REGISTERS_reg_18_6_inst : DFF_X1 port map( D => n1678, CK => net199498, Q =>
                           n566, QN => net245521);
   REGISTERS_reg_18_5_inst : DFF_X1 port map( D => n1700, CK => net199498, Q =>
                           n564, QN => net245520);
   REGISTERS_reg_18_4_inst : DFF_X1 port map( D => n1722, CK => net199498, Q =>
                           n563, QN => net245519);
   REGISTERS_reg_18_3_inst : DFF_X1 port map( D => n1744, CK => net199498, Q =>
                           n562, QN => net245518);
   REGISTERS_reg_18_2_inst : DFF_X1 port map( D => n1766, CK => net199498, Q =>
                           n561, QN => net245517);
   REGISTERS_reg_18_1_inst : DFF_X1 port map( D => n1788, CK => net199498, Q =>
                           n560, QN => net245516);
   REGISTERS_reg_18_0_inst : DFF_X1 port map( D => n1810, CK => net199498, Q =>
                           n559, QN => net245515);
   REGISTERS_reg_19_31_inst : DFF_X1 port map( D => n1094, CK => net199503, Q 
                           => n558, QN => net245514);
   REGISTERS_reg_19_30_inst : DFF_X1 port map( D => n1150, CK => net199503, Q 
                           => n557, QN => net245513);
   REGISTERS_reg_19_29_inst : DFF_X1 port map( D => n1172, CK => net199503, Q 
                           => n556, QN => net245512);
   REGISTERS_reg_19_28_inst : DFF_X1 port map( D => n1194, CK => net199503, Q 
                           => n555, QN => net245511);
   REGISTERS_reg_19_27_inst : DFF_X1 port map( D => n1216, CK => net199503, Q 
                           => n554, QN => net245510);
   REGISTERS_reg_19_26_inst : DFF_X1 port map( D => n1238, CK => net199503, Q 
                           => n553, QN => net245509);
   REGISTERS_reg_19_25_inst : DFF_X1 port map( D => n1260, CK => net199503, Q 
                           => n552, QN => net245508);
   REGISTERS_reg_19_24_inst : DFF_X1 port map( D => n1282, CK => net199503, Q 
                           => n551, QN => net245507);
   REGISTERS_reg_19_23_inst : DFF_X1 port map( D => n1304, CK => net199503, Q 
                           => n550, QN => net245506);
   REGISTERS_reg_19_22_inst : DFF_X1 port map( D => n1326, CK => net199503, Q 
                           => n549, QN => net245505);
   REGISTERS_reg_19_21_inst : DFF_X1 port map( D => n1348, CK => net199503, Q 
                           => n548, QN => net245504);
   REGISTERS_reg_19_20_inst : DFF_X1 port map( D => n1370, CK => net199503, Q 
                           => n547, QN => net245503);
   REGISTERS_reg_19_19_inst : DFF_X1 port map( D => n1392, CK => net199503, Q 
                           => n546, QN => net245502);
   REGISTERS_reg_19_18_inst : DFF_X1 port map( D => n1414, CK => net199503, Q 
                           => n545, QN => net245501);
   REGISTERS_reg_19_17_inst : DFF_X1 port map( D => n1436, CK => net199503, Q 
                           => n543, QN => net245500);
   REGISTERS_reg_19_16_inst : DFF_X1 port map( D => n1458, CK => net199503, Q 
                           => n542, QN => net245499);
   REGISTERS_reg_19_15_inst : DFF_X1 port map( D => n1480, CK => net199503, Q 
                           => n541, QN => net245498);
   REGISTERS_reg_19_14_inst : DFF_X1 port map( D => n1502, CK => net199503, Q 
                           => n540, QN => net245497);
   REGISTERS_reg_19_13_inst : DFF_X1 port map( D => n1524, CK => net199503, Q 
                           => n539, QN => net245496);
   REGISTERS_reg_19_12_inst : DFF_X1 port map( D => n1546, CK => net199503, Q 
                           => n538, QN => net245495);
   REGISTERS_reg_19_11_inst : DFF_X1 port map( D => n1568, CK => net199503, Q 
                           => n537, QN => net245494);
   REGISTERS_reg_19_10_inst : DFF_X1 port map( D => n1590, CK => net199503, Q 
                           => n536, QN => net245493);
   REGISTERS_reg_19_9_inst : DFF_X1 port map( D => n1612, CK => net199503, Q =>
                           n535, QN => net245492);
   REGISTERS_reg_19_8_inst : DFF_X1 port map( D => n1634, CK => net199503, Q =>
                           n534, QN => net245491);
   REGISTERS_reg_19_7_inst : DFF_X1 port map( D => n1656, CK => net199503, Q =>
                           n533, QN => net245490);
   REGISTERS_reg_19_6_inst : DFF_X1 port map( D => n1678, CK => net199503, Q =>
                           n532, QN => net245489);
   REGISTERS_reg_19_5_inst : DFF_X1 port map( D => n1700, CK => net199503, Q =>
                           n531, QN => net245488);
   REGISTERS_reg_19_4_inst : DFF_X1 port map( D => n1722, CK => net199503, Q =>
                           n530, QN => net245487);
   REGISTERS_reg_19_3_inst : DFF_X1 port map( D => n1744, CK => net199503, Q =>
                           n529, QN => net245486);
   REGISTERS_reg_19_2_inst : DFF_X1 port map( D => n1766, CK => net199503, Q =>
                           n528, QN => net245485);
   REGISTERS_reg_19_1_inst : DFF_X1 port map( D => n1788, CK => net199503, Q =>
                           n527, QN => net245484);
   REGISTERS_reg_19_0_inst : DFF_X1 port map( D => n1810, CK => net199503, Q =>
                           n526, QN => net245483);
   REGISTERS_reg_20_31_inst : DFF_X1 port map( D => n1094, CK => net199508, Q 
                           => n525, QN => net245482);
   REGISTERS_reg_20_30_inst : DFF_X1 port map( D => n1150, CK => net199508, Q 
                           => n524, QN => net245481);
   REGISTERS_reg_20_29_inst : DFF_X1 port map( D => n1172, CK => net199508, Q 
                           => n522, QN => net245480);
   REGISTERS_reg_20_28_inst : DFF_X1 port map( D => n1194, CK => net199508, Q 
                           => n521, QN => net245479);
   REGISTERS_reg_20_27_inst : DFF_X1 port map( D => n1216, CK => net199508, Q 
                           => n520, QN => net245478);
   REGISTERS_reg_20_26_inst : DFF_X1 port map( D => n1238, CK => net199508, Q 
                           => n519, QN => net245477);
   REGISTERS_reg_20_25_inst : DFF_X1 port map( D => n1260, CK => net199508, Q 
                           => n518, QN => net245476);
   REGISTERS_reg_20_24_inst : DFF_X1 port map( D => n1282, CK => net199508, Q 
                           => n517, QN => net245475);
   REGISTERS_reg_20_23_inst : DFF_X1 port map( D => n1304, CK => net199508, Q 
                           => n516, QN => net245474);
   REGISTERS_reg_20_22_inst : DFF_X1 port map( D => n1326, CK => net199508, Q 
                           => n515, QN => net245473);
   REGISTERS_reg_20_21_inst : DFF_X1 port map( D => n1348, CK => net199508, Q 
                           => n514, QN => net245472);
   REGISTERS_reg_20_20_inst : DFF_X1 port map( D => n1370, CK => net199508, Q 
                           => n513, QN => net245471);
   REGISTERS_reg_20_19_inst : DFF_X1 port map( D => n1392, CK => net199508, Q 
                           => n512, QN => net245470);
   REGISTERS_reg_20_18_inst : DFF_X1 port map( D => n1414, CK => net199508, Q 
                           => n511, QN => net245469);
   REGISTERS_reg_20_17_inst : DFF_X1 port map( D => n1436, CK => net199508, Q 
                           => n510, QN => net245468);
   REGISTERS_reg_20_16_inst : DFF_X1 port map( D => n1458, CK => net199508, Q 
                           => n509, QN => net245467);
   REGISTERS_reg_20_15_inst : DFF_X1 port map( D => n1480, CK => net199508, Q 
                           => n508, QN => net245466);
   REGISTERS_reg_20_14_inst : DFF_X1 port map( D => n1502, CK => net199508, Q 
                           => n507, QN => net245465);
   REGISTERS_reg_20_13_inst : DFF_X1 port map( D => n1524, CK => net199508, Q 
                           => n506, QN => net245464);
   REGISTERS_reg_20_12_inst : DFF_X1 port map( D => n1546, CK => net199508, Q 
                           => n505, QN => net245463);
   REGISTERS_reg_20_11_inst : DFF_X1 port map( D => n1568, CK => net199508, Q 
                           => n504, QN => net245462);
   REGISTERS_reg_20_10_inst : DFF_X1 port map( D => n1590, CK => net199508, Q 
                           => n503, QN => net245461);
   REGISTERS_reg_20_9_inst : DFF_X1 port map( D => n1612, CK => net199508, Q =>
                           n501, QN => net245460);
   REGISTERS_reg_20_8_inst : DFF_X1 port map( D => n1634, CK => net199508, Q =>
                           n500, QN => net245459);
   REGISTERS_reg_20_7_inst : DFF_X1 port map( D => n1656, CK => net199508, Q =>
                           n499, QN => net245458);
   REGISTERS_reg_20_6_inst : DFF_X1 port map( D => n1678, CK => net199508, Q =>
                           n498, QN => net245457);
   REGISTERS_reg_20_5_inst : DFF_X1 port map( D => n1700, CK => net199508, Q =>
                           n497, QN => net245456);
   REGISTERS_reg_20_4_inst : DFF_X1 port map( D => n1722, CK => net199508, Q =>
                           n496, QN => net245455);
   REGISTERS_reg_20_3_inst : DFF_X1 port map( D => n1744, CK => net199508, Q =>
                           n495, QN => net245454);
   REGISTERS_reg_20_2_inst : DFF_X1 port map( D => n1766, CK => net199508, Q =>
                           n494, QN => net245453);
   REGISTERS_reg_20_1_inst : DFF_X1 port map( D => n1788, CK => net199508, Q =>
                           n493, QN => net245452);
   REGISTERS_reg_20_0_inst : DFF_X1 port map( D => n1810, CK => net199508, Q =>
                           n492, QN => net245451);
   REGISTERS_reg_21_31_inst : DFF_X1 port map( D => n1094, CK => net199513, Q 
                           => n491, QN => net245450);
   REGISTERS_reg_21_30_inst : DFF_X1 port map( D => n1150, CK => net199513, Q 
                           => n490, QN => net245449);
   REGISTERS_reg_21_29_inst : DFF_X1 port map( D => n1172, CK => net199513, Q 
                           => n489, QN => net245448);
   REGISTERS_reg_21_28_inst : DFF_X1 port map( D => n1194, CK => net199513, Q 
                           => n488, QN => net245447);
   REGISTERS_reg_21_27_inst : DFF_X1 port map( D => n1216, CK => net199513, Q 
                           => n487, QN => net245446);
   REGISTERS_reg_21_26_inst : DFF_X1 port map( D => n1238, CK => net199513, Q 
                           => n486, QN => net245445);
   REGISTERS_reg_21_25_inst : DFF_X1 port map( D => n1260, CK => net199513, Q 
                           => n485, QN => net245444);
   REGISTERS_reg_21_24_inst : DFF_X1 port map( D => n1282, CK => net199513, Q 
                           => n484, QN => net245443);
   REGISTERS_reg_21_23_inst : DFF_X1 port map( D => n1304, CK => net199513, Q 
                           => n483, QN => net245442);
   REGISTERS_reg_21_22_inst : DFF_X1 port map( D => n1326, CK => net199513, Q 
                           => n482, QN => net245441);
   REGISTERS_reg_21_21_inst : DFF_X1 port map( D => n1348, CK => net199513, Q 
                           => n480, QN => net245440);
   REGISTERS_reg_21_20_inst : DFF_X1 port map( D => n1370, CK => net199513, Q 
                           => n479, QN => net245439);
   REGISTERS_reg_21_19_inst : DFF_X1 port map( D => n1392, CK => net199513, Q 
                           => n478, QN => net245438);
   REGISTERS_reg_21_18_inst : DFF_X1 port map( D => n1414, CK => net199513, Q 
                           => n477, QN => net245437);
   REGISTERS_reg_21_17_inst : DFF_X1 port map( D => n1436, CK => net199513, Q 
                           => n476, QN => net245436);
   REGISTERS_reg_21_16_inst : DFF_X1 port map( D => n1458, CK => net199513, Q 
                           => n475, QN => net245435);
   REGISTERS_reg_21_15_inst : DFF_X1 port map( D => n1480, CK => net199513, Q 
                           => n474, QN => net245434);
   REGISTERS_reg_21_14_inst : DFF_X1 port map( D => n1502, CK => net199513, Q 
                           => n473, QN => net245433);
   REGISTERS_reg_21_13_inst : DFF_X1 port map( D => n1524, CK => net199513, Q 
                           => n472, QN => net245432);
   REGISTERS_reg_21_12_inst : DFF_X1 port map( D => n1546, CK => net199513, Q 
                           => n471, QN => net245431);
   REGISTERS_reg_21_11_inst : DFF_X1 port map( D => n1568, CK => net199513, Q 
                           => n470, QN => net245430);
   REGISTERS_reg_21_10_inst : DFF_X1 port map( D => n1590, CK => net199513, Q 
                           => n469, QN => net245429);
   REGISTERS_reg_21_9_inst : DFF_X1 port map( D => n1612, CK => net199513, Q =>
                           n468, QN => net245428);
   REGISTERS_reg_21_8_inst : DFF_X1 port map( D => n1634, CK => net199513, Q =>
                           n467, QN => net245427);
   REGISTERS_reg_21_7_inst : DFF_X1 port map( D => n1656, CK => net199513, Q =>
                           n466, QN => net245426);
   REGISTERS_reg_21_6_inst : DFF_X1 port map( D => n1678, CK => net199513, Q =>
                           n465, QN => net245425);
   REGISTERS_reg_21_5_inst : DFF_X1 port map( D => n1700, CK => net199513, Q =>
                           n464, QN => net245424);
   REGISTERS_reg_21_4_inst : DFF_X1 port map( D => n1722, CK => net199513, Q =>
                           n463, QN => net245423);
   REGISTERS_reg_21_3_inst : DFF_X1 port map( D => n1744, CK => net199513, Q =>
                           n462, QN => net245422);
   REGISTERS_reg_21_2_inst : DFF_X1 port map( D => n1766, CK => net199513, Q =>
                           n461, QN => net245421);
   REGISTERS_reg_21_1_inst : DFF_X1 port map( D => n1788, CK => net199513, Q =>
                           n459, QN => net245420);
   REGISTERS_reg_21_0_inst : DFF_X1 port map( D => n1810, CK => net199513, Q =>
                           n458, QN => net245419);
   REGISTERS_reg_22_31_inst : DFF_X1 port map( D => n1094, CK => net199518, Q 
                           => n457, QN => net245418);
   REGISTERS_reg_22_30_inst : DFF_X1 port map( D => n1150, CK => net199518, Q 
                           => n456, QN => net245417);
   REGISTERS_reg_22_29_inst : DFF_X1 port map( D => n1172, CK => net199518, Q 
                           => n455, QN => net245416);
   REGISTERS_reg_22_28_inst : DFF_X1 port map( D => n1194, CK => net199518, Q 
                           => n454, QN => net245415);
   REGISTERS_reg_22_27_inst : DFF_X1 port map( D => n1216, CK => net199518, Q 
                           => n453, QN => net245414);
   REGISTERS_reg_22_26_inst : DFF_X1 port map( D => n1238, CK => net199518, Q 
                           => n452, QN => net245413);
   REGISTERS_reg_22_25_inst : DFF_X1 port map( D => n1260, CK => net199518, Q 
                           => n451, QN => net245412);
   REGISTERS_reg_22_24_inst : DFF_X1 port map( D => n1282, CK => net199518, Q 
                           => n450, QN => net245411);
   REGISTERS_reg_22_23_inst : DFF_X1 port map( D => n1304, CK => net199518, Q 
                           => n449, QN => net245410);
   REGISTERS_reg_22_22_inst : DFF_X1 port map( D => n1326, CK => net199518, Q 
                           => n448, QN => net245409);
   REGISTERS_reg_22_21_inst : DFF_X1 port map( D => n1348, CK => net199518, Q 
                           => n447, QN => net245408);
   REGISTERS_reg_22_20_inst : DFF_X1 port map( D => n1370, CK => net199518, Q 
                           => n446, QN => net245407);
   REGISTERS_reg_22_19_inst : DFF_X1 port map( D => n1392, CK => net199518, Q 
                           => n445, QN => net245406);
   REGISTERS_reg_22_18_inst : DFF_X1 port map( D => n1414, CK => net199518, Q 
                           => n444, QN => net245405);
   REGISTERS_reg_22_17_inst : DFF_X1 port map( D => n1436, CK => net199518, Q 
                           => n443, QN => net245404);
   REGISTERS_reg_22_16_inst : DFF_X1 port map( D => n1458, CK => net199518, Q 
                           => n442, QN => net245403);
   REGISTERS_reg_22_15_inst : DFF_X1 port map( D => n1480, CK => net199518, Q 
                           => n441, QN => net245402);
   REGISTERS_reg_22_14_inst : DFF_X1 port map( D => n1502, CK => net199518, Q 
                           => n440, QN => net245401);
   REGISTERS_reg_22_13_inst : DFF_X1 port map( D => n1524, CK => net199518, Q 
                           => n438, QN => net245400);
   REGISTERS_reg_22_12_inst : DFF_X1 port map( D => n1546, CK => net199518, Q 
                           => n437, QN => net245399);
   REGISTERS_reg_22_11_inst : DFF_X1 port map( D => n1568, CK => net199518, Q 
                           => n436, QN => net245398);
   REGISTERS_reg_22_10_inst : DFF_X1 port map( D => n1590, CK => net199518, Q 
                           => n435, QN => net245397);
   REGISTERS_reg_22_9_inst : DFF_X1 port map( D => n1612, CK => net199518, Q =>
                           n434, QN => net245396);
   REGISTERS_reg_22_8_inst : DFF_X1 port map( D => n1634, CK => net199518, Q =>
                           n433, QN => net245395);
   REGISTERS_reg_22_7_inst : DFF_X1 port map( D => n1656, CK => net199518, Q =>
                           n432, QN => net245394);
   REGISTERS_reg_22_6_inst : DFF_X1 port map( D => n1678, CK => net199518, Q =>
                           n431, QN => net245393);
   REGISTERS_reg_22_5_inst : DFF_X1 port map( D => n1700, CK => net199518, Q =>
                           n430, QN => net245392);
   REGISTERS_reg_22_4_inst : DFF_X1 port map( D => n1722, CK => net199518, Q =>
                           n429, QN => net245391);
   REGISTERS_reg_22_3_inst : DFF_X1 port map( D => n1744, CK => net199518, Q =>
                           n428, QN => net245390);
   REGISTERS_reg_22_2_inst : DFF_X1 port map( D => n1766, CK => net199518, Q =>
                           n427, QN => net245389);
   REGISTERS_reg_22_1_inst : DFF_X1 port map( D => n1788, CK => net199518, Q =>
                           n426, QN => net245388);
   REGISTERS_reg_22_0_inst : DFF_X1 port map( D => n1810, CK => net199518, Q =>
                           n425, QN => net245387);
   REGISTERS_reg_23_31_inst : DFF_X1 port map( D => n1094, CK => net199523, Q 
                           => n424, QN => net245386);
   REGISTERS_reg_23_30_inst : DFF_X1 port map( D => n1150, CK => net199523, Q 
                           => n423, QN => net245385);
   REGISTERS_reg_23_29_inst : DFF_X1 port map( D => n1172, CK => net199523, Q 
                           => n422, QN => net245384);
   REGISTERS_reg_23_28_inst : DFF_X1 port map( D => n1194, CK => net199523, Q 
                           => n421, QN => net245383);
   REGISTERS_reg_23_27_inst : DFF_X1 port map( D => n1216, CK => net199523, Q 
                           => n420, QN => net245382);
   REGISTERS_reg_23_26_inst : DFF_X1 port map( D => n1238, CK => net199523, Q 
                           => n419, QN => net245381);
   REGISTERS_reg_23_25_inst : DFF_X1 port map( D => n1260, CK => net199523, Q 
                           => n418, QN => net245380);
   REGISTERS_reg_23_24_inst : DFF_X1 port map( D => n1282, CK => net199523, Q 
                           => n417, QN => net245379);
   REGISTERS_reg_23_23_inst : DFF_X1 port map( D => n1304, CK => net199523, Q 
                           => n416, QN => net245378);
   REGISTERS_reg_23_22_inst : DFF_X1 port map( D => n1326, CK => net199523, Q 
                           => n415, QN => net245377);
   REGISTERS_reg_23_21_inst : DFF_X1 port map( D => n1348, CK => net199523, Q 
                           => n414, QN => net245376);
   REGISTERS_reg_23_20_inst : DFF_X1 port map( D => n1370, CK => net199523, Q 
                           => n413, QN => net245375);
   REGISTERS_reg_23_19_inst : DFF_X1 port map( D => n1392, CK => net199523, Q 
                           => n412, QN => net245374);
   REGISTERS_reg_23_18_inst : DFF_X1 port map( D => n1414, CK => net199523, Q 
                           => n411, QN => net245373);
   REGISTERS_reg_23_17_inst : DFF_X1 port map( D => n1436, CK => net199523, Q 
                           => n410, QN => net245372);
   REGISTERS_reg_23_16_inst : DFF_X1 port map( D => n1458, CK => net199523, Q 
                           => n409, QN => net245371);
   REGISTERS_reg_23_15_inst : DFF_X1 port map( D => n1480, CK => net199523, Q 
                           => n408, QN => net245370);
   REGISTERS_reg_23_14_inst : DFF_X1 port map( D => n1502, CK => net199523, Q 
                           => n407, QN => net245369);
   REGISTERS_reg_23_13_inst : DFF_X1 port map( D => n1524, CK => net199523, Q 
                           => n406, QN => net245368);
   REGISTERS_reg_23_12_inst : DFF_X1 port map( D => n1546, CK => net199523, Q 
                           => n405, QN => net245367);
   REGISTERS_reg_23_11_inst : DFF_X1 port map( D => n1568, CK => net199523, Q 
                           => n404, QN => net245366);
   REGISTERS_reg_23_10_inst : DFF_X1 port map( D => n1590, CK => net199523, Q 
                           => n403, QN => net245365);
   REGISTERS_reg_23_9_inst : DFF_X1 port map( D => n1612, CK => net199523, Q =>
                           n402, QN => net245364);
   REGISTERS_reg_23_8_inst : DFF_X1 port map( D => n1634, CK => net199523, Q =>
                           n401, QN => net245363);
   REGISTERS_reg_23_7_inst : DFF_X1 port map( D => n1656, CK => net199523, Q =>
                           n400, QN => net245362);
   REGISTERS_reg_23_6_inst : DFF_X1 port map( D => n1678, CK => net199523, Q =>
                           n399, QN => net245361);
   REGISTERS_reg_23_5_inst : DFF_X1 port map( D => n1700, CK => net199523, Q =>
                           n398, QN => net245360);
   REGISTERS_reg_23_4_inst : DFF_X1 port map( D => n1722, CK => net199523, Q =>
                           n397, QN => net245359);
   REGISTERS_reg_23_3_inst : DFF_X1 port map( D => n1744, CK => net199523, Q =>
                           n396, QN => net245358);
   REGISTERS_reg_23_2_inst : DFF_X1 port map( D => n1766, CK => net199523, Q =>
                           n395, QN => net245357);
   REGISTERS_reg_23_1_inst : DFF_X1 port map( D => n1788, CK => net199523, Q =>
                           n394, QN => net245356);
   REGISTERS_reg_23_0_inst : DFF_X1 port map( D => n1810, CK => net199523, Q =>
                           n393, QN => net245355);
   REGISTERS_reg_24_31_inst : DFF_X1 port map( D => n1094, CK => net199528, Q 
                           => n392, QN => net245354);
   REGISTERS_reg_24_30_inst : DFF_X1 port map( D => n1150, CK => net199528, Q 
                           => n391, QN => net245353);
   REGISTERS_reg_24_29_inst : DFF_X1 port map( D => n1172, CK => net199528, Q 
                           => n390, QN => net245352);
   REGISTERS_reg_24_28_inst : DFF_X1 port map( D => n1194, CK => net199528, Q 
                           => n389, QN => net245351);
   REGISTERS_reg_24_27_inst : DFF_X1 port map( D => n1216, CK => net199528, Q 
                           => n388, QN => net245350);
   REGISTERS_reg_24_26_inst : DFF_X1 port map( D => n1238, CK => net199528, Q 
                           => n387, QN => net245349);
   REGISTERS_reg_24_25_inst : DFF_X1 port map( D => n1260, CK => net199528, Q 
                           => n386, QN => net245348);
   REGISTERS_reg_24_24_inst : DFF_X1 port map( D => n1282, CK => net199528, Q 
                           => n385, QN => net245347);
   REGISTERS_reg_24_23_inst : DFF_X1 port map( D => n1304, CK => net199528, Q 
                           => n384, QN => net245346);
   REGISTERS_reg_24_22_inst : DFF_X1 port map( D => n1326, CK => net199528, Q 
                           => n383, QN => net245345);
   REGISTERS_reg_24_21_inst : DFF_X1 port map( D => n1348, CK => net199528, Q 
                           => n382, QN => net245344);
   REGISTERS_reg_24_20_inst : DFF_X1 port map( D => n1370, CK => net199528, Q 
                           => n381, QN => net245343);
   REGISTERS_reg_24_19_inst : DFF_X1 port map( D => n1392, CK => net199528, Q 
                           => n380, QN => net245342);
   REGISTERS_reg_24_18_inst : DFF_X1 port map( D => n1414, CK => net199528, Q 
                           => n379, QN => net245341);
   REGISTERS_reg_24_17_inst : DFF_X1 port map( D => n1436, CK => net199528, Q 
                           => n378, QN => net245340);
   REGISTERS_reg_24_16_inst : DFF_X1 port map( D => n1458, CK => net199528, Q 
                           => n377, QN => net245339);
   REGISTERS_reg_24_15_inst : DFF_X1 port map( D => n1480, CK => net199528, Q 
                           => n376, QN => net245338);
   REGISTERS_reg_24_14_inst : DFF_X1 port map( D => n1502, CK => net199528, Q 
                           => n375, QN => net245337);
   REGISTERS_reg_24_13_inst : DFF_X1 port map( D => n1524, CK => net199528, Q 
                           => n374, QN => net245336);
   REGISTERS_reg_24_12_inst : DFF_X1 port map( D => n1546, CK => net199528, Q 
                           => n373, QN => net245335);
   REGISTERS_reg_24_11_inst : DFF_X1 port map( D => n1568, CK => net199528, Q 
                           => n372, QN => net245334);
   REGISTERS_reg_24_10_inst : DFF_X1 port map( D => n1590, CK => net199528, Q 
                           => n371, QN => net245333);
   REGISTERS_reg_24_9_inst : DFF_X1 port map( D => n1612, CK => net199528, Q =>
                           n370, QN => net245332);
   REGISTERS_reg_24_8_inst : DFF_X1 port map( D => n1634, CK => net199528, Q =>
                           n369, QN => net245331);
   REGISTERS_reg_24_7_inst : DFF_X1 port map( D => n1656, CK => net199528, Q =>
                           n368, QN => net245330);
   REGISTERS_reg_24_6_inst : DFF_X1 port map( D => n1678, CK => net199528, Q =>
                           n367, QN => net245329);
   REGISTERS_reg_24_5_inst : DFF_X1 port map( D => n1700, CK => net199528, Q =>
                           n366, QN => net245328);
   REGISTERS_reg_24_4_inst : DFF_X1 port map( D => n1722, CK => net199528, Q =>
                           n365, QN => net245327);
   REGISTERS_reg_24_3_inst : DFF_X1 port map( D => n1744, CK => net199528, Q =>
                           n364, QN => net245326);
   REGISTERS_reg_24_2_inst : DFF_X1 port map( D => n1766, CK => net199528, Q =>
                           n363, QN => net245325);
   REGISTERS_reg_24_1_inst : DFF_X1 port map( D => n1788, CK => net199528, Q =>
                           n362, QN => net245324);
   REGISTERS_reg_24_0_inst : DFF_X1 port map( D => n1810, CK => net199528, Q =>
                           n361, QN => net245323);
   REGISTERS_reg_25_31_inst : DFF_X1 port map( D => n1094, CK => net199533, Q 
                           => n360, QN => net245322);
   REGISTERS_reg_25_30_inst : DFF_X1 port map( D => n1150, CK => net199533, Q 
                           => n359, QN => net245321);
   REGISTERS_reg_25_29_inst : DFF_X1 port map( D => n1172, CK => net199533, Q 
                           => n358, QN => net245320);
   REGISTERS_reg_25_28_inst : DFF_X1 port map( D => n1194, CK => net199533, Q 
                           => n357, QN => net245319);
   REGISTERS_reg_25_27_inst : DFF_X1 port map( D => n1216, CK => net199533, Q 
                           => n356, QN => net245318);
   REGISTERS_reg_25_26_inst : DFF_X1 port map( D => n1238, CK => net199533, Q 
                           => n355, QN => net245317);
   REGISTERS_reg_25_25_inst : DFF_X1 port map( D => n1260, CK => net199533, Q 
                           => n354, QN => net245316);
   REGISTERS_reg_25_24_inst : DFF_X1 port map( D => n1282, CK => net199533, Q 
                           => n353, QN => net245315);
   REGISTERS_reg_25_23_inst : DFF_X1 port map( D => n1304, CK => net199533, Q 
                           => n352, QN => net245314);
   REGISTERS_reg_25_22_inst : DFF_X1 port map( D => n1326, CK => net199533, Q 
                           => n351, QN => net245313);
   REGISTERS_reg_25_21_inst : DFF_X1 port map( D => n1348, CK => net199533, Q 
                           => n350, QN => net245312);
   REGISTERS_reg_25_20_inst : DFF_X1 port map( D => n1370, CK => net199533, Q 
                           => n349, QN => net245311);
   REGISTERS_reg_25_19_inst : DFF_X1 port map( D => n1392, CK => net199533, Q 
                           => n348, QN => net245310);
   REGISTERS_reg_25_18_inst : DFF_X1 port map( D => n1414, CK => net199533, Q 
                           => n347, QN => net245309);
   REGISTERS_reg_25_17_inst : DFF_X1 port map( D => n1436, CK => net199533, Q 
                           => n346, QN => net245308);
   REGISTERS_reg_25_16_inst : DFF_X1 port map( D => n1458, CK => net199533, Q 
                           => n345, QN => net245307);
   REGISTERS_reg_25_15_inst : DFF_X1 port map( D => n1480, CK => net199533, Q 
                           => n344, QN => net245306);
   REGISTERS_reg_25_14_inst : DFF_X1 port map( D => n1502, CK => net199533, Q 
                           => n343, QN => net245305);
   REGISTERS_reg_25_13_inst : DFF_X1 port map( D => n1524, CK => net199533, Q 
                           => n342, QN => net245304);
   REGISTERS_reg_25_12_inst : DFF_X1 port map( D => n1546, CK => net199533, Q 
                           => n341, QN => net245303);
   REGISTERS_reg_25_11_inst : DFF_X1 port map( D => n1568, CK => net199533, Q 
                           => n340, QN => net245302);
   REGISTERS_reg_25_10_inst : DFF_X1 port map( D => n1590, CK => net199533, Q 
                           => n339, QN => net245301);
   REGISTERS_reg_25_9_inst : DFF_X1 port map( D => n1612, CK => net199533, Q =>
                           n338, QN => net245300);
   REGISTERS_reg_25_8_inst : DFF_X1 port map( D => n1634, CK => net199533, Q =>
                           n337, QN => net245299);
   REGISTERS_reg_25_7_inst : DFF_X1 port map( D => n1656, CK => net199533, Q =>
                           n336, QN => net245298);
   REGISTERS_reg_25_6_inst : DFF_X1 port map( D => n1678, CK => net199533, Q =>
                           n335, QN => net245297);
   REGISTERS_reg_25_5_inst : DFF_X1 port map( D => n1700, CK => net199533, Q =>
                           n334, QN => net245296);
   REGISTERS_reg_25_4_inst : DFF_X1 port map( D => n1722, CK => net199533, Q =>
                           n333, QN => net245295);
   REGISTERS_reg_25_3_inst : DFF_X1 port map( D => n1744, CK => net199533, Q =>
                           n332, QN => net245294);
   REGISTERS_reg_25_2_inst : DFF_X1 port map( D => n1766, CK => net199533, Q =>
                           n331, QN => net245293);
   REGISTERS_reg_25_1_inst : DFF_X1 port map( D => n1788, CK => net199533, Q =>
                           n330, QN => net245292);
   REGISTERS_reg_25_0_inst : DFF_X1 port map( D => n1810, CK => net199533, Q =>
                           n329, QN => net245291);
   REGISTERS_reg_26_31_inst : DFF_X1 port map( D => n1094, CK => net199538, Q 
                           => n328, QN => net245290);
   REGISTERS_reg_26_30_inst : DFF_X1 port map( D => n1150, CK => net199538, Q 
                           => n327, QN => net245289);
   REGISTERS_reg_26_29_inst : DFF_X1 port map( D => n1172, CK => net199538, Q 
                           => n326, QN => net245288);
   REGISTERS_reg_26_28_inst : DFF_X1 port map( D => n1194, CK => net199538, Q 
                           => n325, QN => net245287);
   REGISTERS_reg_26_27_inst : DFF_X1 port map( D => n1216, CK => net199538, Q 
                           => n324, QN => net245286);
   REGISTERS_reg_26_26_inst : DFF_X1 port map( D => n1238, CK => net199538, Q 
                           => n323, QN => net245285);
   REGISTERS_reg_26_25_inst : DFF_X1 port map( D => n1260, CK => net199538, Q 
                           => n322, QN => net245284);
   REGISTERS_reg_26_24_inst : DFF_X1 port map( D => n1282, CK => net199538, Q 
                           => n321, QN => net245283);
   REGISTERS_reg_26_23_inst : DFF_X1 port map( D => n1304, CK => net199538, Q 
                           => n320, QN => net245282);
   REGISTERS_reg_26_22_inst : DFF_X1 port map( D => n1326, CK => net199538, Q 
                           => n319, QN => net245281);
   REGISTERS_reg_26_21_inst : DFF_X1 port map( D => n1348, CK => net199538, Q 
                           => n318, QN => net245280);
   REGISTERS_reg_26_20_inst : DFF_X1 port map( D => n1370, CK => net199538, Q 
                           => n317, QN => net245279);
   REGISTERS_reg_26_19_inst : DFF_X1 port map( D => n1392, CK => net199538, Q 
                           => n316, QN => net245278);
   REGISTERS_reg_26_18_inst : DFF_X1 port map( D => n1414, CK => net199538, Q 
                           => n315, QN => net245277);
   REGISTERS_reg_26_17_inst : DFF_X1 port map( D => n1436, CK => net199538, Q 
                           => n314, QN => net245276);
   REGISTERS_reg_26_16_inst : DFF_X1 port map( D => n1458, CK => net199538, Q 
                           => n313, QN => net245275);
   REGISTERS_reg_26_15_inst : DFF_X1 port map( D => n1480, CK => net199538, Q 
                           => n312, QN => net245274);
   REGISTERS_reg_26_14_inst : DFF_X1 port map( D => n1502, CK => net199538, Q 
                           => n311, QN => net245273);
   REGISTERS_reg_26_13_inst : DFF_X1 port map( D => n1524, CK => net199538, Q 
                           => n310, QN => net245272);
   REGISTERS_reg_26_12_inst : DFF_X1 port map( D => n1546, CK => net199538, Q 
                           => n309, QN => net245271);
   REGISTERS_reg_26_11_inst : DFF_X1 port map( D => n1568, CK => net199538, Q 
                           => n308, QN => net245270);
   REGISTERS_reg_26_10_inst : DFF_X1 port map( D => n1590, CK => net199538, Q 
                           => n307, QN => net245269);
   REGISTERS_reg_26_9_inst : DFF_X1 port map( D => n1612, CK => net199538, Q =>
                           n306, QN => net245268);
   REGISTERS_reg_26_8_inst : DFF_X1 port map( D => n1634, CK => net199538, Q =>
                           n305, QN => net245267);
   REGISTERS_reg_26_7_inst : DFF_X1 port map( D => n1656, CK => net199538, Q =>
                           n304, QN => net245266);
   REGISTERS_reg_26_6_inst : DFF_X1 port map( D => n1678, CK => net199538, Q =>
                           n303, QN => net245265);
   REGISTERS_reg_26_5_inst : DFF_X1 port map( D => n1700, CK => net199538, Q =>
                           n302, QN => net245264);
   REGISTERS_reg_26_4_inst : DFF_X1 port map( D => n1722, CK => net199538, Q =>
                           n301, QN => net245263);
   REGISTERS_reg_26_3_inst : DFF_X1 port map( D => n1744, CK => net199538, Q =>
                           n300, QN => net245262);
   REGISTERS_reg_26_2_inst : DFF_X1 port map( D => n1766, CK => net199538, Q =>
                           n299, QN => net245261);
   REGISTERS_reg_26_1_inst : DFF_X1 port map( D => n1788, CK => net199538, Q =>
                           n298, QN => net245260);
   REGISTERS_reg_26_0_inst : DFF_X1 port map( D => n1810, CK => net199538, Q =>
                           n297, QN => net245259);
   REGISTERS_reg_27_31_inst : DFF_X1 port map( D => n1094, CK => net199543, Q 
                           => n296, QN => net245258);
   REGISTERS_reg_27_30_inst : DFF_X1 port map( D => n1150, CK => net199543, Q 
                           => n295, QN => net245257);
   REGISTERS_reg_27_29_inst : DFF_X1 port map( D => n1172, CK => net199543, Q 
                           => n294, QN => net245256);
   REGISTERS_reg_27_28_inst : DFF_X1 port map( D => n1194, CK => net199543, Q 
                           => n293, QN => net245255);
   REGISTERS_reg_27_27_inst : DFF_X1 port map( D => n1216, CK => net199543, Q 
                           => n292, QN => net245254);
   REGISTERS_reg_27_26_inst : DFF_X1 port map( D => n1238, CK => net199543, Q 
                           => n291, QN => net245253);
   REGISTERS_reg_27_25_inst : DFF_X1 port map( D => n1260, CK => net199543, Q 
                           => n290, QN => net245252);
   REGISTERS_reg_27_24_inst : DFF_X1 port map( D => n1282, CK => net199543, Q 
                           => n289, QN => net245251);
   REGISTERS_reg_27_23_inst : DFF_X1 port map( D => n1304, CK => net199543, Q 
                           => n288, QN => net245250);
   REGISTERS_reg_27_22_inst : DFF_X1 port map( D => n1326, CK => net199543, Q 
                           => n287, QN => net245249);
   REGISTERS_reg_27_21_inst : DFF_X1 port map( D => n1348, CK => net199543, Q 
                           => n286, QN => net245248);
   REGISTERS_reg_27_20_inst : DFF_X1 port map( D => n1370, CK => net199543, Q 
                           => n285, QN => net245247);
   REGISTERS_reg_27_19_inst : DFF_X1 port map( D => n1392, CK => net199543, Q 
                           => n284, QN => net245246);
   REGISTERS_reg_27_18_inst : DFF_X1 port map( D => n1414, CK => net199543, Q 
                           => n283, QN => net245245);
   REGISTERS_reg_27_17_inst : DFF_X1 port map( D => n1436, CK => net199543, Q 
                           => n282, QN => net245244);
   REGISTERS_reg_27_16_inst : DFF_X1 port map( D => n1458, CK => net199543, Q 
                           => n281, QN => net245243);
   REGISTERS_reg_27_15_inst : DFF_X1 port map( D => n1480, CK => net199543, Q 
                           => n280, QN => net245242);
   REGISTERS_reg_27_14_inst : DFF_X1 port map( D => n1502, CK => net199543, Q 
                           => n279, QN => net245241);
   REGISTERS_reg_27_13_inst : DFF_X1 port map( D => n1524, CK => net199543, Q 
                           => n278, QN => net245240);
   REGISTERS_reg_27_12_inst : DFF_X1 port map( D => n1546, CK => net199543, Q 
                           => n277, QN => net245239);
   REGISTERS_reg_27_11_inst : DFF_X1 port map( D => n1568, CK => net199543, Q 
                           => n276, QN => net245238);
   REGISTERS_reg_27_10_inst : DFF_X1 port map( D => n1590, CK => net199543, Q 
                           => n275, QN => net245237);
   REGISTERS_reg_27_9_inst : DFF_X1 port map( D => n1612, CK => net199543, Q =>
                           n274, QN => net245236);
   REGISTERS_reg_27_8_inst : DFF_X1 port map( D => n1634, CK => net199543, Q =>
                           n273, QN => net245235);
   REGISTERS_reg_27_7_inst : DFF_X1 port map( D => n1656, CK => net199543, Q =>
                           n272, QN => net245234);
   REGISTERS_reg_27_6_inst : DFF_X1 port map( D => n1678, CK => net199543, Q =>
                           n271, QN => net245233);
   REGISTERS_reg_27_5_inst : DFF_X1 port map( D => n1700, CK => net199543, Q =>
                           n270, QN => net245232);
   REGISTERS_reg_27_4_inst : DFF_X1 port map( D => n1722, CK => net199543, Q =>
                           n269, QN => net245231);
   REGISTERS_reg_27_3_inst : DFF_X1 port map( D => n1744, CK => net199543, Q =>
                           n268, QN => net245230);
   REGISTERS_reg_27_2_inst : DFF_X1 port map( D => n1766, CK => net199543, Q =>
                           n267, QN => net245229);
   REGISTERS_reg_27_1_inst : DFF_X1 port map( D => n1788, CK => net199543, Q =>
                           n266, QN => net245228);
   REGISTERS_reg_27_0_inst : DFF_X1 port map( D => n1810, CK => net199543, Q =>
                           n265, QN => net245227);
   REGISTERS_reg_28_31_inst : DFF_X1 port map( D => n1094, CK => net199548, Q 
                           => n264, QN => net245226);
   REGISTERS_reg_28_30_inst : DFF_X1 port map( D => n1150, CK => net199548, Q 
                           => n263, QN => net245225);
   REGISTERS_reg_28_29_inst : DFF_X1 port map( D => n1172, CK => net199548, Q 
                           => n262, QN => net245224);
   REGISTERS_reg_28_28_inst : DFF_X1 port map( D => n1194, CK => net199548, Q 
                           => n261, QN => net245223);
   REGISTERS_reg_28_27_inst : DFF_X1 port map( D => n1216, CK => net199548, Q 
                           => n260, QN => net245222);
   REGISTERS_reg_28_26_inst : DFF_X1 port map( D => n1238, CK => net199548, Q 
                           => n259, QN => net245221);
   REGISTERS_reg_28_25_inst : DFF_X1 port map( D => n1260, CK => net199548, Q 
                           => n258, QN => net245220);
   REGISTERS_reg_28_24_inst : DFF_X1 port map( D => n1282, CK => net199548, Q 
                           => n257, QN => net245219);
   REGISTERS_reg_28_23_inst : DFF_X1 port map( D => n1304, CK => net199548, Q 
                           => n256, QN => net245218);
   REGISTERS_reg_28_22_inst : DFF_X1 port map( D => n1326, CK => net199548, Q 
                           => n255, QN => net245217);
   REGISTERS_reg_28_21_inst : DFF_X1 port map( D => n1348, CK => net199548, Q 
                           => n254, QN => net245216);
   REGISTERS_reg_28_20_inst : DFF_X1 port map( D => n1370, CK => net199548, Q 
                           => n253, QN => net245215);
   REGISTERS_reg_28_19_inst : DFF_X1 port map( D => n1392, CK => net199548, Q 
                           => n252, QN => net245214);
   REGISTERS_reg_28_18_inst : DFF_X1 port map( D => n1414, CK => net199548, Q 
                           => n251, QN => net245213);
   REGISTERS_reg_28_17_inst : DFF_X1 port map( D => n1436, CK => net199548, Q 
                           => n250, QN => net245212);
   REGISTERS_reg_28_16_inst : DFF_X1 port map( D => n1458, CK => net199548, Q 
                           => n249, QN => net245211);
   REGISTERS_reg_28_15_inst : DFF_X1 port map( D => n1480, CK => net199548, Q 
                           => n248, QN => net245210);
   REGISTERS_reg_28_14_inst : DFF_X1 port map( D => n1502, CK => net199548, Q 
                           => n247, QN => net245209);
   REGISTERS_reg_28_13_inst : DFF_X1 port map( D => n1524, CK => net199548, Q 
                           => n246, QN => net245208);
   REGISTERS_reg_28_12_inst : DFF_X1 port map( D => n1546, CK => net199548, Q 
                           => n245, QN => net245207);
   REGISTERS_reg_28_11_inst : DFF_X1 port map( D => n1568, CK => net199548, Q 
                           => n244, QN => net245206);
   REGISTERS_reg_28_10_inst : DFF_X1 port map( D => n1590, CK => net199548, Q 
                           => n243, QN => net245205);
   REGISTERS_reg_28_9_inst : DFF_X1 port map( D => n1612, CK => net199548, Q =>
                           n242, QN => net245204);
   REGISTERS_reg_28_8_inst : DFF_X1 port map( D => n1634, CK => net199548, Q =>
                           n241, QN => net245203);
   REGISTERS_reg_28_7_inst : DFF_X1 port map( D => n1656, CK => net199548, Q =>
                           n240, QN => net245202);
   REGISTERS_reg_28_6_inst : DFF_X1 port map( D => n1678, CK => net199548, Q =>
                           n239, QN => net245201);
   REGISTERS_reg_28_5_inst : DFF_X1 port map( D => n1700, CK => net199548, Q =>
                           n238, QN => net245200);
   REGISTERS_reg_28_4_inst : DFF_X1 port map( D => n1722, CK => net199548, Q =>
                           n237, QN => net245199);
   REGISTERS_reg_28_3_inst : DFF_X1 port map( D => n1744, CK => net199548, Q =>
                           n236, QN => net245198);
   REGISTERS_reg_28_2_inst : DFF_X1 port map( D => n1766, CK => net199548, Q =>
                           n235, QN => net245197);
   REGISTERS_reg_28_1_inst : DFF_X1 port map( D => n1788, CK => net199548, Q =>
                           n234, QN => net245196);
   REGISTERS_reg_28_0_inst : DFF_X1 port map( D => n1810, CK => net199548, Q =>
                           n233, QN => net245195);
   REGISTERS_reg_29_31_inst : DFF_X1 port map( D => n1094, CK => net199553, Q 
                           => n232, QN => net245194);
   REGISTERS_reg_29_30_inst : DFF_X1 port map( D => n1150, CK => net199553, Q 
                           => n231, QN => net245193);
   REGISTERS_reg_29_29_inst : DFF_X1 port map( D => n1172, CK => net199553, Q 
                           => n230, QN => net245192);
   REGISTERS_reg_29_28_inst : DFF_X1 port map( D => n1194, CK => net199553, Q 
                           => n229, QN => net245191);
   REGISTERS_reg_29_27_inst : DFF_X1 port map( D => n1216, CK => net199553, Q 
                           => n228, QN => net245190);
   REGISTERS_reg_29_26_inst : DFF_X1 port map( D => n1238, CK => net199553, Q 
                           => n227, QN => net245189);
   REGISTERS_reg_29_25_inst : DFF_X1 port map( D => n1260, CK => net199553, Q 
                           => n226, QN => net245188);
   REGISTERS_reg_29_24_inst : DFF_X1 port map( D => n1282, CK => net199553, Q 
                           => n225, QN => net245187);
   REGISTERS_reg_29_23_inst : DFF_X1 port map( D => n1304, CK => net199553, Q 
                           => n224, QN => net245186);
   REGISTERS_reg_29_22_inst : DFF_X1 port map( D => n1326, CK => net199553, Q 
                           => n223, QN => net245185);
   REGISTERS_reg_29_21_inst : DFF_X1 port map( D => n1348, CK => net199553, Q 
                           => n222, QN => net245184);
   REGISTERS_reg_29_20_inst : DFF_X1 port map( D => n1370, CK => net199553, Q 
                           => n221, QN => net245183);
   REGISTERS_reg_29_19_inst : DFF_X1 port map( D => n1392, CK => net199553, Q 
                           => n220, QN => net245182);
   REGISTERS_reg_29_18_inst : DFF_X1 port map( D => n1414, CK => net199553, Q 
                           => n219, QN => net245181);
   REGISTERS_reg_29_17_inst : DFF_X1 port map( D => n1436, CK => net199553, Q 
                           => n218, QN => net245180);
   REGISTERS_reg_29_16_inst : DFF_X1 port map( D => n1458, CK => net199553, Q 
                           => n217, QN => net245179);
   REGISTERS_reg_29_15_inst : DFF_X1 port map( D => n1480, CK => net199553, Q 
                           => n216, QN => net245178);
   REGISTERS_reg_29_14_inst : DFF_X1 port map( D => n1502, CK => net199553, Q 
                           => n215, QN => net245177);
   REGISTERS_reg_29_13_inst : DFF_X1 port map( D => n1524, CK => net199553, Q 
                           => n214, QN => net245176);
   REGISTERS_reg_29_12_inst : DFF_X1 port map( D => n1546, CK => net199553, Q 
                           => n213, QN => net245175);
   REGISTERS_reg_29_11_inst : DFF_X1 port map( D => n1568, CK => net199553, Q 
                           => n212, QN => net245174);
   REGISTERS_reg_29_10_inst : DFF_X1 port map( D => n1590, CK => net199553, Q 
                           => n211, QN => net245173);
   REGISTERS_reg_29_9_inst : DFF_X1 port map( D => n1612, CK => net199553, Q =>
                           n210, QN => net245172);
   REGISTERS_reg_29_8_inst : DFF_X1 port map( D => n1634, CK => net199553, Q =>
                           n209, QN => net245171);
   REGISTERS_reg_29_7_inst : DFF_X1 port map( D => n1656, CK => net199553, Q =>
                           n208, QN => net245170);
   REGISTERS_reg_29_6_inst : DFF_X1 port map( D => n1678, CK => net199553, Q =>
                           n207, QN => net245169);
   REGISTERS_reg_29_5_inst : DFF_X1 port map( D => n1700, CK => net199553, Q =>
                           n206, QN => net245168);
   REGISTERS_reg_29_4_inst : DFF_X1 port map( D => n1722, CK => net199553, Q =>
                           n205, QN => net245167);
   REGISTERS_reg_29_3_inst : DFF_X1 port map( D => n1744, CK => net199553, Q =>
                           n204, QN => net245166);
   REGISTERS_reg_29_2_inst : DFF_X1 port map( D => n1766, CK => net199553, Q =>
                           n203, QN => net245165);
   REGISTERS_reg_29_1_inst : DFF_X1 port map( D => n1788, CK => net199553, Q =>
                           n202, QN => net245164);
   REGISTERS_reg_29_0_inst : DFF_X1 port map( D => n1810, CK => net199553, Q =>
                           n201, QN => net245163);
   REGISTERS_reg_30_31_inst : DFF_X1 port map( D => n1094, CK => net199558, Q 
                           => n200, QN => net245162);
   REGISTERS_reg_30_30_inst : DFF_X1 port map( D => n1150, CK => net199558, Q 
                           => n199, QN => net245161);
   REGISTERS_reg_30_29_inst : DFF_X1 port map( D => n1172, CK => net199558, Q 
                           => n198, QN => net245160);
   REGISTERS_reg_30_28_inst : DFF_X1 port map( D => n1194, CK => net199558, Q 
                           => n197, QN => net245159);
   REGISTERS_reg_30_27_inst : DFF_X1 port map( D => n1216, CK => net199558, Q 
                           => n196, QN => net245158);
   REGISTERS_reg_30_26_inst : DFF_X1 port map( D => n1238, CK => net199558, Q 
                           => n195, QN => net245157);
   REGISTERS_reg_30_25_inst : DFF_X1 port map( D => n1260, CK => net199558, Q 
                           => n194, QN => net245156);
   REGISTERS_reg_30_24_inst : DFF_X1 port map( D => n1282, CK => net199558, Q 
                           => n193, QN => net245155);
   REGISTERS_reg_30_23_inst : DFF_X1 port map( D => n1304, CK => net199558, Q 
                           => n192, QN => net245154);
   REGISTERS_reg_30_22_inst : DFF_X1 port map( D => n1326, CK => net199558, Q 
                           => n191, QN => net245153);
   REGISTERS_reg_30_21_inst : DFF_X1 port map( D => n1348, CK => net199558, Q 
                           => n190, QN => net245152);
   REGISTERS_reg_30_20_inst : DFF_X1 port map( D => n1370, CK => net199558, Q 
                           => n189, QN => net245151);
   REGISTERS_reg_30_19_inst : DFF_X1 port map( D => n1392, CK => net199558, Q 
                           => n188, QN => net245150);
   REGISTERS_reg_30_18_inst : DFF_X1 port map( D => n1414, CK => net199558, Q 
                           => n187, QN => net245149);
   REGISTERS_reg_30_17_inst : DFF_X1 port map( D => n1436, CK => net199558, Q 
                           => n186, QN => net245148);
   REGISTERS_reg_30_16_inst : DFF_X1 port map( D => n1458, CK => net199558, Q 
                           => n185, QN => net245147);
   REGISTERS_reg_30_15_inst : DFF_X1 port map( D => n1480, CK => net199558, Q 
                           => n184, QN => net245146);
   REGISTERS_reg_30_14_inst : DFF_X1 port map( D => n1502, CK => net199558, Q 
                           => n183, QN => net245145);
   REGISTERS_reg_30_13_inst : DFF_X1 port map( D => n1524, CK => net199558, Q 
                           => n182, QN => net245144);
   REGISTERS_reg_30_12_inst : DFF_X1 port map( D => n1546, CK => net199558, Q 
                           => n181, QN => net245143);
   REGISTERS_reg_30_11_inst : DFF_X1 port map( D => n1568, CK => net199558, Q 
                           => n180, QN => net245142);
   REGISTERS_reg_30_10_inst : DFF_X1 port map( D => n1590, CK => net199558, Q 
                           => n179, QN => net245141);
   REGISTERS_reg_30_9_inst : DFF_X1 port map( D => n1612, CK => net199558, Q =>
                           n176, QN => net245140);
   REGISTERS_reg_30_8_inst : DFF_X1 port map( D => n1634, CK => net199558, Q =>
                           n165, QN => net245139);
   REGISTERS_reg_30_7_inst : DFF_X1 port map( D => n1656, CK => net199558, Q =>
                           n154, QN => net245138);
   REGISTERS_reg_30_6_inst : DFF_X1 port map( D => n1678, CK => net199558, Q =>
                           n143, QN => net245137);
   REGISTERS_reg_30_5_inst : DFF_X1 port map( D => n1700, CK => net199558, Q =>
                           n132, QN => net245136);
   REGISTERS_reg_30_4_inst : DFF_X1 port map( D => n1722, CK => net199558, Q =>
                           n121, QN => net245135);
   REGISTERS_reg_30_3_inst : DFF_X1 port map( D => n1744, CK => net199558, Q =>
                           n110, QN => net245134);
   REGISTERS_reg_30_2_inst : DFF_X1 port map( D => n1766, CK => net199558, Q =>
                           n99, QN => net245133);
   REGISTERS_reg_30_1_inst : DFF_X1 port map( D => n1788, CK => net199558, Q =>
                           n77, QN => net245132);
   REGISTERS_reg_30_0_inst : DFF_X1 port map( D => n1810, CK => net199558, Q =>
                           n55, QN => net245131);
   REGISTERS_reg_31_31_inst : DFF_X1 port map( D => n1094, CK => net199563, Q 
                           => n1090, QN => net245130);
   OUT2_reg_31_inst : DFF_X1 port map( D => N4616, CK => net199403, Q => 
                           OUT2(31), QN => n98);
   REGISTERS_reg_31_30_inst : DFF_X1 port map( D => n1150, CK => net199563, Q 
                           => n1069, QN => net245129);
   OUT2_reg_30_inst : DFF_X1 port map( D => N4614, CK => net199403, Q => 
                           OUT2(30), QN => n96);
   REGISTERS_reg_31_29_inst : DFF_X1 port map( D => n1172, CK => net199563, Q 
                           => n1048, QN => net245128);
   OUT2_reg_29_inst : DFF_X1 port map( D => N4612, CK => net199403, Q => 
                           OUT2(29), QN => n94);
   REGISTERS_reg_31_28_inst : DFF_X1 port map( D => n1194, CK => net199563, Q 
                           => n1027, QN => net245127);
   OUT2_reg_28_inst : DFF_X1 port map( D => N4610, CK => net199403, Q => 
                           OUT2(28), QN => n92);
   REGISTERS_reg_31_27_inst : DFF_X1 port map( D => n1216, CK => net199563, Q 
                           => n1006, QN => net245126);
   OUT2_reg_27_inst : DFF_X1 port map( D => N4608, CK => net199403, Q => 
                           OUT2(27), QN => n90);
   REGISTERS_reg_31_26_inst : DFF_X1 port map( D => n1238, CK => net199563, Q 
                           => n985, QN => net245125);
   OUT2_reg_26_inst : DFF_X1 port map( D => N4606, CK => net199403, Q => 
                           OUT2(26), QN => n88);
   REGISTERS_reg_31_25_inst : DFF_X1 port map( D => n1260, CK => net199563, Q 
                           => n964, QN => net245124);
   OUT2_reg_25_inst : DFF_X1 port map( D => N4604, CK => net199403, Q => 
                           OUT2(25), QN => n86);
   REGISTERS_reg_31_24_inst : DFF_X1 port map( D => n1282, CK => net199563, Q 
                           => n943, QN => net245123);
   OUT2_reg_24_inst : DFF_X1 port map( D => N4602, CK => net199403, Q => 
                           OUT2(24), QN => n84);
   REGISTERS_reg_31_23_inst : DFF_X1 port map( D => n1304, CK => net199563, Q 
                           => n922, QN => net245122);
   OUT2_reg_23_inst : DFF_X1 port map( D => N4600, CK => net199403, Q => 
                           OUT2(23), QN => n82);
   REGISTERS_reg_31_22_inst : DFF_X1 port map( D => n1326, CK => net199563, Q 
                           => n901, QN => net245121);
   OUT2_reg_22_inst : DFF_X1 port map( D => N4598, CK => net199403, Q => 
                           OUT2(22), QN => n80);
   REGISTERS_reg_31_21_inst : DFF_X1 port map( D => n1348, CK => net199563, Q 
                           => n880, QN => net245120);
   OUT2_reg_21_inst : DFF_X1 port map( D => N4596, CK => net199403, Q => 
                           OUT2(21), QN => n78);
   REGISTERS_reg_31_20_inst : DFF_X1 port map( D => n1370, CK => net199563, Q 
                           => n859, QN => net245119);
   OUT2_reg_20_inst : DFF_X1 port map( D => N4594, CK => net199403, Q => 
                           OUT2(20), QN => n76);
   REGISTERS_reg_31_19_inst : DFF_X1 port map( D => n1392, CK => net199563, Q 
                           => n838, QN => net245118);
   OUT2_reg_19_inst : DFF_X1 port map( D => N4592, CK => net199403, Q => 
                           OUT2(19), QN => n74);
   REGISTERS_reg_31_18_inst : DFF_X1 port map( D => n1414, CK => net199563, Q 
                           => n817, QN => net245117);
   OUT2_reg_18_inst : DFF_X1 port map( D => N4590, CK => net199403, Q => 
                           OUT2(18), QN => n72);
   REGISTERS_reg_31_17_inst : DFF_X1 port map( D => n1436, CK => net199563, Q 
                           => n796, QN => net245116);
   OUT2_reg_17_inst : DFF_X1 port map( D => N4588, CK => net199403, Q => 
                           OUT2(17), QN => n70);
   REGISTERS_reg_31_16_inst : DFF_X1 port map( D => n1458, CK => net199563, Q 
                           => n775, QN => net245115);
   OUT2_reg_16_inst : DFF_X1 port map( D => N4586, CK => net199403, Q => 
                           OUT2(16), QN => n68);
   REGISTERS_reg_31_15_inst : DFF_X1 port map( D => n1480, CK => net199563, Q 
                           => n754, QN => net245114);
   OUT2_reg_15_inst : DFF_X1 port map( D => N4584, CK => net199403, Q => 
                           OUT2(15), QN => n66);
   REGISTERS_reg_31_14_inst : DFF_X1 port map( D => n1502, CK => net199563, Q 
                           => n733, QN => net245113);
   OUT2_reg_14_inst : DFF_X1 port map( D => N4582, CK => net199403, Q => 
                           OUT2(14), QN => n64);
   REGISTERS_reg_31_13_inst : DFF_X1 port map( D => n1524, CK => net199563, Q 
                           => n712, QN => net245112);
   OUT2_reg_13_inst : DFF_X1 port map( D => N4580, CK => net199403, Q => 
                           OUT2(13), QN => n62);
   REGISTERS_reg_31_12_inst : DFF_X1 port map( D => n1546, CK => net199563, Q 
                           => n691, QN => net245111);
   OUT2_reg_12_inst : DFF_X1 port map( D => N4578, CK => net199403, Q => 
                           OUT2(12), QN => n60);
   REGISTERS_reg_31_11_inst : DFF_X1 port map( D => n1568, CK => net199563, Q 
                           => n670, QN => net245110);
   OUT2_reg_11_inst : DFF_X1 port map( D => N4576, CK => net199403, Q => 
                           OUT2(11), QN => n58);
   REGISTERS_reg_31_10_inst : DFF_X1 port map( D => n1590, CK => net199563, Q 
                           => n649, QN => net245109);
   OUT2_reg_10_inst : DFF_X1 port map( D => N4574, CK => net199403, Q => 
                           OUT2(10), QN => n56);
   REGISTERS_reg_31_9_inst : DFF_X1 port map( D => n1612, CK => net199563, Q =>
                           n628, QN => net245108);
   OUT2_reg_9_inst : DFF_X1 port map( D => N4572, CK => net199403, Q => OUT2(9)
                           , QN => n54);
   REGISTERS_reg_31_8_inst : DFF_X1 port map( D => n1634, CK => net199563, Q =>
                           n607, QN => net245107);
   OUT2_reg_8_inst : DFF_X1 port map( D => N4570, CK => net199403, Q => OUT2(8)
                           , QN => n52);
   REGISTERS_reg_31_7_inst : DFF_X1 port map( D => n1656, CK => net199563, Q =>
                           n586, QN => net245106);
   OUT2_reg_7_inst : DFF_X1 port map( D => N4568, CK => net199403, Q => OUT2(7)
                           , QN => n50);
   REGISTERS_reg_31_6_inst : DFF_X1 port map( D => n1678, CK => net199563, Q =>
                           n565, QN => net245105);
   OUT2_reg_6_inst : DFF_X1 port map( D => N4566, CK => net199403, Q => OUT2(6)
                           , QN => n48);
   REGISTERS_reg_31_5_inst : DFF_X1 port map( D => n1700, CK => net199563, Q =>
                           n544, QN => net245104);
   OUT2_reg_5_inst : DFF_X1 port map( D => N4564, CK => net199403, Q => OUT2(5)
                           , QN => n46);
   REGISTERS_reg_31_4_inst : DFF_X1 port map( D => n1722, CK => net199563, Q =>
                           n523, QN => net245103);
   OUT2_reg_4_inst : DFF_X1 port map( D => N4562, CK => net199403, Q => OUT2(4)
                           , QN => n44);
   REGISTERS_reg_31_3_inst : DFF_X1 port map( D => n1744, CK => net199563, Q =>
                           n502, QN => net245102);
   OUT2_reg_3_inst : DFF_X1 port map( D => N4560, CK => net199403, Q => OUT2(3)
                           , QN => n42);
   REGISTERS_reg_31_2_inst : DFF_X1 port map( D => n1766, CK => net199563, Q =>
                           n481, QN => net245101);
   OUT2_reg_2_inst : DFF_X1 port map( D => N4558, CK => net199403, Q => OUT2(2)
                           , QN => n40);
   REGISTERS_reg_31_1_inst : DFF_X1 port map( D => n1788, CK => net199563, Q =>
                           n460, QN => net245100);
   OUT2_reg_1_inst : DFF_X1 port map( D => N4556, CK => net199403, Q => OUT2(1)
                           , QN => n38);
   REGISTERS_reg_31_0_inst : DFF_X1 port map( D => n1810, CK => net199563, Q =>
                           n439, QN => net245099);
   OUT2_reg_0_inst : DFF_X1 port map( D => N4554, CK => net199403, Q => OUT2(0)
                           , QN => n36);
   OUT1_reg_31_inst : DFF_X1 port map( D => N4552, CK => net199568, Q => 
                           OUT1(31), QN => n35);
   OUT1_reg_30_inst : DFF_X1 port map( D => N4550, CK => net199568, Q => 
                           OUT1(30), QN => n34);
   OUT1_reg_29_inst : DFF_X1 port map( D => N4548, CK => net199568, Q => 
                           OUT1(29), QN => n33);
   OUT1_reg_28_inst : DFF_X1 port map( D => N4546, CK => net199568, Q => 
                           OUT1(28), QN => n32);
   OUT1_reg_27_inst : DFF_X1 port map( D => N4544, CK => net199568, Q => 
                           OUT1(27), QN => n31);
   OUT1_reg_26_inst : DFF_X1 port map( D => N4542, CK => net199568, Q => 
                           OUT1(26), QN => n30);
   OUT1_reg_25_inst : DFF_X1 port map( D => N4540, CK => net199568, Q => 
                           OUT1(25), QN => n29);
   OUT1_reg_24_inst : DFF_X1 port map( D => N4538, CK => net199568, Q => 
                           OUT1(24), QN => n28);
   OUT1_reg_23_inst : DFF_X1 port map( D => N4536, CK => net199568, Q => 
                           OUT1(23), QN => n27);
   OUT1_reg_22_inst : DFF_X1 port map( D => N4534, CK => net199568, Q => 
                           OUT1(22), QN => n26);
   OUT1_reg_21_inst : DFF_X1 port map( D => N4532, CK => net199568, Q => 
                           OUT1(21), QN => n25);
   OUT1_reg_20_inst : DFF_X1 port map( D => N4530, CK => net199568, Q => 
                           OUT1(20), QN => n24);
   OUT1_reg_19_inst : DFF_X1 port map( D => N4528, CK => net199568, Q => 
                           OUT1(19), QN => n23);
   OUT1_reg_18_inst : DFF_X1 port map( D => N4526, CK => net199568, Q => 
                           OUT1(18), QN => n22);
   OUT1_reg_17_inst : DFF_X1 port map( D => N4524, CK => net199568, Q => 
                           OUT1(17), QN => n21);
   OUT1_reg_16_inst : DFF_X1 port map( D => N4522, CK => net199568, Q => 
                           OUT1(16), QN => n20);
   OUT1_reg_15_inst : DFF_X1 port map( D => N4520, CK => net199568, Q => 
                           OUT1(15), QN => n19);
   OUT1_reg_14_inst : DFF_X1 port map( D => N4518, CK => net199568, Q => 
                           OUT1(14), QN => n18);
   OUT1_reg_13_inst : DFF_X1 port map( D => N4516, CK => net199568, Q => 
                           OUT1(13), QN => n17);
   OUT1_reg_12_inst : DFF_X1 port map( D => N4514, CK => net199568, Q => 
                           OUT1(12), QN => n16);
   OUT1_reg_11_inst : DFF_X1 port map( D => N4512, CK => net199568, Q => 
                           OUT1(11), QN => n15);
   OUT1_reg_10_inst : DFF_X1 port map( D => N4510, CK => net199568, Q => 
                           OUT1(10), QN => n14);
   OUT1_reg_9_inst : DFF_X1 port map( D => N4508, CK => net199568, Q => OUT1(9)
                           , QN => n13);
   OUT1_reg_8_inst : DFF_X1 port map( D => N4506, CK => net199568, Q => OUT1(8)
                           , QN => n12);
   OUT1_reg_7_inst : DFF_X1 port map( D => N4504, CK => net199568, Q => OUT1(7)
                           , QN => n11);
   OUT1_reg_6_inst : DFF_X1 port map( D => N4502, CK => net199568, Q => OUT1(6)
                           , QN => n10);
   OUT1_reg_5_inst : DFF_X1 port map( D => N4500, CK => net199568, Q => OUT1(5)
                           , QN => n9);
   OUT1_reg_4_inst : DFF_X1 port map( D => N4498, CK => net199568, Q => OUT1(4)
                           , QN => n8);
   OUT1_reg_3_inst : DFF_X1 port map( D => N4496, CK => net199568, Q => OUT1(3)
                           , QN => n7);
   OUT1_reg_2_inst : DFF_X1 port map( D => N4494, CK => net199568, Q => OUT1(2)
                           , QN => n6);
   OUT1_reg_1_inst : DFF_X1 port map( D => N4492, CK => net199568, Q => OUT1(1)
                           , QN => n5);
   OUT1_reg_0_inst : DFF_X1 port map( D => N4490, CK => net199568, Q => OUT1(0)
                           , QN => n4);
   clk_gate_OUT2_reg : SNPS_CLOCK_GATE_HIGH_dlx_regfile_0 port map( CLK => Clk,
                           EN => N4615, ENCLK => net199403);
   clk_gate_REGISTERS_reg_0_inst : SNPS_CLOCK_GATE_HIGH_dlx_regfile_33 port 
                           map( CLK => Clk, EN => Rst, ENCLK => net199408);
   clk_gate_REGISTERS_reg_1_inst : SNPS_CLOCK_GATE_HIGH_dlx_regfile_32 port 
                           map( CLK => Clk, EN => N4423, ENCLK => net199413);
   clk_gate_REGISTERS_reg_2_inst : SNPS_CLOCK_GATE_HIGH_dlx_regfile_31 port 
                           map( CLK => Clk, EN => N4359, ENCLK => net199418);
   clk_gate_REGISTERS_reg_3_inst : SNPS_CLOCK_GATE_HIGH_dlx_regfile_30 port 
                           map( CLK => Clk, EN => N4295, ENCLK => net199423);
   clk_gate_REGISTERS_reg_4_inst : SNPS_CLOCK_GATE_HIGH_dlx_regfile_29 port 
                           map( CLK => Clk, EN => N4231, ENCLK => net199428);
   clk_gate_REGISTERS_reg_5_inst : SNPS_CLOCK_GATE_HIGH_dlx_regfile_28 port 
                           map( CLK => Clk, EN => N4167, ENCLK => net199433);
   clk_gate_REGISTERS_reg_6_inst : SNPS_CLOCK_GATE_HIGH_dlx_regfile_27 port 
                           map( CLK => Clk, EN => N4103, ENCLK => net199438);
   clk_gate_REGISTERS_reg_7_inst : SNPS_CLOCK_GATE_HIGH_dlx_regfile_26 port 
                           map( CLK => Clk, EN => N4039, ENCLK => net199443);
   clk_gate_REGISTERS_reg_8_inst : SNPS_CLOCK_GATE_HIGH_dlx_regfile_25 port 
                           map( CLK => Clk, EN => N3975, ENCLK => net199448);
   clk_gate_REGISTERS_reg_9_inst : SNPS_CLOCK_GATE_HIGH_dlx_regfile_24 port 
                           map( CLK => Clk, EN => N3911, ENCLK => net199453);
   clk_gate_REGISTERS_reg_10_inst : SNPS_CLOCK_GATE_HIGH_dlx_regfile_23 port 
                           map( CLK => Clk, EN => N3847, ENCLK => net199458);
   clk_gate_REGISTERS_reg_11_inst : SNPS_CLOCK_GATE_HIGH_dlx_regfile_22 port 
                           map( CLK => Clk, EN => N3783, ENCLK => net199463);
   clk_gate_REGISTERS_reg_12_inst : SNPS_CLOCK_GATE_HIGH_dlx_regfile_21 port 
                           map( CLK => Clk, EN => N3719, ENCLK => net199468);
   clk_gate_REGISTERS_reg_13_inst : SNPS_CLOCK_GATE_HIGH_dlx_regfile_20 port 
                           map( CLK => Clk, EN => N3655, ENCLK => net199473);
   clk_gate_REGISTERS_reg_14_inst : SNPS_CLOCK_GATE_HIGH_dlx_regfile_19 port 
                           map( CLK => Clk, EN => N3591, ENCLK => net199478);
   clk_gate_REGISTERS_reg_15_inst : SNPS_CLOCK_GATE_HIGH_dlx_regfile_18 port 
                           map( CLK => Clk, EN => N3527, ENCLK => net199483);
   clk_gate_REGISTERS_reg_16_inst : SNPS_CLOCK_GATE_HIGH_dlx_regfile_17 port 
                           map( CLK => Clk, EN => N3463, ENCLK => net199488);
   clk_gate_REGISTERS_reg_17_inst : SNPS_CLOCK_GATE_HIGH_dlx_regfile_16 port 
                           map( CLK => Clk, EN => N3399, ENCLK => net199493);
   clk_gate_REGISTERS_reg_18_inst : SNPS_CLOCK_GATE_HIGH_dlx_regfile_15 port 
                           map( CLK => Clk, EN => N3335, ENCLK => net199498);
   clk_gate_REGISTERS_reg_19_inst : SNPS_CLOCK_GATE_HIGH_dlx_regfile_14 port 
                           map( CLK => Clk, EN => N3271, ENCLK => net199503);
   clk_gate_REGISTERS_reg_20_inst : SNPS_CLOCK_GATE_HIGH_dlx_regfile_13 port 
                           map( CLK => Clk, EN => N3207, ENCLK => net199508);
   clk_gate_REGISTERS_reg_21_inst : SNPS_CLOCK_GATE_HIGH_dlx_regfile_12 port 
                           map( CLK => Clk, EN => N3143, ENCLK => net199513);
   clk_gate_REGISTERS_reg_22_inst : SNPS_CLOCK_GATE_HIGH_dlx_regfile_11 port 
                           map( CLK => Clk, EN => N3079, ENCLK => net199518);
   clk_gate_REGISTERS_reg_23_inst : SNPS_CLOCK_GATE_HIGH_dlx_regfile_10 port 
                           map( CLK => Clk, EN => N3015, ENCLK => net199523);
   clk_gate_REGISTERS_reg_24_inst : SNPS_CLOCK_GATE_HIGH_dlx_regfile_9 port 
                           map( CLK => Clk, EN => N2951, ENCLK => net199528);
   clk_gate_REGISTERS_reg_25_inst : SNPS_CLOCK_GATE_HIGH_dlx_regfile_8 port 
                           map( CLK => Clk, EN => N2887, ENCLK => net199533);
   clk_gate_REGISTERS_reg_26_inst : SNPS_CLOCK_GATE_HIGH_dlx_regfile_7 port 
                           map( CLK => Clk, EN => N2823, ENCLK => net199538);
   clk_gate_REGISTERS_reg_27_inst : SNPS_CLOCK_GATE_HIGH_dlx_regfile_6 port 
                           map( CLK => Clk, EN => N2759, ENCLK => net199543);
   clk_gate_REGISTERS_reg_28_inst : SNPS_CLOCK_GATE_HIGH_dlx_regfile_5 port 
                           map( CLK => Clk, EN => N2695, ENCLK => net199548);
   clk_gate_REGISTERS_reg_29_inst : SNPS_CLOCK_GATE_HIGH_dlx_regfile_4 port 
                           map( CLK => Clk, EN => N2631, ENCLK => net199553);
   clk_gate_REGISTERS_reg_30_inst : SNPS_CLOCK_GATE_HIGH_dlx_regfile_3 port 
                           map( CLK => Clk, EN => N2567, ENCLK => net199558);
   clk_gate_REGISTERS_reg_31_inst : SNPS_CLOCK_GATE_HIGH_dlx_regfile_2 port 
                           map( CLK => Clk, EN => N2503, ENCLK => net199563);
   clk_gate_OUT1_reg : SNPS_CLOCK_GATE_HIGH_dlx_regfile_1 port map( CLK => Clk,
                           EN => N4615, ENCLK => net199568);
   U3 : OR2_X1 port map( A1 => Rst, A2 => ENABLE, ZN => N4615);
   U4 : NAND2_X2 port map( A1 => n53, A2 => n1869, ZN => n1868);
   U5 : NAND2_X2 port map( A1 => n53, A2 => n1104, ZN => n1103);
   U6 : NAND3_X2 port map( A1 => n1820, A2 => n2554, A3 => n2555, ZN => n1869);
   U7 : NAND3_X2 port map( A1 => n1820, A2 => n1821, A3 => n1822, ZN => n1104);
   U8 : AND4_X1 port map( A1 => n1665, A2 => n1666, A3 => n1667, A4 => n1668, 
                           ZN => n1664);
   U9 : AND4_X1 port map( A1 => n2154, A2 => n2155, A3 => n2156, A4 => n2157, 
                           ZN => n2153);
   U10 : AND4_X1 port map( A1 => n1489, A2 => n1490, A3 => n1491, A4 => n1492, 
                           ZN => n1488);
   U11 : AND4_X1 port map( A1 => n1291, A2 => n1292, A3 => n1293, A4 => n1294, 
                           ZN => n1290);
   U12 : AND4_X1 port map( A1 => n2175, A2 => n2176, A3 => n2177, A4 => n2178, 
                           ZN => n2174);
   U13 : AND4_X1 port map( A1 => n2469, A2 => n2470, A3 => n2471, A4 => n2472, 
                           ZN => n2468);
   U14 : AND4_X1 port map( A1 => n1643, A2 => n1644, A3 => n1645, A4 => n1646, 
                           ZN => n1642);
   U15 : AND4_X1 port map( A1 => n2091, A2 => n2092, A3 => n2093, A4 => n2094, 
                           ZN => n2090);
   U16 : AND4_X1 port map( A1 => n1687, A2 => n1688, A3 => n1689, A4 => n1690, 
                           ZN => n1686);
   U17 : AND4_X1 port map( A1 => n2112, A2 => n2113, A3 => n2114, A4 => n2115, 
                           ZN => n2111);
   U18 : AND4_X1 port map( A1 => n2133, A2 => n2134, A3 => n2135, A4 => n2136, 
                           ZN => n2132);
   U19 : AND4_X1 port map( A1 => n2280, A2 => n2281, A3 => n2282, A4 => n2283, 
                           ZN => n2279);
   U20 : AND4_X1 port map( A1 => n1335, A2 => n1336, A3 => n1337, A4 => n1338, 
                           ZN => n1334);
   U21 : AND4_X1 port map( A1 => n1599, A2 => n1600, A3 => n1601, A4 => n1602, 
                           ZN => n1598);
   U22 : AND4_X1 port map( A1 => n2427, A2 => n2428, A3 => n2429, A4 => n2430, 
                           ZN => n2426);
   U23 : AND4_X1 port map( A1 => n2301, A2 => n2302, A3 => n2303, A4 => n2304, 
                           ZN => n2300);
   U24 : AND4_X1 port map( A1 => n2322, A2 => n2323, A3 => n2324, A4 => n2325, 
                           ZN => n2321);
   U25 : AND4_X1 port map( A1 => n1577, A2 => n1578, A3 => n1579, A4 => n1580, 
                           ZN => n1576);
   U26 : AND4_X1 port map( A1 => n2343, A2 => n2344, A3 => n2345, A4 => n2346, 
                           ZN => n2342);
   U27 : AND4_X1 port map( A1 => n2364, A2 => n2365, A3 => n2366, A4 => n2367, 
                           ZN => n2363);
   U28 : AND4_X1 port map( A1 => n1555, A2 => n1556, A3 => n1557, A4 => n1558, 
                           ZN => n1554);
   U29 : AND4_X1 port map( A1 => n2406, A2 => n2407, A3 => n2408, A4 => n2409, 
                           ZN => n2405);
   U30 : AND4_X1 port map( A1 => n2385, A2 => n2386, A3 => n2387, A4 => n2388, 
                           ZN => n2384);
   U31 : AND4_X1 port map( A1 => n1533, A2 => n1534, A3 => n1535, A4 => n1536, 
                           ZN => n1532);
   U32 : AND4_X1 port map( A1 => n2196, A2 => n2197, A3 => n2198, A4 => n2199, 
                           ZN => n2195);
   U33 : AND4_X1 port map( A1 => n2217, A2 => n2218, A3 => n2219, A4 => n2220, 
                           ZN => n2216);
   U34 : AND4_X1 port map( A1 => n1313, A2 => n1314, A3 => n1315, A4 => n1316, 
                           ZN => n1312);
   U35 : AND4_X1 port map( A1 => n2448, A2 => n2449, A3 => n2450, A4 => n2451, 
                           ZN => n2447);
   U36 : AND4_X1 port map( A1 => n1621, A2 => n1622, A3 => n1623, A4 => n1624, 
                           ZN => n1620);
   U37 : AND4_X1 port map( A1 => n2238, A2 => n2239, A3 => n2240, A4 => n2241, 
                           ZN => n2237);
   U38 : AND4_X1 port map( A1 => n1379, A2 => n1380, A3 => n1381, A4 => n1382, 
                           ZN => n1378);
   U39 : AND4_X1 port map( A1 => n1511, A2 => n1512, A3 => n1513, A4 => n1514, 
                           ZN => n1510);
   U40 : AND4_X1 port map( A1 => n2259, A2 => n2260, A3 => n2261, A4 => n2262, 
                           ZN => n2258);
   U41 : AND4_X1 port map( A1 => n1776, A2 => n1777, A3 => n1778, A4 => n1779, 
                           ZN => n1775);
   U42 : AND4_X1 port map( A1 => n1965, A2 => n1966, A3 => n1967, A4 => n1968, 
                           ZN => n1964);
   U43 : AND4_X1 port map( A1 => n1423, A2 => n1424, A3 => n1425, A4 => n1426, 
                           ZN => n1422);
   U44 : AND4_X1 port map( A1 => n1247, A2 => n1248, A3 => n1249, A4 => n1250, 
                           ZN => n1246);
   U45 : AND4_X1 port map( A1 => n1986, A2 => n1987, A3 => n1988, A4 => n1989, 
                           ZN => n1985);
   U46 : AND4_X1 port map( A1 => n2565, A2 => n2566, A3 => n2567_port, A4 => 
                           n2568, ZN => n2553);
   U47 : AND4_X1 port map( A1 => n2007, A2 => n2008, A3 => n2009, A4 => n2010, 
                           ZN => n2006);
   U48 : AND4_X1 port map( A1 => n1181, A2 => n1182, A3 => n1183, A4 => n1184, 
                           ZN => n1180);
   U49 : AND4_X1 port map( A1 => n1832, A2 => n1833, A3 => n1834, A4 => n1835, 
                           ZN => n1819);
   U50 : AND4_X1 port map( A1 => n1159, A2 => n1160, A3 => n1161, A4 => n1162, 
                           ZN => n1158);
   U51 : AND4_X1 port map( A1 => n1870, A2 => n1871, A3 => n1872, A4 => n1873, 
                           ZN => n1867);
   U52 : AND4_X1 port map( A1 => n1203, A2 => n1204, A3 => n1205, A4 => n1206, 
                           ZN => n1202);
   U53 : AND4_X1 port map( A1 => n1798, A2 => n1799, A3 => n1800, A4 => n1801, 
                           ZN => n1797);
   U54 : AND4_X1 port map( A1 => n1923, A2 => n1924, A3 => n1925, A4 => n1926, 
                           ZN => n1922);
   U55 : AND4_X1 port map( A1 => n1401, A2 => n1402, A3 => n1403, A4 => n1404, 
                           ZN => n1400);
   U56 : AND4_X1 port map( A1 => n1105, A2 => n1106, A3 => n1107, A4 => n1108, 
                           ZN => n1102);
   U57 : AND4_X1 port map( A1 => n1944, A2 => n1945, A3 => n1946, A4 => n1947, 
                           ZN => n1943);
   U58 : AND4_X1 port map( A1 => n1225, A2 => n1226, A3 => n1227, A4 => n1228, 
                           ZN => n1224);
   U59 : AND4_X1 port map( A1 => n1357, A2 => n1358, A3 => n1359, A4 => n1360, 
                           ZN => n1356);
   U60 : AND4_X1 port map( A1 => n1269, A2 => n1270, A3 => n1271, A4 => n1272, 
                           ZN => n1268);
   U61 : AND4_X1 port map( A1 => n2070, A2 => n2071, A3 => n2072, A4 => n2073, 
                           ZN => n2069);
   U62 : AND4_X1 port map( A1 => n2049, A2 => n2050, A3 => n2051, A4 => n2052, 
                           ZN => n2048);
   U63 : AND4_X1 port map( A1 => n1731, A2 => n1732, A3 => n1733, A4 => n1734, 
                           ZN => n1730);
   U64 : AND4_X1 port map( A1 => n1467, A2 => n1468, A3 => n1469, A4 => n1470, 
                           ZN => n1466);
   U65 : AND4_X1 port map( A1 => n2533, A2 => n2534, A3 => n2535, A4 => n2536, 
                           ZN => n2532);
   U66 : AND4_X1 port map( A1 => n1709, A2 => n1710, A3 => n1711, A4 => n1712, 
                           ZN => n1708);
   U67 : AND4_X1 port map( A1 => n2028, A2 => n2029, A3 => n2030, A4 => n2031, 
                           ZN => n2027);
   U68 : AND4_X1 port map( A1 => n2512, A2 => n2513, A3 => n2514, A4 => n2515, 
                           ZN => n2511);
   U69 : AND4_X1 port map( A1 => n1445, A2 => n1446, A3 => n1447, A4 => n1448, 
                           ZN => n1444);
   U70 : INV_X1 port map( A => n2564, ZN => n2561);
   U71 : INV_X1 port map( A => n1774, ZN => n1768);
   U72 : INV_X1 port map( A => n2510, ZN => n2504);
   U73 : OR3_X1 port map( A1 => n1830, A2 => n2563, A3 => ADD_WR(4), ZN => 
                           n2608);
   U74 : INV_X1 port map( A => ADD_WR(3), ZN => n1830);
   U75 : NAND2_X2 port map( A1 => DATAIN(1), A2 => n53, ZN => n1788);
   U76 : NAND2_X2 port map( A1 => DATAIN(2), A2 => n53, ZN => n1766);
   U77 : NAND2_X2 port map( A1 => DATAIN(3), A2 => n51, ZN => n1744);
   U78 : NAND2_X2 port map( A1 => DATAIN(4), A2 => n51, ZN => n1722);
   U79 : NAND2_X2 port map( A1 => DATAIN(5), A2 => n51, ZN => n1700);
   U80 : NAND2_X2 port map( A1 => DATAIN(6), A2 => n51, ZN => n1678);
   U81 : NAND2_X2 port map( A1 => DATAIN(7), A2 => n51, ZN => n1656);
   U82 : NAND2_X2 port map( A1 => DATAIN(8), A2 => n51, ZN => n1634);
   U83 : NAND2_X2 port map( A1 => DATAIN(0), A2 => n53, ZN => n1810);
   U84 : NAND2_X2 port map( A1 => DATAIN(9), A2 => n51, ZN => n1612);
   U85 : NAND2_X2 port map( A1 => DATAIN(10), A2 => n51, ZN => n1590);
   U86 : NAND2_X2 port map( A1 => DATAIN(11), A2 => n51, ZN => n1568);
   U87 : NAND2_X2 port map( A1 => DATAIN(12), A2 => n51, ZN => n1546);
   U88 : INV_X1 port map( A => ADD_WR(1), ZN => n1824);
   U89 : NAND2_X2 port map( A1 => DATAIN(25), A2 => n49, ZN => n1260);
   U90 : NAND2_X2 port map( A1 => DATAIN(26), A2 => n49, ZN => n1238);
   U91 : NAND2_X2 port map( A1 => DATAIN(27), A2 => n47, ZN => n1216);
   U92 : NAND2_X2 port map( A1 => DATAIN(28), A2 => n47, ZN => n1194);
   U93 : NAND2_X2 port map( A1 => DATAIN(29), A2 => n47, ZN => n1172);
   U94 : NAND2_X2 port map( A1 => DATAIN(30), A2 => n47, ZN => n1150);
   U95 : NAND2_X2 port map( A1 => DATAIN(31), A2 => n47, ZN => n1094);
   U96 : NAND2_X2 port map( A1 => DATAIN(13), A2 => n51, ZN => n1524);
   U97 : NAND2_X2 port map( A1 => DATAIN(14), A2 => n51, ZN => n1502);
   U98 : NAND2_X2 port map( A1 => DATAIN(15), A2 => n49, ZN => n1480);
   U99 : NAND2_X2 port map( A1 => DATAIN(16), A2 => n49, ZN => n1458);
   U100 : NAND2_X2 port map( A1 => DATAIN(17), A2 => n49, ZN => n1436);
   U101 : NAND2_X2 port map( A1 => DATAIN(18), A2 => n49, ZN => n1414);
   U102 : NAND2_X2 port map( A1 => DATAIN(19), A2 => n49, ZN => n1392);
   U103 : NAND2_X2 port map( A1 => DATAIN(20), A2 => n49, ZN => n1370);
   U104 : NAND2_X2 port map( A1 => DATAIN(21), A2 => n49, ZN => n1348);
   U105 : NAND2_X2 port map( A1 => DATAIN(22), A2 => n49, ZN => n1326);
   U106 : NAND2_X2 port map( A1 => DATAIN(23), A2 => n49, ZN => n1304);
   U107 : NAND2_X2 port map( A1 => DATAIN(24), A2 => n49, ZN => n1282);
   U108 : INV_X1 port map( A => ADD_WR(2), ZN => n1826);
   U109 : INV_X1 port map( A => ADD_WR(0), ZN => n1827);
   U110 : NAND2_X2 port map( A1 => n2573, A2 => n2575, ZN => n1878);
   U111 : NAND2_X2 port map( A1 => n2576, A2 => n2574, ZN => n1881);
   U112 : NAND2_X2 port map( A1 => n2576, A2 => n2575, ZN => n1880);
   U113 : NAND2_X2 port map( A1 => n2573, A2 => n2586, ZN => n1891);
   U114 : NAND2_X2 port map( A1 => n2573, A2 => n2574, ZN => n1879);
   U115 : NAND2_X2 port map( A1 => n2573, A2 => n2587, ZN => n1890);
   U116 : NAND2_X2 port map( A1 => n2586, A2 => n2576, ZN => n1893);
   U117 : NAND2_X2 port map( A1 => n2587, A2 => n2576, ZN => n1892);
   U118 : NAND2_X2 port map( A1 => n2577, A2 => n2586, ZN => n1895);
   U119 : NAND2_X2 port map( A1 => n2577, A2 => n2587, ZN => n1894);
   U120 : NAND2_X2 port map( A1 => n2578, A2 => n2586, ZN => n1897);
   U121 : NAND2_X2 port map( A1 => n2578, A2 => n2587, ZN => n1896);
   U122 : NAND2_X2 port map( A1 => n2573, A2 => n2592, ZN => n1903);
   U123 : NAND2_X2 port map( A1 => n2573, A2 => n2593, ZN => n1902);
   U124 : NAND2_X2 port map( A1 => n2592, A2 => n2576, ZN => n1905);
   U125 : NAND2_X2 port map( A1 => n2576, A2 => n2593, ZN => n1904);
   U126 : NAND2_X2 port map( A1 => n2577, A2 => n2592, ZN => n1907);
   U127 : NAND2_X2 port map( A1 => n2577, A2 => n2593, ZN => n1906);
   U128 : NAND2_X2 port map( A1 => n2592, A2 => n2578, ZN => n1909);
   U129 : NAND2_X2 port map( A1 => n2578, A2 => n2593, ZN => n1908);
   U130 : NAND2_X2 port map( A1 => n2573, A2 => n2598, ZN => n1915);
   U131 : NAND2_X2 port map( A1 => n2576, A2 => n2598, ZN => n1917);
   U132 : NAND2_X2 port map( A1 => n2599, A2 => n2576, ZN => n1916);
   U133 : NAND2_X2 port map( A1 => n2577, A2 => n2598, ZN => n1919);
   U134 : NAND2_X2 port map( A1 => n2599, A2 => n2577, ZN => n1918);
   U135 : NAND2_X2 port map( A1 => n2578, A2 => n2598, ZN => n1921);
   U136 : NAND2_X2 port map( A1 => n1843, A2 => n1860, ZN => n1139);
   U137 : NAND2_X2 port map( A1 => n1859, A2 => n1843, ZN => n1140);
   U138 : NAND2_X2 port map( A1 => n1840, A2 => n1860, ZN => n1137);
   U139 : NAND2_X2 port map( A1 => n1840, A2 => n1859, ZN => n1138);
   U140 : NAND2_X2 port map( A1 => n1845, A2 => n1854, ZN => n1131);
   U141 : NAND2_X2 port map( A1 => n1845, A2 => n1853, ZN => n1132);
   U142 : NAND2_X2 port map( A1 => n1844, A2 => n1854, ZN => n1129);
   U143 : NAND2_X2 port map( A1 => n1844, A2 => n1853, ZN => n1130);
   U144 : NAND2_X2 port map( A1 => n1854, A2 => n1843, ZN => n1127);
   U145 : NAND2_X2 port map( A1 => n1853, A2 => n1843, ZN => n1128);
   U146 : NAND2_X2 port map( A1 => n1840, A2 => n1854, ZN => n1125);
   U147 : NAND2_X2 port map( A1 => n1840, A2 => n1853, ZN => n1126);
   U148 : NAND2_X2 port map( A1 => n1845, A2 => n1842, ZN => n1119);
   U149 : NAND2_X2 port map( A1 => n1845, A2 => n1841, ZN => n1120);
   U150 : NAND2_X2 port map( A1 => n1844, A2 => n1842, ZN => n1117);
   U151 : NAND2_X2 port map( A1 => n1844, A2 => n1841, ZN => n1118);
   U152 : NAND2_X2 port map( A1 => n1843, A2 => n1842, ZN => n1115);
   U153 : NAND2_X2 port map( A1 => n1843, A2 => n1841, ZN => n1116);
   U154 : NAND2_X2 port map( A1 => n1840, A2 => n1842, ZN => n1113);
   U155 : NAND2_X2 port map( A1 => n1840, A2 => n1841, ZN => n1114);
   U156 : NAND2_X2 port map( A1 => n1845, A2 => n1865, ZN => n1157);
   U157 : NAND2_X2 port map( A1 => n1866, A2 => n1844, ZN => n1154);
   U158 : NAND2_X2 port map( A1 => n1844, A2 => n1865, ZN => n1155);
   U159 : NAND2_X2 port map( A1 => n1866, A2 => n1843, ZN => n1152);
   U160 : NAND2_X2 port map( A1 => n1843, A2 => n1865, ZN => n1153);
   U161 : NAND2_X2 port map( A1 => n1840, A2 => n1865, ZN => n1151);
   U162 : AND2_X1 port map( A1 => n1823, A2 => ADD_RD2(2), ZN => n1843);
   U163 : NAND2_X2 port map( A1 => n2599, A2 => n2578, ZN => n1920);
   U164 : NAND2_X2 port map( A1 => n2599, A2 => n2573, ZN => n1914);
   U165 : NAND2_X2 port map( A1 => n1866, A2 => n1845, ZN => n1156);
   U166 : AND2_X1 port map( A1 => n2556, A2 => ADD_RD1(2), ZN => n2576);
   U167 : NAND2_X2 port map( A1 => n1866, A2 => n1840, ZN => n1149);
   U168 : INV_X1 port map( A => ADD_RD1(1), ZN => n2556);
   U169 : INV_X1 port map( A => ADD_RD1(4), ZN => n2559);
   U170 : INV_X1 port map( A => ADD_RD1(0), ZN => n2580);
   U171 : INV_X1 port map( A => ADD_RD1(3), ZN => n2579);
   U172 : AND2_X1 port map( A1 => ADD_RD1(1), A2 => ADD_RD1(2), ZN => n2573);
   U173 : AND2_X1 port map( A1 => ADD_RD2(1), A2 => ADD_RD2(2), ZN => n1840);
   U174 : INV_X1 port map( A => ADD_RD2(3), ZN => n1846);
   U175 : INV_X1 port map( A => ADD_RD2(0), ZN => n1847);
   U176 : INV_X1 port map( A => ADD_RD2(4), ZN => n1829);
   U177 : INV_X1 port map( A => Rst, ZN => n53);
   U178 : INV_X1 port map( A => ADD_RD2(1), ZN => n1823);
   U179 : INV_X1 port map( A => Rst, ZN => n51);
   U180 : INV_X1 port map( A => Rst, ZN => n49);
   U181 : INV_X1 port map( A => Rst, ZN => n47);
   U182 : NOR2_X1 port map( A1 => ADD_RD2(2), A2 => n1823, ZN => n1844);
   U183 : AOI21_X1 port map( B1 => n2561, B2 => n2562, A => n2563, ZN => n1820)
                           ;
   U184 : NOR2_X1 port map( A1 => ADD_RD1(2), A2 => n2556, ZN => n2577);
   U185 : NOR2_X1 port map( A1 => ADD_RD2(1), A2 => ADD_RD2(2), ZN => n1845);
   U186 : NOR2_X1 port map( A1 => ADD_RD1(1), A2 => ADD_RD1(2), ZN => n2578);
   U187 : NOR2_X1 port map( A1 => ADD_WR(4), A2 => ADD_WR(3), ZN => n2562);
   U188 : AOI221_X1 port map( B1 => ADD_WR(1), B2 => n1823, C1 => n1824, C2 => 
                           ADD_RD2(1), A => n1825, ZN => n1822);
   U189 : NOR2_X1 port map( A1 => ADD_RD2(0), A2 => n1848, ZN => n1842);
   U190 : AOI221_X1 port map( B1 => ADD_WR(1), B2 => n2556, C1 => n1824, C2 => 
                           ADD_RD1(1), A => n2557, ZN => n2555);
   U191 : NOR2_X1 port map( A1 => ADD_RD1(0), A2 => n2581, ZN => n2575);
   U192 : NAND2_X1 port map( A1 => n2577, A2 => n2575, ZN => n1882);
   U193 : NAND2_X1 port map( A1 => n2578, A2 => n2575, ZN => n1884);
   U194 : NAND3_X1 port map( A1 => n1827, A2 => n1826, A3 => n1824, ZN => n2564
                           );
   U195 : BUF_X1 port map( A => n1142, Z => n2);
   U196 : BUF_X1 port map( A => n1141, Z => n1);
   U197 : BUF_X1 port map( A => n1144, Z => n37);
   U198 : BUF_X1 port map( A => n1143, Z => n3);
   U199 : BUF_X1 port map( A => n1883, Z => n41);
   U200 : BUF_X1 port map( A => n1882, Z => n39);
   U201 : BUF_X1 port map( A => n1885, Z => n45);
   U202 : BUF_X1 port map( A => n1884, Z => n43);
   U203 : OAI22_X1 port map( A1 => n1102, A2 => n1103, B1 => n1104, B2 => n1094
                           , ZN => N4616);
   U204 : NOR4_X1 port map( A1 => n1109, A2 => n1110, A3 => n1111, A4 => n1112,
                           ZN => n1108);
   U205 : OAI22_X1 port map( A1 => n200, A2 => n1113, B1 => n1090, B2 => n1114,
                           ZN => n1112);
   U206 : OAI22_X1 port map( A1 => n264, A2 => n1115, B1 => n232, B2 => n1116, 
                           ZN => n1111);
   U207 : OAI22_X1 port map( A1 => n328, A2 => n1117, B1 => n296, B2 => n1118, 
                           ZN => n1110);
   U208 : OAI22_X1 port map( A1 => n392, A2 => n1119, B1 => n360, B2 => n1120, 
                           ZN => n1109);
   U209 : NOR4_X1 port map( A1 => n1121, A2 => n1122, A3 => n1123, A4 => n1124,
                           ZN => n1107);
   U210 : OAI22_X1 port map( A1 => n457, A2 => n1125, B1 => n424, B2 => n1126, 
                           ZN => n1124);
   U211 : OAI22_X1 port map( A1 => n525, A2 => n1127, B1 => n491, B2 => n1128, 
                           ZN => n1123);
   U212 : OAI22_X1 port map( A1 => n592, A2 => n1129, B1 => n558, B2 => n1130, 
                           ZN => n1122);
   U213 : OAI22_X1 port map( A1 => n659, A2 => n1131, B1 => n625, B2 => n1132, 
                           ZN => n1121);
   U214 : NOR4_X1 port map( A1 => n1133, A2 => n1134, A3 => n1135, A4 => n1136,
                           ZN => n1106);
   U215 : OAI22_X1 port map( A1 => n726, A2 => n1137, B1 => n693, B2 => n1138, 
                           ZN => n1136);
   U216 : OAI22_X1 port map( A1 => n793, A2 => n1139, B1 => n760, B2 => n1140, 
                           ZN => n1135);
   U217 : OAI22_X1 port map( A1 => n861, A2 => n1141, B1 => n827, B2 => n1142, 
                           ZN => n1134);
   U218 : OAI22_X1 port map( A1 => n928, A2 => n1143, B1 => n894, B2 => n1144, 
                           ZN => n1133);
   U219 : NOR4_X1 port map( A1 => n1145, A2 => n1146, A3 => n1147, A4 => n1148,
                           ZN => n1105);
   U220 : OAI22_X1 port map( A1 => n995, A2 => n1149, B1 => n961, B2 => n1151, 
                           ZN => n1148);
   U221 : OAI22_X1 port map( A1 => n1062, A2 => n1152, B1 => n1029, B2 => n1153
                           , ZN => n1147);
   U222 : OAI22_X1 port map( A1 => n107, A2 => n1154, B1 => n1097, B2 => n1155,
                           ZN => n1146);
   U223 : OAI22_X1 port map( A1 => n178, A2 => n1156, B1 => n142, B2 => n1157, 
                           ZN => n1145);
   U224 : OAI22_X1 port map( A1 => n1158, A2 => n1103, B1 => n1104, B2 => n1150
                           , ZN => N4614);
   U225 : NOR4_X1 port map( A1 => n1163, A2 => n1164, A3 => n1165, A4 => n1166,
                           ZN => n1162);
   U226 : OAI22_X1 port map( A1 => n199, A2 => n1113, B1 => n1069, B2 => n1114,
                           ZN => n1166);
   U227 : OAI22_X1 port map( A1 => n263, A2 => n1115, B1 => n231, B2 => n1116, 
                           ZN => n1165);
   U228 : OAI22_X1 port map( A1 => n327, A2 => n1117, B1 => n295, B2 => n1118, 
                           ZN => n1164);
   U229 : OAI22_X1 port map( A1 => n391, A2 => n1119, B1 => n359, B2 => n1120, 
                           ZN => n1163);
   U230 : NOR4_X1 port map( A1 => n1167, A2 => n1168, A3 => n1169, A4 => n1170,
                           ZN => n1161);
   U231 : OAI22_X1 port map( A1 => n456, A2 => n1125, B1 => n423, B2 => n1126, 
                           ZN => n1170);
   U232 : OAI22_X1 port map( A1 => n524, A2 => n1127, B1 => n490, B2 => n1128, 
                           ZN => n1169);
   U233 : OAI22_X1 port map( A1 => n591, A2 => n1129, B1 => n557, B2 => n1130, 
                           ZN => n1168);
   U234 : OAI22_X1 port map( A1 => n658, A2 => n1131, B1 => n624, B2 => n1132, 
                           ZN => n1167);
   U235 : NOR4_X1 port map( A1 => n1171, A2 => n1173, A3 => n1174, A4 => n1175,
                           ZN => n1160);
   U236 : OAI22_X1 port map( A1 => n725, A2 => n1137, B1 => n692, B2 => n1138, 
                           ZN => n1175);
   U237 : OAI22_X1 port map( A1 => n792, A2 => n1139, B1 => n759, B2 => n1140, 
                           ZN => n1174);
   U238 : OAI22_X1 port map( A1 => n860, A2 => n1, B1 => n826, B2 => n1142, ZN 
                           => n1173);
   U239 : OAI22_X1 port map( A1 => n927, A2 => n3, B1 => n893, B2 => n1144, ZN 
                           => n1171);
   U240 : NOR4_X1 port map( A1 => n1176, A2 => n1177, A3 => n1178, A4 => n1179,
                           ZN => n1159);
   U241 : OAI22_X1 port map( A1 => n994, A2 => n1149, B1 => n960, B2 => n1151, 
                           ZN => n1179);
   U242 : OAI22_X1 port map( A1 => n1061, A2 => n1152, B1 => n1028, B2 => n1153
                           , ZN => n1178);
   U243 : OAI22_X1 port map( A1 => n106, A2 => n1154, B1 => n1096, B2 => n1155,
                           ZN => n1177);
   U244 : OAI22_X1 port map( A1 => n177, A2 => n1156, B1 => n141, B2 => n1157, 
                           ZN => n1176);
   U245 : OAI22_X1 port map( A1 => n1180, A2 => n1103, B1 => n1104, B2 => n1172
                           , ZN => N4612);
   U246 : NOR4_X1 port map( A1 => n1185, A2 => n1186, A3 => n1187, A4 => n1188,
                           ZN => n1184);
   U247 : OAI22_X1 port map( A1 => n198, A2 => n1113, B1 => n1048, B2 => n1114,
                           ZN => n1188);
   U248 : OAI22_X1 port map( A1 => n262, A2 => n1115, B1 => n230, B2 => n1116, 
                           ZN => n1187);
   U249 : OAI22_X1 port map( A1 => n326, A2 => n1117, B1 => n294, B2 => n1118, 
                           ZN => n1186);
   U250 : OAI22_X1 port map( A1 => n390, A2 => n1119, B1 => n358, B2 => n1120, 
                           ZN => n1185);
   U251 : NOR4_X1 port map( A1 => n1189, A2 => n1190, A3 => n1191, A4 => n1192,
                           ZN => n1183);
   U252 : OAI22_X1 port map( A1 => n455, A2 => n1125, B1 => n422, B2 => n1126, 
                           ZN => n1192);
   U253 : OAI22_X1 port map( A1 => n522, A2 => n1127, B1 => n489, B2 => n1128, 
                           ZN => n1191);
   U254 : OAI22_X1 port map( A1 => n590, A2 => n1129, B1 => n556, B2 => n1130, 
                           ZN => n1190);
   U255 : OAI22_X1 port map( A1 => n657, A2 => n1131, B1 => n623, B2 => n1132, 
                           ZN => n1189);
   U256 : NOR4_X1 port map( A1 => n1193, A2 => n1195, A3 => n1196, A4 => n1197,
                           ZN => n1182);
   U257 : OAI22_X1 port map( A1 => n724, A2 => n1137, B1 => n690, B2 => n1138, 
                           ZN => n1197);
   U258 : OAI22_X1 port map( A1 => n791, A2 => n1139, B1 => n758, B2 => n1140, 
                           ZN => n1196);
   U259 : OAI22_X1 port map( A1 => n858, A2 => n1141, B1 => n825, B2 => n1142, 
                           ZN => n1195);
   U260 : OAI22_X1 port map( A1 => n926, A2 => n1143, B1 => n892, B2 => n1144, 
                           ZN => n1193);
   U261 : NOR4_X1 port map( A1 => n1198, A2 => n1199, A3 => n1200, A4 => n1201,
                           ZN => n1181);
   U262 : OAI22_X1 port map( A1 => n993, A2 => n1149, B1 => n959, B2 => n1151, 
                           ZN => n1201);
   U263 : OAI22_X1 port map( A1 => n1060, A2 => n1152, B1 => n1026, B2 => n1153
                           , ZN => n1200);
   U264 : OAI22_X1 port map( A1 => n105, A2 => n1154, B1 => n1095, B2 => n1155,
                           ZN => n1199);
   U265 : OAI22_X1 port map( A1 => n175, A2 => n1156, B1 => n140, B2 => n1157, 
                           ZN => n1198);
   U266 : OAI22_X1 port map( A1 => n1202, A2 => n1103, B1 => n1104, B2 => n1194
                           , ZN => N4610);
   U267 : NOR4_X1 port map( A1 => n1207, A2 => n1208, A3 => n1209, A4 => n1210,
                           ZN => n1206);
   U268 : OAI22_X1 port map( A1 => n197, A2 => n1113, B1 => n1027, B2 => n1114,
                           ZN => n1210);
   U269 : OAI22_X1 port map( A1 => n261, A2 => n1115, B1 => n229, B2 => n1116, 
                           ZN => n1209);
   U270 : OAI22_X1 port map( A1 => n325, A2 => n1117, B1 => n293, B2 => n1118, 
                           ZN => n1208);
   U271 : OAI22_X1 port map( A1 => n389, A2 => n1119, B1 => n357, B2 => n1120, 
                           ZN => n1207);
   U272 : NOR4_X1 port map( A1 => n1211, A2 => n1212, A3 => n1213, A4 => n1214,
                           ZN => n1205);
   U273 : OAI22_X1 port map( A1 => n454, A2 => n1125, B1 => n421, B2 => n1126, 
                           ZN => n1214);
   U274 : OAI22_X1 port map( A1 => n521, A2 => n1127, B1 => n488, B2 => n1128, 
                           ZN => n1213);
   U275 : OAI22_X1 port map( A1 => n589, A2 => n1129, B1 => n555, B2 => n1130, 
                           ZN => n1212);
   U276 : OAI22_X1 port map( A1 => n656, A2 => n1131, B1 => n622, B2 => n1132, 
                           ZN => n1211);
   U277 : NOR4_X1 port map( A1 => n1215, A2 => n1217, A3 => n1218, A4 => n1219,
                           ZN => n1204);
   U278 : OAI22_X1 port map( A1 => n723, A2 => n1137, B1 => n689, B2 => n1138, 
                           ZN => n1219);
   U279 : OAI22_X1 port map( A1 => n790, A2 => n1139, B1 => n757, B2 => n1140, 
                           ZN => n1218);
   U280 : OAI22_X1 port map( A1 => n857, A2 => n1141, B1 => n824, B2 => n1142, 
                           ZN => n1217);
   U281 : OAI22_X1 port map( A1 => n925, A2 => n1143, B1 => n891, B2 => n1144, 
                           ZN => n1215);
   U282 : NOR4_X1 port map( A1 => n1220, A2 => n1221, A3 => n1222, A4 => n1223,
                           ZN => n1203);
   U283 : OAI22_X1 port map( A1 => n992, A2 => n1149, B1 => n958, B2 => n1151, 
                           ZN => n1223);
   U284 : OAI22_X1 port map( A1 => n1059, A2 => n1152, B1 => n1025, B2 => n1153
                           , ZN => n1222);
   U285 : OAI22_X1 port map( A1 => n104, A2 => n1154, B1 => n1093, B2 => n1155,
                           ZN => n1221);
   U286 : OAI22_X1 port map( A1 => n174, A2 => n1156, B1 => n139, B2 => n1157, 
                           ZN => n1220);
   U287 : OAI22_X1 port map( A1 => n1224, A2 => n1103, B1 => n1104, B2 => n1216
                           , ZN => N4608);
   U288 : NOR4_X1 port map( A1 => n1229, A2 => n1230, A3 => n1231, A4 => n1232,
                           ZN => n1228);
   U289 : OAI22_X1 port map( A1 => n196, A2 => n1113, B1 => n1006, B2 => n1114,
                           ZN => n1232);
   U290 : OAI22_X1 port map( A1 => n260, A2 => n1115, B1 => n228, B2 => n1116, 
                           ZN => n1231);
   U291 : OAI22_X1 port map( A1 => n324, A2 => n1117, B1 => n292, B2 => n1118, 
                           ZN => n1230);
   U292 : OAI22_X1 port map( A1 => n388, A2 => n1119, B1 => n356, B2 => n1120, 
                           ZN => n1229);
   U293 : NOR4_X1 port map( A1 => n1233, A2 => n1234, A3 => n1235, A4 => n1236,
                           ZN => n1227);
   U294 : OAI22_X1 port map( A1 => n453, A2 => n1125, B1 => n420, B2 => n1126, 
                           ZN => n1236);
   U295 : OAI22_X1 port map( A1 => n520, A2 => n1127, B1 => n487, B2 => n1128, 
                           ZN => n1235);
   U296 : OAI22_X1 port map( A1 => n588, A2 => n1129, B1 => n554, B2 => n1130, 
                           ZN => n1234);
   U297 : OAI22_X1 port map( A1 => n655, A2 => n1131, B1 => n621, B2 => n1132, 
                           ZN => n1233);
   U298 : NOR4_X1 port map( A1 => n1237, A2 => n1239, A3 => n1240, A4 => n1241,
                           ZN => n1226);
   U299 : OAI22_X1 port map( A1 => n722, A2 => n1137, B1 => n688, B2 => n1138, 
                           ZN => n1241);
   U300 : OAI22_X1 port map( A1 => n789, A2 => n1139, B1 => n756, B2 => n1140, 
                           ZN => n1240);
   U301 : OAI22_X1 port map( A1 => n856, A2 => n1141, B1 => n823, B2 => n1142, 
                           ZN => n1239);
   U302 : OAI22_X1 port map( A1 => n924, A2 => n1143, B1 => n890, B2 => n1144, 
                           ZN => n1237);
   U303 : NOR4_X1 port map( A1 => n1242, A2 => n1243, A3 => n1244, A4 => n1245,
                           ZN => n1225);
   U304 : OAI22_X1 port map( A1 => n991, A2 => n1149, B1 => n957, B2 => n1151, 
                           ZN => n1245);
   U305 : OAI22_X1 port map( A1 => n1058, A2 => n1152, B1 => n1024, B2 => n1153
                           , ZN => n1244);
   U306 : OAI22_X1 port map( A1 => n103, A2 => n1154, B1 => n1092, B2 => n1155,
                           ZN => n1243);
   U307 : OAI22_X1 port map( A1 => n173, A2 => n1156, B1 => n138, B2 => n1157, 
                           ZN => n1242);
   U308 : OAI22_X1 port map( A1 => n1246, A2 => n1103, B1 => n1104, B2 => n1238
                           , ZN => N4606);
   U309 : NOR4_X1 port map( A1 => n1251, A2 => n1252, A3 => n1253, A4 => n1254,
                           ZN => n1250);
   U310 : OAI22_X1 port map( A1 => n195, A2 => n1113, B1 => n985, B2 => n1114, 
                           ZN => n1254);
   U311 : OAI22_X1 port map( A1 => n259, A2 => n1115, B1 => n227, B2 => n1116, 
                           ZN => n1253);
   U312 : OAI22_X1 port map( A1 => n323, A2 => n1117, B1 => n291, B2 => n1118, 
                           ZN => n1252);
   U313 : OAI22_X1 port map( A1 => n387, A2 => n1119, B1 => n355, B2 => n1120, 
                           ZN => n1251);
   U314 : NOR4_X1 port map( A1 => n1255, A2 => n1256, A3 => n1257, A4 => n1258,
                           ZN => n1249);
   U315 : OAI22_X1 port map( A1 => n452, A2 => n1125, B1 => n419, B2 => n1126, 
                           ZN => n1258);
   U316 : OAI22_X1 port map( A1 => n519, A2 => n1127, B1 => n486, B2 => n1128, 
                           ZN => n1257);
   U317 : OAI22_X1 port map( A1 => n587, A2 => n1129, B1 => n553, B2 => n1130, 
                           ZN => n1256);
   U318 : OAI22_X1 port map( A1 => n654, A2 => n1131, B1 => n620, B2 => n1132, 
                           ZN => n1255);
   U319 : NOR4_X1 port map( A1 => n1259, A2 => n1261, A3 => n1262, A4 => n1263,
                           ZN => n1248);
   U320 : OAI22_X1 port map( A1 => n721, A2 => n1137, B1 => n687, B2 => n1138, 
                           ZN => n1263);
   U321 : OAI22_X1 port map( A1 => n788, A2 => n1139, B1 => n755, B2 => n1140, 
                           ZN => n1262);
   U322 : OAI22_X1 port map( A1 => n855, A2 => n1141, B1 => n822, B2 => n1142, 
                           ZN => n1261);
   U323 : OAI22_X1 port map( A1 => n923, A2 => n1143, B1 => n889, B2 => n1144, 
                           ZN => n1259);
   U324 : NOR4_X1 port map( A1 => n1264, A2 => n1265, A3 => n1266, A4 => n1267,
                           ZN => n1247);
   U325 : OAI22_X1 port map( A1 => n990, A2 => n1149, B1 => n956, B2 => n1151, 
                           ZN => n1267);
   U326 : OAI22_X1 port map( A1 => n1057, A2 => n1152, B1 => n1023, B2 => n1153
                           , ZN => n1266);
   U327 : OAI22_X1 port map( A1 => n102, A2 => n1154, B1 => n1091, B2 => n1155,
                           ZN => n1265);
   U328 : OAI22_X1 port map( A1 => n172, A2 => n1156, B1 => n137, B2 => n1157, 
                           ZN => n1264);
   U329 : OAI22_X1 port map( A1 => n1268, A2 => n1103, B1 => n1104, B2 => n1260
                           , ZN => N4604);
   U330 : NOR4_X1 port map( A1 => n1273, A2 => n1274, A3 => n1275, A4 => n1276,
                           ZN => n1272);
   U331 : OAI22_X1 port map( A1 => n194, A2 => n1113, B1 => n964, B2 => n1114, 
                           ZN => n1276);
   U332 : OAI22_X1 port map( A1 => n258, A2 => n1115, B1 => n226, B2 => n1116, 
                           ZN => n1275);
   U333 : OAI22_X1 port map( A1 => n322, A2 => n1117, B1 => n290, B2 => n1118, 
                           ZN => n1274);
   U334 : OAI22_X1 port map( A1 => n386, A2 => n1119, B1 => n354, B2 => n1120, 
                           ZN => n1273);
   U335 : NOR4_X1 port map( A1 => n1277, A2 => n1278, A3 => n1279, A4 => n1280,
                           ZN => n1271);
   U336 : OAI22_X1 port map( A1 => n451, A2 => n1125, B1 => n418, B2 => n1126, 
                           ZN => n1280);
   U337 : OAI22_X1 port map( A1 => n518, A2 => n1127, B1 => n485, B2 => n1128, 
                           ZN => n1279);
   U338 : OAI22_X1 port map( A1 => n585, A2 => n1129, B1 => n552, B2 => n1130, 
                           ZN => n1278);
   U339 : OAI22_X1 port map( A1 => n653, A2 => n1131, B1 => n619, B2 => n1132, 
                           ZN => n1277);
   U340 : NOR4_X1 port map( A1 => n1281, A2 => n1283, A3 => n1284, A4 => n1285,
                           ZN => n1270);
   U341 : OAI22_X1 port map( A1 => n720, A2 => n1137, B1 => n686, B2 => n1138, 
                           ZN => n1285);
   U342 : OAI22_X1 port map( A1 => n787, A2 => n1139, B1 => n753, B2 => n1140, 
                           ZN => n1284);
   U343 : OAI22_X1 port map( A1 => n854, A2 => n1141, B1 => n821, B2 => n2, ZN 
                           => n1283);
   U344 : OAI22_X1 port map( A1 => n921, A2 => n1143, B1 => n888, B2 => n37, ZN
                           => n1281);
   U345 : NOR4_X1 port map( A1 => n1286, A2 => n1287, A3 => n1288, A4 => n1289,
                           ZN => n1269);
   U346 : OAI22_X1 port map( A1 => n989, A2 => n1149, B1 => n955, B2 => n1151, 
                           ZN => n1289);
   U347 : OAI22_X1 port map( A1 => n1056, A2 => n1152, B1 => n1022, B2 => n1153
                           , ZN => n1288);
   U348 : OAI22_X1 port map( A1 => n101, A2 => n1154, B1 => n1089, B2 => n1155,
                           ZN => n1287);
   U349 : OAI22_X1 port map( A1 => n171, A2 => n1156, B1 => n136, B2 => n1157, 
                           ZN => n1286);
   U350 : OAI22_X1 port map( A1 => n1290, A2 => n1103, B1 => n1104, B2 => n1282
                           , ZN => N4602);
   U351 : NOR4_X1 port map( A1 => n1295, A2 => n1296, A3 => n1297, A4 => n1298,
                           ZN => n1294);
   U352 : OAI22_X1 port map( A1 => n193, A2 => n1113, B1 => n943, B2 => n1114, 
                           ZN => n1298);
   U353 : OAI22_X1 port map( A1 => n257, A2 => n1115, B1 => n225, B2 => n1116, 
                           ZN => n1297);
   U354 : OAI22_X1 port map( A1 => n321, A2 => n1117, B1 => n289, B2 => n1118, 
                           ZN => n1296);
   U355 : OAI22_X1 port map( A1 => n385, A2 => n1119, B1 => n353, B2 => n1120, 
                           ZN => n1295);
   U356 : NOR4_X1 port map( A1 => n1299, A2 => n1300, A3 => n1301, A4 => n1302,
                           ZN => n1293);
   U357 : OAI22_X1 port map( A1 => n450, A2 => n1125, B1 => n417, B2 => n1126, 
                           ZN => n1302);
   U358 : OAI22_X1 port map( A1 => n517, A2 => n1127, B1 => n484, B2 => n1128, 
                           ZN => n1301);
   U359 : OAI22_X1 port map( A1 => n584, A2 => n1129, B1 => n551, B2 => n1130, 
                           ZN => n1300);
   U360 : OAI22_X1 port map( A1 => n652, A2 => n1131, B1 => n618, B2 => n1132, 
                           ZN => n1299);
   U361 : NOR4_X1 port map( A1 => n1303, A2 => n1305, A3 => n1306, A4 => n1307,
                           ZN => n1292);
   U362 : OAI22_X1 port map( A1 => n719, A2 => n1137, B1 => n685, B2 => n1138, 
                           ZN => n1307);
   U363 : OAI22_X1 port map( A1 => n786, A2 => n1139, B1 => n752, B2 => n1140, 
                           ZN => n1306);
   U364 : OAI22_X1 port map( A1 => n853, A2 => n1141, B1 => n820, B2 => n1142, 
                           ZN => n1305);
   U365 : OAI22_X1 port map( A1 => n920, A2 => n1143, B1 => n887, B2 => n1144, 
                           ZN => n1303);
   U366 : NOR4_X1 port map( A1 => n1308, A2 => n1309, A3 => n1310, A4 => n1311,
                           ZN => n1291);
   U367 : OAI22_X1 port map( A1 => n988, A2 => n1149, B1 => n954, B2 => n1151, 
                           ZN => n1311);
   U368 : OAI22_X1 port map( A1 => n1055, A2 => n1152, B1 => n1021, B2 => n1153
                           , ZN => n1310);
   U369 : OAI22_X1 port map( A1 => n100, A2 => n1154, B1 => n1088, B2 => n1155,
                           ZN => n1309);
   U370 : OAI22_X1 port map( A1 => n170, A2 => n1156, B1 => n135, B2 => n1157, 
                           ZN => n1308);
   U371 : OAI22_X1 port map( A1 => n1312, A2 => n1103, B1 => n1104, B2 => n1304
                           , ZN => N4600);
   U372 : NOR4_X1 port map( A1 => n1317, A2 => n1318, A3 => n1319, A4 => n1320,
                           ZN => n1316);
   U373 : OAI22_X1 port map( A1 => n192, A2 => n1113, B1 => n922, B2 => n1114, 
                           ZN => n1320);
   U374 : OAI22_X1 port map( A1 => n256, A2 => n1115, B1 => n224, B2 => n1116, 
                           ZN => n1319);
   U375 : OAI22_X1 port map( A1 => n320, A2 => n1117, B1 => n288, B2 => n1118, 
                           ZN => n1318);
   U376 : OAI22_X1 port map( A1 => n384, A2 => n1119, B1 => n352, B2 => n1120, 
                           ZN => n1317);
   U377 : NOR4_X1 port map( A1 => n1321, A2 => n1322, A3 => n1323, A4 => n1324,
                           ZN => n1315);
   U378 : OAI22_X1 port map( A1 => n449, A2 => n1125, B1 => n416, B2 => n1126, 
                           ZN => n1324);
   U379 : OAI22_X1 port map( A1 => n516, A2 => n1127, B1 => n483, B2 => n1128, 
                           ZN => n1323);
   U380 : OAI22_X1 port map( A1 => n583, A2 => n1129, B1 => n550, B2 => n1130, 
                           ZN => n1322);
   U381 : OAI22_X1 port map( A1 => n651, A2 => n1131, B1 => n617, B2 => n1132, 
                           ZN => n1321);
   U382 : NOR4_X1 port map( A1 => n1325, A2 => n1327, A3 => n1328, A4 => n1329,
                           ZN => n1314);
   U383 : OAI22_X1 port map( A1 => n718, A2 => n1137, B1 => n684, B2 => n1138, 
                           ZN => n1329);
   U384 : OAI22_X1 port map( A1 => n785, A2 => n1139, B1 => n751, B2 => n1140, 
                           ZN => n1328);
   U385 : OAI22_X1 port map( A1 => n852, A2 => n1141, B1 => n819, B2 => n1142, 
                           ZN => n1327);
   U386 : OAI22_X1 port map( A1 => n919, A2 => n1143, B1 => n886, B2 => n1144, 
                           ZN => n1325);
   U387 : NOR4_X1 port map( A1 => n1330, A2 => n1331, A3 => n1332, A4 => n1333,
                           ZN => n1313);
   U388 : OAI22_X1 port map( A1 => n987, A2 => n1149, B1 => n953, B2 => n1151, 
                           ZN => n1333);
   U389 : OAI22_X1 port map( A1 => n1054, A2 => n1152, B1 => n1020, B2 => n1153
                           , ZN => n1332);
   U390 : OAI22_X1 port map( A1 => n97, A2 => n1154, B1 => n1087, B2 => n1155, 
                           ZN => n1331);
   U391 : OAI22_X1 port map( A1 => n169, A2 => n1156, B1 => n134, B2 => n1157, 
                           ZN => n1330);
   U392 : OAI22_X1 port map( A1 => n1334, A2 => n1103, B1 => n1104, B2 => n1326
                           , ZN => N4598);
   U393 : NOR4_X1 port map( A1 => n1339, A2 => n1340, A3 => n1341, A4 => n1342,
                           ZN => n1338);
   U394 : OAI22_X1 port map( A1 => n191, A2 => n1113, B1 => n901, B2 => n1114, 
                           ZN => n1342);
   U395 : OAI22_X1 port map( A1 => n255, A2 => n1115, B1 => n223, B2 => n1116, 
                           ZN => n1341);
   U396 : OAI22_X1 port map( A1 => n319, A2 => n1117, B1 => n287, B2 => n1118, 
                           ZN => n1340);
   U397 : OAI22_X1 port map( A1 => n383, A2 => n1119, B1 => n351, B2 => n1120, 
                           ZN => n1339);
   U398 : NOR4_X1 port map( A1 => n1343, A2 => n1344, A3 => n1345, A4 => n1346,
                           ZN => n1337);
   U399 : OAI22_X1 port map( A1 => n448, A2 => n1125, B1 => n415, B2 => n1126, 
                           ZN => n1346);
   U400 : OAI22_X1 port map( A1 => n515, A2 => n1127, B1 => n482, B2 => n1128, 
                           ZN => n1345);
   U401 : OAI22_X1 port map( A1 => n582, A2 => n1129, B1 => n549, B2 => n1130, 
                           ZN => n1344);
   U402 : OAI22_X1 port map( A1 => n650, A2 => n1131, B1 => n616, B2 => n1132, 
                           ZN => n1343);
   U403 : NOR4_X1 port map( A1 => n1347, A2 => n1349, A3 => n1350, A4 => n1351,
                           ZN => n1336);
   U404 : OAI22_X1 port map( A1 => n717, A2 => n1137, B1 => n683, B2 => n1138, 
                           ZN => n1351);
   U405 : OAI22_X1 port map( A1 => n784, A2 => n1139, B1 => n750, B2 => n1140, 
                           ZN => n1350);
   U406 : OAI22_X1 port map( A1 => n851, A2 => n1141, B1 => n818, B2 => n1142, 
                           ZN => n1349);
   U407 : OAI22_X1 port map( A1 => n918, A2 => n1143, B1 => n885, B2 => n1144, 
                           ZN => n1347);
   U408 : NOR4_X1 port map( A1 => n1352, A2 => n1353, A3 => n1354, A4 => n1355,
                           ZN => n1335);
   U409 : OAI22_X1 port map( A1 => n986, A2 => n1149, B1 => n952, B2 => n1151, 
                           ZN => n1355);
   U410 : OAI22_X1 port map( A1 => n1053, A2 => n1152, B1 => n1019, B2 => n1153
                           , ZN => n1354);
   U411 : OAI22_X1 port map( A1 => n95, A2 => n1154, B1 => n1086, B2 => n1155, 
                           ZN => n1353);
   U412 : OAI22_X1 port map( A1 => n168, A2 => n1156, B1 => n133, B2 => n1157, 
                           ZN => n1352);
   U413 : OAI22_X1 port map( A1 => n1356, A2 => n1103, B1 => n1104, B2 => n1348
                           , ZN => N4596);
   U414 : NOR4_X1 port map( A1 => n1361, A2 => n1362, A3 => n1363, A4 => n1364,
                           ZN => n1360);
   U415 : OAI22_X1 port map( A1 => n190, A2 => n1113, B1 => n880, B2 => n1114, 
                           ZN => n1364);
   U416 : OAI22_X1 port map( A1 => n254, A2 => n1115, B1 => n222, B2 => n1116, 
                           ZN => n1363);
   U417 : OAI22_X1 port map( A1 => n318, A2 => n1117, B1 => n286, B2 => n1118, 
                           ZN => n1362);
   U418 : OAI22_X1 port map( A1 => n382, A2 => n1119, B1 => n350, B2 => n1120, 
                           ZN => n1361);
   U419 : NOR4_X1 port map( A1 => n1365, A2 => n1366, A3 => n1367, A4 => n1368,
                           ZN => n1359);
   U420 : OAI22_X1 port map( A1 => n447, A2 => n1125, B1 => n414, B2 => n1126, 
                           ZN => n1368);
   U421 : OAI22_X1 port map( A1 => n514, A2 => n1127, B1 => n480, B2 => n1128, 
                           ZN => n1367);
   U422 : OAI22_X1 port map( A1 => n581, A2 => n1129, B1 => n548, B2 => n1130, 
                           ZN => n1366);
   U423 : OAI22_X1 port map( A1 => n648, A2 => n1131, B1 => n615, B2 => n1132, 
                           ZN => n1365);
   U424 : NOR4_X1 port map( A1 => n1369, A2 => n1371, A3 => n1372, A4 => n1373,
                           ZN => n1358);
   U425 : OAI22_X1 port map( A1 => n716, A2 => n1137, B1 => n682, B2 => n1138, 
                           ZN => n1373);
   U426 : OAI22_X1 port map( A1 => n783, A2 => n1139, B1 => n749, B2 => n1140, 
                           ZN => n1372);
   U427 : OAI22_X1 port map( A1 => n850, A2 => n1141, B1 => n816, B2 => n1142, 
                           ZN => n1371);
   U428 : OAI22_X1 port map( A1 => n917, A2 => n1143, B1 => n884, B2 => n1144, 
                           ZN => n1369);
   U429 : NOR4_X1 port map( A1 => n1374, A2 => n1375, A3 => n1376, A4 => n1377,
                           ZN => n1357);
   U430 : OAI22_X1 port map( A1 => n984, A2 => n1149, B1 => n951, B2 => n1151, 
                           ZN => n1377);
   U431 : OAI22_X1 port map( A1 => n1052, A2 => n1152, B1 => n1018, B2 => n1153
                           , ZN => n1376);
   U432 : OAI22_X1 port map( A1 => n93, A2 => n1154, B1 => n1085, B2 => n1155, 
                           ZN => n1375);
   U433 : OAI22_X1 port map( A1 => n167, A2 => n1156, B1 => n131, B2 => n1157, 
                           ZN => n1374);
   U434 : OAI22_X1 port map( A1 => n1378, A2 => n1103, B1 => n1104, B2 => n1370
                           , ZN => N4594);
   U435 : NOR4_X1 port map( A1 => n1383, A2 => n1384, A3 => n1385, A4 => n1386,
                           ZN => n1382);
   U436 : OAI22_X1 port map( A1 => n189, A2 => n1113, B1 => n859, B2 => n1114, 
                           ZN => n1386);
   U437 : OAI22_X1 port map( A1 => n253, A2 => n1115, B1 => n221, B2 => n1116, 
                           ZN => n1385);
   U438 : OAI22_X1 port map( A1 => n317, A2 => n1117, B1 => n285, B2 => n1118, 
                           ZN => n1384);
   U439 : OAI22_X1 port map( A1 => n381, A2 => n1119, B1 => n349, B2 => n1120, 
                           ZN => n1383);
   U440 : NOR4_X1 port map( A1 => n1387, A2 => n1388, A3 => n1389, A4 => n1390,
                           ZN => n1381);
   U441 : OAI22_X1 port map( A1 => n446, A2 => n1125, B1 => n413, B2 => n1126, 
                           ZN => n1390);
   U442 : OAI22_X1 port map( A1 => n513, A2 => n1127, B1 => n479, B2 => n1128, 
                           ZN => n1389);
   U443 : OAI22_X1 port map( A1 => n580, A2 => n1129, B1 => n547, B2 => n1130, 
                           ZN => n1388);
   U444 : OAI22_X1 port map( A1 => n647, A2 => n1131, B1 => n614, B2 => n1132, 
                           ZN => n1387);
   U445 : NOR4_X1 port map( A1 => n1391, A2 => n1393, A3 => n1394, A4 => n1395,
                           ZN => n1380);
   U446 : OAI22_X1 port map( A1 => n715, A2 => n1137, B1 => n681, B2 => n1138, 
                           ZN => n1395);
   U447 : OAI22_X1 port map( A1 => n782, A2 => n1139, B1 => n748, B2 => n1140, 
                           ZN => n1394);
   U448 : OAI22_X1 port map( A1 => n849, A2 => n1141, B1 => n815, B2 => n1142, 
                           ZN => n1393);
   U449 : OAI22_X1 port map( A1 => n916, A2 => n1143, B1 => n883, B2 => n1144, 
                           ZN => n1391);
   U450 : NOR4_X1 port map( A1 => n1396, A2 => n1397, A3 => n1398, A4 => n1399,
                           ZN => n1379);
   U451 : OAI22_X1 port map( A1 => n983, A2 => n1149, B1 => n950, B2 => n1151, 
                           ZN => n1399);
   U452 : OAI22_X1 port map( A1 => n1051, A2 => n1152, B1 => n1017, B2 => n1153
                           , ZN => n1398);
   U453 : OAI22_X1 port map( A1 => n91, A2 => n1154, B1 => n1084, B2 => n1155, 
                           ZN => n1397);
   U454 : OAI22_X1 port map( A1 => n166, A2 => n1156, B1 => n130, B2 => n1157, 
                           ZN => n1396);
   U455 : OAI22_X1 port map( A1 => n1400, A2 => n1103, B1 => n1104, B2 => n1392
                           , ZN => N4592);
   U456 : NOR4_X1 port map( A1 => n1405, A2 => n1406, A3 => n1407, A4 => n1408,
                           ZN => n1404);
   U457 : OAI22_X1 port map( A1 => n188, A2 => n1113, B1 => n838, B2 => n1114, 
                           ZN => n1408);
   U458 : OAI22_X1 port map( A1 => n252, A2 => n1115, B1 => n220, B2 => n1116, 
                           ZN => n1407);
   U459 : OAI22_X1 port map( A1 => n316, A2 => n1117, B1 => n284, B2 => n1118, 
                           ZN => n1406);
   U460 : OAI22_X1 port map( A1 => n380, A2 => n1119, B1 => n348, B2 => n1120, 
                           ZN => n1405);
   U461 : NOR4_X1 port map( A1 => n1409, A2 => n1410, A3 => n1411, A4 => n1412,
                           ZN => n1403);
   U462 : OAI22_X1 port map( A1 => n445, A2 => n1125, B1 => n412, B2 => n1126, 
                           ZN => n1412);
   U463 : OAI22_X1 port map( A1 => n512, A2 => n1127, B1 => n478, B2 => n1128, 
                           ZN => n1411);
   U464 : OAI22_X1 port map( A1 => n579, A2 => n1129, B1 => n546, B2 => n1130, 
                           ZN => n1410);
   U465 : OAI22_X1 port map( A1 => n646, A2 => n1131, B1 => n613, B2 => n1132, 
                           ZN => n1409);
   U466 : NOR4_X1 port map( A1 => n1413, A2 => n1415, A3 => n1416, A4 => n1417,
                           ZN => n1402);
   U467 : OAI22_X1 port map( A1 => n714, A2 => n1137, B1 => n680, B2 => n1138, 
                           ZN => n1417);
   U468 : OAI22_X1 port map( A1 => n781, A2 => n1139, B1 => n747, B2 => n1140, 
                           ZN => n1416);
   U469 : OAI22_X1 port map( A1 => n848, A2 => n1141, B1 => n814, B2 => n1142, 
                           ZN => n1415);
   U470 : OAI22_X1 port map( A1 => n915, A2 => n1143, B1 => n882, B2 => n1144, 
                           ZN => n1413);
   U471 : NOR4_X1 port map( A1 => n1418, A2 => n1419, A3 => n1420, A4 => n1421,
                           ZN => n1401);
   U472 : OAI22_X1 port map( A1 => n982, A2 => n1149, B1 => n949, B2 => n1151, 
                           ZN => n1421);
   U473 : OAI22_X1 port map( A1 => n1050, A2 => n1152, B1 => n1016, B2 => n1153
                           , ZN => n1420);
   U474 : OAI22_X1 port map( A1 => n89, A2 => n1154, B1 => n1083, B2 => n1155, 
                           ZN => n1419);
   U475 : OAI22_X1 port map( A1 => n164, A2 => n1156, B1 => n129, B2 => n1157, 
                           ZN => n1418);
   U476 : OAI22_X1 port map( A1 => n1422, A2 => n1103, B1 => n1104, B2 => n1414
                           , ZN => N4590);
   U477 : NOR4_X1 port map( A1 => n1427, A2 => n1428, A3 => n1429, A4 => n1430,
                           ZN => n1426);
   U478 : OAI22_X1 port map( A1 => n187, A2 => n1113, B1 => n817, B2 => n1114, 
                           ZN => n1430);
   U479 : OAI22_X1 port map( A1 => n251, A2 => n1115, B1 => n219, B2 => n1116, 
                           ZN => n1429);
   U480 : OAI22_X1 port map( A1 => n315, A2 => n1117, B1 => n283, B2 => n1118, 
                           ZN => n1428);
   U481 : OAI22_X1 port map( A1 => n379, A2 => n1119, B1 => n347, B2 => n1120, 
                           ZN => n1427);
   U482 : NOR4_X1 port map( A1 => n1431, A2 => n1432, A3 => n1433, A4 => n1434,
                           ZN => n1425);
   U483 : OAI22_X1 port map( A1 => n444, A2 => n1125, B1 => n411, B2 => n1126, 
                           ZN => n1434);
   U484 : OAI22_X1 port map( A1 => n511, A2 => n1127, B1 => n477, B2 => n1128, 
                           ZN => n1433);
   U485 : OAI22_X1 port map( A1 => n578, A2 => n1129, B1 => n545, B2 => n1130, 
                           ZN => n1432);
   U486 : OAI22_X1 port map( A1 => n645, A2 => n1131, B1 => n612, B2 => n1132, 
                           ZN => n1431);
   U487 : NOR4_X1 port map( A1 => n1435, A2 => n1437, A3 => n1438, A4 => n1439,
                           ZN => n1424);
   U488 : OAI22_X1 port map( A1 => n713, A2 => n1137, B1 => n679, B2 => n1138, 
                           ZN => n1439);
   U489 : OAI22_X1 port map( A1 => n780, A2 => n1139, B1 => n746, B2 => n1140, 
                           ZN => n1438);
   U490 : OAI22_X1 port map( A1 => n847, A2 => n1141, B1 => n813, B2 => n1142, 
                           ZN => n1437);
   U491 : OAI22_X1 port map( A1 => n914, A2 => n1143, B1 => n881, B2 => n1144, 
                           ZN => n1435);
   U492 : NOR4_X1 port map( A1 => n1440, A2 => n1441, A3 => n1442, A4 => n1443,
                           ZN => n1423);
   U493 : OAI22_X1 port map( A1 => n981, A2 => n1149, B1 => n948, B2 => n1151, 
                           ZN => n1443);
   U494 : OAI22_X1 port map( A1 => n1049, A2 => n1152, B1 => n1015, B2 => n1153
                           , ZN => n1442);
   U495 : OAI22_X1 port map( A1 => n87, A2 => n1154, B1 => n1082, B2 => n1155, 
                           ZN => n1441);
   U496 : OAI22_X1 port map( A1 => n163, A2 => n1156, B1 => n128, B2 => n1157, 
                           ZN => n1440);
   U497 : OAI22_X1 port map( A1 => n1444, A2 => n1103, B1 => n1104, B2 => n1436
                           , ZN => N4588);
   U498 : NOR4_X1 port map( A1 => n1449, A2 => n1450, A3 => n1451, A4 => n1452,
                           ZN => n1448);
   U499 : OAI22_X1 port map( A1 => n186, A2 => n1113, B1 => n796, B2 => n1114, 
                           ZN => n1452);
   U500 : OAI22_X1 port map( A1 => n250, A2 => n1115, B1 => n218, B2 => n1116, 
                           ZN => n1451);
   U501 : OAI22_X1 port map( A1 => n314, A2 => n1117, B1 => n282, B2 => n1118, 
                           ZN => n1450);
   U502 : OAI22_X1 port map( A1 => n378, A2 => n1119, B1 => n346, B2 => n1120, 
                           ZN => n1449);
   U503 : NOR4_X1 port map( A1 => n1453, A2 => n1454, A3 => n1455, A4 => n1456,
                           ZN => n1447);
   U504 : OAI22_X1 port map( A1 => n443, A2 => n1125, B1 => n410, B2 => n1126, 
                           ZN => n1456);
   U505 : OAI22_X1 port map( A1 => n510, A2 => n1127, B1 => n476, B2 => n1128, 
                           ZN => n1455);
   U506 : OAI22_X1 port map( A1 => n577, A2 => n1129, B1 => n543, B2 => n1130, 
                           ZN => n1454);
   U507 : OAI22_X1 port map( A1 => n644, A2 => n1131, B1 => n611, B2 => n1132, 
                           ZN => n1453);
   U508 : NOR4_X1 port map( A1 => n1457, A2 => n1459, A3 => n1460, A4 => n1461,
                           ZN => n1446);
   U509 : OAI22_X1 port map( A1 => n711, A2 => n1137, B1 => n678, B2 => n1138, 
                           ZN => n1461);
   U510 : OAI22_X1 port map( A1 => n779, A2 => n1139, B1 => n745, B2 => n1140, 
                           ZN => n1460);
   U511 : OAI22_X1 port map( A1 => n846, A2 => n1141, B1 => n812, B2 => n1142, 
                           ZN => n1459);
   U512 : OAI22_X1 port map( A1 => n913, A2 => n1143, B1 => n879, B2 => n1144, 
                           ZN => n1457);
   U513 : NOR4_X1 port map( A1 => n1462, A2 => n1463, A3 => n1464, A4 => n1465,
                           ZN => n1445);
   U514 : OAI22_X1 port map( A1 => n980, A2 => n1149, B1 => n947, B2 => n1151, 
                           ZN => n1465);
   U515 : OAI22_X1 port map( A1 => n1047, A2 => n1152, B1 => n1014, B2 => n1153
                           , ZN => n1464);
   U516 : OAI22_X1 port map( A1 => n85, A2 => n1154, B1 => n1081, B2 => n1155, 
                           ZN => n1463);
   U517 : OAI22_X1 port map( A1 => n162, A2 => n1156, B1 => n127, B2 => n1157, 
                           ZN => n1462);
   U518 : OAI22_X1 port map( A1 => n1466, A2 => n1103, B1 => n1104, B2 => n1458
                           , ZN => N4586);
   U519 : NOR4_X1 port map( A1 => n1471, A2 => n1472, A3 => n1473, A4 => n1474,
                           ZN => n1470);
   U520 : OAI22_X1 port map( A1 => n185, A2 => n1113, B1 => n775, B2 => n1114, 
                           ZN => n1474);
   U521 : OAI22_X1 port map( A1 => n249, A2 => n1115, B1 => n217, B2 => n1116, 
                           ZN => n1473);
   U522 : OAI22_X1 port map( A1 => n313, A2 => n1117, B1 => n281, B2 => n1118, 
                           ZN => n1472);
   U523 : OAI22_X1 port map( A1 => n377, A2 => n1119, B1 => n345, B2 => n1120, 
                           ZN => n1471);
   U524 : NOR4_X1 port map( A1 => n1475, A2 => n1476, A3 => n1477, A4 => n1478,
                           ZN => n1469);
   U525 : OAI22_X1 port map( A1 => n442, A2 => n1125, B1 => n409, B2 => n1126, 
                           ZN => n1478);
   U526 : OAI22_X1 port map( A1 => n509, A2 => n1127, B1 => n475, B2 => n1128, 
                           ZN => n1477);
   U527 : OAI22_X1 port map( A1 => n576, A2 => n1129, B1 => n542, B2 => n1130, 
                           ZN => n1476);
   U528 : OAI22_X1 port map( A1 => n643, A2 => n1131, B1 => n610, B2 => n1132, 
                           ZN => n1475);
   U529 : NOR4_X1 port map( A1 => n1479, A2 => n1481, A3 => n1482, A4 => n1483,
                           ZN => n1468);
   U530 : OAI22_X1 port map( A1 => n710, A2 => n1137, B1 => n677, B2 => n1138, 
                           ZN => n1483);
   U531 : OAI22_X1 port map( A1 => n778, A2 => n1139, B1 => n744, B2 => n1140, 
                           ZN => n1482);
   U532 : OAI22_X1 port map( A1 => n845, A2 => n1141, B1 => n811, B2 => n1142, 
                           ZN => n1481);
   U533 : OAI22_X1 port map( A1 => n912, A2 => n1143, B1 => n878, B2 => n1144, 
                           ZN => n1479);
   U534 : NOR4_X1 port map( A1 => n1484, A2 => n1485, A3 => n1486, A4 => n1487,
                           ZN => n1467);
   U535 : OAI22_X1 port map( A1 => n979, A2 => n1149, B1 => n946, B2 => n1151, 
                           ZN => n1487);
   U536 : OAI22_X1 port map( A1 => n1046, A2 => n1152, B1 => n1013, B2 => n1153
                           , ZN => n1486);
   U537 : OAI22_X1 port map( A1 => n83, A2 => n1154, B1 => n1080, B2 => n1155, 
                           ZN => n1485);
   U538 : OAI22_X1 port map( A1 => n161, A2 => n1156, B1 => n126, B2 => n1157, 
                           ZN => n1484);
   U539 : OAI22_X1 port map( A1 => n1488, A2 => n1103, B1 => n1104, B2 => n1480
                           , ZN => N4584);
   U540 : NOR4_X1 port map( A1 => n1493, A2 => n1494, A3 => n1495, A4 => n1496,
                           ZN => n1492);
   U541 : OAI22_X1 port map( A1 => n184, A2 => n1113, B1 => n754, B2 => n1114, 
                           ZN => n1496);
   U542 : OAI22_X1 port map( A1 => n248, A2 => n1115, B1 => n216, B2 => n1116, 
                           ZN => n1495);
   U543 : OAI22_X1 port map( A1 => n312, A2 => n1117, B1 => n280, B2 => n1118, 
                           ZN => n1494);
   U544 : OAI22_X1 port map( A1 => n376, A2 => n1119, B1 => n344, B2 => n1120, 
                           ZN => n1493);
   U545 : NOR4_X1 port map( A1 => n1497, A2 => n1498, A3 => n1499, A4 => n1500,
                           ZN => n1491);
   U546 : OAI22_X1 port map( A1 => n441, A2 => n1125, B1 => n408, B2 => n1126, 
                           ZN => n1500);
   U547 : OAI22_X1 port map( A1 => n508, A2 => n1127, B1 => n474, B2 => n1128, 
                           ZN => n1499);
   U548 : OAI22_X1 port map( A1 => n575, A2 => n1129, B1 => n541, B2 => n1130, 
                           ZN => n1498);
   U549 : OAI22_X1 port map( A1 => n642, A2 => n1131, B1 => n609, B2 => n1132, 
                           ZN => n1497);
   U550 : NOR4_X1 port map( A1 => n1501, A2 => n1503, A3 => n1504, A4 => n1505,
                           ZN => n1490);
   U551 : OAI22_X1 port map( A1 => n709, A2 => n1137, B1 => n676, B2 => n1138, 
                           ZN => n1505);
   U552 : OAI22_X1 port map( A1 => n777, A2 => n1139, B1 => n743, B2 => n1140, 
                           ZN => n1504);
   U553 : OAI22_X1 port map( A1 => n844, A2 => n1141, B1 => n810, B2 => n1142, 
                           ZN => n1503);
   U554 : OAI22_X1 port map( A1 => n911, A2 => n1143, B1 => n877, B2 => n1144, 
                           ZN => n1501);
   U555 : NOR4_X1 port map( A1 => n1506, A2 => n1507, A3 => n1508, A4 => n1509,
                           ZN => n1489);
   U556 : OAI22_X1 port map( A1 => n978, A2 => n1149, B1 => n945, B2 => n1151, 
                           ZN => n1509);
   U557 : OAI22_X1 port map( A1 => n1045, A2 => n1152, B1 => n1012, B2 => n1153
                           , ZN => n1508);
   U558 : OAI22_X1 port map( A1 => n81, A2 => n1154, B1 => n1079, B2 => n1155, 
                           ZN => n1507);
   U559 : OAI22_X1 port map( A1 => n160, A2 => n1156, B1 => n125, B2 => n1157, 
                           ZN => n1506);
   U560 : OAI22_X1 port map( A1 => n1510, A2 => n1103, B1 => n1104, B2 => n1502
                           , ZN => N4582);
   U561 : NOR4_X1 port map( A1 => n1515, A2 => n1516, A3 => n1517, A4 => n1518,
                           ZN => n1514);
   U562 : OAI22_X1 port map( A1 => n183, A2 => n1113, B1 => n733, B2 => n1114, 
                           ZN => n1518);
   U563 : OAI22_X1 port map( A1 => n247, A2 => n1115, B1 => n215, B2 => n1116, 
                           ZN => n1517);
   U564 : OAI22_X1 port map( A1 => n311, A2 => n1117, B1 => n279, B2 => n1118, 
                           ZN => n1516);
   U565 : OAI22_X1 port map( A1 => n375, A2 => n1119, B1 => n343, B2 => n1120, 
                           ZN => n1515);
   U566 : NOR4_X1 port map( A1 => n1519, A2 => n1520, A3 => n1521, A4 => n1522,
                           ZN => n1513);
   U567 : OAI22_X1 port map( A1 => n440, A2 => n1125, B1 => n407, B2 => n1126, 
                           ZN => n1522);
   U568 : OAI22_X1 port map( A1 => n507, A2 => n1127, B1 => n473, B2 => n1128, 
                           ZN => n1521);
   U569 : OAI22_X1 port map( A1 => n574, A2 => n1129, B1 => n540, B2 => n1130, 
                           ZN => n1520);
   U570 : OAI22_X1 port map( A1 => n641, A2 => n1131, B1 => n608, B2 => n1132, 
                           ZN => n1519);
   U571 : NOR4_X1 port map( A1 => n1523, A2 => n1525, A3 => n1526, A4 => n1527,
                           ZN => n1512);
   U572 : OAI22_X1 port map( A1 => n708, A2 => n1137, B1 => n675, B2 => n1138, 
                           ZN => n1527);
   U573 : OAI22_X1 port map( A1 => n776, A2 => n1139, B1 => n742, B2 => n1140, 
                           ZN => n1526);
   U574 : OAI22_X1 port map( A1 => n843, A2 => n1141, B1 => n809, B2 => n1142, 
                           ZN => n1525);
   U575 : OAI22_X1 port map( A1 => n910, A2 => n1143, B1 => n876, B2 => n1144, 
                           ZN => n1523);
   U576 : NOR4_X1 port map( A1 => n1528, A2 => n1529, A3 => n1530, A4 => n1531,
                           ZN => n1511);
   U577 : OAI22_X1 port map( A1 => n977, A2 => n1149, B1 => n944, B2 => n1151, 
                           ZN => n1531);
   U578 : OAI22_X1 port map( A1 => n1044, A2 => n1152, B1 => n1011, B2 => n1153
                           , ZN => n1530);
   U579 : OAI22_X1 port map( A1 => n79, A2 => n1154, B1 => n1078, B2 => n1155, 
                           ZN => n1529);
   U580 : OAI22_X1 port map( A1 => n159, A2 => n1156, B1 => n124, B2 => n1157, 
                           ZN => n1528);
   U581 : OAI22_X1 port map( A1 => n1532, A2 => n1103, B1 => n1104, B2 => n1524
                           , ZN => N4580);
   U582 : NOR4_X1 port map( A1 => n1537, A2 => n1538, A3 => n1539, A4 => n1540,
                           ZN => n1536);
   U583 : OAI22_X1 port map( A1 => n182, A2 => n1113, B1 => n712, B2 => n1114, 
                           ZN => n1540);
   U584 : OAI22_X1 port map( A1 => n246, A2 => n1115, B1 => n214, B2 => n1116, 
                           ZN => n1539);
   U585 : OAI22_X1 port map( A1 => n310, A2 => n1117, B1 => n278, B2 => n1118, 
                           ZN => n1538);
   U586 : OAI22_X1 port map( A1 => n374, A2 => n1119, B1 => n342, B2 => n1120, 
                           ZN => n1537);
   U587 : NOR4_X1 port map( A1 => n1541, A2 => n1542, A3 => n1543, A4 => n1544,
                           ZN => n1535);
   U588 : OAI22_X1 port map( A1 => n438, A2 => n1125, B1 => n406, B2 => n1126, 
                           ZN => n1544);
   U589 : OAI22_X1 port map( A1 => n506, A2 => n1127, B1 => n472, B2 => n1128, 
                           ZN => n1543);
   U590 : OAI22_X1 port map( A1 => n573, A2 => n1129, B1 => n539, B2 => n1130, 
                           ZN => n1542);
   U591 : OAI22_X1 port map( A1 => n640, A2 => n1131, B1 => n606, B2 => n1132, 
                           ZN => n1541);
   U592 : NOR4_X1 port map( A1 => n1545, A2 => n1547, A3 => n1548, A4 => n1549,
                           ZN => n1534);
   U593 : OAI22_X1 port map( A1 => n707, A2 => n1137, B1 => n674, B2 => n1138, 
                           ZN => n1549);
   U594 : OAI22_X1 port map( A1 => n774, A2 => n1139, B1 => n741, B2 => n1140, 
                           ZN => n1548);
   U595 : OAI22_X1 port map( A1 => n842, A2 => n1141, B1 => n808, B2 => n1142, 
                           ZN => n1547);
   U596 : OAI22_X1 port map( A1 => n909, A2 => n1143, B1 => n875, B2 => n1144, 
                           ZN => n1545);
   U597 : NOR4_X1 port map( A1 => n1550, A2 => n1551, A3 => n1552, A4 => n1553,
                           ZN => n1533);
   U598 : OAI22_X1 port map( A1 => n976, A2 => n1149, B1 => n942, B2 => n1151, 
                           ZN => n1553);
   U599 : OAI22_X1 port map( A1 => n1043, A2 => n1152, B1 => n1010, B2 => n1153
                           , ZN => n1552);
   U600 : OAI22_X1 port map( A1 => n75, A2 => n1154, B1 => n1077, B2 => n1155, 
                           ZN => n1551);
   U601 : OAI22_X1 port map( A1 => n158, A2 => n1156, B1 => n123, B2 => n1157, 
                           ZN => n1550);
   U602 : OAI22_X1 port map( A1 => n1554, A2 => n1103, B1 => n1104, B2 => n1546
                           , ZN => N4578);
   U603 : NOR4_X1 port map( A1 => n1559, A2 => n1560, A3 => n1561, A4 => n1562,
                           ZN => n1558);
   U604 : OAI22_X1 port map( A1 => n181, A2 => n1113, B1 => n691, B2 => n1114, 
                           ZN => n1562);
   U605 : OAI22_X1 port map( A1 => n245, A2 => n1115, B1 => n213, B2 => n1116, 
                           ZN => n1561);
   U606 : OAI22_X1 port map( A1 => n309, A2 => n1117, B1 => n277, B2 => n1118, 
                           ZN => n1560);
   U607 : OAI22_X1 port map( A1 => n373, A2 => n1119, B1 => n341, B2 => n1120, 
                           ZN => n1559);
   U608 : NOR4_X1 port map( A1 => n1563, A2 => n1564, A3 => n1565, A4 => n1566,
                           ZN => n1557);
   U609 : OAI22_X1 port map( A1 => n437, A2 => n1125, B1 => n405, B2 => n1126, 
                           ZN => n1566);
   U610 : OAI22_X1 port map( A1 => n505, A2 => n1127, B1 => n471, B2 => n1128, 
                           ZN => n1565);
   U611 : OAI22_X1 port map( A1 => n572, A2 => n1129, B1 => n538, B2 => n1130, 
                           ZN => n1564);
   U612 : OAI22_X1 port map( A1 => n639, A2 => n1131, B1 => n605, B2 => n1132, 
                           ZN => n1563);
   U613 : NOR4_X1 port map( A1 => n1567, A2 => n1569, A3 => n1570, A4 => n1571,
                           ZN => n1556);
   U614 : OAI22_X1 port map( A1 => n706, A2 => n1137, B1 => n673, B2 => n1138, 
                           ZN => n1571);
   U615 : OAI22_X1 port map( A1 => n773, A2 => n1139, B1 => n740, B2 => n1140, 
                           ZN => n1570);
   U616 : OAI22_X1 port map( A1 => n841, A2 => n1141, B1 => n807, B2 => n1142, 
                           ZN => n1569);
   U617 : OAI22_X1 port map( A1 => n908, A2 => n1143, B1 => n874, B2 => n1144, 
                           ZN => n1567);
   U618 : NOR4_X1 port map( A1 => n1572, A2 => n1573, A3 => n1574, A4 => n1575,
                           ZN => n1555);
   U619 : OAI22_X1 port map( A1 => n975, A2 => n1149, B1 => n941, B2 => n1151, 
                           ZN => n1575);
   U620 : OAI22_X1 port map( A1 => n1042, A2 => n1152, B1 => n1009, B2 => n1153
                           , ZN => n1574);
   U621 : OAI22_X1 port map( A1 => n73, A2 => n1154, B1 => n1076, B2 => n1155, 
                           ZN => n1573);
   U622 : OAI22_X1 port map( A1 => n157, A2 => n1156, B1 => n122, B2 => n1157, 
                           ZN => n1572);
   U623 : OAI22_X1 port map( A1 => n1576, A2 => n1103, B1 => n1104, B2 => n1568
                           , ZN => N4576);
   U624 : NOR4_X1 port map( A1 => n1581, A2 => n1582, A3 => n1583, A4 => n1584,
                           ZN => n1580);
   U625 : OAI22_X1 port map( A1 => n180, A2 => n1113, B1 => n670, B2 => n1114, 
                           ZN => n1584);
   U626 : OAI22_X1 port map( A1 => n244, A2 => n1115, B1 => n212, B2 => n1116, 
                           ZN => n1583);
   U627 : OAI22_X1 port map( A1 => n308, A2 => n1117, B1 => n276, B2 => n1118, 
                           ZN => n1582);
   U628 : OAI22_X1 port map( A1 => n372, A2 => n1119, B1 => n340, B2 => n1120, 
                           ZN => n1581);
   U629 : NOR4_X1 port map( A1 => n1585, A2 => n1586, A3 => n1587, A4 => n1588,
                           ZN => n1579);
   U630 : OAI22_X1 port map( A1 => n436, A2 => n1125, B1 => n404, B2 => n1126, 
                           ZN => n1588);
   U631 : OAI22_X1 port map( A1 => n504, A2 => n1127, B1 => n470, B2 => n1128, 
                           ZN => n1587);
   U632 : OAI22_X1 port map( A1 => n571, A2 => n1129, B1 => n537, B2 => n1130, 
                           ZN => n1586);
   U633 : OAI22_X1 port map( A1 => n638, A2 => n1131, B1 => n604, B2 => n1132, 
                           ZN => n1585);
   U634 : NOR4_X1 port map( A1 => n1589, A2 => n1591, A3 => n1592, A4 => n1593,
                           ZN => n1578);
   U635 : OAI22_X1 port map( A1 => n705, A2 => n1137, B1 => n672, B2 => n1138, 
                           ZN => n1593);
   U636 : OAI22_X1 port map( A1 => n772, A2 => n1139, B1 => n739, B2 => n1140, 
                           ZN => n1592);
   U637 : OAI22_X1 port map( A1 => n840, A2 => n1, B1 => n806, B2 => n2, ZN => 
                           n1591);
   U638 : OAI22_X1 port map( A1 => n907, A2 => n3, B1 => n873, B2 => n37, ZN =>
                           n1589);
   U639 : NOR4_X1 port map( A1 => n1594, A2 => n1595, A3 => n1596, A4 => n1597,
                           ZN => n1577);
   U640 : OAI22_X1 port map( A1 => n974, A2 => n1149, B1 => n940, B2 => n1151, 
                           ZN => n1597);
   U641 : OAI22_X1 port map( A1 => n1041, A2 => n1152, B1 => n1008, B2 => n1153
                           , ZN => n1596);
   U642 : OAI22_X1 port map( A1 => n71, A2 => n1154, B1 => n1075, B2 => n1155, 
                           ZN => n1595);
   U643 : OAI22_X1 port map( A1 => n156, A2 => n1156, B1 => n120, B2 => n1157, 
                           ZN => n1594);
   U644 : OAI22_X1 port map( A1 => n1598, A2 => n1103, B1 => n1104, B2 => n1590
                           , ZN => N4574);
   U645 : NOR4_X1 port map( A1 => n1603, A2 => n1604, A3 => n1605, A4 => n1606,
                           ZN => n1602);
   U646 : OAI22_X1 port map( A1 => n179, A2 => n1113, B1 => n649, B2 => n1114, 
                           ZN => n1606);
   U647 : OAI22_X1 port map( A1 => n243, A2 => n1115, B1 => n211, B2 => n1116, 
                           ZN => n1605);
   U648 : OAI22_X1 port map( A1 => n307, A2 => n1117, B1 => n275, B2 => n1118, 
                           ZN => n1604);
   U649 : OAI22_X1 port map( A1 => n371, A2 => n1119, B1 => n339, B2 => n1120, 
                           ZN => n1603);
   U650 : NOR4_X1 port map( A1 => n1607, A2 => n1608, A3 => n1609, A4 => n1610,
                           ZN => n1601);
   U651 : OAI22_X1 port map( A1 => n435, A2 => n1125, B1 => n403, B2 => n1126, 
                           ZN => n1610);
   U652 : OAI22_X1 port map( A1 => n503, A2 => n1127, B1 => n469, B2 => n1128, 
                           ZN => n1609);
   U653 : OAI22_X1 port map( A1 => n570, A2 => n1129, B1 => n536, B2 => n1130, 
                           ZN => n1608);
   U654 : OAI22_X1 port map( A1 => n637, A2 => n1131, B1 => n603, B2 => n1132, 
                           ZN => n1607);
   U655 : NOR4_X1 port map( A1 => n1611, A2 => n1613, A3 => n1614, A4 => n1615,
                           ZN => n1600);
   U656 : OAI22_X1 port map( A1 => n704, A2 => n1137, B1 => n671, B2 => n1138, 
                           ZN => n1615);
   U657 : OAI22_X1 port map( A1 => n771, A2 => n1139, B1 => n738, B2 => n1140, 
                           ZN => n1614);
   U658 : OAI22_X1 port map( A1 => n839, A2 => n1, B1 => n805, B2 => n2, ZN => 
                           n1613);
   U659 : OAI22_X1 port map( A1 => n906, A2 => n3, B1 => n872, B2 => n37, ZN =>
                           n1611);
   U660 : NOR4_X1 port map( A1 => n1616, A2 => n1617, A3 => n1618, A4 => n1619,
                           ZN => n1599);
   U661 : OAI22_X1 port map( A1 => n973, A2 => n1149, B1 => n939, B2 => n1151, 
                           ZN => n1619);
   U662 : OAI22_X1 port map( A1 => n1040, A2 => n1152, B1 => n1007, B2 => n1153
                           , ZN => n1618);
   U663 : OAI22_X1 port map( A1 => n69, A2 => n1154, B1 => n1074, B2 => n1155, 
                           ZN => n1617);
   U664 : OAI22_X1 port map( A1 => n155, A2 => n1156, B1 => n119, B2 => n1157, 
                           ZN => n1616);
   U665 : OAI22_X1 port map( A1 => n1620, A2 => n1103, B1 => n1104, B2 => n1612
                           , ZN => N4572);
   U666 : NOR4_X1 port map( A1 => n1625, A2 => n1626, A3 => n1627, A4 => n1628,
                           ZN => n1624);
   U667 : OAI22_X1 port map( A1 => n176, A2 => n1113, B1 => n628, B2 => n1114, 
                           ZN => n1628);
   U668 : OAI22_X1 port map( A1 => n242, A2 => n1115, B1 => n210, B2 => n1116, 
                           ZN => n1627);
   U669 : OAI22_X1 port map( A1 => n306, A2 => n1117, B1 => n274, B2 => n1118, 
                           ZN => n1626);
   U670 : OAI22_X1 port map( A1 => n370, A2 => n1119, B1 => n338, B2 => n1120, 
                           ZN => n1625);
   U671 : NOR4_X1 port map( A1 => n1629, A2 => n1630, A3 => n1631, A4 => n1632,
                           ZN => n1623);
   U672 : OAI22_X1 port map( A1 => n434, A2 => n1125, B1 => n402, B2 => n1126, 
                           ZN => n1632);
   U673 : OAI22_X1 port map( A1 => n501, A2 => n1127, B1 => n468, B2 => n1128, 
                           ZN => n1631);
   U674 : OAI22_X1 port map( A1 => n569, A2 => n1129, B1 => n535, B2 => n1130, 
                           ZN => n1630);
   U675 : OAI22_X1 port map( A1 => n636, A2 => n1131, B1 => n602, B2 => n1132, 
                           ZN => n1629);
   U676 : NOR4_X1 port map( A1 => n1633, A2 => n1635, A3 => n1636, A4 => n1637,
                           ZN => n1622);
   U677 : OAI22_X1 port map( A1 => n703, A2 => n1137, B1 => n669, B2 => n1138, 
                           ZN => n1637);
   U678 : OAI22_X1 port map( A1 => n770, A2 => n1139, B1 => n737, B2 => n1140, 
                           ZN => n1636);
   U679 : OAI22_X1 port map( A1 => n837, A2 => n1, B1 => n804, B2 => n2, ZN => 
                           n1635);
   U680 : OAI22_X1 port map( A1 => n905, A2 => n3, B1 => n871, B2 => n37, ZN =>
                           n1633);
   U681 : NOR4_X1 port map( A1 => n1638, A2 => n1639, A3 => n1640, A4 => n1641,
                           ZN => n1621);
   U682 : OAI22_X1 port map( A1 => n972, A2 => n1149, B1 => n938, B2 => n1151, 
                           ZN => n1641);
   U683 : OAI22_X1 port map( A1 => n1039, A2 => n1152, B1 => n1005, B2 => n1153
                           , ZN => n1640);
   U684 : OAI22_X1 port map( A1 => n67, A2 => n1154, B1 => n1073, B2 => n1155, 
                           ZN => n1639);
   U685 : OAI22_X1 port map( A1 => n153, A2 => n1156, B1 => n118, B2 => n1157, 
                           ZN => n1638);
   U686 : OAI22_X1 port map( A1 => n1642, A2 => n1103, B1 => n1104, B2 => n1634
                           , ZN => N4570);
   U687 : NOR4_X1 port map( A1 => n1647, A2 => n1648, A3 => n1649, A4 => n1650,
                           ZN => n1646);
   U688 : OAI22_X1 port map( A1 => n165, A2 => n1113, B1 => n607, B2 => n1114, 
                           ZN => n1650);
   U689 : OAI22_X1 port map( A1 => n241, A2 => n1115, B1 => n209, B2 => n1116, 
                           ZN => n1649);
   U690 : OAI22_X1 port map( A1 => n305, A2 => n1117, B1 => n273, B2 => n1118, 
                           ZN => n1648);
   U691 : OAI22_X1 port map( A1 => n369, A2 => n1119, B1 => n337, B2 => n1120, 
                           ZN => n1647);
   U692 : NOR4_X1 port map( A1 => n1651, A2 => n1652, A3 => n1653, A4 => n1654,
                           ZN => n1645);
   U693 : OAI22_X1 port map( A1 => n433, A2 => n1125, B1 => n401, B2 => n1126, 
                           ZN => n1654);
   U694 : OAI22_X1 port map( A1 => n500, A2 => n1127, B1 => n467, B2 => n1128, 
                           ZN => n1653);
   U695 : OAI22_X1 port map( A1 => n568, A2 => n1129, B1 => n534, B2 => n1130, 
                           ZN => n1652);
   U696 : OAI22_X1 port map( A1 => n635, A2 => n1131, B1 => n601, B2 => n1132, 
                           ZN => n1651);
   U697 : NOR4_X1 port map( A1 => n1655, A2 => n1657, A3 => n1658, A4 => n1659,
                           ZN => n1644);
   U698 : OAI22_X1 port map( A1 => n702, A2 => n1137, B1 => n668, B2 => n1138, 
                           ZN => n1659);
   U699 : OAI22_X1 port map( A1 => n769, A2 => n1139, B1 => n736, B2 => n1140, 
                           ZN => n1658);
   U700 : OAI22_X1 port map( A1 => n836, A2 => n1, B1 => n803, B2 => n2, ZN => 
                           n1657);
   U701 : OAI22_X1 port map( A1 => n904, A2 => n3, B1 => n870, B2 => n37, ZN =>
                           n1655);
   U702 : NOR4_X1 port map( A1 => n1660, A2 => n1661, A3 => n1662, A4 => n1663,
                           ZN => n1643);
   U703 : OAI22_X1 port map( A1 => n971, A2 => n1149, B1 => n937, B2 => n1151, 
                           ZN => n1663);
   U704 : OAI22_X1 port map( A1 => n1038, A2 => n1152, B1 => n1004, B2 => n1153
                           , ZN => n1662);
   U705 : OAI22_X1 port map( A1 => n65, A2 => n1154, B1 => n1072, B2 => n1155, 
                           ZN => n1661);
   U706 : OAI22_X1 port map( A1 => n152, A2 => n1156, B1 => n117, B2 => n1157, 
                           ZN => n1660);
   U707 : OAI22_X1 port map( A1 => n1664, A2 => n1103, B1 => n1104, B2 => n1656
                           , ZN => N4568);
   U708 : NOR4_X1 port map( A1 => n1669, A2 => n1670, A3 => n1671, A4 => n1672,
                           ZN => n1668);
   U709 : OAI22_X1 port map( A1 => n154, A2 => n1113, B1 => n586, B2 => n1114, 
                           ZN => n1672);
   U710 : OAI22_X1 port map( A1 => n240, A2 => n1115, B1 => n208, B2 => n1116, 
                           ZN => n1671);
   U711 : OAI22_X1 port map( A1 => n304, A2 => n1117, B1 => n272, B2 => n1118, 
                           ZN => n1670);
   U712 : OAI22_X1 port map( A1 => n368, A2 => n1119, B1 => n336, B2 => n1120, 
                           ZN => n1669);
   U713 : NOR4_X1 port map( A1 => n1673, A2 => n1674, A3 => n1675, A4 => n1676,
                           ZN => n1667);
   U714 : OAI22_X1 port map( A1 => n432, A2 => n1125, B1 => n400, B2 => n1126, 
                           ZN => n1676);
   U715 : OAI22_X1 port map( A1 => n499, A2 => n1127, B1 => n466, B2 => n1128, 
                           ZN => n1675);
   U716 : OAI22_X1 port map( A1 => n567, A2 => n1129, B1 => n533, B2 => n1130, 
                           ZN => n1674);
   U717 : OAI22_X1 port map( A1 => n634, A2 => n1131, B1 => n600, B2 => n1132, 
                           ZN => n1673);
   U718 : NOR4_X1 port map( A1 => n1677, A2 => n1679, A3 => n1680, A4 => n1681,
                           ZN => n1666);
   U719 : OAI22_X1 port map( A1 => n701, A2 => n1137, B1 => n667, B2 => n1138, 
                           ZN => n1681);
   U720 : OAI22_X1 port map( A1 => n768, A2 => n1139, B1 => n735, B2 => n1140, 
                           ZN => n1680);
   U721 : OAI22_X1 port map( A1 => n835, A2 => n1, B1 => n802, B2 => n2, ZN => 
                           n1679);
   U722 : OAI22_X1 port map( A1 => n903, A2 => n3, B1 => n869, B2 => n37, ZN =>
                           n1677);
   U723 : NOR4_X1 port map( A1 => n1682, A2 => n1683, A3 => n1684, A4 => n1685,
                           ZN => n1665);
   U724 : OAI22_X1 port map( A1 => n970, A2 => n1149, B1 => n936, B2 => n1151, 
                           ZN => n1685);
   U725 : OAI22_X1 port map( A1 => n1037, A2 => n1152, B1 => n1003, B2 => n1153
                           , ZN => n1684);
   U726 : OAI22_X1 port map( A1 => n63, A2 => n1154, B1 => n1071, B2 => n1155, 
                           ZN => n1683);
   U727 : OAI22_X1 port map( A1 => n151, A2 => n1156, B1 => n116, B2 => n1157, 
                           ZN => n1682);
   U728 : OAI22_X1 port map( A1 => n1686, A2 => n1103, B1 => n1104, B2 => n1678
                           , ZN => N4566);
   U729 : NOR4_X1 port map( A1 => n1691, A2 => n1692, A3 => n1693, A4 => n1694,
                           ZN => n1690);
   U730 : OAI22_X1 port map( A1 => n143, A2 => n1113, B1 => n565, B2 => n1114, 
                           ZN => n1694);
   U731 : OAI22_X1 port map( A1 => n239, A2 => n1115, B1 => n207, B2 => n1116, 
                           ZN => n1693);
   U732 : OAI22_X1 port map( A1 => n303, A2 => n1117, B1 => n271, B2 => n1118, 
                           ZN => n1692);
   U733 : OAI22_X1 port map( A1 => n367, A2 => n1119, B1 => n335, B2 => n1120, 
                           ZN => n1691);
   U734 : NOR4_X1 port map( A1 => n1695, A2 => n1696, A3 => n1697, A4 => n1698,
                           ZN => n1689);
   U735 : OAI22_X1 port map( A1 => n431, A2 => n1125, B1 => n399, B2 => n1126, 
                           ZN => n1698);
   U736 : OAI22_X1 port map( A1 => n498, A2 => n1127, B1 => n465, B2 => n1128, 
                           ZN => n1697);
   U737 : OAI22_X1 port map( A1 => n566, A2 => n1129, B1 => n532, B2 => n1130, 
                           ZN => n1696);
   U738 : OAI22_X1 port map( A1 => n633, A2 => n1131, B1 => n599, B2 => n1132, 
                           ZN => n1695);
   U739 : NOR4_X1 port map( A1 => n1699, A2 => n1701, A3 => n1702, A4 => n1703,
                           ZN => n1688);
   U740 : OAI22_X1 port map( A1 => n700, A2 => n1137, B1 => n666, B2 => n1138, 
                           ZN => n1703);
   U741 : OAI22_X1 port map( A1 => n767, A2 => n1139, B1 => n734, B2 => n1140, 
                           ZN => n1702);
   U742 : OAI22_X1 port map( A1 => n834, A2 => n1, B1 => n801, B2 => n2, ZN => 
                           n1701);
   U743 : OAI22_X1 port map( A1 => n902, A2 => n3, B1 => n868, B2 => n37, ZN =>
                           n1699);
   U744 : NOR4_X1 port map( A1 => n1704, A2 => n1705, A3 => n1706, A4 => n1707,
                           ZN => n1687);
   U745 : OAI22_X1 port map( A1 => n969, A2 => n1149, B1 => n935, B2 => n1151, 
                           ZN => n1707);
   U746 : OAI22_X1 port map( A1 => n1036, A2 => n1152, B1 => n1002, B2 => n1153
                           , ZN => n1706);
   U747 : OAI22_X1 port map( A1 => n61, A2 => n1154, B1 => n1070, B2 => n1155, 
                           ZN => n1705);
   U748 : OAI22_X1 port map( A1 => n150, A2 => n1156, B1 => n115, B2 => n1157, 
                           ZN => n1704);
   U749 : OAI22_X1 port map( A1 => n1708, A2 => n1103, B1 => n1104, B2 => n1700
                           , ZN => N4564);
   U750 : NOR4_X1 port map( A1 => n1713, A2 => n1714, A3 => n1715, A4 => n1716,
                           ZN => n1712);
   U751 : OAI22_X1 port map( A1 => n132, A2 => n1113, B1 => n544, B2 => n1114, 
                           ZN => n1716);
   U752 : OAI22_X1 port map( A1 => n238, A2 => n1115, B1 => n206, B2 => n1116, 
                           ZN => n1715);
   U753 : OAI22_X1 port map( A1 => n302, A2 => n1117, B1 => n270, B2 => n1118, 
                           ZN => n1714);
   U754 : OAI22_X1 port map( A1 => n366, A2 => n1119, B1 => n334, B2 => n1120, 
                           ZN => n1713);
   U755 : NOR4_X1 port map( A1 => n1717, A2 => n1718, A3 => n1719, A4 => n1720,
                           ZN => n1711);
   U756 : OAI22_X1 port map( A1 => n430, A2 => n1125, B1 => n398, B2 => n1126, 
                           ZN => n1720);
   U757 : OAI22_X1 port map( A1 => n497, A2 => n1127, B1 => n464, B2 => n1128, 
                           ZN => n1719);
   U758 : OAI22_X1 port map( A1 => n564, A2 => n1129, B1 => n531, B2 => n1130, 
                           ZN => n1718);
   U759 : OAI22_X1 port map( A1 => n632, A2 => n1131, B1 => n598, B2 => n1132, 
                           ZN => n1717);
   U760 : NOR4_X1 port map( A1 => n1721, A2 => n1723, A3 => n1724, A4 => n1725,
                           ZN => n1710);
   U761 : OAI22_X1 port map( A1 => n699, A2 => n1137, B1 => n665, B2 => n1138, 
                           ZN => n1725);
   U762 : OAI22_X1 port map( A1 => n766, A2 => n1139, B1 => n732, B2 => n1140, 
                           ZN => n1724);
   U763 : OAI22_X1 port map( A1 => n833, A2 => n1, B1 => n800, B2 => n2, ZN => 
                           n1723);
   U764 : OAI22_X1 port map( A1 => n900, A2 => n3, B1 => n867, B2 => n37, ZN =>
                           n1721);
   U765 : NOR4_X1 port map( A1 => n1726, A2 => n1727, A3 => n1728, A4 => n1729,
                           ZN => n1709);
   U766 : OAI22_X1 port map( A1 => n968, A2 => n1149, B1 => n934, B2 => n1151, 
                           ZN => n1729);
   U767 : OAI22_X1 port map( A1 => n1035, A2 => n1152, B1 => n1001, B2 => n1153
                           , ZN => n1728);
   U768 : OAI22_X1 port map( A1 => n59, A2 => n1154, B1 => n1068, B2 => n1155, 
                           ZN => n1727);
   U769 : OAI22_X1 port map( A1 => n149, A2 => n1156, B1 => n114, B2 => n1157, 
                           ZN => n1726);
   U770 : OAI22_X1 port map( A1 => n1730, A2 => n1103, B1 => n1104, B2 => n1722
                           , ZN => N4562);
   U771 : NOR4_X1 port map( A1 => n1735, A2 => n1736, A3 => n1737, A4 => n1738,
                           ZN => n1734);
   U772 : OAI22_X1 port map( A1 => n121, A2 => n1113, B1 => n523, B2 => n1114, 
                           ZN => n1738);
   U773 : OAI22_X1 port map( A1 => n237, A2 => n1115, B1 => n205, B2 => n1116, 
                           ZN => n1737);
   U774 : OAI22_X1 port map( A1 => n301, A2 => n1117, B1 => n269, B2 => n1118, 
                           ZN => n1736);
   U775 : OAI22_X1 port map( A1 => n365, A2 => n1119, B1 => n333, B2 => n1120, 
                           ZN => n1735);
   U776 : NOR4_X1 port map( A1 => n1739, A2 => n1740, A3 => n1741, A4 => n1742,
                           ZN => n1733);
   U777 : OAI22_X1 port map( A1 => n429, A2 => n1125, B1 => n397, B2 => n1126, 
                           ZN => n1742);
   U778 : OAI22_X1 port map( A1 => n496, A2 => n1127, B1 => n463, B2 => n1128, 
                           ZN => n1741);
   U779 : OAI22_X1 port map( A1 => n563, A2 => n1129, B1 => n530, B2 => n1130, 
                           ZN => n1740);
   U780 : OAI22_X1 port map( A1 => n631, A2 => n1131, B1 => n597, B2 => n1132, 
                           ZN => n1739);
   U781 : NOR4_X1 port map( A1 => n1743, A2 => n1745, A3 => n1746, A4 => n1747,
                           ZN => n1732);
   U782 : OAI22_X1 port map( A1 => n698, A2 => n1137, B1 => n664, B2 => n1138, 
                           ZN => n1747);
   U783 : OAI22_X1 port map( A1 => n765, A2 => n1139, B1 => n731, B2 => n1140, 
                           ZN => n1746);
   U784 : OAI22_X1 port map( A1 => n832, A2 => n1, B1 => n799, B2 => n2, ZN => 
                           n1745);
   U785 : OAI22_X1 port map( A1 => n899, A2 => n3, B1 => n866, B2 => n37, ZN =>
                           n1743);
   U786 : NOR4_X1 port map( A1 => n1748, A2 => n1749, A3 => n1750, A4 => n1751,
                           ZN => n1731);
   U787 : OAI22_X1 port map( A1 => n967, A2 => n1149, B1 => n933, B2 => n1151, 
                           ZN => n1751);
   U788 : OAI22_X1 port map( A1 => n1034, A2 => n1152, B1 => n1000, B2 => n1153
                           , ZN => n1750);
   U789 : OAI22_X1 port map( A1 => n57, A2 => n1154, B1 => n1067, B2 => n1155, 
                           ZN => n1749);
   U790 : OAI22_X1 port map( A1 => n148, A2 => n1156, B1 => n113, B2 => n1157, 
                           ZN => n1748);
   U791 : OAI22_X1 port map( A1 => n1752, A2 => n1103, B1 => n1744, B2 => n1104
                           , ZN => N4560);
   U792 : NOR4_X1 port map( A1 => n1753, A2 => n1754, A3 => n1755, A4 => n1756,
                           ZN => n1752);
   U793 : OAI211_X1 port map( C1 => n1101, C2 => n1154, A => n1757, B => n1758,
                           ZN => n1756);
   U794 : NOR4_X1 port map( A1 => n1759, A2 => n1760, A3 => n1761, A4 => n1762,
                           ZN => n1758);
   U795 : OAI22_X1 port map( A1 => n110, A2 => n1113, B1 => n204, B2 => n1116, 
                           ZN => n1762);
   U796 : OAI22_X1 port map( A1 => n236, A2 => n1115, B1 => n268, B2 => n1118, 
                           ZN => n1761);
   U797 : OAI22_X1 port map( A1 => n300, A2 => n1117, B1 => n332, B2 => n1120, 
                           ZN => n1760);
   U798 : OAI22_X1 port map( A1 => n364, A2 => n1119, B1 => n396, B2 => n1126, 
                           ZN => n1759);
   U799 : NOR4_X1 port map( A1 => n1763, A2 => n1764, A3 => n1765, A4 => n1767,
                           ZN => n1757);
   U800 : OAI22_X1 port map( A1 => n428, A2 => n1125, B1 => n462, B2 => n1128, 
                           ZN => n1767);
   U801 : OAI22_X1 port map( A1 => n495, A2 => n1127, B1 => n529, B2 => n1130, 
                           ZN => n1765);
   U802 : OAI22_X1 port map( A1 => n562, A2 => n1129, B1 => n596, B2 => n1132, 
                           ZN => n1764);
   U803 : OAI22_X1 port map( A1 => n630, A2 => n1131, B1 => n663, B2 => n1138, 
                           ZN => n1763);
   U804 : OAI211_X1 port map( C1 => n147, C2 => n1156, A => n1768, B => n1769, 
                           ZN => n1755);
   U805 : NOR4_X1 port map( A1 => n1770, A2 => n1771, A3 => n1772, A4 => n1773,
                           ZN => n1769);
   U806 : OAI22_X1 port map( A1 => n764, A2 => n1139, B1 => n798, B2 => n2, ZN 
                           => n1773);
   U807 : OAI22_X1 port map( A1 => n697, A2 => n1137, B1 => n730, B2 => n1140, 
                           ZN => n1772);
   U808 : OAI22_X1 port map( A1 => n898, A2 => n3, B1 => n932, B2 => n1151, ZN 
                           => n1771);
   U809 : OAI22_X1 port map( A1 => n831, A2 => n1, B1 => n865, B2 => n37, ZN =>
                           n1770);
   U810 : OAI22_X1 port map( A1 => n1114, A2 => n502, B1 => n1157, B2 => n112, 
                           ZN => n1774);
   U811 : OAI22_X1 port map( A1 => n1033, A2 => n1152, B1 => n1066, B2 => n1155
                           , ZN => n1754);
   U812 : OAI22_X1 port map( A1 => n966, A2 => n1149, B1 => n999, B2 => n1153, 
                           ZN => n1753);
   U813 : OAI22_X1 port map( A1 => n1775, A2 => n1103, B1 => n1104, B2 => n1766
                           , ZN => N4558);
   U814 : NOR4_X1 port map( A1 => n1780, A2 => n1781, A3 => n1782, A4 => n1783,
                           ZN => n1779);
   U815 : OAI22_X1 port map( A1 => n99, A2 => n1113, B1 => n481, B2 => n1114, 
                           ZN => n1783);
   U816 : OAI22_X1 port map( A1 => n235, A2 => n1115, B1 => n203, B2 => n1116, 
                           ZN => n1782);
   U817 : OAI22_X1 port map( A1 => n299, A2 => n1117, B1 => n267, B2 => n1118, 
                           ZN => n1781);
   U818 : OAI22_X1 port map( A1 => n363, A2 => n1119, B1 => n331, B2 => n1120, 
                           ZN => n1780);
   U819 : NOR4_X1 port map( A1 => n1784, A2 => n1785, A3 => n1786, A4 => n1787,
                           ZN => n1778);
   U820 : OAI22_X1 port map( A1 => n427, A2 => n1125, B1 => n395, B2 => n1126, 
                           ZN => n1787);
   U821 : OAI22_X1 port map( A1 => n494, A2 => n1127, B1 => n461, B2 => n1128, 
                           ZN => n1786);
   U822 : OAI22_X1 port map( A1 => n561, A2 => n1129, B1 => n528, B2 => n1130, 
                           ZN => n1785);
   U823 : OAI22_X1 port map( A1 => n629, A2 => n1131, B1 => n595, B2 => n1132, 
                           ZN => n1784);
   U824 : NOR4_X1 port map( A1 => n1789, A2 => n1790, A3 => n1791, A4 => n1792,
                           ZN => n1777);
   U825 : OAI22_X1 port map( A1 => n696, A2 => n1137, B1 => n662, B2 => n1138, 
                           ZN => n1792);
   U826 : OAI22_X1 port map( A1 => n763, A2 => n1139, B1 => n729, B2 => n1140, 
                           ZN => n1791);
   U827 : OAI22_X1 port map( A1 => n830, A2 => n1, B1 => n797, B2 => n2, ZN => 
                           n1790);
   U828 : OAI22_X1 port map( A1 => n897, A2 => n3, B1 => n864, B2 => n37, ZN =>
                           n1789);
   U829 : NOR4_X1 port map( A1 => n1793, A2 => n1794, A3 => n1795, A4 => n1796,
                           ZN => n1776);
   U830 : OAI22_X1 port map( A1 => n965, A2 => n1149, B1 => n931, B2 => n1151, 
                           ZN => n1796);
   U831 : OAI22_X1 port map( A1 => n1032, A2 => n1152, B1 => n998, B2 => n1153,
                           ZN => n1795);
   U832 : OAI22_X1 port map( A1 => n1100, A2 => n1154, B1 => n1065, B2 => n1155
                           , ZN => n1794);
   U833 : OAI22_X1 port map( A1 => n146, A2 => n1156, B1 => n111, B2 => n1157, 
                           ZN => n1793);
   U834 : OAI22_X1 port map( A1 => n1797, A2 => n1103, B1 => n1104, B2 => n1788
                           , ZN => N4556);
   U835 : NOR4_X1 port map( A1 => n1802, A2 => n1803, A3 => n1804, A4 => n1805,
                           ZN => n1801);
   U836 : OAI22_X1 port map( A1 => n77, A2 => n1113, B1 => n460, B2 => n1114, 
                           ZN => n1805);
   U837 : OAI22_X1 port map( A1 => n234, A2 => n1115, B1 => n202, B2 => n1116, 
                           ZN => n1804);
   U838 : OAI22_X1 port map( A1 => n298, A2 => n1117, B1 => n266, B2 => n1118, 
                           ZN => n1803);
   U839 : OAI22_X1 port map( A1 => n362, A2 => n1119, B1 => n330, B2 => n1120, 
                           ZN => n1802);
   U840 : NOR4_X1 port map( A1 => n1806, A2 => n1807, A3 => n1808, A4 => n1809,
                           ZN => n1800);
   U841 : OAI22_X1 port map( A1 => n426, A2 => n1125, B1 => n394, B2 => n1126, 
                           ZN => n1809);
   U842 : OAI22_X1 port map( A1 => n493, A2 => n1127, B1 => n459, B2 => n1128, 
                           ZN => n1808);
   U843 : OAI22_X1 port map( A1 => n560, A2 => n1129, B1 => n527, B2 => n1130, 
                           ZN => n1807);
   U844 : OAI22_X1 port map( A1 => n627, A2 => n1131, B1 => n594, B2 => n1132, 
                           ZN => n1806);
   U845 : NOR4_X1 port map( A1 => n1811, A2 => n1812, A3 => n1813, A4 => n1814,
                           ZN => n1799);
   U846 : OAI22_X1 port map( A1 => n695, A2 => n1137, B1 => n661, B2 => n1138, 
                           ZN => n1814);
   U847 : OAI22_X1 port map( A1 => n762, A2 => n1139, B1 => n728, B2 => n1140, 
                           ZN => n1813);
   U848 : OAI22_X1 port map( A1 => n829, A2 => n1, B1 => n795, B2 => n2, ZN => 
                           n1812);
   U849 : OAI22_X1 port map( A1 => n896, A2 => n3, B1 => n863, B2 => n37, ZN =>
                           n1811);
   U850 : NOR4_X1 port map( A1 => n1815, A2 => n1816, A3 => n1817, A4 => n1818,
                           ZN => n1798);
   U851 : OAI22_X1 port map( A1 => n963, A2 => n1149, B1 => n930, B2 => n1151, 
                           ZN => n1818);
   U852 : OAI22_X1 port map( A1 => n1031, A2 => n1152, B1 => n997, B2 => n1153,
                           ZN => n1817);
   U853 : OAI22_X1 port map( A1 => n1099, A2 => n1154, B1 => n1064, B2 => n1155
                           , ZN => n1816);
   U854 : OAI22_X1 port map( A1 => n145, A2 => n1156, B1 => n109, B2 => n1157, 
                           ZN => n1815);
   U855 : OAI22_X1 port map( A1 => n1819, A2 => n1103, B1 => n1104, B2 => n1810
                           , ZN => N4554);
   U856 : OAI221_X1 port map( B1 => n1826, B2 => ADD_RD2(2), C1 => n1827, C2 =>
                           ADD_RD2(0), A => n1828, ZN => n1825);
   U857 : AOI22_X1 port map( A1 => n1826, A2 => ADD_RD2(2), B1 => n1827, B2 => 
                           ADD_RD2(0), ZN => n1828);
   U858 : AOI221_X1 port map( B1 => n1829, B2 => ADD_WR(4), C1 => n1830, C2 => 
                           ADD_RD2(3), A => n1831, ZN => n1821);
   U859 : OAI22_X1 port map( A1 => ADD_WR(4), A2 => n1829, B1 => n1830, B2 => 
                           ADD_RD2(3), ZN => n1831);
   U860 : NOR4_X1 port map( A1 => n1836, A2 => n1837, A3 => n1838, A4 => n1839,
                           ZN => n1835);
   U861 : OAI22_X1 port map( A1 => n55, A2 => n1113, B1 => n439, B2 => n1114, 
                           ZN => n1839);
   U862 : OAI22_X1 port map( A1 => n233, A2 => n1115, B1 => n201, B2 => n1116, 
                           ZN => n1838);
   U863 : OAI22_X1 port map( A1 => n297, A2 => n1117, B1 => n265, B2 => n1118, 
                           ZN => n1837);
   U864 : OAI22_X1 port map( A1 => n361, A2 => n1119, B1 => n329, B2 => n1120, 
                           ZN => n1836);
   U865 : NOR3_X1 port map( A1 => n1829, A2 => n1846, A3 => n1847, ZN => n1841)
                           ;
   U866 : NAND2_X1 port map( A1 => ADD_RD2(4), A2 => ADD_RD2(3), ZN => n1848);
   U867 : NOR4_X1 port map( A1 => n1849, A2 => n1850, A3 => n1851, A4 => n1852,
                           ZN => n1834);
   U868 : OAI22_X1 port map( A1 => n425, A2 => n1125, B1 => n393, B2 => n1126, 
                           ZN => n1852);
   U869 : OAI22_X1 port map( A1 => n492, A2 => n1127, B1 => n458, B2 => n1128, 
                           ZN => n1851);
   U870 : OAI22_X1 port map( A1 => n559, A2 => n1129, B1 => n526, B2 => n1130, 
                           ZN => n1850);
   U871 : OAI22_X1 port map( A1 => n626, A2 => n1131, B1 => n593, B2 => n1132, 
                           ZN => n1849);
   U872 : NOR3_X1 port map( A1 => ADD_RD2(3), A2 => n1829, A3 => n1847, ZN => 
                           n1853);
   U873 : NOR3_X1 port map( A1 => ADD_RD2(3), A2 => ADD_RD2(0), A3 => n1829, ZN
                           => n1854);
   U874 : NOR4_X1 port map( A1 => n1855, A2 => n1856, A3 => n1857, A4 => n1858,
                           ZN => n1833);
   U875 : OAI22_X1 port map( A1 => n694, A2 => n1137, B1 => n660, B2 => n1138, 
                           ZN => n1858);
   U876 : OAI22_X1 port map( A1 => n761, A2 => n1139, B1 => n727, B2 => n1140, 
                           ZN => n1857);
   U877 : OAI22_X1 port map( A1 => n828, A2 => n1, B1 => n794, B2 => n2, ZN => 
                           n1856);
   U878 : NAND2_X1 port map( A1 => n1844, A2 => n1859, ZN => n1142);
   U879 : NAND2_X1 port map( A1 => n1844, A2 => n1860, ZN => n1141);
   U880 : OAI22_X1 port map( A1 => n895, A2 => n3, B1 => n862, B2 => n37, ZN =>
                           n1855);
   U881 : NAND2_X1 port map( A1 => n1859, A2 => n1845, ZN => n1144);
   U882 : NOR3_X1 port map( A1 => ADD_RD2(4), A2 => n1846, A3 => n1847, ZN => 
                           n1859);
   U883 : NAND2_X1 port map( A1 => n1845, A2 => n1860, ZN => n1143);
   U884 : NOR3_X1 port map( A1 => ADD_RD2(4), A2 => ADD_RD2(0), A3 => n1846, ZN
                           => n1860);
   U885 : NOR4_X1 port map( A1 => n1861, A2 => n1862, A3 => n1863, A4 => n1864,
                           ZN => n1832);
   U886 : OAI22_X1 port map( A1 => n962, A2 => n1149, B1 => n929, B2 => n1151, 
                           ZN => n1864);
   U887 : OAI22_X1 port map( A1 => n1030, A2 => n1152, B1 => n996, B2 => n1153,
                           ZN => n1863);
   U888 : OAI22_X1 port map( A1 => n1098, A2 => n1154, B1 => n1063, B2 => n1155
                           , ZN => n1862);
   U889 : OAI22_X1 port map( A1 => n144, A2 => n1156, B1 => n108, B2 => n1157, 
                           ZN => n1861);
   U890 : NOR3_X1 port map( A1 => ADD_RD2(4), A2 => ADD_RD2(3), A3 => n1847, ZN
                           => n1865);
   U891 : NOR3_X1 port map( A1 => ADD_RD2(4), A2 => ADD_RD2(3), A3 => 
                           ADD_RD2(0), ZN => n1866);
   U892 : OAI22_X1 port map( A1 => n1867, A2 => n1868, B1 => n1869, B2 => n1094
                           , ZN => N4552);
   U893 : NOR4_X1 port map( A1 => n1874, A2 => n1875, A3 => n1876, A4 => n1877,
                           ZN => n1873);
   U894 : OAI22_X1 port map( A1 => n200, A2 => n1878, B1 => n1090, B2 => n1879,
                           ZN => n1877);
   U895 : OAI22_X1 port map( A1 => n264, A2 => n1880, B1 => n232, B2 => n1881, 
                           ZN => n1876);
   U896 : OAI22_X1 port map( A1 => n328, A2 => n1882, B1 => n296, B2 => n1883, 
                           ZN => n1875);
   U897 : OAI22_X1 port map( A1 => n392, A2 => n1884, B1 => n360, B2 => n1885, 
                           ZN => n1874);
   U898 : NOR4_X1 port map( A1 => n1886, A2 => n1887, A3 => n1888, A4 => n1889,
                           ZN => n1872);
   U899 : OAI22_X1 port map( A1 => n457, A2 => n1890, B1 => n424, B2 => n1891, 
                           ZN => n1889);
   U900 : OAI22_X1 port map( A1 => n525, A2 => n1892, B1 => n491, B2 => n1893, 
                           ZN => n1888);
   U901 : OAI22_X1 port map( A1 => n592, A2 => n1894, B1 => n558, B2 => n1895, 
                           ZN => n1887);
   U902 : OAI22_X1 port map( A1 => n659, A2 => n1896, B1 => n625, B2 => n1897, 
                           ZN => n1886);
   U903 : NOR4_X1 port map( A1 => n1898, A2 => n1899, A3 => n1900, A4 => n1901,
                           ZN => n1871);
   U904 : OAI22_X1 port map( A1 => n726, A2 => n1902, B1 => n693, B2 => n1903, 
                           ZN => n1901);
   U905 : OAI22_X1 port map( A1 => n793, A2 => n1904, B1 => n760, B2 => n1905, 
                           ZN => n1900);
   U906 : OAI22_X1 port map( A1 => n861, A2 => n1906, B1 => n827, B2 => n1907, 
                           ZN => n1899);
   U907 : OAI22_X1 port map( A1 => n928, A2 => n1908, B1 => n894, B2 => n1909, 
                           ZN => n1898);
   U908 : NOR4_X1 port map( A1 => n1910, A2 => n1911, A3 => n1912, A4 => n1913,
                           ZN => n1870);
   U909 : OAI22_X1 port map( A1 => n995, A2 => n1914, B1 => n961, B2 => n1915, 
                           ZN => n1913);
   U910 : OAI22_X1 port map( A1 => n1062, A2 => n1916, B1 => n1029, B2 => n1917
                           , ZN => n1912);
   U911 : OAI22_X1 port map( A1 => n107, A2 => n1918, B1 => n1097, B2 => n1919,
                           ZN => n1911);
   U912 : OAI22_X1 port map( A1 => n178, A2 => n1920, B1 => n142, B2 => n1921, 
                           ZN => n1910);
   U913 : OAI22_X1 port map( A1 => n1922, A2 => n1868, B1 => n1869, B2 => n1150
                           , ZN => N4550);
   U914 : NOR4_X1 port map( A1 => n1927, A2 => n1928, A3 => n1929, A4 => n1930,
                           ZN => n1926);
   U915 : OAI22_X1 port map( A1 => n199, A2 => n1878, B1 => n1069, B2 => n1879,
                           ZN => n1930);
   U916 : OAI22_X1 port map( A1 => n263, A2 => n1880, B1 => n231, B2 => n1881, 
                           ZN => n1929);
   U917 : OAI22_X1 port map( A1 => n327, A2 => n39, B1 => n295, B2 => n1883, ZN
                           => n1928);
   U918 : OAI22_X1 port map( A1 => n391, A2 => n43, B1 => n359, B2 => n1885, ZN
                           => n1927);
   U919 : NOR4_X1 port map( A1 => n1931, A2 => n1932, A3 => n1933, A4 => n1934,
                           ZN => n1925);
   U920 : OAI22_X1 port map( A1 => n456, A2 => n1890, B1 => n423, B2 => n1891, 
                           ZN => n1934);
   U921 : OAI22_X1 port map( A1 => n524, A2 => n1892, B1 => n490, B2 => n1893, 
                           ZN => n1933);
   U922 : OAI22_X1 port map( A1 => n591, A2 => n1894, B1 => n557, B2 => n1895, 
                           ZN => n1932);
   U923 : OAI22_X1 port map( A1 => n658, A2 => n1896, B1 => n624, B2 => n1897, 
                           ZN => n1931);
   U924 : NOR4_X1 port map( A1 => n1935, A2 => n1936, A3 => n1937, A4 => n1938,
                           ZN => n1924);
   U925 : OAI22_X1 port map( A1 => n725, A2 => n1902, B1 => n692, B2 => n1903, 
                           ZN => n1938);
   U926 : OAI22_X1 port map( A1 => n792, A2 => n1904, B1 => n759, B2 => n1905, 
                           ZN => n1937);
   U927 : OAI22_X1 port map( A1 => n860, A2 => n1906, B1 => n826, B2 => n1907, 
                           ZN => n1936);
   U928 : OAI22_X1 port map( A1 => n927, A2 => n1908, B1 => n893, B2 => n1909, 
                           ZN => n1935);
   U929 : NOR4_X1 port map( A1 => n1939, A2 => n1940, A3 => n1941, A4 => n1942,
                           ZN => n1923);
   U930 : OAI22_X1 port map( A1 => n994, A2 => n1914, B1 => n960, B2 => n1915, 
                           ZN => n1942);
   U931 : OAI22_X1 port map( A1 => n1061, A2 => n1916, B1 => n1028, B2 => n1917
                           , ZN => n1941);
   U932 : OAI22_X1 port map( A1 => n106, A2 => n1918, B1 => n1096, B2 => n1919,
                           ZN => n1940);
   U933 : OAI22_X1 port map( A1 => n177, A2 => n1920, B1 => n141, B2 => n1921, 
                           ZN => n1939);
   U934 : OAI22_X1 port map( A1 => n1943, A2 => n1868, B1 => n1869, B2 => n1172
                           , ZN => N4548);
   U935 : NOR4_X1 port map( A1 => n1948, A2 => n1949, A3 => n1950, A4 => n1951,
                           ZN => n1947);
   U936 : OAI22_X1 port map( A1 => n198, A2 => n1878, B1 => n1048, B2 => n1879,
                           ZN => n1951);
   U937 : OAI22_X1 port map( A1 => n262, A2 => n1880, B1 => n230, B2 => n1881, 
                           ZN => n1950);
   U938 : OAI22_X1 port map( A1 => n326, A2 => n1882, B1 => n294, B2 => n1883, 
                           ZN => n1949);
   U939 : OAI22_X1 port map( A1 => n390, A2 => n1884, B1 => n358, B2 => n1885, 
                           ZN => n1948);
   U940 : NOR4_X1 port map( A1 => n1952, A2 => n1953, A3 => n1954, A4 => n1955,
                           ZN => n1946);
   U941 : OAI22_X1 port map( A1 => n455, A2 => n1890, B1 => n422, B2 => n1891, 
                           ZN => n1955);
   U942 : OAI22_X1 port map( A1 => n522, A2 => n1892, B1 => n489, B2 => n1893, 
                           ZN => n1954);
   U943 : OAI22_X1 port map( A1 => n590, A2 => n1894, B1 => n556, B2 => n1895, 
                           ZN => n1953);
   U944 : OAI22_X1 port map( A1 => n657, A2 => n1896, B1 => n623, B2 => n1897, 
                           ZN => n1952);
   U945 : NOR4_X1 port map( A1 => n1956, A2 => n1957, A3 => n1958, A4 => n1959,
                           ZN => n1945);
   U946 : OAI22_X1 port map( A1 => n724, A2 => n1902, B1 => n690, B2 => n1903, 
                           ZN => n1959);
   U947 : OAI22_X1 port map( A1 => n791, A2 => n1904, B1 => n758, B2 => n1905, 
                           ZN => n1958);
   U948 : OAI22_X1 port map( A1 => n858, A2 => n1906, B1 => n825, B2 => n1907, 
                           ZN => n1957);
   U949 : OAI22_X1 port map( A1 => n926, A2 => n1908, B1 => n892, B2 => n1909, 
                           ZN => n1956);
   U950 : NOR4_X1 port map( A1 => n1960, A2 => n1961, A3 => n1962, A4 => n1963,
                           ZN => n1944);
   U951 : OAI22_X1 port map( A1 => n993, A2 => n1914, B1 => n959, B2 => n1915, 
                           ZN => n1963);
   U952 : OAI22_X1 port map( A1 => n1060, A2 => n1916, B1 => n1026, B2 => n1917
                           , ZN => n1962);
   U953 : OAI22_X1 port map( A1 => n105, A2 => n1918, B1 => n1095, B2 => n1919,
                           ZN => n1961);
   U954 : OAI22_X1 port map( A1 => n175, A2 => n1920, B1 => n140, B2 => n1921, 
                           ZN => n1960);
   U955 : OAI22_X1 port map( A1 => n1964, A2 => n1868, B1 => n1869, B2 => n1194
                           , ZN => N4546);
   U956 : NOR4_X1 port map( A1 => n1969, A2 => n1970, A3 => n1971, A4 => n1972,
                           ZN => n1968);
   U957 : OAI22_X1 port map( A1 => n197, A2 => n1878, B1 => n1027, B2 => n1879,
                           ZN => n1972);
   U958 : OAI22_X1 port map( A1 => n261, A2 => n1880, B1 => n229, B2 => n1881, 
                           ZN => n1971);
   U959 : OAI22_X1 port map( A1 => n325, A2 => n1882, B1 => n293, B2 => n1883, 
                           ZN => n1970);
   U960 : OAI22_X1 port map( A1 => n389, A2 => n1884, B1 => n357, B2 => n1885, 
                           ZN => n1969);
   U961 : NOR4_X1 port map( A1 => n1973, A2 => n1974, A3 => n1975, A4 => n1976,
                           ZN => n1967);
   U962 : OAI22_X1 port map( A1 => n454, A2 => n1890, B1 => n421, B2 => n1891, 
                           ZN => n1976);
   U963 : OAI22_X1 port map( A1 => n521, A2 => n1892, B1 => n488, B2 => n1893, 
                           ZN => n1975);
   U964 : OAI22_X1 port map( A1 => n589, A2 => n1894, B1 => n555, B2 => n1895, 
                           ZN => n1974);
   U965 : OAI22_X1 port map( A1 => n656, A2 => n1896, B1 => n622, B2 => n1897, 
                           ZN => n1973);
   U966 : NOR4_X1 port map( A1 => n1977, A2 => n1978, A3 => n1979, A4 => n1980,
                           ZN => n1966);
   U967 : OAI22_X1 port map( A1 => n723, A2 => n1902, B1 => n689, B2 => n1903, 
                           ZN => n1980);
   U968 : OAI22_X1 port map( A1 => n790, A2 => n1904, B1 => n757, B2 => n1905, 
                           ZN => n1979);
   U969 : OAI22_X1 port map( A1 => n857, A2 => n1906, B1 => n824, B2 => n1907, 
                           ZN => n1978);
   U970 : OAI22_X1 port map( A1 => n925, A2 => n1908, B1 => n891, B2 => n1909, 
                           ZN => n1977);
   U971 : NOR4_X1 port map( A1 => n1981, A2 => n1982, A3 => n1983, A4 => n1984,
                           ZN => n1965);
   U972 : OAI22_X1 port map( A1 => n992, A2 => n1914, B1 => n958, B2 => n1915, 
                           ZN => n1984);
   U973 : OAI22_X1 port map( A1 => n1059, A2 => n1916, B1 => n1025, B2 => n1917
                           , ZN => n1983);
   U974 : OAI22_X1 port map( A1 => n104, A2 => n1918, B1 => n1093, B2 => n1919,
                           ZN => n1982);
   U975 : OAI22_X1 port map( A1 => n174, A2 => n1920, B1 => n139, B2 => n1921, 
                           ZN => n1981);
   U976 : OAI22_X1 port map( A1 => n1985, A2 => n1868, B1 => n1869, B2 => n1216
                           , ZN => N4544);
   U977 : NOR4_X1 port map( A1 => n1990, A2 => n1991, A3 => n1992, A4 => n1993,
                           ZN => n1989);
   U978 : OAI22_X1 port map( A1 => n196, A2 => n1878, B1 => n1006, B2 => n1879,
                           ZN => n1993);
   U979 : OAI22_X1 port map( A1 => n260, A2 => n1880, B1 => n228, B2 => n1881, 
                           ZN => n1992);
   U980 : OAI22_X1 port map( A1 => n324, A2 => n1882, B1 => n292, B2 => n1883, 
                           ZN => n1991);
   U981 : OAI22_X1 port map( A1 => n388, A2 => n1884, B1 => n356, B2 => n1885, 
                           ZN => n1990);
   U982 : NOR4_X1 port map( A1 => n1994, A2 => n1995, A3 => n1996, A4 => n1997,
                           ZN => n1988);
   U983 : OAI22_X1 port map( A1 => n453, A2 => n1890, B1 => n420, B2 => n1891, 
                           ZN => n1997);
   U984 : OAI22_X1 port map( A1 => n520, A2 => n1892, B1 => n487, B2 => n1893, 
                           ZN => n1996);
   U985 : OAI22_X1 port map( A1 => n588, A2 => n1894, B1 => n554, B2 => n1895, 
                           ZN => n1995);
   U986 : OAI22_X1 port map( A1 => n655, A2 => n1896, B1 => n621, B2 => n1897, 
                           ZN => n1994);
   U987 : NOR4_X1 port map( A1 => n1998, A2 => n1999, A3 => n2000, A4 => n2001,
                           ZN => n1987);
   U988 : OAI22_X1 port map( A1 => n722, A2 => n1902, B1 => n688, B2 => n1903, 
                           ZN => n2001);
   U989 : OAI22_X1 port map( A1 => n789, A2 => n1904, B1 => n756, B2 => n1905, 
                           ZN => n2000);
   U990 : OAI22_X1 port map( A1 => n856, A2 => n1906, B1 => n823, B2 => n1907, 
                           ZN => n1999);
   U991 : OAI22_X1 port map( A1 => n924, A2 => n1908, B1 => n890, B2 => n1909, 
                           ZN => n1998);
   U992 : NOR4_X1 port map( A1 => n2002, A2 => n2003, A3 => n2004, A4 => n2005,
                           ZN => n1986);
   U993 : OAI22_X1 port map( A1 => n991, A2 => n1914, B1 => n957, B2 => n1915, 
                           ZN => n2005);
   U994 : OAI22_X1 port map( A1 => n1058, A2 => n1916, B1 => n1024, B2 => n1917
                           , ZN => n2004);
   U995 : OAI22_X1 port map( A1 => n103, A2 => n1918, B1 => n1092, B2 => n1919,
                           ZN => n2003);
   U996 : OAI22_X1 port map( A1 => n173, A2 => n1920, B1 => n138, B2 => n1921, 
                           ZN => n2002);
   U997 : OAI22_X1 port map( A1 => n2006, A2 => n1868, B1 => n1869, B2 => n1238
                           , ZN => N4542);
   U998 : NOR4_X1 port map( A1 => n2011, A2 => n2012, A3 => n2013, A4 => n2014,
                           ZN => n2010);
   U999 : OAI22_X1 port map( A1 => n195, A2 => n1878, B1 => n985, B2 => n1879, 
                           ZN => n2014);
   U1000 : OAI22_X1 port map( A1 => n259, A2 => n1880, B1 => n227, B2 => n1881,
                           ZN => n2013);
   U1001 : OAI22_X1 port map( A1 => n323, A2 => n1882, B1 => n291, B2 => n1883,
                           ZN => n2012);
   U1002 : OAI22_X1 port map( A1 => n387, A2 => n1884, B1 => n355, B2 => n1885,
                           ZN => n2011);
   U1003 : NOR4_X1 port map( A1 => n2015, A2 => n2016, A3 => n2017, A4 => n2018
                           , ZN => n2009);
   U1004 : OAI22_X1 port map( A1 => n452, A2 => n1890, B1 => n419, B2 => n1891,
                           ZN => n2018);
   U1005 : OAI22_X1 port map( A1 => n519, A2 => n1892, B1 => n486, B2 => n1893,
                           ZN => n2017);
   U1006 : OAI22_X1 port map( A1 => n587, A2 => n1894, B1 => n553, B2 => n1895,
                           ZN => n2016);
   U1007 : OAI22_X1 port map( A1 => n654, A2 => n1896, B1 => n620, B2 => n1897,
                           ZN => n2015);
   U1008 : NOR4_X1 port map( A1 => n2019, A2 => n2020, A3 => n2021, A4 => n2022
                           , ZN => n2008);
   U1009 : OAI22_X1 port map( A1 => n721, A2 => n1902, B1 => n687, B2 => n1903,
                           ZN => n2022);
   U1010 : OAI22_X1 port map( A1 => n788, A2 => n1904, B1 => n755, B2 => n1905,
                           ZN => n2021);
   U1011 : OAI22_X1 port map( A1 => n855, A2 => n1906, B1 => n822, B2 => n1907,
                           ZN => n2020);
   U1012 : OAI22_X1 port map( A1 => n923, A2 => n1908, B1 => n889, B2 => n1909,
                           ZN => n2019);
   U1013 : NOR4_X1 port map( A1 => n2023, A2 => n2024, A3 => n2025, A4 => n2026
                           , ZN => n2007);
   U1014 : OAI22_X1 port map( A1 => n990, A2 => n1914, B1 => n956, B2 => n1915,
                           ZN => n2026);
   U1015 : OAI22_X1 port map( A1 => n1057, A2 => n1916, B1 => n1023, B2 => 
                           n1917, ZN => n2025);
   U1016 : OAI22_X1 port map( A1 => n102, A2 => n1918, B1 => n1091, B2 => n1919
                           , ZN => n2024);
   U1017 : OAI22_X1 port map( A1 => n172, A2 => n1920, B1 => n137, B2 => n1921,
                           ZN => n2023);
   U1018 : OAI22_X1 port map( A1 => n2027, A2 => n1868, B1 => n1869, B2 => 
                           n1260, ZN => N4540);
   U1019 : NOR4_X1 port map( A1 => n2032, A2 => n2033, A3 => n2034, A4 => n2035
                           , ZN => n2031);
   U1020 : OAI22_X1 port map( A1 => n194, A2 => n1878, B1 => n964, B2 => n1879,
                           ZN => n2035);
   U1021 : OAI22_X1 port map( A1 => n258, A2 => n1880, B1 => n226, B2 => n1881,
                           ZN => n2034);
   U1022 : OAI22_X1 port map( A1 => n322, A2 => n1882, B1 => n290, B2 => n41, 
                           ZN => n2033);
   U1023 : OAI22_X1 port map( A1 => n386, A2 => n1884, B1 => n354, B2 => n45, 
                           ZN => n2032);
   U1024 : NOR4_X1 port map( A1 => n2036, A2 => n2037, A3 => n2038, A4 => n2039
                           , ZN => n2030);
   U1025 : OAI22_X1 port map( A1 => n451, A2 => n1890, B1 => n418, B2 => n1891,
                           ZN => n2039);
   U1026 : OAI22_X1 port map( A1 => n518, A2 => n1892, B1 => n485, B2 => n1893,
                           ZN => n2038);
   U1027 : OAI22_X1 port map( A1 => n585, A2 => n1894, B1 => n552, B2 => n1895,
                           ZN => n2037);
   U1028 : OAI22_X1 port map( A1 => n653, A2 => n1896, B1 => n619, B2 => n1897,
                           ZN => n2036);
   U1029 : NOR4_X1 port map( A1 => n2040, A2 => n2041, A3 => n2042, A4 => n2043
                           , ZN => n2029);
   U1030 : OAI22_X1 port map( A1 => n720, A2 => n1902, B1 => n686, B2 => n1903,
                           ZN => n2043);
   U1031 : OAI22_X1 port map( A1 => n787, A2 => n1904, B1 => n753, B2 => n1905,
                           ZN => n2042);
   U1032 : OAI22_X1 port map( A1 => n854, A2 => n1906, B1 => n821, B2 => n1907,
                           ZN => n2041);
   U1033 : OAI22_X1 port map( A1 => n921, A2 => n1908, B1 => n888, B2 => n1909,
                           ZN => n2040);
   U1034 : NOR4_X1 port map( A1 => n2044, A2 => n2045, A3 => n2046, A4 => n2047
                           , ZN => n2028);
   U1035 : OAI22_X1 port map( A1 => n989, A2 => n1914, B1 => n955, B2 => n1915,
                           ZN => n2047);
   U1036 : OAI22_X1 port map( A1 => n1056, A2 => n1916, B1 => n1022, B2 => 
                           n1917, ZN => n2046);
   U1037 : OAI22_X1 port map( A1 => n101, A2 => n1918, B1 => n1089, B2 => n1919
                           , ZN => n2045);
   U1038 : OAI22_X1 port map( A1 => n171, A2 => n1920, B1 => n136, B2 => n1921,
                           ZN => n2044);
   U1039 : OAI22_X1 port map( A1 => n2048, A2 => n1868, B1 => n1869, B2 => 
                           n1282, ZN => N4538);
   U1040 : NOR4_X1 port map( A1 => n2053, A2 => n2054, A3 => n2055, A4 => n2056
                           , ZN => n2052);
   U1041 : OAI22_X1 port map( A1 => n193, A2 => n1878, B1 => n943, B2 => n1879,
                           ZN => n2056);
   U1042 : OAI22_X1 port map( A1 => n257, A2 => n1880, B1 => n225, B2 => n1881,
                           ZN => n2055);
   U1043 : OAI22_X1 port map( A1 => n321, A2 => n1882, B1 => n289, B2 => n1883,
                           ZN => n2054);
   U1044 : OAI22_X1 port map( A1 => n385, A2 => n1884, B1 => n353, B2 => n1885,
                           ZN => n2053);
   U1045 : NOR4_X1 port map( A1 => n2057, A2 => n2058, A3 => n2059, A4 => n2060
                           , ZN => n2051);
   U1046 : OAI22_X1 port map( A1 => n450, A2 => n1890, B1 => n417, B2 => n1891,
                           ZN => n2060);
   U1047 : OAI22_X1 port map( A1 => n517, A2 => n1892, B1 => n484, B2 => n1893,
                           ZN => n2059);
   U1048 : OAI22_X1 port map( A1 => n584, A2 => n1894, B1 => n551, B2 => n1895,
                           ZN => n2058);
   U1049 : OAI22_X1 port map( A1 => n652, A2 => n1896, B1 => n618, B2 => n1897,
                           ZN => n2057);
   U1050 : NOR4_X1 port map( A1 => n2061, A2 => n2062, A3 => n2063, A4 => n2064
                           , ZN => n2050);
   U1051 : OAI22_X1 port map( A1 => n719, A2 => n1902, B1 => n685, B2 => n1903,
                           ZN => n2064);
   U1052 : OAI22_X1 port map( A1 => n786, A2 => n1904, B1 => n752, B2 => n1905,
                           ZN => n2063);
   U1053 : OAI22_X1 port map( A1 => n853, A2 => n1906, B1 => n820, B2 => n1907,
                           ZN => n2062);
   U1054 : OAI22_X1 port map( A1 => n920, A2 => n1908, B1 => n887, B2 => n1909,
                           ZN => n2061);
   U1055 : NOR4_X1 port map( A1 => n2065, A2 => n2066, A3 => n2067, A4 => n2068
                           , ZN => n2049);
   U1056 : OAI22_X1 port map( A1 => n988, A2 => n1914, B1 => n954, B2 => n1915,
                           ZN => n2068);
   U1057 : OAI22_X1 port map( A1 => n1055, A2 => n1916, B1 => n1021, B2 => 
                           n1917, ZN => n2067);
   U1058 : OAI22_X1 port map( A1 => n100, A2 => n1918, B1 => n1088, B2 => n1919
                           , ZN => n2066);
   U1059 : OAI22_X1 port map( A1 => n170, A2 => n1920, B1 => n135, B2 => n1921,
                           ZN => n2065);
   U1060 : OAI22_X1 port map( A1 => n2069, A2 => n1868, B1 => n1869, B2 => 
                           n1304, ZN => N4536);
   U1061 : NOR4_X1 port map( A1 => n2074, A2 => n2075, A3 => n2076, A4 => n2077
                           , ZN => n2073);
   U1062 : OAI22_X1 port map( A1 => n192, A2 => n1878, B1 => n922, B2 => n1879,
                           ZN => n2077);
   U1063 : OAI22_X1 port map( A1 => n256, A2 => n1880, B1 => n224, B2 => n1881,
                           ZN => n2076);
   U1064 : OAI22_X1 port map( A1 => n320, A2 => n1882, B1 => n288, B2 => n1883,
                           ZN => n2075);
   U1065 : OAI22_X1 port map( A1 => n384, A2 => n1884, B1 => n352, B2 => n1885,
                           ZN => n2074);
   U1066 : NOR4_X1 port map( A1 => n2078, A2 => n2079, A3 => n2080, A4 => n2081
                           , ZN => n2072);
   U1067 : OAI22_X1 port map( A1 => n449, A2 => n1890, B1 => n416, B2 => n1891,
                           ZN => n2081);
   U1068 : OAI22_X1 port map( A1 => n516, A2 => n1892, B1 => n483, B2 => n1893,
                           ZN => n2080);
   U1069 : OAI22_X1 port map( A1 => n583, A2 => n1894, B1 => n550, B2 => n1895,
                           ZN => n2079);
   U1070 : OAI22_X1 port map( A1 => n651, A2 => n1896, B1 => n617, B2 => n1897,
                           ZN => n2078);
   U1071 : NOR4_X1 port map( A1 => n2082, A2 => n2083, A3 => n2084, A4 => n2085
                           , ZN => n2071);
   U1072 : OAI22_X1 port map( A1 => n718, A2 => n1902, B1 => n684, B2 => n1903,
                           ZN => n2085);
   U1073 : OAI22_X1 port map( A1 => n785, A2 => n1904, B1 => n751, B2 => n1905,
                           ZN => n2084);
   U1074 : OAI22_X1 port map( A1 => n852, A2 => n1906, B1 => n819, B2 => n1907,
                           ZN => n2083);
   U1075 : OAI22_X1 port map( A1 => n919, A2 => n1908, B1 => n886, B2 => n1909,
                           ZN => n2082);
   U1076 : NOR4_X1 port map( A1 => n2086, A2 => n2087, A3 => n2088, A4 => n2089
                           , ZN => n2070);
   U1077 : OAI22_X1 port map( A1 => n987, A2 => n1914, B1 => n953, B2 => n1915,
                           ZN => n2089);
   U1078 : OAI22_X1 port map( A1 => n1054, A2 => n1916, B1 => n1020, B2 => 
                           n1917, ZN => n2088);
   U1079 : OAI22_X1 port map( A1 => n97, A2 => n1918, B1 => n1087, B2 => n1919,
                           ZN => n2087);
   U1080 : OAI22_X1 port map( A1 => n169, A2 => n1920, B1 => n134, B2 => n1921,
                           ZN => n2086);
   U1081 : OAI22_X1 port map( A1 => n2090, A2 => n1868, B1 => n1869, B2 => 
                           n1326, ZN => N4534);
   U1082 : NOR4_X1 port map( A1 => n2095, A2 => n2096, A3 => n2097, A4 => n2098
                           , ZN => n2094);
   U1083 : OAI22_X1 port map( A1 => n191, A2 => n1878, B1 => n901, B2 => n1879,
                           ZN => n2098);
   U1084 : OAI22_X1 port map( A1 => n255, A2 => n1880, B1 => n223, B2 => n1881,
                           ZN => n2097);
   U1085 : OAI22_X1 port map( A1 => n319, A2 => n1882, B1 => n287, B2 => n1883,
                           ZN => n2096);
   U1086 : OAI22_X1 port map( A1 => n383, A2 => n1884, B1 => n351, B2 => n1885,
                           ZN => n2095);
   U1087 : NOR4_X1 port map( A1 => n2099, A2 => n2100, A3 => n2101, A4 => n2102
                           , ZN => n2093);
   U1088 : OAI22_X1 port map( A1 => n448, A2 => n1890, B1 => n415, B2 => n1891,
                           ZN => n2102);
   U1089 : OAI22_X1 port map( A1 => n515, A2 => n1892, B1 => n482, B2 => n1893,
                           ZN => n2101);
   U1090 : OAI22_X1 port map( A1 => n582, A2 => n1894, B1 => n549, B2 => n1895,
                           ZN => n2100);
   U1091 : OAI22_X1 port map( A1 => n650, A2 => n1896, B1 => n616, B2 => n1897,
                           ZN => n2099);
   U1092 : NOR4_X1 port map( A1 => n2103, A2 => n2104, A3 => n2105, A4 => n2106
                           , ZN => n2092);
   U1093 : OAI22_X1 port map( A1 => n717, A2 => n1902, B1 => n683, B2 => n1903,
                           ZN => n2106);
   U1094 : OAI22_X1 port map( A1 => n784, A2 => n1904, B1 => n750, B2 => n1905,
                           ZN => n2105);
   U1095 : OAI22_X1 port map( A1 => n851, A2 => n1906, B1 => n818, B2 => n1907,
                           ZN => n2104);
   U1096 : OAI22_X1 port map( A1 => n918, A2 => n1908, B1 => n885, B2 => n1909,
                           ZN => n2103);
   U1097 : NOR4_X1 port map( A1 => n2107, A2 => n2108, A3 => n2109, A4 => n2110
                           , ZN => n2091);
   U1098 : OAI22_X1 port map( A1 => n986, A2 => n1914, B1 => n952, B2 => n1915,
                           ZN => n2110);
   U1099 : OAI22_X1 port map( A1 => n1053, A2 => n1916, B1 => n1019, B2 => 
                           n1917, ZN => n2109);
   U1100 : OAI22_X1 port map( A1 => n95, A2 => n1918, B1 => n1086, B2 => n1919,
                           ZN => n2108);
   U1101 : OAI22_X1 port map( A1 => n168, A2 => n1920, B1 => n133, B2 => n1921,
                           ZN => n2107);
   U1102 : OAI22_X1 port map( A1 => n2111, A2 => n1868, B1 => n1869, B2 => 
                           n1348, ZN => N4532);
   U1103 : NOR4_X1 port map( A1 => n2116, A2 => n2117, A3 => n2118, A4 => n2119
                           , ZN => n2115);
   U1104 : OAI22_X1 port map( A1 => n190, A2 => n1878, B1 => n880, B2 => n1879,
                           ZN => n2119);
   U1105 : OAI22_X1 port map( A1 => n254, A2 => n1880, B1 => n222, B2 => n1881,
                           ZN => n2118);
   U1106 : OAI22_X1 port map( A1 => n318, A2 => n1882, B1 => n286, B2 => n1883,
                           ZN => n2117);
   U1107 : OAI22_X1 port map( A1 => n382, A2 => n1884, B1 => n350, B2 => n1885,
                           ZN => n2116);
   U1108 : NOR4_X1 port map( A1 => n2120, A2 => n2121, A3 => n2122, A4 => n2123
                           , ZN => n2114);
   U1109 : OAI22_X1 port map( A1 => n447, A2 => n1890, B1 => n414, B2 => n1891,
                           ZN => n2123);
   U1110 : OAI22_X1 port map( A1 => n514, A2 => n1892, B1 => n480, B2 => n1893,
                           ZN => n2122);
   U1111 : OAI22_X1 port map( A1 => n581, A2 => n1894, B1 => n548, B2 => n1895,
                           ZN => n2121);
   U1112 : OAI22_X1 port map( A1 => n648, A2 => n1896, B1 => n615, B2 => n1897,
                           ZN => n2120);
   U1113 : NOR4_X1 port map( A1 => n2124, A2 => n2125, A3 => n2126, A4 => n2127
                           , ZN => n2113);
   U1114 : OAI22_X1 port map( A1 => n716, A2 => n1902, B1 => n682, B2 => n1903,
                           ZN => n2127);
   U1115 : OAI22_X1 port map( A1 => n783, A2 => n1904, B1 => n749, B2 => n1905,
                           ZN => n2126);
   U1116 : OAI22_X1 port map( A1 => n850, A2 => n1906, B1 => n816, B2 => n1907,
                           ZN => n2125);
   U1117 : OAI22_X1 port map( A1 => n917, A2 => n1908, B1 => n884, B2 => n1909,
                           ZN => n2124);
   U1118 : NOR4_X1 port map( A1 => n2128, A2 => n2129, A3 => n2130, A4 => n2131
                           , ZN => n2112);
   U1119 : OAI22_X1 port map( A1 => n984, A2 => n1914, B1 => n951, B2 => n1915,
                           ZN => n2131);
   U1120 : OAI22_X1 port map( A1 => n1052, A2 => n1916, B1 => n1018, B2 => 
                           n1917, ZN => n2130);
   U1121 : OAI22_X1 port map( A1 => n93, A2 => n1918, B1 => n1085, B2 => n1919,
                           ZN => n2129);
   U1122 : OAI22_X1 port map( A1 => n167, A2 => n1920, B1 => n131, B2 => n1921,
                           ZN => n2128);
   U1123 : OAI22_X1 port map( A1 => n2132, A2 => n1868, B1 => n1869, B2 => 
                           n1370, ZN => N4530);
   U1124 : NOR4_X1 port map( A1 => n2137, A2 => n2138, A3 => n2139, A4 => n2140
                           , ZN => n2136);
   U1125 : OAI22_X1 port map( A1 => n189, A2 => n1878, B1 => n859, B2 => n1879,
                           ZN => n2140);
   U1126 : OAI22_X1 port map( A1 => n253, A2 => n1880, B1 => n221, B2 => n1881,
                           ZN => n2139);
   U1127 : OAI22_X1 port map( A1 => n317, A2 => n1882, B1 => n285, B2 => n1883,
                           ZN => n2138);
   U1128 : OAI22_X1 port map( A1 => n381, A2 => n1884, B1 => n349, B2 => n1885,
                           ZN => n2137);
   U1129 : NOR4_X1 port map( A1 => n2141, A2 => n2142, A3 => n2143, A4 => n2144
                           , ZN => n2135);
   U1130 : OAI22_X1 port map( A1 => n446, A2 => n1890, B1 => n413, B2 => n1891,
                           ZN => n2144);
   U1131 : OAI22_X1 port map( A1 => n513, A2 => n1892, B1 => n479, B2 => n1893,
                           ZN => n2143);
   U1132 : OAI22_X1 port map( A1 => n580, A2 => n1894, B1 => n547, B2 => n1895,
                           ZN => n2142);
   U1133 : OAI22_X1 port map( A1 => n647, A2 => n1896, B1 => n614, B2 => n1897,
                           ZN => n2141);
   U1134 : NOR4_X1 port map( A1 => n2145, A2 => n2146, A3 => n2147, A4 => n2148
                           , ZN => n2134);
   U1135 : OAI22_X1 port map( A1 => n715, A2 => n1902, B1 => n681, B2 => n1903,
                           ZN => n2148);
   U1136 : OAI22_X1 port map( A1 => n782, A2 => n1904, B1 => n748, B2 => n1905,
                           ZN => n2147);
   U1137 : OAI22_X1 port map( A1 => n849, A2 => n1906, B1 => n815, B2 => n1907,
                           ZN => n2146);
   U1138 : OAI22_X1 port map( A1 => n916, A2 => n1908, B1 => n883, B2 => n1909,
                           ZN => n2145);
   U1139 : NOR4_X1 port map( A1 => n2149, A2 => n2150, A3 => n2151, A4 => n2152
                           , ZN => n2133);
   U1140 : OAI22_X1 port map( A1 => n983, A2 => n1914, B1 => n950, B2 => n1915,
                           ZN => n2152);
   U1141 : OAI22_X1 port map( A1 => n1051, A2 => n1916, B1 => n1017, B2 => 
                           n1917, ZN => n2151);
   U1142 : OAI22_X1 port map( A1 => n91, A2 => n1918, B1 => n1084, B2 => n1919,
                           ZN => n2150);
   U1143 : OAI22_X1 port map( A1 => n166, A2 => n1920, B1 => n130, B2 => n1921,
                           ZN => n2149);
   U1144 : OAI22_X1 port map( A1 => n2153, A2 => n1868, B1 => n1869, B2 => 
                           n1392, ZN => N4528);
   U1145 : NOR4_X1 port map( A1 => n2158, A2 => n2159, A3 => n2160, A4 => n2161
                           , ZN => n2157);
   U1146 : OAI22_X1 port map( A1 => n188, A2 => n1878, B1 => n838, B2 => n1879,
                           ZN => n2161);
   U1147 : OAI22_X1 port map( A1 => n252, A2 => n1880, B1 => n220, B2 => n1881,
                           ZN => n2160);
   U1148 : OAI22_X1 port map( A1 => n316, A2 => n1882, B1 => n284, B2 => n1883,
                           ZN => n2159);
   U1149 : OAI22_X1 port map( A1 => n380, A2 => n1884, B1 => n348, B2 => n1885,
                           ZN => n2158);
   U1150 : NOR4_X1 port map( A1 => n2162, A2 => n2163, A3 => n2164, A4 => n2165
                           , ZN => n2156);
   U1151 : OAI22_X1 port map( A1 => n445, A2 => n1890, B1 => n412, B2 => n1891,
                           ZN => n2165);
   U1152 : OAI22_X1 port map( A1 => n512, A2 => n1892, B1 => n478, B2 => n1893,
                           ZN => n2164);
   U1153 : OAI22_X1 port map( A1 => n579, A2 => n1894, B1 => n546, B2 => n1895,
                           ZN => n2163);
   U1154 : OAI22_X1 port map( A1 => n646, A2 => n1896, B1 => n613, B2 => n1897,
                           ZN => n2162);
   U1155 : NOR4_X1 port map( A1 => n2166, A2 => n2167, A3 => n2168, A4 => n2169
                           , ZN => n2155);
   U1156 : OAI22_X1 port map( A1 => n714, A2 => n1902, B1 => n680, B2 => n1903,
                           ZN => n2169);
   U1157 : OAI22_X1 port map( A1 => n781, A2 => n1904, B1 => n747, B2 => n1905,
                           ZN => n2168);
   U1158 : OAI22_X1 port map( A1 => n848, A2 => n1906, B1 => n814, B2 => n1907,
                           ZN => n2167);
   U1159 : OAI22_X1 port map( A1 => n915, A2 => n1908, B1 => n882, B2 => n1909,
                           ZN => n2166);
   U1160 : NOR4_X1 port map( A1 => n2170, A2 => n2171, A3 => n2172, A4 => n2173
                           , ZN => n2154);
   U1161 : OAI22_X1 port map( A1 => n982, A2 => n1914, B1 => n949, B2 => n1915,
                           ZN => n2173);
   U1162 : OAI22_X1 port map( A1 => n1050, A2 => n1916, B1 => n1016, B2 => 
                           n1917, ZN => n2172);
   U1163 : OAI22_X1 port map( A1 => n89, A2 => n1918, B1 => n1083, B2 => n1919,
                           ZN => n2171);
   U1164 : OAI22_X1 port map( A1 => n164, A2 => n1920, B1 => n129, B2 => n1921,
                           ZN => n2170);
   U1165 : OAI22_X1 port map( A1 => n2174, A2 => n1868, B1 => n1869, B2 => 
                           n1414, ZN => N4526);
   U1166 : NOR4_X1 port map( A1 => n2179, A2 => n2180, A3 => n2181, A4 => n2182
                           , ZN => n2178);
   U1167 : OAI22_X1 port map( A1 => n187, A2 => n1878, B1 => n817, B2 => n1879,
                           ZN => n2182);
   U1168 : OAI22_X1 port map( A1 => n251, A2 => n1880, B1 => n219, B2 => n1881,
                           ZN => n2181);
   U1169 : OAI22_X1 port map( A1 => n315, A2 => n1882, B1 => n283, B2 => n1883,
                           ZN => n2180);
   U1170 : OAI22_X1 port map( A1 => n379, A2 => n1884, B1 => n347, B2 => n1885,
                           ZN => n2179);
   U1171 : NOR4_X1 port map( A1 => n2183, A2 => n2184, A3 => n2185, A4 => n2186
                           , ZN => n2177);
   U1172 : OAI22_X1 port map( A1 => n444, A2 => n1890, B1 => n411, B2 => n1891,
                           ZN => n2186);
   U1173 : OAI22_X1 port map( A1 => n511, A2 => n1892, B1 => n477, B2 => n1893,
                           ZN => n2185);
   U1174 : OAI22_X1 port map( A1 => n578, A2 => n1894, B1 => n545, B2 => n1895,
                           ZN => n2184);
   U1175 : OAI22_X1 port map( A1 => n645, A2 => n1896, B1 => n612, B2 => n1897,
                           ZN => n2183);
   U1176 : NOR4_X1 port map( A1 => n2187, A2 => n2188, A3 => n2189, A4 => n2190
                           , ZN => n2176);
   U1177 : OAI22_X1 port map( A1 => n713, A2 => n1902, B1 => n679, B2 => n1903,
                           ZN => n2190);
   U1178 : OAI22_X1 port map( A1 => n780, A2 => n1904, B1 => n746, B2 => n1905,
                           ZN => n2189);
   U1179 : OAI22_X1 port map( A1 => n847, A2 => n1906, B1 => n813, B2 => n1907,
                           ZN => n2188);
   U1180 : OAI22_X1 port map( A1 => n914, A2 => n1908, B1 => n881, B2 => n1909,
                           ZN => n2187);
   U1181 : NOR4_X1 port map( A1 => n2191, A2 => n2192, A3 => n2193, A4 => n2194
                           , ZN => n2175);
   U1182 : OAI22_X1 port map( A1 => n981, A2 => n1914, B1 => n948, B2 => n1915,
                           ZN => n2194);
   U1183 : OAI22_X1 port map( A1 => n1049, A2 => n1916, B1 => n1015, B2 => 
                           n1917, ZN => n2193);
   U1184 : OAI22_X1 port map( A1 => n87, A2 => n1918, B1 => n1082, B2 => n1919,
                           ZN => n2192);
   U1185 : OAI22_X1 port map( A1 => n163, A2 => n1920, B1 => n128, B2 => n1921,
                           ZN => n2191);
   U1186 : OAI22_X1 port map( A1 => n2195, A2 => n1868, B1 => n1869, B2 => 
                           n1436, ZN => N4524);
   U1187 : NOR4_X1 port map( A1 => n2200, A2 => n2201, A3 => n2202, A4 => n2203
                           , ZN => n2199);
   U1188 : OAI22_X1 port map( A1 => n186, A2 => n1878, B1 => n796, B2 => n1879,
                           ZN => n2203);
   U1189 : OAI22_X1 port map( A1 => n250, A2 => n1880, B1 => n218, B2 => n1881,
                           ZN => n2202);
   U1190 : OAI22_X1 port map( A1 => n314, A2 => n1882, B1 => n282, B2 => n1883,
                           ZN => n2201);
   U1191 : OAI22_X1 port map( A1 => n378, A2 => n1884, B1 => n346, B2 => n1885,
                           ZN => n2200);
   U1192 : NOR4_X1 port map( A1 => n2204, A2 => n2205, A3 => n2206, A4 => n2207
                           , ZN => n2198);
   U1193 : OAI22_X1 port map( A1 => n443, A2 => n1890, B1 => n410, B2 => n1891,
                           ZN => n2207);
   U1194 : OAI22_X1 port map( A1 => n510, A2 => n1892, B1 => n476, B2 => n1893,
                           ZN => n2206);
   U1195 : OAI22_X1 port map( A1 => n577, A2 => n1894, B1 => n543, B2 => n1895,
                           ZN => n2205);
   U1196 : OAI22_X1 port map( A1 => n644, A2 => n1896, B1 => n611, B2 => n1897,
                           ZN => n2204);
   U1197 : NOR4_X1 port map( A1 => n2208, A2 => n2209, A3 => n2210, A4 => n2211
                           , ZN => n2197);
   U1198 : OAI22_X1 port map( A1 => n711, A2 => n1902, B1 => n678, B2 => n1903,
                           ZN => n2211);
   U1199 : OAI22_X1 port map( A1 => n779, A2 => n1904, B1 => n745, B2 => n1905,
                           ZN => n2210);
   U1200 : OAI22_X1 port map( A1 => n846, A2 => n1906, B1 => n812, B2 => n1907,
                           ZN => n2209);
   U1201 : OAI22_X1 port map( A1 => n913, A2 => n1908, B1 => n879, B2 => n1909,
                           ZN => n2208);
   U1202 : NOR4_X1 port map( A1 => n2212, A2 => n2213, A3 => n2214, A4 => n2215
                           , ZN => n2196);
   U1203 : OAI22_X1 port map( A1 => n980, A2 => n1914, B1 => n947, B2 => n1915,
                           ZN => n2215);
   U1204 : OAI22_X1 port map( A1 => n1047, A2 => n1916, B1 => n1014, B2 => 
                           n1917, ZN => n2214);
   U1205 : OAI22_X1 port map( A1 => n85, A2 => n1918, B1 => n1081, B2 => n1919,
                           ZN => n2213);
   U1206 : OAI22_X1 port map( A1 => n162, A2 => n1920, B1 => n127, B2 => n1921,
                           ZN => n2212);
   U1207 : OAI22_X1 port map( A1 => n2216, A2 => n1868, B1 => n1869, B2 => 
                           n1458, ZN => N4522);
   U1208 : NOR4_X1 port map( A1 => n2221, A2 => n2222, A3 => n2223, A4 => n2224
                           , ZN => n2220);
   U1209 : OAI22_X1 port map( A1 => n185, A2 => n1878, B1 => n775, B2 => n1879,
                           ZN => n2224);
   U1210 : OAI22_X1 port map( A1 => n249, A2 => n1880, B1 => n217, B2 => n1881,
                           ZN => n2223);
   U1211 : OAI22_X1 port map( A1 => n313, A2 => n1882, B1 => n281, B2 => n1883,
                           ZN => n2222);
   U1212 : OAI22_X1 port map( A1 => n377, A2 => n1884, B1 => n345, B2 => n1885,
                           ZN => n2221);
   U1213 : NOR4_X1 port map( A1 => n2225, A2 => n2226, A3 => n2227, A4 => n2228
                           , ZN => n2219);
   U1214 : OAI22_X1 port map( A1 => n442, A2 => n1890, B1 => n409, B2 => n1891,
                           ZN => n2228);
   U1215 : OAI22_X1 port map( A1 => n509, A2 => n1892, B1 => n475, B2 => n1893,
                           ZN => n2227);
   U1216 : OAI22_X1 port map( A1 => n576, A2 => n1894, B1 => n542, B2 => n1895,
                           ZN => n2226);
   U1217 : OAI22_X1 port map( A1 => n643, A2 => n1896, B1 => n610, B2 => n1897,
                           ZN => n2225);
   U1218 : NOR4_X1 port map( A1 => n2229, A2 => n2230, A3 => n2231, A4 => n2232
                           , ZN => n2218);
   U1219 : OAI22_X1 port map( A1 => n710, A2 => n1902, B1 => n677, B2 => n1903,
                           ZN => n2232);
   U1220 : OAI22_X1 port map( A1 => n778, A2 => n1904, B1 => n744, B2 => n1905,
                           ZN => n2231);
   U1221 : OAI22_X1 port map( A1 => n845, A2 => n1906, B1 => n811, B2 => n1907,
                           ZN => n2230);
   U1222 : OAI22_X1 port map( A1 => n912, A2 => n1908, B1 => n878, B2 => n1909,
                           ZN => n2229);
   U1223 : NOR4_X1 port map( A1 => n2233, A2 => n2234, A3 => n2235, A4 => n2236
                           , ZN => n2217);
   U1224 : OAI22_X1 port map( A1 => n979, A2 => n1914, B1 => n946, B2 => n1915,
                           ZN => n2236);
   U1225 : OAI22_X1 port map( A1 => n1046, A2 => n1916, B1 => n1013, B2 => 
                           n1917, ZN => n2235);
   U1226 : OAI22_X1 port map( A1 => n83, A2 => n1918, B1 => n1080, B2 => n1919,
                           ZN => n2234);
   U1227 : OAI22_X1 port map( A1 => n161, A2 => n1920, B1 => n126, B2 => n1921,
                           ZN => n2233);
   U1228 : OAI22_X1 port map( A1 => n2237, A2 => n1868, B1 => n1869, B2 => 
                           n1480, ZN => N4520);
   U1229 : NOR4_X1 port map( A1 => n2242, A2 => n2243, A3 => n2244, A4 => n2245
                           , ZN => n2241);
   U1230 : OAI22_X1 port map( A1 => n184, A2 => n1878, B1 => n754, B2 => n1879,
                           ZN => n2245);
   U1231 : OAI22_X1 port map( A1 => n248, A2 => n1880, B1 => n216, B2 => n1881,
                           ZN => n2244);
   U1232 : OAI22_X1 port map( A1 => n312, A2 => n1882, B1 => n280, B2 => n1883,
                           ZN => n2243);
   U1233 : OAI22_X1 port map( A1 => n376, A2 => n1884, B1 => n344, B2 => n1885,
                           ZN => n2242);
   U1234 : NOR4_X1 port map( A1 => n2246, A2 => n2247, A3 => n2248, A4 => n2249
                           , ZN => n2240);
   U1235 : OAI22_X1 port map( A1 => n441, A2 => n1890, B1 => n408, B2 => n1891,
                           ZN => n2249);
   U1236 : OAI22_X1 port map( A1 => n508, A2 => n1892, B1 => n474, B2 => n1893,
                           ZN => n2248);
   U1237 : OAI22_X1 port map( A1 => n575, A2 => n1894, B1 => n541, B2 => n1895,
                           ZN => n2247);
   U1238 : OAI22_X1 port map( A1 => n642, A2 => n1896, B1 => n609, B2 => n1897,
                           ZN => n2246);
   U1239 : NOR4_X1 port map( A1 => n2250, A2 => n2251, A3 => n2252, A4 => n2253
                           , ZN => n2239);
   U1240 : OAI22_X1 port map( A1 => n709, A2 => n1902, B1 => n676, B2 => n1903,
                           ZN => n2253);
   U1241 : OAI22_X1 port map( A1 => n777, A2 => n1904, B1 => n743, B2 => n1905,
                           ZN => n2252);
   U1242 : OAI22_X1 port map( A1 => n844, A2 => n1906, B1 => n810, B2 => n1907,
                           ZN => n2251);
   U1243 : OAI22_X1 port map( A1 => n911, A2 => n1908, B1 => n877, B2 => n1909,
                           ZN => n2250);
   U1244 : NOR4_X1 port map( A1 => n2254, A2 => n2255, A3 => n2256, A4 => n2257
                           , ZN => n2238);
   U1245 : OAI22_X1 port map( A1 => n978, A2 => n1914, B1 => n945, B2 => n1915,
                           ZN => n2257);
   U1246 : OAI22_X1 port map( A1 => n1045, A2 => n1916, B1 => n1012, B2 => 
                           n1917, ZN => n2256);
   U1247 : OAI22_X1 port map( A1 => n81, A2 => n1918, B1 => n1079, B2 => n1919,
                           ZN => n2255);
   U1248 : OAI22_X1 port map( A1 => n160, A2 => n1920, B1 => n125, B2 => n1921,
                           ZN => n2254);
   U1249 : OAI22_X1 port map( A1 => n2258, A2 => n1868, B1 => n1869, B2 => 
                           n1502, ZN => N4518);
   U1250 : NOR4_X1 port map( A1 => n2263, A2 => n2264, A3 => n2265, A4 => n2266
                           , ZN => n2262);
   U1251 : OAI22_X1 port map( A1 => n183, A2 => n1878, B1 => n733, B2 => n1879,
                           ZN => n2266);
   U1252 : OAI22_X1 port map( A1 => n247, A2 => n1880, B1 => n215, B2 => n1881,
                           ZN => n2265);
   U1253 : OAI22_X1 port map( A1 => n311, A2 => n1882, B1 => n279, B2 => n1883,
                           ZN => n2264);
   U1254 : OAI22_X1 port map( A1 => n375, A2 => n1884, B1 => n343, B2 => n1885,
                           ZN => n2263);
   U1255 : NOR4_X1 port map( A1 => n2267, A2 => n2268, A3 => n2269, A4 => n2270
                           , ZN => n2261);
   U1256 : OAI22_X1 port map( A1 => n440, A2 => n1890, B1 => n407, B2 => n1891,
                           ZN => n2270);
   U1257 : OAI22_X1 port map( A1 => n507, A2 => n1892, B1 => n473, B2 => n1893,
                           ZN => n2269);
   U1258 : OAI22_X1 port map( A1 => n574, A2 => n1894, B1 => n540, B2 => n1895,
                           ZN => n2268);
   U1259 : OAI22_X1 port map( A1 => n641, A2 => n1896, B1 => n608, B2 => n1897,
                           ZN => n2267);
   U1260 : NOR4_X1 port map( A1 => n2271, A2 => n2272, A3 => n2273, A4 => n2274
                           , ZN => n2260);
   U1261 : OAI22_X1 port map( A1 => n708, A2 => n1902, B1 => n675, B2 => n1903,
                           ZN => n2274);
   U1262 : OAI22_X1 port map( A1 => n776, A2 => n1904, B1 => n742, B2 => n1905,
                           ZN => n2273);
   U1263 : OAI22_X1 port map( A1 => n843, A2 => n1906, B1 => n809, B2 => n1907,
                           ZN => n2272);
   U1264 : OAI22_X1 port map( A1 => n910, A2 => n1908, B1 => n876, B2 => n1909,
                           ZN => n2271);
   U1265 : NOR4_X1 port map( A1 => n2275, A2 => n2276, A3 => n2277, A4 => n2278
                           , ZN => n2259);
   U1266 : OAI22_X1 port map( A1 => n977, A2 => n1914, B1 => n944, B2 => n1915,
                           ZN => n2278);
   U1267 : OAI22_X1 port map( A1 => n1044, A2 => n1916, B1 => n1011, B2 => 
                           n1917, ZN => n2277);
   U1268 : OAI22_X1 port map( A1 => n79, A2 => n1918, B1 => n1078, B2 => n1919,
                           ZN => n2276);
   U1269 : OAI22_X1 port map( A1 => n159, A2 => n1920, B1 => n124, B2 => n1921,
                           ZN => n2275);
   U1270 : OAI22_X1 port map( A1 => n2279, A2 => n1868, B1 => n1869, B2 => 
                           n1524, ZN => N4516);
   U1271 : NOR4_X1 port map( A1 => n2284, A2 => n2285, A3 => n2286, A4 => n2287
                           , ZN => n2283);
   U1272 : OAI22_X1 port map( A1 => n182, A2 => n1878, B1 => n712, B2 => n1879,
                           ZN => n2287);
   U1273 : OAI22_X1 port map( A1 => n246, A2 => n1880, B1 => n214, B2 => n1881,
                           ZN => n2286);
   U1274 : OAI22_X1 port map( A1 => n310, A2 => n1882, B1 => n278, B2 => n1883,
                           ZN => n2285);
   U1275 : OAI22_X1 port map( A1 => n374, A2 => n1884, B1 => n342, B2 => n1885,
                           ZN => n2284);
   U1276 : NOR4_X1 port map( A1 => n2288, A2 => n2289, A3 => n2290, A4 => n2291
                           , ZN => n2282);
   U1277 : OAI22_X1 port map( A1 => n438, A2 => n1890, B1 => n406, B2 => n1891,
                           ZN => n2291);
   U1278 : OAI22_X1 port map( A1 => n506, A2 => n1892, B1 => n472, B2 => n1893,
                           ZN => n2290);
   U1279 : OAI22_X1 port map( A1 => n573, A2 => n1894, B1 => n539, B2 => n1895,
                           ZN => n2289);
   U1280 : OAI22_X1 port map( A1 => n640, A2 => n1896, B1 => n606, B2 => n1897,
                           ZN => n2288);
   U1281 : NOR4_X1 port map( A1 => n2292, A2 => n2293, A3 => n2294, A4 => n2295
                           , ZN => n2281);
   U1282 : OAI22_X1 port map( A1 => n707, A2 => n1902, B1 => n674, B2 => n1903,
                           ZN => n2295);
   U1283 : OAI22_X1 port map( A1 => n774, A2 => n1904, B1 => n741, B2 => n1905,
                           ZN => n2294);
   U1284 : OAI22_X1 port map( A1 => n842, A2 => n1906, B1 => n808, B2 => n1907,
                           ZN => n2293);
   U1285 : OAI22_X1 port map( A1 => n909, A2 => n1908, B1 => n875, B2 => n1909,
                           ZN => n2292);
   U1286 : NOR4_X1 port map( A1 => n2296, A2 => n2297, A3 => n2298, A4 => n2299
                           , ZN => n2280);
   U1287 : OAI22_X1 port map( A1 => n976, A2 => n1914, B1 => n942, B2 => n1915,
                           ZN => n2299);
   U1288 : OAI22_X1 port map( A1 => n1043, A2 => n1916, B1 => n1010, B2 => 
                           n1917, ZN => n2298);
   U1289 : OAI22_X1 port map( A1 => n75, A2 => n1918, B1 => n1077, B2 => n1919,
                           ZN => n2297);
   U1290 : OAI22_X1 port map( A1 => n158, A2 => n1920, B1 => n123, B2 => n1921,
                           ZN => n2296);
   U1291 : OAI22_X1 port map( A1 => n2300, A2 => n1868, B1 => n1869, B2 => 
                           n1546, ZN => N4514);
   U1292 : NOR4_X1 port map( A1 => n2305, A2 => n2306, A3 => n2307, A4 => n2308
                           , ZN => n2304);
   U1293 : OAI22_X1 port map( A1 => n181, A2 => n1878, B1 => n691, B2 => n1879,
                           ZN => n2308);
   U1294 : OAI22_X1 port map( A1 => n245, A2 => n1880, B1 => n213, B2 => n1881,
                           ZN => n2307);
   U1295 : OAI22_X1 port map( A1 => n309, A2 => n1882, B1 => n277, B2 => n1883,
                           ZN => n2306);
   U1296 : OAI22_X1 port map( A1 => n373, A2 => n1884, B1 => n341, B2 => n1885,
                           ZN => n2305);
   U1297 : NOR4_X1 port map( A1 => n2309, A2 => n2310, A3 => n2311, A4 => n2312
                           , ZN => n2303);
   U1298 : OAI22_X1 port map( A1 => n437, A2 => n1890, B1 => n405, B2 => n1891,
                           ZN => n2312);
   U1299 : OAI22_X1 port map( A1 => n505, A2 => n1892, B1 => n471, B2 => n1893,
                           ZN => n2311);
   U1300 : OAI22_X1 port map( A1 => n572, A2 => n1894, B1 => n538, B2 => n1895,
                           ZN => n2310);
   U1301 : OAI22_X1 port map( A1 => n639, A2 => n1896, B1 => n605, B2 => n1897,
                           ZN => n2309);
   U1302 : NOR4_X1 port map( A1 => n2313, A2 => n2314, A3 => n2315, A4 => n2316
                           , ZN => n2302);
   U1303 : OAI22_X1 port map( A1 => n706, A2 => n1902, B1 => n673, B2 => n1903,
                           ZN => n2316);
   U1304 : OAI22_X1 port map( A1 => n773, A2 => n1904, B1 => n740, B2 => n1905,
                           ZN => n2315);
   U1305 : OAI22_X1 port map( A1 => n841, A2 => n1906, B1 => n807, B2 => n1907,
                           ZN => n2314);
   U1306 : OAI22_X1 port map( A1 => n908, A2 => n1908, B1 => n874, B2 => n1909,
                           ZN => n2313);
   U1307 : NOR4_X1 port map( A1 => n2317, A2 => n2318, A3 => n2319, A4 => n2320
                           , ZN => n2301);
   U1308 : OAI22_X1 port map( A1 => n975, A2 => n1914, B1 => n941, B2 => n1915,
                           ZN => n2320);
   U1309 : OAI22_X1 port map( A1 => n1042, A2 => n1916, B1 => n1009, B2 => 
                           n1917, ZN => n2319);
   U1310 : OAI22_X1 port map( A1 => n73, A2 => n1918, B1 => n1076, B2 => n1919,
                           ZN => n2318);
   U1311 : OAI22_X1 port map( A1 => n157, A2 => n1920, B1 => n122, B2 => n1921,
                           ZN => n2317);
   U1312 : OAI22_X1 port map( A1 => n2321, A2 => n1868, B1 => n1869, B2 => 
                           n1568, ZN => N4512);
   U1313 : NOR4_X1 port map( A1 => n2326, A2 => n2327, A3 => n2328, A4 => n2329
                           , ZN => n2325);
   U1314 : OAI22_X1 port map( A1 => n180, A2 => n1878, B1 => n670, B2 => n1879,
                           ZN => n2329);
   U1315 : OAI22_X1 port map( A1 => n244, A2 => n1880, B1 => n212, B2 => n1881,
                           ZN => n2328);
   U1316 : OAI22_X1 port map( A1 => n308, A2 => n39, B1 => n276, B2 => n41, ZN 
                           => n2327);
   U1317 : OAI22_X1 port map( A1 => n372, A2 => n43, B1 => n340, B2 => n45, ZN 
                           => n2326);
   U1318 : NOR4_X1 port map( A1 => n2330, A2 => n2331, A3 => n2332, A4 => n2333
                           , ZN => n2324);
   U1319 : OAI22_X1 port map( A1 => n436, A2 => n1890, B1 => n404, B2 => n1891,
                           ZN => n2333);
   U1320 : OAI22_X1 port map( A1 => n504, A2 => n1892, B1 => n470, B2 => n1893,
                           ZN => n2332);
   U1321 : OAI22_X1 port map( A1 => n571, A2 => n1894, B1 => n537, B2 => n1895,
                           ZN => n2331);
   U1322 : OAI22_X1 port map( A1 => n638, A2 => n1896, B1 => n604, B2 => n1897,
                           ZN => n2330);
   U1323 : NOR4_X1 port map( A1 => n2334, A2 => n2335, A3 => n2336, A4 => n2337
                           , ZN => n2323);
   U1324 : OAI22_X1 port map( A1 => n705, A2 => n1902, B1 => n672, B2 => n1903,
                           ZN => n2337);
   U1325 : OAI22_X1 port map( A1 => n772, A2 => n1904, B1 => n739, B2 => n1905,
                           ZN => n2336);
   U1326 : OAI22_X1 port map( A1 => n840, A2 => n1906, B1 => n806, B2 => n1907,
                           ZN => n2335);
   U1327 : OAI22_X1 port map( A1 => n907, A2 => n1908, B1 => n873, B2 => n1909,
                           ZN => n2334);
   U1328 : NOR4_X1 port map( A1 => n2338, A2 => n2339, A3 => n2340, A4 => n2341
                           , ZN => n2322);
   U1329 : OAI22_X1 port map( A1 => n974, A2 => n1914, B1 => n940, B2 => n1915,
                           ZN => n2341);
   U1330 : OAI22_X1 port map( A1 => n1041, A2 => n1916, B1 => n1008, B2 => 
                           n1917, ZN => n2340);
   U1331 : OAI22_X1 port map( A1 => n71, A2 => n1918, B1 => n1075, B2 => n1919,
                           ZN => n2339);
   U1332 : OAI22_X1 port map( A1 => n156, A2 => n1920, B1 => n120, B2 => n1921,
                           ZN => n2338);
   U1333 : OAI22_X1 port map( A1 => n2342, A2 => n1868, B1 => n1869, B2 => 
                           n1590, ZN => N4510);
   U1334 : NOR4_X1 port map( A1 => n2347, A2 => n2348, A3 => n2349, A4 => n2350
                           , ZN => n2346);
   U1335 : OAI22_X1 port map( A1 => n179, A2 => n1878, B1 => n649, B2 => n1879,
                           ZN => n2350);
   U1336 : OAI22_X1 port map( A1 => n243, A2 => n1880, B1 => n211, B2 => n1881,
                           ZN => n2349);
   U1337 : OAI22_X1 port map( A1 => n307, A2 => n39, B1 => n275, B2 => n41, ZN 
                           => n2348);
   U1338 : OAI22_X1 port map( A1 => n371, A2 => n43, B1 => n339, B2 => n45, ZN 
                           => n2347);
   U1339 : NOR4_X1 port map( A1 => n2351, A2 => n2352, A3 => n2353, A4 => n2354
                           , ZN => n2345);
   U1340 : OAI22_X1 port map( A1 => n435, A2 => n1890, B1 => n403, B2 => n1891,
                           ZN => n2354);
   U1341 : OAI22_X1 port map( A1 => n503, A2 => n1892, B1 => n469, B2 => n1893,
                           ZN => n2353);
   U1342 : OAI22_X1 port map( A1 => n570, A2 => n1894, B1 => n536, B2 => n1895,
                           ZN => n2352);
   U1343 : OAI22_X1 port map( A1 => n637, A2 => n1896, B1 => n603, B2 => n1897,
                           ZN => n2351);
   U1344 : NOR4_X1 port map( A1 => n2355, A2 => n2356, A3 => n2357, A4 => n2358
                           , ZN => n2344);
   U1345 : OAI22_X1 port map( A1 => n704, A2 => n1902, B1 => n671, B2 => n1903,
                           ZN => n2358);
   U1346 : OAI22_X1 port map( A1 => n771, A2 => n1904, B1 => n738, B2 => n1905,
                           ZN => n2357);
   U1347 : OAI22_X1 port map( A1 => n839, A2 => n1906, B1 => n805, B2 => n1907,
                           ZN => n2356);
   U1348 : OAI22_X1 port map( A1 => n906, A2 => n1908, B1 => n872, B2 => n1909,
                           ZN => n2355);
   U1349 : NOR4_X1 port map( A1 => n2359, A2 => n2360, A3 => n2361, A4 => n2362
                           , ZN => n2343);
   U1350 : OAI22_X1 port map( A1 => n973, A2 => n1914, B1 => n939, B2 => n1915,
                           ZN => n2362);
   U1351 : OAI22_X1 port map( A1 => n1040, A2 => n1916, B1 => n1007, B2 => 
                           n1917, ZN => n2361);
   U1352 : OAI22_X1 port map( A1 => n69, A2 => n1918, B1 => n1074, B2 => n1919,
                           ZN => n2360);
   U1353 : OAI22_X1 port map( A1 => n155, A2 => n1920, B1 => n119, B2 => n1921,
                           ZN => n2359);
   U1354 : OAI22_X1 port map( A1 => n2363, A2 => n1868, B1 => n1869, B2 => 
                           n1612, ZN => N4508);
   U1355 : NOR4_X1 port map( A1 => n2368, A2 => n2369, A3 => n2370, A4 => n2371
                           , ZN => n2367);
   U1356 : OAI22_X1 port map( A1 => n176, A2 => n1878, B1 => n628, B2 => n1879,
                           ZN => n2371);
   U1357 : OAI22_X1 port map( A1 => n242, A2 => n1880, B1 => n210, B2 => n1881,
                           ZN => n2370);
   U1358 : OAI22_X1 port map( A1 => n306, A2 => n39, B1 => n274, B2 => n41, ZN 
                           => n2369);
   U1359 : OAI22_X1 port map( A1 => n370, A2 => n43, B1 => n338, B2 => n45, ZN 
                           => n2368);
   U1360 : NOR4_X1 port map( A1 => n2372, A2 => n2373, A3 => n2374, A4 => n2375
                           , ZN => n2366);
   U1361 : OAI22_X1 port map( A1 => n434, A2 => n1890, B1 => n402, B2 => n1891,
                           ZN => n2375);
   U1362 : OAI22_X1 port map( A1 => n501, A2 => n1892, B1 => n468, B2 => n1893,
                           ZN => n2374);
   U1363 : OAI22_X1 port map( A1 => n569, A2 => n1894, B1 => n535, B2 => n1895,
                           ZN => n2373);
   U1364 : OAI22_X1 port map( A1 => n636, A2 => n1896, B1 => n602, B2 => n1897,
                           ZN => n2372);
   U1365 : NOR4_X1 port map( A1 => n2376, A2 => n2377, A3 => n2378, A4 => n2379
                           , ZN => n2365);
   U1366 : OAI22_X1 port map( A1 => n703, A2 => n1902, B1 => n669, B2 => n1903,
                           ZN => n2379);
   U1367 : OAI22_X1 port map( A1 => n770, A2 => n1904, B1 => n737, B2 => n1905,
                           ZN => n2378);
   U1368 : OAI22_X1 port map( A1 => n837, A2 => n1906, B1 => n804, B2 => n1907,
                           ZN => n2377);
   U1369 : OAI22_X1 port map( A1 => n905, A2 => n1908, B1 => n871, B2 => n1909,
                           ZN => n2376);
   U1370 : NOR4_X1 port map( A1 => n2380, A2 => n2381, A3 => n2382, A4 => n2383
                           , ZN => n2364);
   U1371 : OAI22_X1 port map( A1 => n972, A2 => n1914, B1 => n938, B2 => n1915,
                           ZN => n2383);
   U1372 : OAI22_X1 port map( A1 => n1039, A2 => n1916, B1 => n1005, B2 => 
                           n1917, ZN => n2382);
   U1373 : OAI22_X1 port map( A1 => n67, A2 => n1918, B1 => n1073, B2 => n1919,
                           ZN => n2381);
   U1374 : OAI22_X1 port map( A1 => n153, A2 => n1920, B1 => n118, B2 => n1921,
                           ZN => n2380);
   U1375 : OAI22_X1 port map( A1 => n2384, A2 => n1868, B1 => n1869, B2 => 
                           n1634, ZN => N4506);
   U1376 : NOR4_X1 port map( A1 => n2389, A2 => n2390, A3 => n2391, A4 => n2392
                           , ZN => n2388);
   U1377 : OAI22_X1 port map( A1 => n165, A2 => n1878, B1 => n607, B2 => n1879,
                           ZN => n2392);
   U1378 : OAI22_X1 port map( A1 => n241, A2 => n1880, B1 => n209, B2 => n1881,
                           ZN => n2391);
   U1379 : OAI22_X1 port map( A1 => n305, A2 => n39, B1 => n273, B2 => n41, ZN 
                           => n2390);
   U1380 : OAI22_X1 port map( A1 => n369, A2 => n43, B1 => n337, B2 => n45, ZN 
                           => n2389);
   U1381 : NOR4_X1 port map( A1 => n2393, A2 => n2394, A3 => n2395, A4 => n2396
                           , ZN => n2387);
   U1382 : OAI22_X1 port map( A1 => n433, A2 => n1890, B1 => n401, B2 => n1891,
                           ZN => n2396);
   U1383 : OAI22_X1 port map( A1 => n500, A2 => n1892, B1 => n467, B2 => n1893,
                           ZN => n2395);
   U1384 : OAI22_X1 port map( A1 => n568, A2 => n1894, B1 => n534, B2 => n1895,
                           ZN => n2394);
   U1385 : OAI22_X1 port map( A1 => n635, A2 => n1896, B1 => n601, B2 => n1897,
                           ZN => n2393);
   U1386 : NOR4_X1 port map( A1 => n2397, A2 => n2398, A3 => n2399, A4 => n2400
                           , ZN => n2386);
   U1387 : OAI22_X1 port map( A1 => n702, A2 => n1902, B1 => n668, B2 => n1903,
                           ZN => n2400);
   U1388 : OAI22_X1 port map( A1 => n769, A2 => n1904, B1 => n736, B2 => n1905,
                           ZN => n2399);
   U1389 : OAI22_X1 port map( A1 => n836, A2 => n1906, B1 => n803, B2 => n1907,
                           ZN => n2398);
   U1390 : OAI22_X1 port map( A1 => n904, A2 => n1908, B1 => n870, B2 => n1909,
                           ZN => n2397);
   U1391 : NOR4_X1 port map( A1 => n2401, A2 => n2402, A3 => n2403, A4 => n2404
                           , ZN => n2385);
   U1392 : OAI22_X1 port map( A1 => n971, A2 => n1914, B1 => n937, B2 => n1915,
                           ZN => n2404);
   U1393 : OAI22_X1 port map( A1 => n1038, A2 => n1916, B1 => n1004, B2 => 
                           n1917, ZN => n2403);
   U1394 : OAI22_X1 port map( A1 => n65, A2 => n1918, B1 => n1072, B2 => n1919,
                           ZN => n2402);
   U1395 : OAI22_X1 port map( A1 => n152, A2 => n1920, B1 => n117, B2 => n1921,
                           ZN => n2401);
   U1396 : OAI22_X1 port map( A1 => n2405, A2 => n1868, B1 => n1869, B2 => 
                           n1656, ZN => N4504);
   U1397 : NOR4_X1 port map( A1 => n2410, A2 => n2411, A3 => n2412, A4 => n2413
                           , ZN => n2409);
   U1398 : OAI22_X1 port map( A1 => n154, A2 => n1878, B1 => n586, B2 => n1879,
                           ZN => n2413);
   U1399 : OAI22_X1 port map( A1 => n240, A2 => n1880, B1 => n208, B2 => n1881,
                           ZN => n2412);
   U1400 : OAI22_X1 port map( A1 => n304, A2 => n39, B1 => n272, B2 => n41, ZN 
                           => n2411);
   U1401 : OAI22_X1 port map( A1 => n368, A2 => n43, B1 => n336, B2 => n45, ZN 
                           => n2410);
   U1402 : NOR4_X1 port map( A1 => n2414, A2 => n2415, A3 => n2416, A4 => n2417
                           , ZN => n2408);
   U1403 : OAI22_X1 port map( A1 => n432, A2 => n1890, B1 => n400, B2 => n1891,
                           ZN => n2417);
   U1404 : OAI22_X1 port map( A1 => n499, A2 => n1892, B1 => n466, B2 => n1893,
                           ZN => n2416);
   U1405 : OAI22_X1 port map( A1 => n567, A2 => n1894, B1 => n533, B2 => n1895,
                           ZN => n2415);
   U1406 : OAI22_X1 port map( A1 => n634, A2 => n1896, B1 => n600, B2 => n1897,
                           ZN => n2414);
   U1407 : NOR4_X1 port map( A1 => n2418, A2 => n2419, A3 => n2420, A4 => n2421
                           , ZN => n2407);
   U1408 : OAI22_X1 port map( A1 => n701, A2 => n1902, B1 => n667, B2 => n1903,
                           ZN => n2421);
   U1409 : OAI22_X1 port map( A1 => n768, A2 => n1904, B1 => n735, B2 => n1905,
                           ZN => n2420);
   U1410 : OAI22_X1 port map( A1 => n835, A2 => n1906, B1 => n802, B2 => n1907,
                           ZN => n2419);
   U1411 : OAI22_X1 port map( A1 => n903, A2 => n1908, B1 => n869, B2 => n1909,
                           ZN => n2418);
   U1412 : NOR4_X1 port map( A1 => n2422, A2 => n2423, A3 => n2424, A4 => n2425
                           , ZN => n2406);
   U1413 : OAI22_X1 port map( A1 => n970, A2 => n1914, B1 => n936, B2 => n1915,
                           ZN => n2425);
   U1414 : OAI22_X1 port map( A1 => n1037, A2 => n1916, B1 => n1003, B2 => 
                           n1917, ZN => n2424);
   U1415 : OAI22_X1 port map( A1 => n63, A2 => n1918, B1 => n1071, B2 => n1919,
                           ZN => n2423);
   U1416 : OAI22_X1 port map( A1 => n151, A2 => n1920, B1 => n116, B2 => n1921,
                           ZN => n2422);
   U1417 : OAI22_X1 port map( A1 => n2426, A2 => n1868, B1 => n1869, B2 => 
                           n1678, ZN => N4502);
   U1418 : NOR4_X1 port map( A1 => n2431, A2 => n2432, A3 => n2433, A4 => n2434
                           , ZN => n2430);
   U1419 : OAI22_X1 port map( A1 => n143, A2 => n1878, B1 => n565, B2 => n1879,
                           ZN => n2434);
   U1420 : OAI22_X1 port map( A1 => n239, A2 => n1880, B1 => n207, B2 => n1881,
                           ZN => n2433);
   U1421 : OAI22_X1 port map( A1 => n303, A2 => n39, B1 => n271, B2 => n41, ZN 
                           => n2432);
   U1422 : OAI22_X1 port map( A1 => n367, A2 => n43, B1 => n335, B2 => n45, ZN 
                           => n2431);
   U1423 : NOR4_X1 port map( A1 => n2435, A2 => n2436, A3 => n2437, A4 => n2438
                           , ZN => n2429);
   U1424 : OAI22_X1 port map( A1 => n431, A2 => n1890, B1 => n399, B2 => n1891,
                           ZN => n2438);
   U1425 : OAI22_X1 port map( A1 => n498, A2 => n1892, B1 => n465, B2 => n1893,
                           ZN => n2437);
   U1426 : OAI22_X1 port map( A1 => n566, A2 => n1894, B1 => n532, B2 => n1895,
                           ZN => n2436);
   U1427 : OAI22_X1 port map( A1 => n633, A2 => n1896, B1 => n599, B2 => n1897,
                           ZN => n2435);
   U1428 : NOR4_X1 port map( A1 => n2439, A2 => n2440, A3 => n2441, A4 => n2442
                           , ZN => n2428);
   U1429 : OAI22_X1 port map( A1 => n700, A2 => n1902, B1 => n666, B2 => n1903,
                           ZN => n2442);
   U1430 : OAI22_X1 port map( A1 => n767, A2 => n1904, B1 => n734, B2 => n1905,
                           ZN => n2441);
   U1431 : OAI22_X1 port map( A1 => n834, A2 => n1906, B1 => n801, B2 => n1907,
                           ZN => n2440);
   U1432 : OAI22_X1 port map( A1 => n902, A2 => n1908, B1 => n868, B2 => n1909,
                           ZN => n2439);
   U1433 : NOR4_X1 port map( A1 => n2443, A2 => n2444, A3 => n2445, A4 => n2446
                           , ZN => n2427);
   U1434 : OAI22_X1 port map( A1 => n969, A2 => n1914, B1 => n935, B2 => n1915,
                           ZN => n2446);
   U1435 : OAI22_X1 port map( A1 => n1036, A2 => n1916, B1 => n1002, B2 => 
                           n1917, ZN => n2445);
   U1436 : OAI22_X1 port map( A1 => n61, A2 => n1918, B1 => n1070, B2 => n1919,
                           ZN => n2444);
   U1437 : OAI22_X1 port map( A1 => n150, A2 => n1920, B1 => n115, B2 => n1921,
                           ZN => n2443);
   U1438 : OAI22_X1 port map( A1 => n2447, A2 => n1868, B1 => n1869, B2 => 
                           n1700, ZN => N4500);
   U1439 : NOR4_X1 port map( A1 => n2452, A2 => n2453, A3 => n2454, A4 => n2455
                           , ZN => n2451);
   U1440 : OAI22_X1 port map( A1 => n132, A2 => n1878, B1 => n544, B2 => n1879,
                           ZN => n2455);
   U1441 : OAI22_X1 port map( A1 => n238, A2 => n1880, B1 => n206, B2 => n1881,
                           ZN => n2454);
   U1442 : OAI22_X1 port map( A1 => n302, A2 => n39, B1 => n270, B2 => n41, ZN 
                           => n2453);
   U1443 : OAI22_X1 port map( A1 => n366, A2 => n43, B1 => n334, B2 => n45, ZN 
                           => n2452);
   U1444 : NOR4_X1 port map( A1 => n2456, A2 => n2457, A3 => n2458, A4 => n2459
                           , ZN => n2450);
   U1445 : OAI22_X1 port map( A1 => n430, A2 => n1890, B1 => n398, B2 => n1891,
                           ZN => n2459);
   U1446 : OAI22_X1 port map( A1 => n497, A2 => n1892, B1 => n464, B2 => n1893,
                           ZN => n2458);
   U1447 : OAI22_X1 port map( A1 => n564, A2 => n1894, B1 => n531, B2 => n1895,
                           ZN => n2457);
   U1448 : OAI22_X1 port map( A1 => n632, A2 => n1896, B1 => n598, B2 => n1897,
                           ZN => n2456);
   U1449 : NOR4_X1 port map( A1 => n2460, A2 => n2461, A3 => n2462, A4 => n2463
                           , ZN => n2449);
   U1450 : OAI22_X1 port map( A1 => n699, A2 => n1902, B1 => n665, B2 => n1903,
                           ZN => n2463);
   U1451 : OAI22_X1 port map( A1 => n766, A2 => n1904, B1 => n732, B2 => n1905,
                           ZN => n2462);
   U1452 : OAI22_X1 port map( A1 => n833, A2 => n1906, B1 => n800, B2 => n1907,
                           ZN => n2461);
   U1453 : OAI22_X1 port map( A1 => n900, A2 => n1908, B1 => n867, B2 => n1909,
                           ZN => n2460);
   U1454 : NOR4_X1 port map( A1 => n2464, A2 => n2465, A3 => n2466, A4 => n2467
                           , ZN => n2448);
   U1455 : OAI22_X1 port map( A1 => n968, A2 => n1914, B1 => n934, B2 => n1915,
                           ZN => n2467);
   U1456 : OAI22_X1 port map( A1 => n1035, A2 => n1916, B1 => n1001, B2 => 
                           n1917, ZN => n2466);
   U1457 : OAI22_X1 port map( A1 => n59, A2 => n1918, B1 => n1068, B2 => n1919,
                           ZN => n2465);
   U1458 : OAI22_X1 port map( A1 => n149, A2 => n1920, B1 => n114, B2 => n1921,
                           ZN => n2464);
   U1459 : OAI22_X1 port map( A1 => n2468, A2 => n1868, B1 => n1869, B2 => 
                           n1722, ZN => N4498);
   U1460 : NOR4_X1 port map( A1 => n2473, A2 => n2474, A3 => n2475, A4 => n2476
                           , ZN => n2472);
   U1461 : OAI22_X1 port map( A1 => n121, A2 => n1878, B1 => n523, B2 => n1879,
                           ZN => n2476);
   U1462 : OAI22_X1 port map( A1 => n237, A2 => n1880, B1 => n205, B2 => n1881,
                           ZN => n2475);
   U1463 : OAI22_X1 port map( A1 => n301, A2 => n39, B1 => n269, B2 => n41, ZN 
                           => n2474);
   U1464 : OAI22_X1 port map( A1 => n365, A2 => n43, B1 => n333, B2 => n45, ZN 
                           => n2473);
   U1465 : NOR4_X1 port map( A1 => n2477, A2 => n2478, A3 => n2479, A4 => n2480
                           , ZN => n2471);
   U1466 : OAI22_X1 port map( A1 => n429, A2 => n1890, B1 => n397, B2 => n1891,
                           ZN => n2480);
   U1467 : OAI22_X1 port map( A1 => n496, A2 => n1892, B1 => n463, B2 => n1893,
                           ZN => n2479);
   U1468 : OAI22_X1 port map( A1 => n563, A2 => n1894, B1 => n530, B2 => n1895,
                           ZN => n2478);
   U1469 : OAI22_X1 port map( A1 => n631, A2 => n1896, B1 => n597, B2 => n1897,
                           ZN => n2477);
   U1470 : NOR4_X1 port map( A1 => n2481, A2 => n2482, A3 => n2483, A4 => n2484
                           , ZN => n2470);
   U1471 : OAI22_X1 port map( A1 => n698, A2 => n1902, B1 => n664, B2 => n1903,
                           ZN => n2484);
   U1472 : OAI22_X1 port map( A1 => n765, A2 => n1904, B1 => n731, B2 => n1905,
                           ZN => n2483);
   U1473 : OAI22_X1 port map( A1 => n832, A2 => n1906, B1 => n799, B2 => n1907,
                           ZN => n2482);
   U1474 : OAI22_X1 port map( A1 => n899, A2 => n1908, B1 => n866, B2 => n1909,
                           ZN => n2481);
   U1475 : NOR4_X1 port map( A1 => n2485, A2 => n2486, A3 => n2487, A4 => n2488
                           , ZN => n2469);
   U1476 : OAI22_X1 port map( A1 => n967, A2 => n1914, B1 => n933, B2 => n1915,
                           ZN => n2488);
   U1477 : OAI22_X1 port map( A1 => n1034, A2 => n1916, B1 => n1000, B2 => 
                           n1917, ZN => n2487);
   U1478 : OAI22_X1 port map( A1 => n57, A2 => n1918, B1 => n1067, B2 => n1919,
                           ZN => n2486);
   U1479 : OAI22_X1 port map( A1 => n148, A2 => n1920, B1 => n113, B2 => n1921,
                           ZN => n2485);
   U1480 : OAI22_X1 port map( A1 => n2489, A2 => n1868, B1 => n1869, B2 => 
                           n1744, ZN => N4496);
   U1481 : NOR4_X1 port map( A1 => n2490, A2 => n2491, A3 => n2492, A4 => n2493
                           , ZN => n2489);
   U1482 : OAI211_X1 port map( C1 => n1101, C2 => n1918, A => n2494, B => n2495
                           , ZN => n2493);
   U1483 : NOR4_X1 port map( A1 => n2496, A2 => n2497, A3 => n2498, A4 => n2499
                           , ZN => n2495);
   U1484 : OAI22_X1 port map( A1 => n110, A2 => n1878, B1 => n204, B2 => n1881,
                           ZN => n2499);
   U1485 : OAI22_X1 port map( A1 => n236, A2 => n1880, B1 => n268, B2 => n41, 
                           ZN => n2498);
   U1486 : OAI22_X1 port map( A1 => n300, A2 => n39, B1 => n332, B2 => n45, ZN 
                           => n2497);
   U1487 : OAI22_X1 port map( A1 => n364, A2 => n43, B1 => n396, B2 => n1891, 
                           ZN => n2496);
   U1488 : NOR4_X1 port map( A1 => n2500, A2 => n2501, A3 => n2502, A4 => 
                           n2503_port, ZN => n2494);
   U1489 : OAI22_X1 port map( A1 => n428, A2 => n1890, B1 => n462, B2 => n1893,
                           ZN => n2503_port);
   U1490 : OAI22_X1 port map( A1 => n495, A2 => n1892, B1 => n529, B2 => n1895,
                           ZN => n2502);
   U1491 : OAI22_X1 port map( A1 => n562, A2 => n1894, B1 => n596, B2 => n1897,
                           ZN => n2501);
   U1492 : OAI22_X1 port map( A1 => n630, A2 => n1896, B1 => n663, B2 => n1903,
                           ZN => n2500);
   U1493 : OAI211_X1 port map( C1 => n147, C2 => n1920, A => n2504, B => n2505,
                           ZN => n2492);
   U1494 : NOR4_X1 port map( A1 => n2506, A2 => n2507, A3 => n2508, A4 => n2509
                           , ZN => n2505);
   U1495 : OAI22_X1 port map( A1 => n764, A2 => n1904, B1 => n798, B2 => n1907,
                           ZN => n2509);
   U1496 : OAI22_X1 port map( A1 => n697, A2 => n1902, B1 => n730, B2 => n1905,
                           ZN => n2508);
   U1497 : OAI22_X1 port map( A1 => n898, A2 => n1908, B1 => n932, B2 => n1915,
                           ZN => n2507);
   U1498 : OAI22_X1 port map( A1 => n831, A2 => n1906, B1 => n865, B2 => n1909,
                           ZN => n2506);
   U1499 : OAI22_X1 port map( A1 => n1879, A2 => n502, B1 => n1921, B2 => n112,
                           ZN => n2510);
   U1500 : OAI22_X1 port map( A1 => n1033, A2 => n1916, B1 => n1066, B2 => 
                           n1919, ZN => n2491);
   U1501 : OAI22_X1 port map( A1 => n966, A2 => n1914, B1 => n999, B2 => n1917,
                           ZN => n2490);
   U1502 : OAI22_X1 port map( A1 => n2511, A2 => n1868, B1 => n1869, B2 => 
                           n1766, ZN => N4494);
   U1503 : NOR4_X1 port map( A1 => n2516, A2 => n2517, A3 => n2518, A4 => n2519
                           , ZN => n2515);
   U1504 : OAI22_X1 port map( A1 => n99, A2 => n1878, B1 => n481, B2 => n1879, 
                           ZN => n2519);
   U1505 : OAI22_X1 port map( A1 => n235, A2 => n1880, B1 => n203, B2 => n1881,
                           ZN => n2518);
   U1506 : OAI22_X1 port map( A1 => n299, A2 => n39, B1 => n267, B2 => n41, ZN 
                           => n2517);
   U1507 : OAI22_X1 port map( A1 => n363, A2 => n43, B1 => n331, B2 => n45, ZN 
                           => n2516);
   U1508 : NOR4_X1 port map( A1 => n2520, A2 => n2521, A3 => n2522, A4 => n2523
                           , ZN => n2514);
   U1509 : OAI22_X1 port map( A1 => n427, A2 => n1890, B1 => n395, B2 => n1891,
                           ZN => n2523);
   U1510 : OAI22_X1 port map( A1 => n494, A2 => n1892, B1 => n461, B2 => n1893,
                           ZN => n2522);
   U1511 : OAI22_X1 port map( A1 => n561, A2 => n1894, B1 => n528, B2 => n1895,
                           ZN => n2521);
   U1512 : OAI22_X1 port map( A1 => n629, A2 => n1896, B1 => n595, B2 => n1897,
                           ZN => n2520);
   U1513 : NOR4_X1 port map( A1 => n2524, A2 => n2525, A3 => n2526, A4 => n2527
                           , ZN => n2513);
   U1514 : OAI22_X1 port map( A1 => n696, A2 => n1902, B1 => n662, B2 => n1903,
                           ZN => n2527);
   U1515 : OAI22_X1 port map( A1 => n763, A2 => n1904, B1 => n729, B2 => n1905,
                           ZN => n2526);
   U1516 : OAI22_X1 port map( A1 => n830, A2 => n1906, B1 => n797, B2 => n1907,
                           ZN => n2525);
   U1517 : OAI22_X1 port map( A1 => n897, A2 => n1908, B1 => n864, B2 => n1909,
                           ZN => n2524);
   U1518 : NOR4_X1 port map( A1 => n2528, A2 => n2529, A3 => n2530, A4 => n2531
                           , ZN => n2512);
   U1519 : OAI22_X1 port map( A1 => n965, A2 => n1914, B1 => n931, B2 => n1915,
                           ZN => n2531);
   U1520 : OAI22_X1 port map( A1 => n1032, A2 => n1916, B1 => n998, B2 => n1917
                           , ZN => n2530);
   U1521 : OAI22_X1 port map( A1 => n1100, A2 => n1918, B1 => n1065, B2 => 
                           n1919, ZN => n2529);
   U1522 : OAI22_X1 port map( A1 => n146, A2 => n1920, B1 => n111, B2 => n1921,
                           ZN => n2528);
   U1523 : OAI22_X1 port map( A1 => n2532, A2 => n1868, B1 => n1869, B2 => 
                           n1788, ZN => N4492);
   U1524 : NOR4_X1 port map( A1 => n2537, A2 => n2538, A3 => n2539, A4 => n2540
                           , ZN => n2536);
   U1525 : OAI22_X1 port map( A1 => n77, A2 => n1878, B1 => n460, B2 => n1879, 
                           ZN => n2540);
   U1526 : OAI22_X1 port map( A1 => n234, A2 => n1880, B1 => n202, B2 => n1881,
                           ZN => n2539);
   U1527 : OAI22_X1 port map( A1 => n298, A2 => n39, B1 => n266, B2 => n41, ZN 
                           => n2538);
   U1528 : OAI22_X1 port map( A1 => n362, A2 => n43, B1 => n330, B2 => n45, ZN 
                           => n2537);
   U1529 : NOR4_X1 port map( A1 => n2541, A2 => n2542, A3 => n2543, A4 => n2544
                           , ZN => n2535);
   U1530 : OAI22_X1 port map( A1 => n426, A2 => n1890, B1 => n394, B2 => n1891,
                           ZN => n2544);
   U1531 : OAI22_X1 port map( A1 => n493, A2 => n1892, B1 => n459, B2 => n1893,
                           ZN => n2543);
   U1532 : OAI22_X1 port map( A1 => n560, A2 => n1894, B1 => n527, B2 => n1895,
                           ZN => n2542);
   U1533 : OAI22_X1 port map( A1 => n627, A2 => n1896, B1 => n594, B2 => n1897,
                           ZN => n2541);
   U1534 : NOR4_X1 port map( A1 => n2545, A2 => n2546, A3 => n2547, A4 => n2548
                           , ZN => n2534);
   U1535 : OAI22_X1 port map( A1 => n695, A2 => n1902, B1 => n661, B2 => n1903,
                           ZN => n2548);
   U1536 : OAI22_X1 port map( A1 => n762, A2 => n1904, B1 => n728, B2 => n1905,
                           ZN => n2547);
   U1537 : OAI22_X1 port map( A1 => n829, A2 => n1906, B1 => n795, B2 => n1907,
                           ZN => n2546);
   U1538 : OAI22_X1 port map( A1 => n896, A2 => n1908, B1 => n863, B2 => n1909,
                           ZN => n2545);
   U1539 : NOR4_X1 port map( A1 => n2549, A2 => n2550, A3 => n2551, A4 => n2552
                           , ZN => n2533);
   U1540 : OAI22_X1 port map( A1 => n963, A2 => n1914, B1 => n930, B2 => n1915,
                           ZN => n2552);
   U1541 : OAI22_X1 port map( A1 => n1031, A2 => n1916, B1 => n997, B2 => n1917
                           , ZN => n2551);
   U1542 : OAI22_X1 port map( A1 => n1099, A2 => n1918, B1 => n1064, B2 => 
                           n1919, ZN => n2550);
   U1543 : OAI22_X1 port map( A1 => n145, A2 => n1920, B1 => n109, B2 => n1921,
                           ZN => n2549);
   U1544 : OAI22_X1 port map( A1 => n2553, A2 => n1868, B1 => n1869, B2 => 
                           n1810, ZN => N4490);
   U1545 : OAI221_X1 port map( B1 => n1826, B2 => ADD_RD1(2), C1 => n1827, C2 
                           => ADD_RD1(0), A => n2558, ZN => n2557);
   U1546 : AOI22_X1 port map( A1 => n1826, A2 => ADD_RD1(2), B1 => n1827, B2 =>
                           ADD_RD1(0), ZN => n2558);
   U1547 : AOI221_X1 port map( B1 => n2559, B2 => ADD_WR(4), C1 => n1830, C2 =>
                           ADD_RD1(3), A => n2560, ZN => n2554);
   U1548 : OAI22_X1 port map( A1 => ADD_WR(4), A2 => n2559, B1 => n1830, B2 => 
                           ADD_RD1(3), ZN => n2560);
   U1549 : NOR4_X1 port map( A1 => n2569, A2 => n2570, A3 => n2571, A4 => n2572
                           , ZN => n2568);
   U1550 : OAI22_X1 port map( A1 => n55, A2 => n1878, B1 => n439, B2 => n1879, 
                           ZN => n2572);
   U1551 : OAI22_X1 port map( A1 => n233, A2 => n1880, B1 => n201, B2 => n1881,
                           ZN => n2571);
   U1552 : OAI22_X1 port map( A1 => n297, A2 => n39, B1 => n265, B2 => n41, ZN 
                           => n2570);
   U1553 : NAND2_X1 port map( A1 => n2577, A2 => n2574, ZN => n1883);
   U1554 : OAI22_X1 port map( A1 => n361, A2 => n43, B1 => n329, B2 => n45, ZN 
                           => n2569);
   U1555 : NAND2_X1 port map( A1 => n2578, A2 => n2574, ZN => n1885);
   U1556 : NOR3_X1 port map( A1 => n2559, A2 => n2579, A3 => n2580, ZN => n2574
                           );
   U1557 : NAND2_X1 port map( A1 => ADD_RD1(4), A2 => ADD_RD1(3), ZN => n2581);
   U1558 : NOR4_X1 port map( A1 => n2582, A2 => n2583, A3 => n2584, A4 => n2585
                           , ZN => n2567_port);
   U1559 : OAI22_X1 port map( A1 => n425, A2 => n1890, B1 => n393, B2 => n1891,
                           ZN => n2585);
   U1560 : OAI22_X1 port map( A1 => n492, A2 => n1892, B1 => n458, B2 => n1893,
                           ZN => n2584);
   U1561 : OAI22_X1 port map( A1 => n559, A2 => n1894, B1 => n526, B2 => n1895,
                           ZN => n2583);
   U1562 : OAI22_X1 port map( A1 => n626, A2 => n1896, B1 => n593, B2 => n1897,
                           ZN => n2582);
   U1563 : NOR3_X1 port map( A1 => ADD_RD1(3), A2 => n2559, A3 => n2580, ZN => 
                           n2586);
   U1564 : NOR3_X1 port map( A1 => ADD_RD1(3), A2 => ADD_RD1(0), A3 => n2559, 
                           ZN => n2587);
   U1565 : NOR4_X1 port map( A1 => n2588, A2 => n2589, A3 => n2590, A4 => n2591
                           , ZN => n2566);
   U1566 : OAI22_X1 port map( A1 => n694, A2 => n1902, B1 => n660, B2 => n1903,
                           ZN => n2591);
   U1567 : OAI22_X1 port map( A1 => n761, A2 => n1904, B1 => n727, B2 => n1905,
                           ZN => n2590);
   U1568 : OAI22_X1 port map( A1 => n828, A2 => n1906, B1 => n794, B2 => n1907,
                           ZN => n2589);
   U1569 : OAI22_X1 port map( A1 => n895, A2 => n1908, B1 => n862, B2 => n1909,
                           ZN => n2588);
   U1570 : NOR3_X1 port map( A1 => ADD_RD1(4), A2 => n2579, A3 => n2580, ZN => 
                           n2592);
   U1571 : NOR3_X1 port map( A1 => ADD_RD1(4), A2 => ADD_RD1(0), A3 => n2579, 
                           ZN => n2593);
   U1572 : NOR4_X1 port map( A1 => n2594, A2 => n2595, A3 => n2596, A4 => n2597
                           , ZN => n2565);
   U1573 : OAI22_X1 port map( A1 => n962, A2 => n1914, B1 => n929, B2 => n1915,
                           ZN => n2597);
   U1574 : OAI22_X1 port map( A1 => n1030, A2 => n1916, B1 => n996, B2 => n1917
                           , ZN => n2596);
   U1575 : OAI22_X1 port map( A1 => n1098, A2 => n1918, B1 => n1063, B2 => 
                           n1919, ZN => n2595);
   U1576 : OAI22_X1 port map( A1 => n144, A2 => n1920, B1 => n108, B2 => n1921,
                           ZN => n2594);
   U1577 : NOR3_X1 port map( A1 => ADD_RD1(4), A2 => ADD_RD1(3), A3 => n2580, 
                           ZN => n2598);
   U1578 : NOR3_X1 port map( A1 => ADD_RD1(4), A2 => ADD_RD1(3), A3 => 
                           ADD_RD1(0), ZN => n2599);
   U1579 : OAI21_X1 port map( B1 => n2600, B2 => n2601, A => n47, ZN => N4423);
   U1580 : OAI21_X1 port map( B1 => n2601, B2 => n2602, A => n47, ZN => N4359);
   U1581 : OAI21_X1 port map( B1 => n2601, B2 => n2603, A => n47, ZN => N4295);
   U1582 : OAI21_X1 port map( B1 => n2601, B2 => n2604, A => n47, ZN => N4231);
   U1583 : OAI21_X1 port map( B1 => n2601, B2 => n2605, A => n47, ZN => N4167);
   U1584 : OAI21_X1 port map( B1 => n2601, B2 => n2606, A => n47, ZN => N4103);
   U1585 : OAI21_X1 port map( B1 => n2601, B2 => n2607, A => n47, ZN => N4039);
   U1586 : NAND2_X1 port map( A1 => n2562, A2 => WR, ZN => n2601);
   U1587 : OAI21_X1 port map( B1 => n2564, B2 => n2608, A => n53, ZN => N3975);
   U1588 : OAI21_X1 port map( B1 => n2600, B2 => n2608, A => n47, ZN => N3911);
   U1589 : OAI21_X1 port map( B1 => n2608, B2 => n2602, A => n53, ZN => N3847);
   U1590 : OAI21_X1 port map( B1 => n2608, B2 => n2603, A => n53, ZN => N3783);
   U1591 : OAI21_X1 port map( B1 => n2608, B2 => n2604, A => n53, ZN => N3719);
   U1592 : OAI21_X1 port map( B1 => n2608, B2 => n2605, A => n53, ZN => N3655);
   U1593 : OAI21_X1 port map( B1 => n2608, B2 => n2606, A => n53, ZN => N3591);
   U1594 : OAI21_X1 port map( B1 => n2608, B2 => n2607, A => n53, ZN => N3527);
   U1595 : INV_X1 port map( A => WR, ZN => n2563);
   U1596 : OAI21_X1 port map( B1 => n2564, B2 => n2609, A => n53, ZN => N3463);
   U1597 : OAI21_X1 port map( B1 => n2600, B2 => n2609, A => n53, ZN => N3399);
   U1598 : OAI21_X1 port map( B1 => n2609, B2 => n2602, A => n53, ZN => N3335);
   U1599 : OAI21_X1 port map( B1 => n2609, B2 => n2603, A => n49, ZN => N3271);
   U1600 : OAI21_X1 port map( B1 => n2609, B2 => n2604, A => n53, ZN => N3207);
   U1601 : OAI21_X1 port map( B1 => n2609, B2 => n2605, A => n47, ZN => N3143);
   U1602 : OAI21_X1 port map( B1 => n2609, B2 => n2606, A => n51, ZN => N3079);
   U1603 : OAI21_X1 port map( B1 => n2609, B2 => n2607, A => n49, ZN => N3015);
   U1604 : NAND3_X1 port map( A1 => ADD_WR(4), A2 => WR, A3 => n1830, ZN => 
                           n2609);
   U1605 : OAI21_X1 port map( B1 => n2564, B2 => n2610, A => n53, ZN => N2951);
   U1606 : OAI21_X1 port map( B1 => n2600, B2 => n2610, A => n47, ZN => N2887);
   U1607 : NAND3_X1 port map( A1 => ADD_WR(0), A2 => n1826, A3 => n1824, ZN => 
                           n2600);
   U1608 : OAI21_X1 port map( B1 => n2610, B2 => n2602, A => n53, ZN => N2823);
   U1609 : NAND3_X1 port map( A1 => ADD_WR(1), A2 => n1827, A3 => n1826, ZN => 
                           n2602);
   U1610 : OAI21_X1 port map( B1 => n2610, B2 => n2603, A => n47, ZN => N2759);
   U1611 : NAND3_X1 port map( A1 => ADD_WR(0), A2 => ADD_WR(1), A3 => n1826, ZN
                           => n2603);
   U1612 : OAI21_X1 port map( B1 => n2610, B2 => n2604, A => n53, ZN => N2695);
   U1613 : NAND3_X1 port map( A1 => ADD_WR(2), A2 => n1827, A3 => n1824, ZN => 
                           n2604);
   U1614 : OAI21_X1 port map( B1 => n2610, B2 => n2605, A => n47, ZN => N2631);
   U1615 : NAND3_X1 port map( A1 => ADD_WR(2), A2 => ADD_WR(0), A3 => n1824, ZN
                           => n2605);
   U1616 : OAI21_X1 port map( B1 => n2610, B2 => n2606, A => n53, ZN => N2567);
   U1617 : NAND3_X1 port map( A1 => ADD_WR(2), A2 => ADD_WR(1), A3 => n1827, ZN
                           => n2606);
   U1618 : OAI21_X1 port map( B1 => n2610, B2 => n2607, A => n47, ZN => N2503);
   U1619 : NAND3_X1 port map( A1 => ADD_WR(0), A2 => ADD_WR(2), A3 => ADD_WR(1)
                           , ZN => n2607);
   U1620 : NAND3_X1 port map( A1 => ADD_WR(4), A2 => ADD_WR(3), A3 => WR, ZN =>
                           n2610);

end SYN_A;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity 
   dlx_cu_MICROCODE_MEM_SIZE64_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE13 is

   port( Clk, Rst : in std_logic;  IR_IN : in std_logic_vector (31 downto 0);  
         stall_exe_i, mispredict_i : in std_logic;  D1_i, D2_i : in 
         std_logic_vector (4 downto 0);  S1_LATCH_EN, S2_LATCH_EN, S3_LATCH_EN 
         : out std_logic;  S_MUX_PC_BUS : out std_logic_vector (1 downto 0);  
         S_EXT, S_EXT_SIGN, S_EQ_NEQ : out std_logic;  S_MUX_DEST : out 
         std_logic_vector (1 downto 0);  S_MUX_LINK, S_MUX_MEM, S_MEM_W_R, 
         S_MEM_EN, S_RF_W_wb, S_RF_W_mem, S_RF_W_exe, S_MUX_ALUIN, stall_exe_o,
         stall_dec_o, stall_fetch_o, stall_btb_o, was_branch_o, was_jmp_o : out
         std_logic;  ALU_WORD_o : out std_logic_vector (12 downto 0);  
         ALU_OPCODE : out std_logic_vector (0 to 4));

end dlx_cu_MICROCODE_MEM_SIZE64_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE13;

architecture SYN_dlx_cu_hw of 
   dlx_cu_MICROCODE_MEM_SIZE64_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE13 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X2
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component 
      SNPS_CLOCK_GATE_HIGH_dlx_cu_MICROCODE_MEM_SIZE64_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE13_0
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component alu_ctrl
      port( OP : in std_logic_vector (0 to 4);  ALU_WORD : out std_logic_vector
            (12 downto 0));
   end component;
   
   component cw_mem_MICROCODE_MEM_SIZE64_OP_CODE_SIZE6_CW_SIZE13
      port( OPCODE_IN : in std_logic_vector (5 downto 0);  CW_OUT : out 
            std_logic_vector (12 downto 0));
   end component;
   
   component stall_logic_FUNC_SIZE11_OP_CODE_SIZE6
      port( OPCODE_i : in std_logic_vector (5 downto 0);  FUNC_i : in 
            std_logic_vector (10 downto 0);  rA_i, rB_i, D1_i, D2_i : in 
            std_logic_vector (4 downto 0);  S_mem_LOAD_i, S_exe_LOAD_i, 
            S_exe_WRITE_i : in std_logic;  S_MUX_PC_BUS_i : in std_logic_vector
            (1 downto 0);  mispredict_i : in std_logic;  bubble_dec_o, 
            bubble_exe_o, stall_exe_o, stall_dec_o, stall_btb_o, stall_fetch_o 
            : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFS_X1
      port( D, CK, SN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal S_MUX_PC_BUS_1_port, S_MUX_PC_BUS_0_port, S_MEM_W_R_port, n122, 
      S_MEM_LOAD, S_EXE_LOAD, next_bubble_dec, stall_dec_o_TEMP, 
      stall_btb_o_TEMP, stall_fetch_o_TEMP, cw_from_mem_12_port, 
      cw_from_mem_11_port, cw_from_mem_10_port, cw_from_mem_9_port, 
      cw_from_mem_8_port, cw_from_mem_7_port, cw_from_mem_6_port, 
      cw_from_mem_5_port, cw_from_mem_4_port, cw_from_mem_3_port, 
      cw_from_mem_2_port, cw_from_mem_1_port, cw_from_mem_0_port, 
      aluOpcode_d_4_port, aluOpcode_d_3_port, aluOpcode_d_2_port, 
      aluOpcode_d_1_port, aluOpcode_d_0_port, N20, N21, N22, N23, N24, N25, N26
      , N27, N29, N30, N31, N32, net199583, n2, n3, n4, n5, n8, n9, n10, n11, 
      n12, n13, n14, n15, n16, n17, n18, n19, n20_port, n21_port, n22_port, 
      n23_port, n24_port, n25_port, n26_port, n27_port, n28, n29_port, n30_port
      , n31_port, n32_port, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, 
      n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57
      , n58, n59, n60, n61, n65, n70, n71, n72, n74, n75, n76, n77, n78, n79, 
      n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94
      , n95, n96, n97, n98, n99, n101, n102, n103, n110, n111, n113, n114, n115
      , n1, n6, n7, n62, n63, n64, n66, n67, n68, n69, n73, n100, n104, n105, 
      n106, n107, n108, n109, n112, n116, n117, n118, n119, n120, n121, 
      net245093, net245094, net245095, net245096, net245097, net245098 : 
      std_logic;

begin
   S_MUX_PC_BUS <= ( S_MUX_PC_BUS_1_port, S_MUX_PC_BUS_0_port );
   S_MEM_W_R <= S_MEM_W_R_port;
   stall_exe_o <= stall_exe_i;
   
   bubble_dec_reg : DFF_X1 port map( D => n113, CK => Clk, Q => n73, QN => n114
                           );
   cw_e_reg_0_inst : DFFR_X1 port map( D => N21, CK => net199583, RN => n100, Q
                           => n122, QN => n2);
   cw_e_reg_5_inst : DFFR_X1 port map( D => N26, CK => net199583, RN => n100, Q
                           => S_MUX_DEST(1), QN => n111);
   cw_e_reg_4_inst : DFFR_X1 port map( D => N25, CK => net199583, RN => n100, Q
                           => S_MUX_DEST(0), QN => n110);
   cw_e_reg_3_inst : DFFR_X1 port map( D => N24, CK => net199583, RN => n100, Q
                           => n3, QN => net245098);
   cw_e_reg_2_inst : DFFR_X1 port map( D => N23, CK => net199583, RN => n100, Q
                           => net245097, QN => n4);
   cw_e_reg_1_inst : DFFR_X1 port map( D => N22, CK => net199583, RN => n100, Q
                           => net245096, QN => n5);
   cw_m_reg_2_inst : DFFR_X1 port map( D => N31, CK => Clk, RN => n100, Q => 
                           S_MEM_W_R_port, QN => net245095);
   cw_m_reg_3_inst : DFFR_X1 port map( D => N32, CK => Clk, RN => n100, Q => 
                           S_MEM_EN, QN => n115);
   cw_m_reg_0_inst : DFFR_X1 port map( D => N29, CK => Clk, RN => n100, Q => 
                           S_RF_W_mem, QN => n103);
   cw_w_reg_0_inst : DFFS_X1 port map( D => n103, CK => Clk, SN => n100, Q => 
                           n102, QN => S_RF_W_wb);
   U3 : XOR2_X1 port map( A => S_MUX_PC_BUS_1_port, B => S_MUX_PC_BUS_0_port, Z
                           => was_jmp_o);
   U8 : MUX2_X1 port map( A => n73, B => next_bubble_dec, S => n100, Z => n113)
                           ;
   U13 : NAND3_X1 port map( A1 => n19, A2 => IR_IN(28), A3 => n20_port, ZN => 
                           n18);
   U24 : NAND3_X1 port map( A1 => n34, A2 => n43, A3 => n21_port, ZN => n42);
   U60 : NAND3_X1 port map( A1 => IR_IN(30), A2 => IR_IN(29), A3 => n72, ZN => 
                           n58);
   U78 : NAND3_X1 port map( A1 => IR_IN(5), A2 => IR_IN(4), A3 => n61, ZN => 
                           n54);
   U92 : NAND3_X1 port map( A1 => n97, A2 => n93, A3 => n21_port, ZN => n41);
   STALL_L : stall_logic_FUNC_SIZE11_OP_CODE_SIZE6 port map( OPCODE_i(5) => 
                           IR_IN(31), OPCODE_i(4) => IR_IN(30), OPCODE_i(3) => 
                           IR_IN(29), OPCODE_i(2) => IR_IN(28), OPCODE_i(1) => 
                           IR_IN(27), OPCODE_i(0) => IR_IN(26), FUNC_i(10) => 
                           n104, FUNC_i(9) => n105, FUNC_i(8) => n106, 
                           FUNC_i(7) => n107, FUNC_i(6) => n108, FUNC_i(5) => 
                           n109, FUNC_i(4) => n112, FUNC_i(3) => n116, 
                           FUNC_i(2) => n117, FUNC_i(1) => n118, FUNC_i(0) => 
                           n119, rA_i(4) => IR_IN(25), rA_i(3) => IR_IN(24), 
                           rA_i(2) => IR_IN(23), rA_i(1) => IR_IN(22), rA_i(0) 
                           => IR_IN(21), rB_i(4) => IR_IN(20), rB_i(3) => 
                           IR_IN(19), rB_i(2) => IR_IN(18), rB_i(1) => 
                           IR_IN(17), rB_i(0) => IR_IN(16), D1_i(4) => D1_i(4),
                           D1_i(3) => D1_i(3), D1_i(2) => D1_i(2), D1_i(1) => 
                           D1_i(1), D1_i(0) => D1_i(0), D2_i(4) => D2_i(4), 
                           D2_i(3) => D2_i(3), D2_i(2) => D2_i(2), D2_i(1) => 
                           D2_i(1), D2_i(0) => D2_i(0), S_mem_LOAD_i => 
                           S_MEM_LOAD, S_exe_LOAD_i => S_EXE_LOAD, 
                           S_exe_WRITE_i => n122, S_MUX_PC_BUS_i(1) => n120, 
                           S_MUX_PC_BUS_i(0) => n121, mispredict_i => 
                           mispredict_i, bubble_dec_o => next_bubble_dec, 
                           bubble_exe_o => net245093, stall_exe_o => net245094,
                           stall_dec_o => stall_dec_o_TEMP, stall_btb_o => 
                           stall_btb_o_TEMP, stall_fetch_o => 
                           stall_fetch_o_TEMP);
   CWM : cw_mem_MICROCODE_MEM_SIZE64_OP_CODE_SIZE6_CW_SIZE13 port map( 
                           OPCODE_IN(5) => IR_IN(31), OPCODE_IN(4) => IR_IN(30)
                           , OPCODE_IN(3) => IR_IN(29), OPCODE_IN(2) => 
                           IR_IN(28), OPCODE_IN(1) => IR_IN(27), OPCODE_IN(0) 
                           => IR_IN(26), CW_OUT(12) => cw_from_mem_12_port, 
                           CW_OUT(11) => cw_from_mem_11_port, CW_OUT(10) => 
                           cw_from_mem_10_port, CW_OUT(9) => cw_from_mem_9_port
                           , CW_OUT(8) => cw_from_mem_8_port, CW_OUT(7) => 
                           cw_from_mem_7_port, CW_OUT(6) => cw_from_mem_6_port,
                           CW_OUT(5) => cw_from_mem_5_port, CW_OUT(4) => 
                           cw_from_mem_4_port, CW_OUT(3) => cw_from_mem_3_port,
                           CW_OUT(2) => cw_from_mem_2_port, CW_OUT(1) => 
                           cw_from_mem_1_port, CW_OUT(0) => cw_from_mem_0_port)
                           ;
   ALU_C : alu_ctrl port map( OP(0) => aluOpcode_d_4_port, OP(1) => 
                           aluOpcode_d_3_port, OP(2) => aluOpcode_d_2_port, 
                           OP(3) => aluOpcode_d_1_port, OP(4) => 
                           aluOpcode_d_0_port, ALU_WORD(12) => ALU_WORD_o(12), 
                           ALU_WORD(11) => ALU_WORD_o(11), ALU_WORD(10) => 
                           ALU_WORD_o(10), ALU_WORD(9) => ALU_WORD_o(9), 
                           ALU_WORD(8) => ALU_WORD_o(8), ALU_WORD(7) => 
                           ALU_WORD_o(7), ALU_WORD(6) => ALU_WORD_o(6), 
                           ALU_WORD(5) => ALU_WORD_o(5), ALU_WORD(4) => 
                           ALU_WORD_o(4), ALU_WORD(3) => ALU_WORD_o(3), 
                           ALU_WORD(2) => ALU_WORD_o(2), ALU_WORD(1) => 
                           ALU_WORD_o(1), ALU_WORD(0) => ALU_WORD_o(0));
   clk_gate_cw_e_reg : 
                           SNPS_CLOCK_GATE_HIGH_dlx_cu_MICROCODE_MEM_SIZE64_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE13_0 
                           port map( CLK => Clk, EN => N20, ENCLK => net199583)
                           ;
   U114 : AND2_X1 port map( A1 => n114, A2 => cw_from_mem_8_port, ZN => 
                           S_EQ_NEQ);
   U109 : NOR2_X1 port map( A1 => n115, A2 => S_MEM_W_R_port, ZN => S_MEM_LOAD)
                           ;
   U47 : NAND2_X1 port map( A1 => IR_IN(4), A2 => IR_IN(5), ZN => n8);
   U96 : NAND2_X1 port map( A1 => n89, A2 => n99, ZN => n98);
   U95 : NOR4_X1 port map( A1 => IR_IN(9), A2 => IR_IN(8), A3 => IR_IN(29), A4 
                           => n98, ZN => n92);
   U94 : NAND2_X1 port map( A1 => n44, A2 => n92, ZN => n49);
   U74 : NOR3_X1 port map( A1 => IR_IN(5), A2 => n39, A3 => n75, ZN => n82);
   U73 : NAND4_X1 port map( A1 => n92, A2 => IR_IN(26), A3 => n82, A4 => n61, 
                           ZN => n47);
   U26 : AOI221_X1 port map( B1 => IR_IN(4), B2 => IR_IN(3), C1 => n45, C2 => 
                           n46, A => n47, ZN => n29_port);
   U70 : NOR2_X1 port map( A1 => n39, A2 => IR_IN(1), ZN => n60);
   U68 : NOR2_X1 port map( A1 => n46, A2 => n25_port, ZN => n34);
   U20 : NAND2_X1 port map( A1 => n21_port, A2 => n34, ZN => n15);
   U100 : NOR3_X1 port map( A1 => IR_IN(2), A2 => n46, A3 => n75, ZN => n93);
   U77 : NAND2_X1 port map( A1 => n21_port, A2 => n93, ZN => n31_port);
   U85 : NAND2_X1 port map( A1 => IR_IN(30), A2 => IR_IN(29), ZN => n96);
   U19 : OAI21_X1 port map( B1 => n12, B2 => n33, A => IR_IN(31), ZN => 
                           n32_port);
   U18 : OAI221_X1 port map( B1 => n8, B2 => n15, C1 => n8, C2 => n31_port, A 
                           => n32_port, ZN => n30_port);
   U17 : NOR2_X1 port map( A1 => n29_port, A2 => n30_port, ZN => n10);
   U56 : NOR2_X1 port map( A1 => n61, A2 => n26_port, ZN => n14);
   U10 : AOI22_X1 port map( A1 => IR_IN(26), A2 => n12, B1 => n13, B2 => n14, 
                           ZN => n11);
   U9 : OAI211_X1 port map( C1 => n8, C2 => n9, A => n10, B => n11, ZN => 
                           aluOpcode_d_4_port);
   U91 : INV_X1 port map( A => IR_IN(31), ZN => n55);
   U90 : NAND2_X1 port map( A1 => IR_IN(29), A2 => n55, ZN => n56);
   U48 : NOR2_X1 port map( A1 => IR_IN(0), A2 => n26_port, ZN => n43);
   U46 : NOR2_X1 port map( A1 => n8, A2 => n61, ZN => n50);
   U28 : OAI221_X1 port map( B1 => n43, B2 => IR_IN(1), C1 => n43, C2 => n50, A
                           => n46, ZN => n48);
   U27 : NOR2_X1 port map( A1 => n48, A2 => n49, ZN => n28);
   U16 : AOI22_X1 port map( A1 => IR_IN(30), A2 => n27_port, B1 => IR_IN(2), B2
                           => n28, ZN => n16);
   U71 : NOR4_X1 port map( A1 => IR_IN(1), A2 => IR_IN(2), A3 => n46, A4 => 
                           n26_port, ZN => n22_port);
   U15 : NOR3_X1 port map( A1 => n25_port, A2 => n26_port, A3 => n9, ZN => 
                           n23_port);
   U25 : AOI21_X1 port map( B1 => n12, B2 => n44, A => n33, ZN => n40);
   U23 : OAI211_X1 port map( C1 => n40, C2 => IR_IN(31), A => n41, B => n42, ZN
                           => n24_port);
   U14 : AOI211_X1 port map( C1 => n21_port, C2 => n22_port, A => n23_port, B 
                           => n24_port, ZN => n17);
   U89 : NOR2_X1 port map( A1 => IR_IN(30), A2 => n56, ZN => n19);
   U12 : NAND4_X1 port map( A1 => n10, A2 => n16, A3 => n17, A4 => n18, ZN => 
                           aluOpcode_d_3_port);
   U65 : NOR3_X1 port map( A1 => IR_IN(2), A2 => n61, A3 => n26_port, ZN => n59
                           );
   U36 : OAI221_X1 port map( B1 => n59, B2 => n60, C1 => n59, C2 => n50, A => 
                           n21_port, ZN => n35);
   U33 : OAI221_X1 port map( B1 => n27_port, B2 => IR_IN(31), C1 => n27_port, 
                           C2 => n12, A => IR_IN(26), ZN => n36);
   U31 : OAI21_X1 port map( B1 => n55, B2 => n20_port, A => n56, ZN => n52);
   U30 : NOR3_X1 port map( A1 => n39, A2 => n54, A3 => n9, ZN => n53);
   U29 : AOI21_X1 port map( B1 => n51, B2 => n52, A => n53, ZN => n37);
   U22 : AOI211_X1 port map( C1 => n28, C2 => n39, A => n29_port, B => n24_port
                           , ZN => n38);
   U83 : INV_X1 port map( A => IR_IN(29), ZN => n91);
   U80 : AOI221_X1 port map( B1 => n94, B2 => IR_IN(26), C1 => n33, C2 => n44, 
                           A => n95, ZN => n76);
   U76 : NOR2_X1 port map( A1 => n54, A2 => n31_port, ZN => n78);
   U72 : NOR3_X1 port map( A1 => IR_IN(3), A2 => n45, A3 => n47, ZN => n79);
   U67 : OAI221_X1 port map( B1 => n22_port, B2 => n34, C1 => n22_port, C2 => 
                           IR_IN(5), A => n61, ZN => n85);
   U64 : OAI211_X1 port map( C1 => n84, C2 => n59, A => IR_IN(1), B => n46, ZN 
                           => n86);
   U62 : NOR2_X1 port map( A1 => n91, A2 => n20_port, ZN => n88);
   U59 : AOI211_X1 port map( C1 => IR_IN(31), C2 => n57, A => IR_IN(26), B => 
                           n58, ZN => n90);
   U58 : AOI21_X1 port map( B1 => n88, B2 => n89, A => n90, ZN => n87);
   U57 : OAI221_X1 port map( B1 => n49, B2 => n85, C1 => n49, C2 => n86, A => 
                           n87, ZN => n65);
   U55 : NOR4_X1 port map( A1 => IR_IN(4), A2 => IR_IN(5), A3 => IR_IN(0), A4 
                           => n25_port, ZN => n83);
   U54 : AOI211_X1 port map( C1 => n14, C2 => n75, A => n83, B => n84, ZN => 
                           n81);
   U53 : NAND2_X1 port map( A1 => n82, A2 => n45, ZN => n74);
   U51 : AOI221_X1 port map( B1 => n61, B2 => n81, C1 => n74, C2 => n81, A => 
                           n9, ZN => n80);
   U50 : NOR4_X1 port map( A1 => n78, A2 => n79, A3 => n65, A4 => n80, ZN => 
                           n77);
   U49 : OAI211_X1 port map( C1 => IR_IN(0), C2 => n41, A => n76, B => n77, ZN 
                           => aluOpcode_d_0_port);
   U119 : NOR2_X1 port map( A1 => n2, A2 => stall_exe_i, ZN => N29);
   U117 : NOR2_X1 port map( A1 => n4, A2 => stall_exe_i, ZN => N31);
   U118 : NOR2_X1 port map( A1 => n5, A2 => stall_exe_i, ZN => N30);
   U52 : NAND2_X1 port map( A1 => n21_port, A2 => n46, ZN => n9);
   U34 : NOR2_X1 port map( A1 => n57, A2 => n58, ZN => n12);
   U104 : NAND2_X1 port map( A1 => IR_IN(5), A2 => n45, ZN => n26_port);
   U21 : NAND4_X1 port map( A1 => n35, A2 => n36, A3 => n37, A4 => n38, ZN => 
                           aluOpcode_d_2_port);
   U99 : INV_X1 port map( A => IR_IN(26), ZN => n44);
   U127 : NOR2_X1 port map( A1 => stall_dec_o_TEMP, A2 => n73, ZN => n101);
   U107 : AND2_X1 port map( A1 => n114, A2 => cw_from_mem_11_port, ZN => 
                           S_MUX_PC_BUS_0_port);
   U106 : AND2_X1 port map( A1 => cw_from_mem_12_port, A2 => n114, ZN => 
                           S_MUX_PC_BUS_1_port);
   cw_e_reg_6_inst : DFFR_X2 port map( D => N27, CK => net199583, RN => n100, Q
                           => S_MUX_ALUIN, QN => n69);
   U75 : INV_X1 port map( A => IR_IN(2), ZN => n39);
   U113 : AND2_X1 port map( A1 => n4, A2 => n3, ZN => S_EXE_LOAD);
   U101 : INV_X1 port map( A => IR_IN(1), ZN => n75);
   U79 : INV_X1 port map( A => IR_IN(0), ZN => n61);
   U105 : INV_X1 port map( A => IR_IN(4), ZN => n45);
   U102 : INV_X1 port map( A => IR_IN(3), ZN => n46);
   U66 : INV_X1 port map( A => n54, ZN => n84);
   U103 : INV_X1 port map( A => n26_port, ZN => n97);
   U69 : INV_X1 port map( A => n60, ZN => n25_port);
   U88 : INV_X1 port map( A => n19, ZN => n71);
   U93 : INV_X1 port map( A => n49, ZN => n21_port);
   U116 : AND2_X1 port map( A1 => N20, A2 => n3, ZN => N32);
   U11 : INV_X1 port map( A => n15, ZN => n13);
   U4 : AND2_X1 port map( A1 => S_MUX_PC_BUS_1_port, A2 => S_MUX_PC_BUS_0_port,
                           ZN => was_branch_o);
   U5 : OR2_X1 port map( A1 => stall_exe_i, A2 => stall_fetch_o_TEMP, ZN => 
                           stall_fetch_o);
   U6 : OR2_X1 port map( A1 => stall_exe_i, A2 => stall_dec_o_TEMP, ZN => 
                           stall_dec_o);
   U7 : OR2_X1 port map( A1 => stall_exe_i, A2 => stall_btb_o_TEMP, ZN => 
                           stall_btb_o);
   U125 : AND2_X1 port map( A1 => n101, A2 => cw_from_mem_1_port, ZN => N22);
   U124 : AND2_X1 port map( A1 => n101, A2 => cw_from_mem_2_port, ZN => N23);
   U121 : AND2_X1 port map( A1 => n101, A2 => cw_from_mem_5_port, ZN => N26);
   U122 : AND2_X1 port map( A1 => n101, A2 => cw_from_mem_4_port, ZN => N25);
   U126 : AND2_X1 port map( A1 => n101, A2 => cw_from_mem_0_port, ZN => N21);
   U123 : AND2_X1 port map( A1 => n101, A2 => cw_from_mem_3_port, ZN => N24);
   cw_m_reg_1_inst : DFFR_X2 port map( D => N30, CK => Clk, RN => n100, Q => 
                           S_MUX_MEM, QN => n68);
   U32 : OAI21_X1 port map( B1 => IR_IN(26), B2 => n71, A => n70, ZN => n1);
   U35 : INV_X1 port map( A => n72, ZN => n6);
   U37 : INV_X1 port map( A => n31_port, ZN => n7);
   U38 : AOI222_X1 port map( A1 => n1, A2 => n6, B1 => IR_IN(26), B2 => n33, C1
                           => n7, C2 => n50, ZN => n62);
   U39 : AOI22_X1 port map( A1 => IR_IN(1), A2 => n43, B1 => n50, B2 => n75, ZN
                           => n63);
   U40 : AOI21_X1 port map( B1 => n74, B2 => n63, A => n9, ZN => n64);
   U41 : NOR3_X1 port map( A1 => n46, A2 => n47, A3 => IR_IN(4), ZN => n66);
   U42 : NOR3_X1 port map( A1 => n65, A2 => n64, A3 => n66, ZN => n67);
   U43 : OAI211_X1 port map( C1 => n61, C2 => n41, A => n62, B => n67, ZN => 
                           aluOpcode_d_1_port);
   U44 : INV_X1 port map( A => stall_exe_i, ZN => N20);
   U45 : AND2_X2 port map( A1 => n114, A2 => cw_from_mem_7_port, ZN => 
                           S_MUX_LINK);
   U61 : INV_X1 port map( A => Rst, ZN => n100);
   U63 : AND2_X1 port map( A1 => n101, A2 => cw_from_mem_6_port, ZN => N27);
   U81 : INV_X1 port map( A => IR_IN(27), ZN => n72);
   U82 : NOR2_X1 port map( A1 => IR_IN(28), A2 => n56, ZN => n27_port);
   U84 : AND2_X2 port map( A1 => cw_from_mem_10_port, A2 => n114, ZN => S_EXT);
   U86 : AOI221_X1 port map( B1 => IR_IN(27), B2 => n44, C1 => n72, C2 => 
                           IR_IN(26), A => n70, ZN => n95);
   U87 : AND2_X1 port map( A1 => cw_from_mem_9_port, A2 => n114, ZN => 
                           S_EXT_SIGN);
   U97 : NOR2_X1 port map( A1 => IR_IN(27), A2 => n71, ZN => n94);
   U98 : NAND2_X1 port map( A1 => IR_IN(26), A2 => IR_IN(27), ZN => n20_port);
   U108 : NOR4_X1 port map( A1 => IR_IN(7), A2 => IR_IN(6), A3 => IR_IN(27), A4
                           => IR_IN(10), ZN => n99);
   U110 : NOR3_X1 port map( A1 => IR_IN(31), A2 => IR_IN(28), A3 => IR_IN(30), 
                           ZN => n89);
   U111 : NOR3_X1 port map( A1 => IR_IN(28), A2 => n72, A3 => n96, ZN => n33);
   U112 : NAND4_X1 port map( A1 => IR_IN(28), A2 => IR_IN(30), A3 => n55, A4 =>
                           n91, ZN => n70);
   U115 : INV_X1 port map( A => IR_IN(28), ZN => n57);
   U120 : NOR2_X1 port map( A1 => IR_IN(28), A2 => IR_IN(30), ZN => n51);
   n104 <= '0';
   n105 <= '0';
   n106 <= '0';
   n107 <= '0';
   n108 <= '0';
   n109 <= '0';
   n112 <= '0';
   n116 <= '0';
   n117 <= '0';
   n118 <= '0';
   n119 <= '0';
   n120 <= '0';
   n121 <= '0';

end SYN_dlx_cu_hw;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity jump_logic is

   port( NPCF_i, IR_i, A_i : in std_logic_vector (31 downto 0);  A_o : out 
         std_logic_vector (31 downto 0);  rA_o, rB_o, rC_o : out 
         std_logic_vector (4 downto 0);  branch_target_o, sum_addr_o, 
         extended_imm : out std_logic_vector (31 downto 0);  taken_o : out 
         std_logic;  FW_X_i, FW_W_i : in std_logic_vector (31 downto 0);  
         S_FW_Adec_i : in std_logic_vector (1 downto 0);  S_EXT_i, S_EXT_SIGN_i
         , S_MUX_LINK_i, S_EQ_NEQ_i : in std_logic);

end jump_logic;

architecture SYN_struct of jump_logic is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component mux41_MUX_SIZE32_0
      port( IN0, IN1, IN2, IN3 : in std_logic_vector (31 downto 0);  CTRL : in 
            std_logic_vector (1 downto 0);  OUT1 : out std_logic_vector (31 
            downto 0));
   end component;
   
   component mux21_4
      port( IN0, IN1 : in std_logic_vector (31 downto 0);  CTRL : in std_logic;
            OUT1 : out std_logic_vector (31 downto 0));
   end component;
   
   component zerocheck
      port( IN0 : in std_logic_vector (31 downto 0);  CTRL : in std_logic;  
            OUT1 : out std_logic);
   end component;
   
   component mux21_0
      port( IN0, IN1 : in std_logic_vector (31 downto 0);  CTRL : in std_logic;
            OUT1 : out std_logic_vector (31 downto 0));
   end component;
   
   component p4add_N32_logN5_0
      port( A, B : in std_logic_vector (31 downto 0);  Cin, sign : in std_logic
            ;  S : out std_logic_vector (31 downto 0);  Cout : out std_logic);
   end component;
   
   component extender_32
      port( IN1 : in std_logic_vector (31 downto 0);  CTRL, SIGN : in std_logic
            ;  OUT1 : out std_logic_vector (31 downto 0));
   end component;
   
   signal X_Logic0_port, A_o_31_port, A_o_30_port, A_o_29_port, A_o_28_port, 
      A_o_27_port, A_o_26_port, A_o_25_port, A_o_24_port, A_o_23_port, 
      A_o_22_port, A_o_21_port, A_o_20_port, A_o_19_port, A_o_18_port, 
      A_o_17_port, A_o_16_port, A_o_15_port, A_o_14_port, A_o_13_port, 
      A_o_12_port, A_o_11_port, A_o_10_port, A_o_9_port, A_o_8_port, A_o_7_port
      , A_o_6_port, A_o_5_port, A_o_4_port, A_o_3_port, A_o_2_port, A_o_1_port,
      A_o_0_port, sum_addr_o_31_port, sum_addr_o_30_port, sum_addr_o_29_port, 
      sum_addr_o_28_port, sum_addr_o_27_port, sum_addr_o_26_port, 
      sum_addr_o_25_port, sum_addr_o_24_port, sum_addr_o_23_port, 
      sum_addr_o_22_port, sum_addr_o_21_port, sum_addr_o_20_port, 
      sum_addr_o_19_port, sum_addr_o_18_port, sum_addr_o_17_port, 
      sum_addr_o_16_port, sum_addr_o_15_port, sum_addr_o_14_port, 
      sum_addr_o_13_port, sum_addr_o_12_port, sum_addr_o_11_port, 
      sum_addr_o_10_port, sum_addr_o_9_port, sum_addr_o_8_port, 
      sum_addr_o_7_port, sum_addr_o_6_port, sum_addr_o_5_port, 
      sum_addr_o_4_port, sum_addr_o_3_port, sum_addr_o_2_port, 
      sum_addr_o_1_port, sum_addr_o_0_port, ext_imm_31_port, ext_imm_30_port, 
      ext_imm_28_port, ext_imm_26_port, ext_imm_24_port, ext_imm_23_port, 
      ext_imm_22_port, ext_imm_21_port, ext_imm_20_port, ext_imm_19_port, 
      ext_imm_18_port, ext_imm_17_port, ext_imm_16_port, ext_imm_15_port, 
      ext_imm_14_port, ext_imm_13_port, ext_imm_12_port, ext_imm_11_port, 
      ext_imm_10_port, ext_imm_9_port, ext_imm_8_port, ext_imm_7_port, 
      ext_imm_6_port, ext_imm_5_port, ext_imm_4_port, ext_imm_3_port, 
      ext_imm_2_port, ext_imm_1_port, ext_imm_0_port, branch_sel, n1, n2, n3, 
      n6, n7, n8, n9, n10, n11, net245092 : std_logic;

begin
   A_o <= ( A_o_31_port, A_o_30_port, A_o_29_port, A_o_28_port, A_o_27_port, 
      A_o_26_port, A_o_25_port, A_o_24_port, A_o_23_port, A_o_22_port, 
      A_o_21_port, A_o_20_port, A_o_19_port, A_o_18_port, A_o_17_port, 
      A_o_16_port, A_o_15_port, A_o_14_port, A_o_13_port, A_o_12_port, 
      A_o_11_port, A_o_10_port, A_o_9_port, A_o_8_port, A_o_7_port, A_o_6_port,
      A_o_5_port, A_o_4_port, A_o_3_port, A_o_2_port, A_o_1_port, A_o_0_port );
   rA_o <= ( IR_i(25), IR_i(24), IR_i(23), IR_i(22), IR_i(21) );
   rB_o <= ( IR_i(20), IR_i(19), IR_i(18), IR_i(17), IR_i(16) );
   rC_o <= ( IR_i(15), IR_i(14), IR_i(13), IR_i(12), IR_i(11) );
   sum_addr_o <= ( sum_addr_o_31_port, sum_addr_o_30_port, sum_addr_o_29_port, 
      sum_addr_o_28_port, sum_addr_o_27_port, sum_addr_o_26_port, 
      sum_addr_o_25_port, sum_addr_o_24_port, sum_addr_o_23_port, 
      sum_addr_o_22_port, sum_addr_o_21_port, sum_addr_o_20_port, 
      sum_addr_o_19_port, sum_addr_o_18_port, sum_addr_o_17_port, 
      sum_addr_o_16_port, sum_addr_o_15_port, sum_addr_o_14_port, 
      sum_addr_o_13_port, sum_addr_o_12_port, sum_addr_o_11_port, 
      sum_addr_o_10_port, sum_addr_o_9_port, sum_addr_o_8_port, 
      sum_addr_o_7_port, sum_addr_o_6_port, sum_addr_o_5_port, 
      sum_addr_o_4_port, sum_addr_o_3_port, sum_addr_o_2_port, 
      sum_addr_o_1_port, sum_addr_o_0_port );
   
   X_Logic0_port <= '0';
   EXTENDER : extender_32 port map( IN1(31) => n6, IN1(30) => n7, IN1(29) => n8
                           , IN1(28) => n9, IN1(27) => n10, IN1(26) => n11, 
                           IN1(25) => IR_i(25), IN1(24) => IR_i(24), IN1(23) =>
                           IR_i(23), IN1(22) => IR_i(22), IN1(21) => IR_i(21), 
                           IN1(20) => IR_i(20), IN1(19) => IR_i(19), IN1(18) =>
                           IR_i(18), IN1(17) => IR_i(17), IN1(16) => IR_i(16), 
                           IN1(15) => IR_i(15), IN1(14) => IR_i(14), IN1(13) =>
                           IR_i(13), IN1(12) => IR_i(12), IN1(11) => IR_i(11), 
                           IN1(10) => IR_i(10), IN1(9) => IR_i(9), IN1(8) => 
                           IR_i(8), IN1(7) => IR_i(7), IN1(6) => IR_i(6), 
                           IN1(5) => IR_i(5), IN1(4) => IR_i(4), IN1(3) => 
                           IR_i(3), IN1(2) => IR_i(2), IN1(1) => IR_i(1), 
                           IN1(0) => IR_i(0), CTRL => S_EXT_i, SIGN => 
                           S_EXT_SIGN_i, OUT1(31) => ext_imm_31_port, OUT1(30) 
                           => ext_imm_30_port, OUT1(29) => n3, OUT1(28) => 
                           ext_imm_28_port, OUT1(27) => n2, OUT1(26) => 
                           ext_imm_26_port, OUT1(25) => n1, OUT1(24) => 
                           ext_imm_24_port, OUT1(23) => ext_imm_23_port, 
                           OUT1(22) => ext_imm_22_port, OUT1(21) => 
                           ext_imm_21_port, OUT1(20) => ext_imm_20_port, 
                           OUT1(19) => ext_imm_19_port, OUT1(18) => 
                           ext_imm_18_port, OUT1(17) => ext_imm_17_port, 
                           OUT1(16) => ext_imm_16_port, OUT1(15) => 
                           ext_imm_15_port, OUT1(14) => ext_imm_14_port, 
                           OUT1(13) => ext_imm_13_port, OUT1(12) => 
                           ext_imm_12_port, OUT1(11) => ext_imm_11_port, 
                           OUT1(10) => ext_imm_10_port, OUT1(9) => 
                           ext_imm_9_port, OUT1(8) => ext_imm_8_port, OUT1(7) 
                           => ext_imm_7_port, OUT1(6) => ext_imm_6_port, 
                           OUT1(5) => ext_imm_5_port, OUT1(4) => ext_imm_4_port
                           , OUT1(3) => ext_imm_3_port, OUT1(2) => 
                           ext_imm_2_port, OUT1(1) => ext_imm_1_port, OUT1(0) 
                           => ext_imm_0_port);
   JUMPADDER : p4add_N32_logN5_0 port map( A(31) => NPCF_i(31), A(30) => 
                           NPCF_i(30), A(29) => NPCF_i(29), A(28) => NPCF_i(28)
                           , A(27) => NPCF_i(27), A(26) => NPCF_i(26), A(25) =>
                           NPCF_i(25), A(24) => NPCF_i(24), A(23) => NPCF_i(23)
                           , A(22) => NPCF_i(22), A(21) => NPCF_i(21), A(20) =>
                           NPCF_i(20), A(19) => NPCF_i(19), A(18) => NPCF_i(18)
                           , A(17) => NPCF_i(17), A(16) => NPCF_i(16), A(15) =>
                           NPCF_i(15), A(14) => NPCF_i(14), A(13) => NPCF_i(13)
                           , A(12) => NPCF_i(12), A(11) => NPCF_i(11), A(10) =>
                           NPCF_i(10), A(9) => NPCF_i(9), A(8) => NPCF_i(8), 
                           A(7) => NPCF_i(7), A(6) => NPCF_i(6), A(5) => 
                           NPCF_i(5), A(4) => NPCF_i(4), A(3) => NPCF_i(3), 
                           A(2) => NPCF_i(2), A(1) => NPCF_i(1), A(0) => 
                           NPCF_i(0), B(31) => ext_imm_31_port, B(30) => 
                           ext_imm_30_port, B(29) => n3, B(28) => 
                           ext_imm_28_port, B(27) => n2, B(26) => 
                           ext_imm_26_port, B(25) => n1, B(24) => 
                           ext_imm_24_port, B(23) => ext_imm_23_port, B(22) => 
                           ext_imm_22_port, B(21) => ext_imm_21_port, B(20) => 
                           ext_imm_20_port, B(19) => ext_imm_19_port, B(18) => 
                           ext_imm_18_port, B(17) => ext_imm_17_port, B(16) => 
                           ext_imm_16_port, B(15) => ext_imm_15_port, B(14) => 
                           ext_imm_14_port, B(13) => ext_imm_13_port, B(12) => 
                           ext_imm_12_port, B(11) => ext_imm_11_port, B(10) => 
                           ext_imm_10_port, B(9) => ext_imm_9_port, B(8) => 
                           ext_imm_8_port, B(7) => ext_imm_7_port, B(6) => 
                           ext_imm_6_port, B(5) => ext_imm_5_port, B(4) => 
                           ext_imm_4_port, B(3) => ext_imm_3_port, B(2) => 
                           ext_imm_2_port, B(1) => ext_imm_1_port, B(0) => 
                           ext_imm_0_port, Cin => X_Logic0_port, sign => 
                           X_Logic0_port, S(31) => sum_addr_o_31_port, S(30) =>
                           sum_addr_o_30_port, S(29) => sum_addr_o_29_port, 
                           S(28) => sum_addr_o_28_port, S(27) => 
                           sum_addr_o_27_port, S(26) => sum_addr_o_26_port, 
                           S(25) => sum_addr_o_25_port, S(24) => 
                           sum_addr_o_24_port, S(23) => sum_addr_o_23_port, 
                           S(22) => sum_addr_o_22_port, S(21) => 
                           sum_addr_o_21_port, S(20) => sum_addr_o_20_port, 
                           S(19) => sum_addr_o_19_port, S(18) => 
                           sum_addr_o_18_port, S(17) => sum_addr_o_17_port, 
                           S(16) => sum_addr_o_16_port, S(15) => 
                           sum_addr_o_15_port, S(14) => sum_addr_o_14_port, 
                           S(13) => sum_addr_o_13_port, S(12) => 
                           sum_addr_o_12_port, S(11) => sum_addr_o_11_port, 
                           S(10) => sum_addr_o_10_port, S(9) => 
                           sum_addr_o_9_port, S(8) => sum_addr_o_8_port, S(7) 
                           => sum_addr_o_7_port, S(6) => sum_addr_o_6_port, 
                           S(5) => sum_addr_o_5_port, S(4) => sum_addr_o_4_port
                           , S(3) => sum_addr_o_3_port, S(2) => 
                           sum_addr_o_2_port, S(1) => sum_addr_o_1_port, S(0) 
                           => sum_addr_o_0_port, Cout => net245092);
   BRANCHMUX : mux21_0 port map( IN0(31) => sum_addr_o_31_port, IN0(30) => 
                           sum_addr_o_30_port, IN0(29) => sum_addr_o_29_port, 
                           IN0(28) => sum_addr_o_28_port, IN0(27) => 
                           sum_addr_o_27_port, IN0(26) => sum_addr_o_26_port, 
                           IN0(25) => sum_addr_o_25_port, IN0(24) => 
                           sum_addr_o_24_port, IN0(23) => sum_addr_o_23_port, 
                           IN0(22) => sum_addr_o_22_port, IN0(21) => 
                           sum_addr_o_21_port, IN0(20) => sum_addr_o_20_port, 
                           IN0(19) => sum_addr_o_19_port, IN0(18) => 
                           sum_addr_o_18_port, IN0(17) => sum_addr_o_17_port, 
                           IN0(16) => sum_addr_o_16_port, IN0(15) => 
                           sum_addr_o_15_port, IN0(14) => sum_addr_o_14_port, 
                           IN0(13) => sum_addr_o_13_port, IN0(12) => 
                           sum_addr_o_12_port, IN0(11) => sum_addr_o_11_port, 
                           IN0(10) => sum_addr_o_10_port, IN0(9) => 
                           sum_addr_o_9_port, IN0(8) => sum_addr_o_8_port, 
                           IN0(7) => sum_addr_o_7_port, IN0(6) => 
                           sum_addr_o_6_port, IN0(5) => sum_addr_o_5_port, 
                           IN0(4) => sum_addr_o_4_port, IN0(3) => 
                           sum_addr_o_3_port, IN0(2) => sum_addr_o_2_port, 
                           IN0(1) => sum_addr_o_1_port, IN0(0) => 
                           sum_addr_o_0_port, IN1(31) => NPCF_i(31), IN1(30) =>
                           NPCF_i(30), IN1(29) => NPCF_i(29), IN1(28) => 
                           NPCF_i(28), IN1(27) => NPCF_i(27), IN1(26) => 
                           NPCF_i(26), IN1(25) => NPCF_i(25), IN1(24) => 
                           NPCF_i(24), IN1(23) => NPCF_i(23), IN1(22) => 
                           NPCF_i(22), IN1(21) => NPCF_i(21), IN1(20) => 
                           NPCF_i(20), IN1(19) => NPCF_i(19), IN1(18) => 
                           NPCF_i(18), IN1(17) => NPCF_i(17), IN1(16) => 
                           NPCF_i(16), IN1(15) => NPCF_i(15), IN1(14) => 
                           NPCF_i(14), IN1(13) => NPCF_i(13), IN1(12) => 
                           NPCF_i(12), IN1(11) => NPCF_i(11), IN1(10) => 
                           NPCF_i(10), IN1(9) => NPCF_i(9), IN1(8) => NPCF_i(8)
                           , IN1(7) => NPCF_i(7), IN1(6) => NPCF_i(6), IN1(5) 
                           => NPCF_i(5), IN1(4) => NPCF_i(4), IN1(3) => 
                           NPCF_i(3), IN1(2) => NPCF_i(2), IN1(1) => NPCF_i(1),
                           IN1(0) => NPCF_i(0), CTRL => branch_sel, OUT1(31) =>
                           branch_target_o(31), OUT1(30) => branch_target_o(30)
                           , OUT1(29) => branch_target_o(29), OUT1(28) => 
                           branch_target_o(28), OUT1(27) => branch_target_o(27)
                           , OUT1(26) => branch_target_o(26), OUT1(25) => 
                           branch_target_o(25), OUT1(24) => branch_target_o(24)
                           , OUT1(23) => branch_target_o(23), OUT1(22) => 
                           branch_target_o(22), OUT1(21) => branch_target_o(21)
                           , OUT1(20) => branch_target_o(20), OUT1(19) => 
                           branch_target_o(19), OUT1(18) => branch_target_o(18)
                           , OUT1(17) => branch_target_o(17), OUT1(16) => 
                           branch_target_o(16), OUT1(15) => branch_target_o(15)
                           , OUT1(14) => branch_target_o(14), OUT1(13) => 
                           branch_target_o(13), OUT1(12) => branch_target_o(12)
                           , OUT1(11) => branch_target_o(11), OUT1(10) => 
                           branch_target_o(10), OUT1(9) => branch_target_o(9), 
                           OUT1(8) => branch_target_o(8), OUT1(7) => 
                           branch_target_o(7), OUT1(6) => branch_target_o(6), 
                           OUT1(5) => branch_target_o(5), OUT1(4) => 
                           branch_target_o(4), OUT1(3) => branch_target_o(3), 
                           OUT1(2) => branch_target_o(2), OUT1(1) => 
                           branch_target_o(1), OUT1(0) => branch_target_o(0));
   ZC : zerocheck port map( IN0(31) => A_o_31_port, IN0(30) => A_o_30_port, 
                           IN0(29) => A_o_29_port, IN0(28) => A_o_28_port, 
                           IN0(27) => A_o_27_port, IN0(26) => A_o_26_port, 
                           IN0(25) => A_o_25_port, IN0(24) => A_o_24_port, 
                           IN0(23) => A_o_23_port, IN0(22) => A_o_22_port, 
                           IN0(21) => A_o_21_port, IN0(20) => A_o_20_port, 
                           IN0(19) => A_o_19_port, IN0(18) => A_o_18_port, 
                           IN0(17) => A_o_17_port, IN0(16) => A_o_16_port, 
                           IN0(15) => A_o_15_port, IN0(14) => A_o_14_port, 
                           IN0(13) => A_o_13_port, IN0(12) => A_o_12_port, 
                           IN0(11) => A_o_11_port, IN0(10) => A_o_10_port, 
                           IN0(9) => A_o_9_port, IN0(8) => A_o_8_port, IN0(7) 
                           => A_o_7_port, IN0(6) => A_o_6_port, IN0(5) => 
                           A_o_5_port, IN0(4) => A_o_4_port, IN0(3) => 
                           A_o_3_port, IN0(2) => A_o_2_port, IN0(1) => 
                           A_o_1_port, IN0(0) => A_o_0_port, CTRL => S_EQ_NEQ_i
                           , OUT1 => branch_sel);
   MUXLINK : mux21_4 port map( IN0(31) => ext_imm_31_port, IN0(30) => 
                           ext_imm_30_port, IN0(29) => n3, IN0(28) => 
                           ext_imm_28_port, IN0(27) => n2, IN0(26) => 
                           ext_imm_26_port, IN0(25) => n1, IN0(24) => 
                           ext_imm_24_port, IN0(23) => ext_imm_23_port, IN0(22)
                           => ext_imm_22_port, IN0(21) => ext_imm_21_port, 
                           IN0(20) => ext_imm_20_port, IN0(19) => 
                           ext_imm_19_port, IN0(18) => ext_imm_18_port, IN0(17)
                           => ext_imm_17_port, IN0(16) => ext_imm_16_port, 
                           IN0(15) => ext_imm_15_port, IN0(14) => 
                           ext_imm_14_port, IN0(13) => ext_imm_13_port, IN0(12)
                           => ext_imm_12_port, IN0(11) => ext_imm_11_port, 
                           IN0(10) => ext_imm_10_port, IN0(9) => ext_imm_9_port
                           , IN0(8) => ext_imm_8_port, IN0(7) => ext_imm_7_port
                           , IN0(6) => ext_imm_6_port, IN0(5) => ext_imm_5_port
                           , IN0(4) => ext_imm_4_port, IN0(3) => ext_imm_3_port
                           , IN0(2) => ext_imm_2_port, IN0(1) => ext_imm_1_port
                           , IN0(0) => ext_imm_0_port, IN1(31) => NPCF_i(31), 
                           IN1(30) => NPCF_i(30), IN1(29) => NPCF_i(29), 
                           IN1(28) => NPCF_i(28), IN1(27) => NPCF_i(27), 
                           IN1(26) => NPCF_i(26), IN1(25) => NPCF_i(25), 
                           IN1(24) => NPCF_i(24), IN1(23) => NPCF_i(23), 
                           IN1(22) => NPCF_i(22), IN1(21) => NPCF_i(21), 
                           IN1(20) => NPCF_i(20), IN1(19) => NPCF_i(19), 
                           IN1(18) => NPCF_i(18), IN1(17) => NPCF_i(17), 
                           IN1(16) => NPCF_i(16), IN1(15) => NPCF_i(15), 
                           IN1(14) => NPCF_i(14), IN1(13) => NPCF_i(13), 
                           IN1(12) => NPCF_i(12), IN1(11) => NPCF_i(11), 
                           IN1(10) => NPCF_i(10), IN1(9) => NPCF_i(9), IN1(8) 
                           => NPCF_i(8), IN1(7) => NPCF_i(7), IN1(6) => 
                           NPCF_i(6), IN1(5) => NPCF_i(5), IN1(4) => NPCF_i(4),
                           IN1(3) => NPCF_i(3), IN1(2) => NPCF_i(2), IN1(1) => 
                           NPCF_i(1), IN1(0) => NPCF_i(0), CTRL => S_MUX_LINK_i
                           , OUT1(31) => extended_imm(31), OUT1(30) => 
                           extended_imm(30), OUT1(29) => extended_imm(29), 
                           OUT1(28) => extended_imm(28), OUT1(27) => 
                           extended_imm(27), OUT1(26) => extended_imm(26), 
                           OUT1(25) => extended_imm(25), OUT1(24) => 
                           extended_imm(24), OUT1(23) => extended_imm(23), 
                           OUT1(22) => extended_imm(22), OUT1(21) => 
                           extended_imm(21), OUT1(20) => extended_imm(20), 
                           OUT1(19) => extended_imm(19), OUT1(18) => 
                           extended_imm(18), OUT1(17) => extended_imm(17), 
                           OUT1(16) => extended_imm(16), OUT1(15) => 
                           extended_imm(15), OUT1(14) => extended_imm(14), 
                           OUT1(13) => extended_imm(13), OUT1(12) => 
                           extended_imm(12), OUT1(11) => extended_imm(11), 
                           OUT1(10) => extended_imm(10), OUT1(9) => 
                           extended_imm(9), OUT1(8) => extended_imm(8), OUT1(7)
                           => extended_imm(7), OUT1(6) => extended_imm(6), 
                           OUT1(5) => extended_imm(5), OUT1(4) => 
                           extended_imm(4), OUT1(3) => extended_imm(3), OUT1(2)
                           => extended_imm(2), OUT1(1) => extended_imm(1), 
                           OUT1(0) => extended_imm(0));
   MUX_FWA : mux41_MUX_SIZE32_0 port map( IN0(31) => A_i(31), IN0(30) => 
                           A_i(30), IN0(29) => A_i(29), IN0(28) => A_i(28), 
                           IN0(27) => A_i(27), IN0(26) => A_i(26), IN0(25) => 
                           A_i(25), IN0(24) => A_i(24), IN0(23) => A_i(23), 
                           IN0(22) => A_i(22), IN0(21) => A_i(21), IN0(20) => 
                           A_i(20), IN0(19) => A_i(19), IN0(18) => A_i(18), 
                           IN0(17) => A_i(17), IN0(16) => A_i(16), IN0(15) => 
                           A_i(15), IN0(14) => A_i(14), IN0(13) => A_i(13), 
                           IN0(12) => A_i(12), IN0(11) => A_i(11), IN0(10) => 
                           A_i(10), IN0(9) => A_i(9), IN0(8) => A_i(8), IN0(7) 
                           => A_i(7), IN0(6) => A_i(6), IN0(5) => A_i(5), 
                           IN0(4) => A_i(4), IN0(3) => A_i(3), IN0(2) => A_i(2)
                           , IN0(1) => A_i(1), IN0(0) => A_i(0), IN1(31) => 
                           FW_X_i(31), IN1(30) => FW_X_i(30), IN1(29) => 
                           FW_X_i(29), IN1(28) => FW_X_i(28), IN1(27) => 
                           FW_X_i(27), IN1(26) => FW_X_i(26), IN1(25) => 
                           FW_X_i(25), IN1(24) => FW_X_i(24), IN1(23) => 
                           FW_X_i(23), IN1(22) => FW_X_i(22), IN1(21) => 
                           FW_X_i(21), IN1(20) => FW_X_i(20), IN1(19) => 
                           FW_X_i(19), IN1(18) => FW_X_i(18), IN1(17) => 
                           FW_X_i(17), IN1(16) => FW_X_i(16), IN1(15) => 
                           FW_X_i(15), IN1(14) => FW_X_i(14), IN1(13) => 
                           FW_X_i(13), IN1(12) => FW_X_i(12), IN1(11) => 
                           FW_X_i(11), IN1(10) => FW_X_i(10), IN1(9) => 
                           FW_X_i(9), IN1(8) => FW_X_i(8), IN1(7) => FW_X_i(7),
                           IN1(6) => FW_X_i(6), IN1(5) => FW_X_i(5), IN1(4) => 
                           FW_X_i(4), IN1(3) => FW_X_i(3), IN1(2) => FW_X_i(2),
                           IN1(1) => FW_X_i(1), IN1(0) => FW_X_i(0), IN2(31) =>
                           FW_W_i(31), IN2(30) => FW_W_i(30), IN2(29) => 
                           FW_W_i(29), IN2(28) => FW_W_i(28), IN2(27) => 
                           FW_W_i(27), IN2(26) => FW_W_i(26), IN2(25) => 
                           FW_W_i(25), IN2(24) => FW_W_i(24), IN2(23) => 
                           FW_W_i(23), IN2(22) => FW_W_i(22), IN2(21) => 
                           FW_W_i(21), IN2(20) => FW_W_i(20), IN2(19) => 
                           FW_W_i(19), IN2(18) => FW_W_i(18), IN2(17) => 
                           FW_W_i(17), IN2(16) => FW_W_i(16), IN2(15) => 
                           FW_W_i(15), IN2(14) => FW_W_i(14), IN2(13) => 
                           FW_W_i(13), IN2(12) => FW_W_i(12), IN2(11) => 
                           FW_W_i(11), IN2(10) => FW_W_i(10), IN2(9) => 
                           FW_W_i(9), IN2(8) => FW_W_i(8), IN2(7) => FW_W_i(7),
                           IN2(6) => FW_W_i(6), IN2(5) => FW_W_i(5), IN2(4) => 
                           FW_W_i(4), IN2(3) => FW_W_i(3), IN2(2) => FW_W_i(2),
                           IN2(1) => FW_W_i(1), IN2(0) => FW_W_i(0), IN3(31) =>
                           X_Logic0_port, IN3(30) => X_Logic0_port, IN3(29) => 
                           X_Logic0_port, IN3(28) => X_Logic0_port, IN3(27) => 
                           X_Logic0_port, IN3(26) => X_Logic0_port, IN3(25) => 
                           X_Logic0_port, IN3(24) => X_Logic0_port, IN3(23) => 
                           X_Logic0_port, IN3(22) => X_Logic0_port, IN3(21) => 
                           X_Logic0_port, IN3(20) => X_Logic0_port, IN3(19) => 
                           X_Logic0_port, IN3(18) => X_Logic0_port, IN3(17) => 
                           X_Logic0_port, IN3(16) => X_Logic0_port, IN3(15) => 
                           X_Logic0_port, IN3(14) => X_Logic0_port, IN3(13) => 
                           X_Logic0_port, IN3(12) => X_Logic0_port, IN3(11) => 
                           X_Logic0_port, IN3(10) => X_Logic0_port, IN3(9) => 
                           X_Logic0_port, IN3(8) => X_Logic0_port, IN3(7) => 
                           X_Logic0_port, IN3(6) => X_Logic0_port, IN3(5) => 
                           X_Logic0_port, IN3(4) => X_Logic0_port, IN3(3) => 
                           X_Logic0_port, IN3(2) => X_Logic0_port, IN3(1) => 
                           X_Logic0_port, IN3(0) => X_Logic0_port, CTRL(1) => 
                           S_FW_Adec_i(1), CTRL(0) => S_FW_Adec_i(0), OUT1(31) 
                           => A_o_31_port, OUT1(30) => A_o_30_port, OUT1(29) =>
                           A_o_29_port, OUT1(28) => A_o_28_port, OUT1(27) => 
                           A_o_27_port, OUT1(26) => A_o_26_port, OUT1(25) => 
                           A_o_25_port, OUT1(24) => A_o_24_port, OUT1(23) => 
                           A_o_23_port, OUT1(22) => A_o_22_port, OUT1(21) => 
                           A_o_21_port, OUT1(20) => A_o_20_port, OUT1(19) => 
                           A_o_19_port, OUT1(18) => A_o_18_port, OUT1(17) => 
                           A_o_17_port, OUT1(16) => A_o_16_port, OUT1(15) => 
                           A_o_15_port, OUT1(14) => A_o_14_port, OUT1(13) => 
                           A_o_13_port, OUT1(12) => A_o_12_port, OUT1(11) => 
                           A_o_11_port, OUT1(10) => A_o_10_port, OUT1(9) => 
                           A_o_9_port, OUT1(8) => A_o_8_port, OUT1(7) => 
                           A_o_7_port, OUT1(6) => A_o_6_port, OUT1(5) => 
                           A_o_5_port, OUT1(4) => A_o_4_port, OUT1(3) => 
                           A_o_3_port, OUT1(2) => A_o_2_port, OUT1(1) => 
                           A_o_1_port, OUT1(0) => A_o_0_port);
   U2 : INV_X1 port map( A => branch_sel, ZN => taken_o);
   n6 <= '0';
   n7 <= '0';
   n8 <= '0';
   n9 <= '0';
   n10 <= '0';
   n11 <= '0';

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity fetch_regs is

   port( NPCF_i, IR_i : in std_logic_vector (31 downto 0);  NPCF_o, IR_o : out 
         std_logic_vector (31 downto 0);  stall_i, clk, rst : in std_logic);

end fetch_regs;

architecture SYN_struct of fetch_regs is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component ff32_en_IR
      port( D : in std_logic_vector (31 downto 0);  en, clk, rst : in std_logic
            ;  Q : out std_logic_vector (31 downto 0));
   end component;
   
   component ff32_en_1
      port( D : in std_logic_vector (31 downto 0);  en, clk, rst : in std_logic
            ;  Q : out std_logic_vector (31 downto 0));
   end component;
   
   signal enable : std_logic;

begin
   
   NPCF : ff32_en_1 port map( D(31) => NPCF_i(31), D(30) => NPCF_i(30), D(29) 
                           => NPCF_i(29), D(28) => NPCF_i(28), D(27) => 
                           NPCF_i(27), D(26) => NPCF_i(26), D(25) => NPCF_i(25)
                           , D(24) => NPCF_i(24), D(23) => NPCF_i(23), D(22) =>
                           NPCF_i(22), D(21) => NPCF_i(21), D(20) => NPCF_i(20)
                           , D(19) => NPCF_i(19), D(18) => NPCF_i(18), D(17) =>
                           NPCF_i(17), D(16) => NPCF_i(16), D(15) => NPCF_i(15)
                           , D(14) => NPCF_i(14), D(13) => NPCF_i(13), D(12) =>
                           NPCF_i(12), D(11) => NPCF_i(11), D(10) => NPCF_i(10)
                           , D(9) => NPCF_i(9), D(8) => NPCF_i(8), D(7) => 
                           NPCF_i(7), D(6) => NPCF_i(6), D(5) => NPCF_i(5), 
                           D(4) => NPCF_i(4), D(3) => NPCF_i(3), D(2) => 
                           NPCF_i(2), D(1) => NPCF_i(1), D(0) => NPCF_i(0), en 
                           => enable, clk => clk, rst => rst, Q(31) => 
                           NPCF_o(31), Q(30) => NPCF_o(30), Q(29) => NPCF_o(29)
                           , Q(28) => NPCF_o(28), Q(27) => NPCF_o(27), Q(26) =>
                           NPCF_o(26), Q(25) => NPCF_o(25), Q(24) => NPCF_o(24)
                           , Q(23) => NPCF_o(23), Q(22) => NPCF_o(22), Q(21) =>
                           NPCF_o(21), Q(20) => NPCF_o(20), Q(19) => NPCF_o(19)
                           , Q(18) => NPCF_o(18), Q(17) => NPCF_o(17), Q(16) =>
                           NPCF_o(16), Q(15) => NPCF_o(15), Q(14) => NPCF_o(14)
                           , Q(13) => NPCF_o(13), Q(12) => NPCF_o(12), Q(11) =>
                           NPCF_o(11), Q(10) => NPCF_o(10), Q(9) => NPCF_o(9), 
                           Q(8) => NPCF_o(8), Q(7) => NPCF_o(7), Q(6) => 
                           NPCF_o(6), Q(5) => NPCF_o(5), Q(4) => NPCF_o(4), 
                           Q(3) => NPCF_o(3), Q(2) => NPCF_o(2), Q(1) => 
                           NPCF_o(1), Q(0) => NPCF_o(0));
   IR : ff32_en_IR port map( D(31) => IR_i(31), D(30) => IR_i(30), D(29) => 
                           IR_i(29), D(28) => IR_i(28), D(27) => IR_i(27), 
                           D(26) => IR_i(26), D(25) => IR_i(25), D(24) => 
                           IR_i(24), D(23) => IR_i(23), D(22) => IR_i(22), 
                           D(21) => IR_i(21), D(20) => IR_i(20), D(19) => 
                           IR_i(19), D(18) => IR_i(18), D(17) => IR_i(17), 
                           D(16) => IR_i(16), D(15) => IR_i(15), D(14) => 
                           IR_i(14), D(13) => IR_i(13), D(12) => IR_i(12), 
                           D(11) => IR_i(11), D(10) => IR_i(10), D(9) => 
                           IR_i(9), D(8) => IR_i(8), D(7) => IR_i(7), D(6) => 
                           IR_i(6), D(5) => IR_i(5), D(4) => IR_i(4), D(3) => 
                           IR_i(3), D(2) => IR_i(2), D(1) => IR_i(1), D(0) => 
                           IR_i(0), en => enable, clk => clk, rst => rst, Q(31)
                           => IR_o(31), Q(30) => IR_o(30), Q(29) => IR_o(29), 
                           Q(28) => IR_o(28), Q(27) => IR_o(27), Q(26) => 
                           IR_o(26), Q(25) => IR_o(25), Q(24) => IR_o(24), 
                           Q(23) => IR_o(23), Q(22) => IR_o(22), Q(21) => 
                           IR_o(21), Q(20) => IR_o(20), Q(19) => IR_o(19), 
                           Q(18) => IR_o(18), Q(17) => IR_o(17), Q(16) => 
                           IR_o(16), Q(15) => IR_o(15), Q(14) => IR_o(14), 
                           Q(13) => IR_o(13), Q(12) => IR_o(12), Q(11) => 
                           IR_o(11), Q(10) => IR_o(10), Q(9) => IR_o(9), Q(8) 
                           => IR_o(8), Q(7) => IR_o(7), Q(6) => IR_o(6), Q(5) 
                           => IR_o(5), Q(4) => IR_o(4), Q(3) => IR_o(3), Q(2) 
                           => IR_o(2), Q(1) => IR_o(1), Q(0) => IR_o(0));
   U1 : INV_X1 port map( A => stall_i, ZN => enable);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity btb_N_LINES4_SIZE32 is

   port( clock, reset, stall_i : in std_logic;  TAG_i : in std_logic_vector (3 
         downto 0);  target_PC_i : in std_logic_vector (31 downto 0);  
         was_taken_i : in std_logic;  predicted_next_PC_o : out 
         std_logic_vector (31 downto 0);  taken_o, mispredict_o : out std_logic
         );

end btb_N_LINES4_SIZE32;

architecture SYN_bhe of btb_N_LINES4_SIZE32 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_1
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_2
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_3
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_4
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_5
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_6
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_7
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_8
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_9
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_10
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_11
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_12
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_13
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_14
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_15
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_16
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_0
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component predictor_2_1
      port( clock, reset, enable, taken_i : in std_logic;  prediction_o : out 
            std_logic);
   end component;
   
   component predictor_2_2
      port( clock, reset, enable, taken_i : in std_logic;  prediction_o : out 
            std_logic);
   end component;
   
   component predictor_2_3
      port( clock, reset, enable, taken_i : in std_logic;  prediction_o : out 
            std_logic);
   end component;
   
   component predictor_2_4
      port( clock, reset, enable, taken_i : in std_logic;  prediction_o : out 
            std_logic);
   end component;
   
   component predictor_2_5
      port( clock, reset, enable, taken_i : in std_logic;  prediction_o : out 
            std_logic);
   end component;
   
   component predictor_2_6
      port( clock, reset, enable, taken_i : in std_logic;  prediction_o : out 
            std_logic);
   end component;
   
   component predictor_2_7
      port( clock, reset, enable, taken_i : in std_logic;  prediction_o : out 
            std_logic);
   end component;
   
   component predictor_2_8
      port( clock, reset, enable, taken_i : in std_logic;  prediction_o : out 
            std_logic);
   end component;
   
   component predictor_2_9
      port( clock, reset, enable, taken_i : in std_logic;  prediction_o : out 
            std_logic);
   end component;
   
   component predictor_2_10
      port( clock, reset, enable, taken_i : in std_logic;  prediction_o : out 
            std_logic);
   end component;
   
   component predictor_2_11
      port( clock, reset, enable, taken_i : in std_logic;  prediction_o : out 
            std_logic);
   end component;
   
   component predictor_2_12
      port( clock, reset, enable, taken_i : in std_logic;  prediction_o : out 
            std_logic);
   end component;
   
   component predictor_2_13
      port( clock, reset, enable, taken_i : in std_logic;  prediction_o : out 
            std_logic);
   end component;
   
   component predictor_2_14
      port( clock, reset, enable, taken_i : in std_logic;  prediction_o : out 
            std_logic);
   end component;
   
   component predictor_2_15
      port( clock, reset, enable, taken_i : in std_logic;  prediction_o : out 
            std_logic);
   end component;
   
   component predictor_2_0
      port( clock, reset, enable, taken_i : in std_logic;  prediction_o : out 
            std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFS_X1
      port( D, CK, SN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal predicted_next_PC_o_31_port, predicted_next_PC_o_30_port, 
      predicted_next_PC_o_29_port, predicted_next_PC_o_28_port, 
      predicted_next_PC_o_27_port, predicted_next_PC_o_26_port, 
      predicted_next_PC_o_25_port, predicted_next_PC_o_24_port, 
      predicted_next_PC_o_23_port, predicted_next_PC_o_22_port, 
      predicted_next_PC_o_21_port, predicted_next_PC_o_20_port, 
      predicted_next_PC_o_19_port, predicted_next_PC_o_18_port, 
      predicted_next_PC_o_17_port, predicted_next_PC_o_16_port, 
      predicted_next_PC_o_15_port, predicted_next_PC_o_14_port, 
      predicted_next_PC_o_13_port, predicted_next_PC_o_12_port, 
      predicted_next_PC_o_11_port, predicted_next_PC_o_10_port, 
      predicted_next_PC_o_9_port, predicted_next_PC_o_8_port, 
      predicted_next_PC_o_7_port, predicted_next_PC_o_6_port, 
      predicted_next_PC_o_5_port, predicted_next_PC_o_4_port, 
      predicted_next_PC_o_3_port, predicted_next_PC_o_2_port, 
      predicted_next_PC_o_1_port, predicted_next_PC_o_0_port, taken_o_port, 
      mispredict_o_port, taken_15_port, taken_14_port, taken_13_port, 
      taken_12_port, taken_11_port, taken_10_port, taken_9_port, taken_8_port, 
      taken_7_port, taken_6_port, taken_5_port, taken_4_port, taken_3_port, 
      taken_2_port, taken_1_port, taken_0_port, write_enable_15_port, 
      write_enable_14_port, write_enable_13_port, write_enable_12_port, 
      write_enable_11_port, write_enable_10_port, write_enable_9_port, 
      write_enable_8_port, write_enable_7_port, write_enable_6_port, 
      write_enable_5_port, write_enable_4_port, write_enable_3_port, 
      write_enable_2_port, write_enable_1_port, write_enable_0_port, 
      predict_PC_0_31_port, predict_PC_0_30_port, predict_PC_0_29_port, 
      predict_PC_0_28_port, predict_PC_0_27_port, predict_PC_0_26_port, 
      predict_PC_0_25_port, predict_PC_0_24_port, predict_PC_0_23_port, 
      predict_PC_0_22_port, predict_PC_0_21_port, predict_PC_0_20_port, 
      predict_PC_0_19_port, predict_PC_0_18_port, predict_PC_0_17_port, 
      predict_PC_0_16_port, predict_PC_0_15_port, predict_PC_0_14_port, 
      predict_PC_0_13_port, predict_PC_0_12_port, predict_PC_0_11_port, 
      predict_PC_0_10_port, predict_PC_0_9_port, predict_PC_0_8_port, 
      predict_PC_0_7_port, predict_PC_0_6_port, predict_PC_0_5_port, 
      predict_PC_0_4_port, predict_PC_0_3_port, predict_PC_0_2_port, 
      predict_PC_0_1_port, predict_PC_0_0_port, predict_PC_1_31_port, 
      predict_PC_1_30_port, predict_PC_1_29_port, predict_PC_1_28_port, 
      predict_PC_1_27_port, predict_PC_1_26_port, predict_PC_1_25_port, 
      predict_PC_1_24_port, predict_PC_1_23_port, predict_PC_1_22_port, 
      predict_PC_1_21_port, predict_PC_1_20_port, predict_PC_1_19_port, 
      predict_PC_1_18_port, predict_PC_1_17_port, predict_PC_1_16_port, 
      predict_PC_1_15_port, predict_PC_1_14_port, predict_PC_1_13_port, 
      predict_PC_1_12_port, predict_PC_1_11_port, predict_PC_1_10_port, 
      predict_PC_1_9_port, predict_PC_1_8_port, predict_PC_1_7_port, 
      predict_PC_1_6_port, predict_PC_1_5_port, predict_PC_1_4_port, 
      predict_PC_1_3_port, predict_PC_1_2_port, predict_PC_1_1_port, 
      predict_PC_1_0_port, predict_PC_2_31_port, predict_PC_2_30_port, 
      predict_PC_2_29_port, predict_PC_2_28_port, predict_PC_2_27_port, 
      predict_PC_2_26_port, predict_PC_2_25_port, predict_PC_2_24_port, 
      predict_PC_2_23_port, predict_PC_2_22_port, predict_PC_2_21_port, 
      predict_PC_2_20_port, predict_PC_2_19_port, predict_PC_2_18_port, 
      predict_PC_2_17_port, predict_PC_2_16_port, predict_PC_2_15_port, 
      predict_PC_2_14_port, predict_PC_2_13_port, predict_PC_2_12_port, 
      predict_PC_2_11_port, predict_PC_2_10_port, predict_PC_2_9_port, 
      predict_PC_2_8_port, predict_PC_2_7_port, predict_PC_2_6_port, 
      predict_PC_2_5_port, predict_PC_2_4_port, predict_PC_2_3_port, 
      predict_PC_2_2_port, predict_PC_2_1_port, predict_PC_2_0_port, 
      predict_PC_3_31_port, predict_PC_3_30_port, predict_PC_3_29_port, 
      predict_PC_3_28_port, predict_PC_3_27_port, predict_PC_3_26_port, 
      predict_PC_3_25_port, predict_PC_3_24_port, predict_PC_3_23_port, 
      predict_PC_3_22_port, predict_PC_3_21_port, predict_PC_3_20_port, 
      predict_PC_3_19_port, predict_PC_3_18_port, predict_PC_3_17_port, 
      predict_PC_3_16_port, predict_PC_3_15_port, predict_PC_3_14_port, 
      predict_PC_3_13_port, predict_PC_3_12_port, predict_PC_3_11_port, 
      predict_PC_3_10_port, predict_PC_3_9_port, predict_PC_3_8_port, 
      predict_PC_3_7_port, predict_PC_3_6_port, predict_PC_3_5_port, 
      predict_PC_3_4_port, predict_PC_3_3_port, predict_PC_3_2_port, 
      predict_PC_3_1_port, predict_PC_3_0_port, predict_PC_4_31_port, 
      predict_PC_4_30_port, predict_PC_4_29_port, predict_PC_4_28_port, 
      predict_PC_4_27_port, predict_PC_4_26_port, predict_PC_4_25_port, 
      predict_PC_4_24_port, predict_PC_4_23_port, predict_PC_4_22_port, 
      predict_PC_4_21_port, predict_PC_4_20_port, predict_PC_4_19_port, 
      predict_PC_4_18_port, predict_PC_4_17_port, predict_PC_4_16_port, 
      predict_PC_4_15_port, predict_PC_4_14_port, predict_PC_4_13_port, 
      predict_PC_4_12_port, predict_PC_4_11_port, predict_PC_4_10_port, 
      predict_PC_4_9_port, predict_PC_4_8_port, predict_PC_4_7_port, 
      predict_PC_4_6_port, predict_PC_4_5_port, predict_PC_4_4_port, 
      predict_PC_4_3_port, predict_PC_4_2_port, predict_PC_4_1_port, 
      predict_PC_4_0_port, predict_PC_5_31_port, predict_PC_5_30_port, 
      predict_PC_5_29_port, predict_PC_5_28_port, predict_PC_5_27_port, 
      predict_PC_5_26_port, predict_PC_5_25_port, predict_PC_5_24_port, 
      predict_PC_5_23_port, predict_PC_5_22_port, predict_PC_5_21_port, 
      predict_PC_5_20_port, predict_PC_5_19_port, predict_PC_5_18_port, 
      predict_PC_5_17_port, predict_PC_5_16_port, predict_PC_5_15_port, 
      predict_PC_5_14_port, predict_PC_5_13_port, predict_PC_5_12_port, 
      predict_PC_5_11_port, predict_PC_5_10_port, predict_PC_5_9_port, 
      predict_PC_5_8_port, predict_PC_5_7_port, predict_PC_5_6_port, 
      predict_PC_5_5_port, predict_PC_5_4_port, predict_PC_5_3_port, 
      predict_PC_5_2_port, predict_PC_5_1_port, predict_PC_5_0_port, 
      predict_PC_6_31_port, predict_PC_6_30_port, predict_PC_6_29_port, 
      predict_PC_6_28_port, predict_PC_6_27_port, predict_PC_6_26_port, 
      predict_PC_6_25_port, predict_PC_6_24_port, predict_PC_6_23_port, 
      predict_PC_6_22_port, predict_PC_6_21_port, predict_PC_6_20_port, 
      predict_PC_6_19_port, predict_PC_6_18_port, predict_PC_6_17_port, 
      predict_PC_6_16_port, predict_PC_6_15_port, predict_PC_6_14_port, 
      predict_PC_6_13_port, predict_PC_6_12_port, predict_PC_6_11_port, 
      predict_PC_6_10_port, predict_PC_6_9_port, predict_PC_6_8_port, 
      predict_PC_6_7_port, predict_PC_6_6_port, predict_PC_6_5_port, 
      predict_PC_6_4_port, predict_PC_6_3_port, predict_PC_6_2_port, 
      predict_PC_6_1_port, predict_PC_6_0_port, predict_PC_7_31_port, 
      predict_PC_7_30_port, predict_PC_7_29_port, predict_PC_7_28_port, 
      predict_PC_7_27_port, predict_PC_7_26_port, predict_PC_7_25_port, 
      predict_PC_7_24_port, predict_PC_7_23_port, predict_PC_7_22_port, 
      predict_PC_7_21_port, predict_PC_7_20_port, predict_PC_7_19_port, 
      predict_PC_7_18_port, predict_PC_7_17_port, predict_PC_7_16_port, 
      predict_PC_7_15_port, predict_PC_7_14_port, predict_PC_7_13_port, 
      predict_PC_7_12_port, predict_PC_7_11_port, predict_PC_7_10_port, 
      predict_PC_7_9_port, predict_PC_7_8_port, predict_PC_7_7_port, 
      predict_PC_7_6_port, predict_PC_7_5_port, predict_PC_7_4_port, 
      predict_PC_7_3_port, predict_PC_7_2_port, predict_PC_7_1_port, 
      predict_PC_7_0_port, predict_PC_8_31_port, predict_PC_8_30_port, 
      predict_PC_8_29_port, predict_PC_8_28_port, predict_PC_8_27_port, 
      predict_PC_8_26_port, predict_PC_8_25_port, predict_PC_8_24_port, 
      predict_PC_8_23_port, predict_PC_8_22_port, predict_PC_8_21_port, 
      predict_PC_8_20_port, predict_PC_8_19_port, predict_PC_8_18_port, 
      predict_PC_8_17_port, predict_PC_8_16_port, predict_PC_8_15_port, 
      predict_PC_8_14_port, predict_PC_8_13_port, predict_PC_8_12_port, 
      predict_PC_8_11_port, predict_PC_8_10_port, predict_PC_8_9_port, 
      predict_PC_8_8_port, predict_PC_8_7_port, predict_PC_8_6_port, 
      predict_PC_8_5_port, predict_PC_8_4_port, predict_PC_8_3_port, 
      predict_PC_8_2_port, predict_PC_8_1_port, predict_PC_8_0_port, 
      predict_PC_9_31_port, predict_PC_9_30_port, predict_PC_9_29_port, 
      predict_PC_9_28_port, predict_PC_9_27_port, predict_PC_9_26_port, 
      predict_PC_9_25_port, predict_PC_9_24_port, predict_PC_9_23_port, 
      predict_PC_9_22_port, predict_PC_9_21_port, predict_PC_9_20_port, 
      predict_PC_9_19_port, predict_PC_9_18_port, predict_PC_9_17_port, 
      predict_PC_9_16_port, predict_PC_9_15_port, predict_PC_9_14_port, 
      predict_PC_9_13_port, predict_PC_9_12_port, predict_PC_9_11_port, 
      predict_PC_9_10_port, predict_PC_9_9_port, predict_PC_9_8_port, 
      predict_PC_9_7_port, predict_PC_9_6_port, predict_PC_9_5_port, 
      predict_PC_9_4_port, predict_PC_9_3_port, predict_PC_9_2_port, 
      predict_PC_9_1_port, predict_PC_9_0_port, predict_PC_10_31_port, 
      predict_PC_10_30_port, predict_PC_10_29_port, predict_PC_10_28_port, 
      predict_PC_10_27_port, predict_PC_10_26_port, predict_PC_10_25_port, 
      predict_PC_10_24_port, predict_PC_10_23_port, predict_PC_10_22_port, 
      predict_PC_10_21_port, predict_PC_10_20_port, predict_PC_10_19_port, 
      predict_PC_10_18_port, predict_PC_10_17_port, predict_PC_10_16_port, 
      predict_PC_10_15_port, predict_PC_10_14_port, predict_PC_10_13_port, 
      predict_PC_10_12_port, predict_PC_10_11_port, predict_PC_10_10_port, 
      predict_PC_10_9_port, predict_PC_10_8_port, predict_PC_10_7_port, 
      predict_PC_10_6_port, predict_PC_10_5_port, predict_PC_10_4_port, 
      predict_PC_10_3_port, predict_PC_10_2_port, predict_PC_10_1_port, 
      predict_PC_10_0_port, predict_PC_11_31_port, predict_PC_11_30_port, 
      predict_PC_11_29_port, predict_PC_11_28_port, predict_PC_11_27_port, 
      predict_PC_11_26_port, predict_PC_11_25_port, predict_PC_11_24_port, 
      predict_PC_11_23_port, predict_PC_11_22_port, predict_PC_11_21_port, 
      predict_PC_11_20_port, predict_PC_11_19_port, predict_PC_11_18_port, 
      predict_PC_11_17_port, predict_PC_11_16_port, predict_PC_11_15_port, 
      predict_PC_11_14_port, predict_PC_11_13_port, predict_PC_11_12_port, 
      predict_PC_11_11_port, predict_PC_11_10_port, predict_PC_11_9_port, 
      predict_PC_11_8_port, predict_PC_11_7_port, predict_PC_11_6_port, 
      predict_PC_11_5_port, predict_PC_11_4_port, predict_PC_11_3_port, 
      predict_PC_11_2_port, predict_PC_11_1_port, predict_PC_11_0_port, 
      predict_PC_12_31_port, predict_PC_12_30_port, predict_PC_12_29_port, 
      predict_PC_12_28_port, predict_PC_12_27_port, predict_PC_12_26_port, 
      predict_PC_12_25_port, predict_PC_12_24_port, predict_PC_12_23_port, 
      predict_PC_12_22_port, predict_PC_12_21_port, predict_PC_12_20_port, 
      predict_PC_12_19_port, predict_PC_12_18_port, predict_PC_12_17_port, 
      predict_PC_12_16_port, predict_PC_12_15_port, predict_PC_12_14_port, 
      predict_PC_12_13_port, predict_PC_12_12_port, predict_PC_12_11_port, 
      predict_PC_12_10_port, predict_PC_12_9_port, predict_PC_12_8_port, 
      predict_PC_12_7_port, predict_PC_12_6_port, predict_PC_12_5_port, 
      predict_PC_12_4_port, predict_PC_12_3_port, predict_PC_12_2_port, 
      predict_PC_12_1_port, predict_PC_12_0_port, predict_PC_13_31_port, 
      predict_PC_13_30_port, predict_PC_13_29_port, predict_PC_13_28_port, 
      predict_PC_13_27_port, predict_PC_13_26_port, predict_PC_13_25_port, 
      predict_PC_13_24_port, predict_PC_13_23_port, predict_PC_13_22_port, 
      predict_PC_13_21_port, predict_PC_13_20_port, predict_PC_13_19_port, 
      predict_PC_13_18_port, predict_PC_13_17_port, predict_PC_13_16_port, 
      predict_PC_13_15_port, predict_PC_13_14_port, predict_PC_13_13_port, 
      predict_PC_13_12_port, predict_PC_13_11_port, predict_PC_13_10_port, 
      predict_PC_13_9_port, predict_PC_13_8_port, predict_PC_13_7_port, 
      predict_PC_13_6_port, predict_PC_13_5_port, predict_PC_13_4_port, 
      predict_PC_13_3_port, predict_PC_13_2_port, predict_PC_13_1_port, 
      predict_PC_13_0_port, predict_PC_14_31_port, predict_PC_14_30_port, 
      predict_PC_14_29_port, predict_PC_14_28_port, predict_PC_14_27_port, 
      predict_PC_14_26_port, predict_PC_14_25_port, predict_PC_14_24_port, 
      predict_PC_14_23_port, predict_PC_14_22_port, predict_PC_14_21_port, 
      predict_PC_14_20_port, predict_PC_14_19_port, predict_PC_14_18_port, 
      predict_PC_14_17_port, predict_PC_14_16_port, predict_PC_14_15_port, 
      predict_PC_14_14_port, predict_PC_14_13_port, predict_PC_14_12_port, 
      predict_PC_14_11_port, predict_PC_14_10_port, predict_PC_14_9_port, 
      predict_PC_14_8_port, predict_PC_14_7_port, predict_PC_14_6_port, 
      predict_PC_14_5_port, predict_PC_14_4_port, predict_PC_14_3_port, 
      predict_PC_14_2_port, predict_PC_14_1_port, predict_PC_14_0_port, 
      predict_PC_15_31_port, predict_PC_15_30_port, predict_PC_15_29_port, 
      predict_PC_15_28_port, predict_PC_15_27_port, predict_PC_15_26_port, 
      predict_PC_15_25_port, predict_PC_15_24_port, predict_PC_15_23_port, 
      predict_PC_15_22_port, predict_PC_15_21_port, predict_PC_15_20_port, 
      predict_PC_15_19_port, predict_PC_15_18_port, predict_PC_15_17_port, 
      predict_PC_15_16_port, predict_PC_15_15_port, predict_PC_15_14_port, 
      predict_PC_15_13_port, predict_PC_15_12_port, predict_PC_15_11_port, 
      predict_PC_15_10_port, predict_PC_15_9_port, predict_PC_15_8_port, 
      predict_PC_15_7_port, predict_PC_15_6_port, predict_PC_15_5_port, 
      predict_PC_15_4_port, predict_PC_15_3_port, predict_PC_15_2_port, 
      predict_PC_15_1_port, predict_PC_15_0_port, N38, N39, N40, N41, N42, N43,
      N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N86, N118, N150, N182, 
      N214, N246, N278, N310, N342, N374, N406, N438, N470, N502, N534, N566, 
      N567, net199633, net199638, net199643, net199648, net199653, net199658, 
      net199663, net199668, net199673, net199678, net199683, net199688, 
      net199693, net199698, net199703, net199708, net199713, n483, n485, n487, 
      n489, n491, n493, n495, n497, n499, n501, n503, n505, n507, n509, n511, 
      n513, n515, n517, n519, n521, n523, n525, n527, n529, n531, n533, n535, 
      n537, n539, n541, n543, n545, n546, n547, n548, n549, n550, n551, n552, 
      n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, 
      n565, n566_port, n567_port, n568, n569, n570, n571, n572, n573, n574, 
      n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, 
      n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, 
      n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, 
      n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, 
      n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, 
      n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, 
      n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, 
      n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, 
      n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, 
      n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, 
      n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, 
      n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, 
      n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, 
      n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, 
      n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, 
      n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, 
      n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, 
      n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, 
      n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, 
      n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, 
      n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, 
      n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, 
      n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, 
      n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, 
      n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, 
      n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, 
      n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, 
      n899, n900, n901, n902, n903, n943, n944, n945, n946, n947, n948, n949, 
      n951, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, 
      n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, 
      n978, n979, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, 
      n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29
      , n30, n31, n32, n33, n34, n35, n36, n37, n38_port, n39_port, n40_port, 
      n41_port, n42_port, n43_port, n44_port, n45_port, n46_port, n47_port, 
      n48_port, n49_port, n50_port, n51_port, n52_port, n53_port, n54, n55, n56
      , n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, 
      n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85
      , n86_port, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, 
      n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, 
      n111, n112, n113, net244547, net244548, net244549, net244550, net244551, 
      net244552, net244553, net244554, net244555, net244556, net244557, 
      net244558, net244559, net244560, net244561, net244562, net244563, 
      net244564, net244565, net244566, net244567, net244568, net244569, 
      net244570, net244571, net244572, net244573, net244574, net244575, 
      net244576, net244577, net244578, net244579, net244580, net244581, 
      net244582, net244583, net244584, net244585, net244586, net244587, 
      net244588, net244589, net244590, net244591, net244592, net244593, 
      net244594, net244595, net244596, net244597, net244598, net244599, 
      net244600, net244601, net244602, net244603, net244604, net244605, 
      net244606, net244607, net244608, net244609, net244610, net244611, 
      net244612, net244613, net244614, net244615, net244616, net244617, 
      net244618, net244619, net244620, net244621, net244622, net244623, 
      net244624, net244625, net244626, net244627, net244628, net244629, 
      net244630, net244631, net244632, net244633, net244634, net244635, 
      net244636, net244637, net244638, net244639, net244640, net244641, 
      net244642, net244643, net244644, net244645, net244646, net244647, 
      net244648, net244649, net244650, net244651, net244652, net244653, 
      net244654, net244655, net244656, net244657, net244658, net244659, 
      net244660, net244661, net244662, net244663, net244664, net244665, 
      net244666, net244667, net244668, net244669, net244670, net244671, 
      net244672, net244673, net244674, net244675, net244676, net244677, 
      net244678, net244679, net244680, net244681, net244682, net244683, 
      net244684, net244685, net244686, net244687, net244688, net244689, 
      net244690, net244691, net244692, net244693, net244694, net244695, 
      net244696, net244697, net244698, net244699, net244700, net244701, 
      net244702, net244703, net244704, net244705, net244706, net244707, 
      net244708, net244709, net244710, net244711, net244712, net244713, 
      net244714, net244715, net244716, net244717, net244718, net244719, 
      net244720, net244721, net244722, net244723, net244724, net244725, 
      net244726, net244727, net244728, net244729, net244730, net244731, 
      net244732, net244733, net244734, net244735, net244736, net244737, 
      net244738, net244739, net244740, net244741, net244742, net244743, 
      net244744, net244745, net244746, net244747, net244748, net244749, 
      net244750, net244751, net244752, net244753, net244754, net244755, 
      net244756, net244757, net244758, net244759, net244760, net244761, 
      net244762, net244763, net244764, net244765, net244766, net244767, 
      net244768, net244769, net244770, net244771, net244772, net244773, 
      net244774, net244775, net244776, net244777, net244778, net244779, 
      net244780, net244781, net244782, net244783, net244784, net244785, 
      net244786, net244787, net244788, net244789, net244790, net244791, 
      net244792, net244793, net244794, net244795, net244796, net244797, 
      net244798, net244799, net244800, net244801, net244802, net244803, 
      net244804, net244805, net244806, net244807, net244808, net244809, 
      net244810, net244811, net244812, net244813, net244814, net244815, 
      net244816, net244817, net244818, net244819, net244820, net244821, 
      net244822, net244823, net244824, net244825, net244826, net244827, 
      net244828, net244829, net244830, net244831, net244832, net244833, 
      net244834, net244835, net244836, net244837, net244838, net244839, 
      net244840, net244841, net244842, net244843, net244844, net244845, 
      net244846, net244847, net244848, net244849, net244850, net244851, 
      net244852, net244853, net244854, net244855, net244856, net244857, 
      net244858, net244859, net244860, net244861, net244862, net244863, 
      net244864, net244865, net244866, net244867, net244868, net244869, 
      net244870, net244871, net244872, net244873, net244874, net244875, 
      net244876, net244877, net244878, net244879, net244880, net244881, 
      net244882, net244883, net244884, net244885, net244886, net244887, 
      net244888, net244889, net244890, net244891, net244892, net244893, 
      net244894, net244895, net244896, net244897, net244898, net244899, 
      net244900, net244901, net244902, net244903, net244904, net244905, 
      net244906, net244907, net244908, net244909, net244910, net244911, 
      net244912, net244913, net244914, net244915, net244916, net244917, 
      net244918, net244919, net244920, net244921, net244922, net244923, 
      net244924, net244925, net244926, net244927, net244928, net244929, 
      net244930, net244931, net244932, net244933, net244934, net244935, 
      net244936, net244937, net244938, net244939, net244940, net244941, 
      net244942, net244943, net244944, net244945, net244946, net244947, 
      net244948, net244949, net244950, net244951, net244952, net244953, 
      net244954, net244955, net244956, net244957, net244958, net244959, 
      net244960, net244961, net244962, net244963, net244964, net244965, 
      net244966, net244967, net244968, net244969, net244970, net244971, 
      net244972, net244973, net244974, net244975, net244976, net244977, 
      net244978, net244979, net244980, net244981, net244982, net244983, 
      net244984, net244985, net244986, net244987, net244988, net244989, 
      net244990, net244991, net244992, net244993, net244994, net244995, 
      net244996, net244997, net244998, net244999, net245000, net245001, 
      net245002, net245003, net245004, net245005, net245006, net245007, 
      net245008, net245009, net245010, net245011, net245012, net245013, 
      net245014, net245015, net245016, net245017, net245018, net245019, 
      net245020, net245021, net245022, net245023, net245024, net245025, 
      net245026, net245027, net245028, net245029, net245030, net245031, 
      net245032, net245033, net245034, net245035, net245036, net245037, 
      net245038, net245039, net245040, net245041, net245042, net245043, 
      net245044, net245045, net245046, net245047, net245048, net245049, 
      net245050, net245051, net245052, net245053, net245054, net245055, 
      net245056, net245057, net245058, net245059, net245060, net245061, 
      net245062, net245063, net245064, net245065, net245066, net245067, 
      net245068, net245069, net245070, net245071, net245072, net245073, 
      net245074, net245075, net245076, net245077, net245078, net245079, 
      net245080, net245081, net245082, net245083, net245084, net245085, 
      net245086, net245087, net245088, net245089, net245090, net245091 : 
      std_logic;

begin
   predicted_next_PC_o <= ( predicted_next_PC_o_31_port, 
      predicted_next_PC_o_30_port, predicted_next_PC_o_29_port, 
      predicted_next_PC_o_28_port, predicted_next_PC_o_27_port, 
      predicted_next_PC_o_26_port, predicted_next_PC_o_25_port, 
      predicted_next_PC_o_24_port, predicted_next_PC_o_23_port, 
      predicted_next_PC_o_22_port, predicted_next_PC_o_21_port, 
      predicted_next_PC_o_20_port, predicted_next_PC_o_19_port, 
      predicted_next_PC_o_18_port, predicted_next_PC_o_17_port, 
      predicted_next_PC_o_16_port, predicted_next_PC_o_15_port, 
      predicted_next_PC_o_14_port, predicted_next_PC_o_13_port, 
      predicted_next_PC_o_12_port, predicted_next_PC_o_11_port, 
      predicted_next_PC_o_10_port, predicted_next_PC_o_9_port, 
      predicted_next_PC_o_8_port, predicted_next_PC_o_7_port, 
      predicted_next_PC_o_6_port, predicted_next_PC_o_5_port, 
      predicted_next_PC_o_4_port, predicted_next_PC_o_3_port, 
      predicted_next_PC_o_2_port, predicted_next_PC_o_1_port, 
      predicted_next_PC_o_0_port );
   taken_o <= taken_o_port;
   mispredict_o <= mispredict_o_port;
   
   last_TAG_reg_3_inst : DFFS_X1 port map( D => n972, CK => net199633, SN => 
                           n99, Q => n977, QN => n12);
   last_TAG_reg_2_inst : DFFS_X1 port map( D => n973, CK => net199633, SN => 
                           n90, Q => n976, QN => n10);
   last_TAG_reg_1_inst : DFFS_X1 port map( D => n974, CK => net199633, SN => 
                           n92, Q => n979, QN => n11);
   last_TAG_reg_0_inst : DFFR_X1 port map( D => TAG_i(0), CK => net199633, RN 
                           => n100, Q => n9, QN => n978);
   write_enable_reg_15_inst : DFFR_X1 port map( D => N53, CK => net199633, RN 
                           => n94, Q => write_enable_15_port, QN => n971);
   write_enable_reg_14_inst : DFFR_X1 port map( D => N52, CK => net199633, RN 
                           => n92, Q => write_enable_14_port, QN => n970);
   write_enable_reg_13_inst : DFFR_X1 port map( D => N51, CK => net199633, RN 
                           => n95, Q => write_enable_13_port, QN => n969);
   write_enable_reg_12_inst : DFFR_X1 port map( D => N50, CK => net199633, RN 
                           => n96, Q => write_enable_12_port, QN => n968);
   write_enable_reg_11_inst : DFFR_X1 port map( D => N49, CK => net199633, RN 
                           => n98, Q => write_enable_11_port, QN => n967);
   write_enable_reg_10_inst : DFFR_X1 port map( D => N48, CK => net199633, RN 
                           => n99, Q => write_enable_10_port, QN => n966);
   write_enable_reg_9_inst : DFFR_X1 port map( D => N47, CK => net199633, RN =>
                           n98, Q => write_enable_9_port, QN => n965);
   write_enable_reg_8_inst : DFFR_X1 port map( D => N46, CK => net199633, RN =>
                           n97, Q => write_enable_8_port, QN => n964);
   write_enable_reg_7_inst : DFFR_X1 port map( D => N45, CK => net199633, RN =>
                           n100, Q => write_enable_7_port, QN => n963);
   write_enable_reg_6_inst : DFFR_X1 port map( D => N44, CK => net199633, RN =>
                           n97, Q => write_enable_6_port, QN => n962);
   write_enable_reg_5_inst : DFFR_X1 port map( D => N43, CK => net199633, RN =>
                           n99, Q => write_enable_5_port, QN => n961);
   write_enable_reg_4_inst : DFFR_X1 port map( D => N42, CK => net199633, RN =>
                           n98, Q => write_enable_4_port, QN => n960);
   write_enable_reg_3_inst : DFFR_X1 port map( D => N41, CK => net199633, RN =>
                           n97, Q => write_enable_3_port, QN => n959);
   write_enable_reg_2_inst : DFFR_X1 port map( D => N40, CK => net199633, RN =>
                           n100, Q => write_enable_2_port, QN => n958);
   write_enable_reg_1_inst : DFFR_X1 port map( D => N39, CK => net199633, RN =>
                           n100, Q => write_enable_1_port, QN => n957);
   write_enable_reg_0_inst : DFFR_X1 port map( D => N38, CK => net199633, RN =>
                           n99, Q => write_enable_0_port, QN => n956);
   last_taken_reg : DFF_X1 port map( D => n955, CK => clock, Q => n13, QN => 
                           n975);
   predict_PC_reg_0_31_inst : DFFR_X1 port map( D => target_PC_i(31), CK => 
                           net199638, RN => n100, Q => predict_PC_0_31_port, QN
                           => net245091);
   predict_PC_reg_0_30_inst : DFFR_X1 port map( D => target_PC_i(30), CK => 
                           net199638, RN => n97, Q => predict_PC_0_30_port, QN 
                           => net245090);
   predict_PC_reg_0_29_inst : DFFR_X1 port map( D => target_PC_i(29), CK => 
                           net199638, RN => n98, Q => predict_PC_0_29_port, QN 
                           => net245089);
   predict_PC_reg_0_28_inst : DFFR_X1 port map( D => target_PC_i(28), CK => 
                           net199638, RN => n99, Q => predict_PC_0_28_port, QN 
                           => net245088);
   predict_PC_reg_0_27_inst : DFFR_X1 port map( D => target_PC_i(27), CK => 
                           net199638, RN => n100, Q => predict_PC_0_27_port, QN
                           => net245087);
   predict_PC_reg_0_26_inst : DFFR_X1 port map( D => target_PC_i(26), CK => 
                           net199638, RN => n97, Q => predict_PC_0_26_port, QN 
                           => net245086);
   predict_PC_reg_0_25_inst : DFFR_X1 port map( D => target_PC_i(25), CK => 
                           net199638, RN => n98, Q => predict_PC_0_25_port, QN 
                           => net245085);
   predict_PC_reg_0_24_inst : DFFR_X1 port map( D => target_PC_i(24), CK => 
                           net199638, RN => n99, Q => predict_PC_0_24_port, QN 
                           => net245084);
   predict_PC_reg_0_23_inst : DFFR_X1 port map( D => target_PC_i(23), CK => 
                           net199638, RN => n100, Q => predict_PC_0_23_port, QN
                           => net245083);
   predict_PC_reg_0_22_inst : DFFR_X1 port map( D => target_PC_i(22), CK => 
                           net199638, RN => n97, Q => predict_PC_0_22_port, QN 
                           => net245082);
   predict_PC_reg_0_21_inst : DFFR_X1 port map( D => target_PC_i(21), CK => 
                           net199638, RN => n98, Q => predict_PC_0_21_port, QN 
                           => net245081);
   predict_PC_reg_0_20_inst : DFFR_X1 port map( D => target_PC_i(20), CK => 
                           net199638, RN => n99, Q => predict_PC_0_20_port, QN 
                           => net245080);
   predict_PC_reg_0_19_inst : DFFR_X1 port map( D => target_PC_i(19), CK => 
                           net199638, RN => n97, Q => predict_PC_0_19_port, QN 
                           => net245079);
   predict_PC_reg_0_18_inst : DFFR_X1 port map( D => target_PC_i(18), CK => 
                           net199638, RN => n97, Q => predict_PC_0_18_port, QN 
                           => net245078);
   predict_PC_reg_0_17_inst : DFFR_X1 port map( D => target_PC_i(17), CK => 
                           net199638, RN => n97, Q => predict_PC_0_17_port, QN 
                           => net245077);
   predict_PC_reg_0_16_inst : DFFR_X1 port map( D => target_PC_i(16), CK => 
                           net199638, RN => n97, Q => predict_PC_0_16_port, QN 
                           => net245076);
   predict_PC_reg_0_15_inst : DFFR_X1 port map( D => target_PC_i(15), CK => 
                           net199638, RN => n97, Q => predict_PC_0_15_port, QN 
                           => net245075);
   predict_PC_reg_0_14_inst : DFFR_X1 port map( D => target_PC_i(14), CK => 
                           net199638, RN => n97, Q => predict_PC_0_14_port, QN 
                           => net245074);
   predict_PC_reg_0_13_inst : DFFR_X1 port map( D => target_PC_i(13), CK => 
                           net199638, RN => n97, Q => predict_PC_0_13_port, QN 
                           => net245073);
   predict_PC_reg_0_12_inst : DFFR_X1 port map( D => target_PC_i(12), CK => 
                           net199638, RN => n97, Q => predict_PC_0_12_port, QN 
                           => net245072);
   predict_PC_reg_0_11_inst : DFFR_X1 port map( D => target_PC_i(11), CK => 
                           net199638, RN => n97, Q => predict_PC_0_11_port, QN 
                           => net245071);
   predict_PC_reg_0_10_inst : DFFR_X1 port map( D => target_PC_i(10), CK => 
                           net199638, RN => n97, Q => predict_PC_0_10_port, QN 
                           => net245070);
   predict_PC_reg_0_9_inst : DFFR_X1 port map( D => target_PC_i(9), CK => 
                           net199638, RN => n97, Q => predict_PC_0_9_port, QN 
                           => net245069);
   predict_PC_reg_0_8_inst : DFFR_X1 port map( D => target_PC_i(8), CK => 
                           net199638, RN => n97, Q => predict_PC_0_8_port, QN 
                           => net245068);
   predict_PC_reg_0_7_inst : DFFR_X1 port map( D => target_PC_i(7), CK => 
                           net199638, RN => n98, Q => predict_PC_0_7_port, QN 
                           => net245067);
   predict_PC_reg_0_6_inst : DFFR_X1 port map( D => target_PC_i(6), CK => 
                           net199638, RN => n98, Q => predict_PC_0_6_port, QN 
                           => net245066);
   predict_PC_reg_0_5_inst : DFFR_X1 port map( D => target_PC_i(5), CK => 
                           net199638, RN => n98, Q => predict_PC_0_5_port, QN 
                           => net245065);
   predict_PC_reg_0_4_inst : DFFR_X1 port map( D => target_PC_i(4), CK => 
                           net199638, RN => n98, Q => predict_PC_0_4_port, QN 
                           => net245064);
   predict_PC_reg_0_3_inst : DFFR_X1 port map( D => target_PC_i(3), CK => 
                           net199638, RN => n98, Q => predict_PC_0_3_port, QN 
                           => net245063);
   predict_PC_reg_0_2_inst : DFFR_X1 port map( D => target_PC_i(2), CK => 
                           net199638, RN => n98, Q => predict_PC_0_2_port, QN 
                           => net245062);
   predict_PC_reg_0_1_inst : DFFR_X1 port map( D => target_PC_i(1), CK => 
                           net199638, RN => n98, Q => predict_PC_0_1_port, QN 
                           => net245061);
   predict_PC_reg_0_0_inst : DFFR_X1 port map( D => target_PC_i(0), CK => 
                           net199638, RN => n98, Q => predict_PC_0_0_port, QN 
                           => net245060);
   predict_PC_reg_1_31_inst : DFFR_X1 port map( D => target_PC_i(31), CK => 
                           net199643, RN => n98, Q => predict_PC_1_31_port, QN 
                           => net245059);
   predict_PC_reg_1_30_inst : DFFR_X1 port map( D => target_PC_i(30), CK => 
                           net199643, RN => n98, Q => predict_PC_1_30_port, QN 
                           => net245058);
   predict_PC_reg_1_29_inst : DFFR_X1 port map( D => target_PC_i(29), CK => 
                           net199643, RN => n98, Q => predict_PC_1_29_port, QN 
                           => net245057);
   predict_PC_reg_1_28_inst : DFFR_X1 port map( D => target_PC_i(28), CK => 
                           net199643, RN => n98, Q => predict_PC_1_28_port, QN 
                           => net245056);
   predict_PC_reg_1_27_inst : DFFR_X1 port map( D => target_PC_i(27), CK => 
                           net199643, RN => n99, Q => predict_PC_1_27_port, QN 
                           => net245055);
   predict_PC_reg_1_26_inst : DFFR_X1 port map( D => target_PC_i(26), CK => 
                           net199643, RN => n99, Q => predict_PC_1_26_port, QN 
                           => net245054);
   predict_PC_reg_1_25_inst : DFFR_X1 port map( D => target_PC_i(25), CK => 
                           net199643, RN => n99, Q => predict_PC_1_25_port, QN 
                           => net245053);
   predict_PC_reg_1_24_inst : DFFR_X1 port map( D => target_PC_i(24), CK => 
                           net199643, RN => n99, Q => predict_PC_1_24_port, QN 
                           => net245052);
   predict_PC_reg_1_23_inst : DFFR_X1 port map( D => target_PC_i(23), CK => 
                           net199643, RN => n99, Q => predict_PC_1_23_port, QN 
                           => net245051);
   predict_PC_reg_1_22_inst : DFFR_X1 port map( D => target_PC_i(22), CK => 
                           net199643, RN => n99, Q => predict_PC_1_22_port, QN 
                           => net245050);
   predict_PC_reg_1_21_inst : DFFR_X1 port map( D => target_PC_i(21), CK => 
                           net199643, RN => n99, Q => predict_PC_1_21_port, QN 
                           => net245049);
   predict_PC_reg_1_20_inst : DFFR_X1 port map( D => target_PC_i(20), CK => 
                           net199643, RN => n99, Q => predict_PC_1_20_port, QN 
                           => net245048);
   predict_PC_reg_1_19_inst : DFFR_X1 port map( D => target_PC_i(19), CK => 
                           net199643, RN => n99, Q => predict_PC_1_19_port, QN 
                           => net245047);
   predict_PC_reg_1_18_inst : DFFR_X1 port map( D => target_PC_i(18), CK => 
                           net199643, RN => n99, Q => predict_PC_1_18_port, QN 
                           => net245046);
   predict_PC_reg_1_17_inst : DFFR_X1 port map( D => target_PC_i(17), CK => 
                           net199643, RN => n99, Q => predict_PC_1_17_port, QN 
                           => net245045);
   predict_PC_reg_1_16_inst : DFFR_X1 port map( D => target_PC_i(16), CK => 
                           net199643, RN => n99, Q => predict_PC_1_16_port, QN 
                           => net245044);
   predict_PC_reg_1_15_inst : DFFR_X1 port map( D => target_PC_i(15), CK => 
                           net199643, RN => n100, Q => predict_PC_1_15_port, QN
                           => net245043);
   predict_PC_reg_1_14_inst : DFFR_X1 port map( D => target_PC_i(14), CK => 
                           net199643, RN => n100, Q => predict_PC_1_14_port, QN
                           => net245042);
   predict_PC_reg_1_13_inst : DFFR_X1 port map( D => target_PC_i(13), CK => 
                           net199643, RN => n100, Q => predict_PC_1_13_port, QN
                           => net245041);
   predict_PC_reg_1_12_inst : DFFR_X1 port map( D => target_PC_i(12), CK => 
                           net199643, RN => n100, Q => predict_PC_1_12_port, QN
                           => net245040);
   predict_PC_reg_1_11_inst : DFFR_X1 port map( D => target_PC_i(11), CK => 
                           net199643, RN => n100, Q => predict_PC_1_11_port, QN
                           => net245039);
   predict_PC_reg_1_10_inst : DFFR_X1 port map( D => target_PC_i(10), CK => 
                           net199643, RN => n100, Q => predict_PC_1_10_port, QN
                           => net245038);
   predict_PC_reg_1_9_inst : DFFR_X1 port map( D => target_PC_i(9), CK => 
                           net199643, RN => n100, Q => predict_PC_1_9_port, QN 
                           => net245037);
   predict_PC_reg_1_8_inst : DFFR_X1 port map( D => target_PC_i(8), CK => 
                           net199643, RN => n100, Q => predict_PC_1_8_port, QN 
                           => net245036);
   predict_PC_reg_1_7_inst : DFFR_X1 port map( D => target_PC_i(7), CK => 
                           net199643, RN => n100, Q => predict_PC_1_7_port, QN 
                           => net245035);
   predict_PC_reg_1_6_inst : DFFR_X1 port map( D => target_PC_i(6), CK => 
                           net199643, RN => n100, Q => predict_PC_1_6_port, QN 
                           => net245034);
   predict_PC_reg_1_5_inst : DFFR_X1 port map( D => target_PC_i(5), CK => 
                           net199643, RN => n100, Q => predict_PC_1_5_port, QN 
                           => net245033);
   predict_PC_reg_1_4_inst : DFFR_X1 port map( D => target_PC_i(4), CK => 
                           net199643, RN => n98, Q => predict_PC_1_4_port, QN 
                           => net245032);
   predict_PC_reg_1_3_inst : DFFR_X1 port map( D => target_PC_i(3), CK => 
                           net199643, RN => n111, Q => predict_PC_1_3_port, QN 
                           => net245031);
   predict_PC_reg_1_2_inst : DFFR_X1 port map( D => target_PC_i(2), CK => 
                           net199643, RN => n99, Q => predict_PC_1_2_port, QN 
                           => net245030);
   predict_PC_reg_1_1_inst : DFFR_X1 port map( D => target_PC_i(1), CK => 
                           net199643, RN => n99, Q => predict_PC_1_1_port, QN 
                           => net245029);
   predict_PC_reg_1_0_inst : DFFR_X1 port map( D => target_PC_i(0), CK => 
                           net199643, RN => n101, Q => predict_PC_1_0_port, QN 
                           => net245028);
   predict_PC_reg_2_31_inst : DFFR_X1 port map( D => target_PC_i(31), CK => 
                           net199648, RN => n103, Q => predict_PC_2_31_port, QN
                           => net245027);
   predict_PC_reg_2_30_inst : DFFR_X1 port map( D => target_PC_i(30), CK => 
                           net199648, RN => n112, Q => predict_PC_2_30_port, QN
                           => net245026);
   predict_PC_reg_2_29_inst : DFFR_X1 port map( D => target_PC_i(29), CK => 
                           net199648, RN => n113, Q => predict_PC_2_29_port, QN
                           => net245025);
   predict_PC_reg_2_28_inst : DFFR_X1 port map( D => target_PC_i(28), CK => 
                           net199648, RN => n112, Q => predict_PC_2_28_port, QN
                           => net245024);
   predict_PC_reg_2_27_inst : DFFR_X1 port map( D => target_PC_i(27), CK => 
                           net199648, RN => n98, Q => predict_PC_2_27_port, QN 
                           => net245023);
   predict_PC_reg_2_26_inst : DFFR_X1 port map( D => target_PC_i(26), CK => 
                           net199648, RN => n105, Q => predict_PC_2_26_port, QN
                           => net245022);
   predict_PC_reg_2_25_inst : DFFR_X1 port map( D => target_PC_i(25), CK => 
                           net199648, RN => n109, Q => predict_PC_2_25_port, QN
                           => net245021);
   predict_PC_reg_2_24_inst : DFFR_X1 port map( D => target_PC_i(24), CK => 
                           net199648, RN => n106, Q => predict_PC_2_24_port, QN
                           => net245020);
   predict_PC_reg_2_23_inst : DFFR_X1 port map( D => target_PC_i(23), CK => 
                           net199648, RN => n95, Q => predict_PC_2_23_port, QN 
                           => net245019);
   predict_PC_reg_2_22_inst : DFFR_X1 port map( D => target_PC_i(22), CK => 
                           net199648, RN => n106, Q => predict_PC_2_22_port, QN
                           => net245018);
   predict_PC_reg_2_21_inst : DFFR_X1 port map( D => target_PC_i(21), CK => 
                           net199648, RN => n101, Q => predict_PC_2_21_port, QN
                           => net245017);
   predict_PC_reg_2_20_inst : DFFR_X1 port map( D => target_PC_i(20), CK => 
                           net199648, RN => n102, Q => predict_PC_2_20_port, QN
                           => net245016);
   predict_PC_reg_2_19_inst : DFFR_X1 port map( D => target_PC_i(19), CK => 
                           net199648, RN => n103, Q => predict_PC_2_19_port, QN
                           => net245015);
   predict_PC_reg_2_18_inst : DFFR_X1 port map( D => target_PC_i(18), CK => 
                           net199648, RN => n110, Q => predict_PC_2_18_port, QN
                           => net245014);
   predict_PC_reg_2_17_inst : DFFR_X1 port map( D => target_PC_i(17), CK => 
                           net199648, RN => n107, Q => predict_PC_2_17_port, QN
                           => net245013);
   predict_PC_reg_2_16_inst : DFFR_X1 port map( D => target_PC_i(16), CK => 
                           net199648, RN => n103, Q => predict_PC_2_16_port, QN
                           => net245012);
   predict_PC_reg_2_15_inst : DFFR_X1 port map( D => target_PC_i(15), CK => 
                           net199648, RN => n108, Q => predict_PC_2_15_port, QN
                           => net245011);
   predict_PC_reg_2_14_inst : DFFR_X1 port map( D => target_PC_i(14), CK => 
                           net199648, RN => n109, Q => predict_PC_2_14_port, QN
                           => net245010);
   predict_PC_reg_2_13_inst : DFFR_X1 port map( D => target_PC_i(13), CK => 
                           net199648, RN => n105, Q => predict_PC_2_13_port, QN
                           => net245009);
   predict_PC_reg_2_12_inst : DFFR_X1 port map( D => target_PC_i(12), CK => 
                           net199648, RN => n106, Q => predict_PC_2_12_port, QN
                           => net245008);
   predict_PC_reg_2_11_inst : DFFR_X1 port map( D => target_PC_i(11), CK => 
                           net199648, RN => n104, Q => predict_PC_2_11_port, QN
                           => net245007);
   predict_PC_reg_2_10_inst : DFFR_X1 port map( D => target_PC_i(10), CK => 
                           net199648, RN => n102, Q => predict_PC_2_10_port, QN
                           => net245006);
   predict_PC_reg_2_9_inst : DFFR_X1 port map( D => target_PC_i(9), CK => 
                           net199648, RN => n111, Q => predict_PC_2_9_port, QN 
                           => net245005);
   predict_PC_reg_2_8_inst : DFFR_X1 port map( D => target_PC_i(8), CK => 
                           net199648, RN => n111, Q => predict_PC_2_8_port, QN 
                           => net245004);
   predict_PC_reg_2_7_inst : DFFR_X1 port map( D => target_PC_i(7), CK => 
                           net199648, RN => n111, Q => predict_PC_2_7_port, QN 
                           => net245003);
   predict_PC_reg_2_6_inst : DFFR_X1 port map( D => target_PC_i(6), CK => 
                           net199648, RN => n104, Q => predict_PC_2_6_port, QN 
                           => net245002);
   predict_PC_reg_2_5_inst : DFFR_X1 port map( D => target_PC_i(5), CK => 
                           net199648, RN => n103, Q => predict_PC_2_5_port, QN 
                           => net245001);
   predict_PC_reg_2_4_inst : DFFR_X1 port map( D => target_PC_i(4), CK => 
                           net199648, RN => n112, Q => predict_PC_2_4_port, QN 
                           => net245000);
   predict_PC_reg_2_3_inst : DFFR_X1 port map( D => target_PC_i(3), CK => 
                           net199648, RN => n113, Q => predict_PC_2_3_port, QN 
                           => net244999);
   predict_PC_reg_2_2_inst : DFFR_X1 port map( D => target_PC_i(2), CK => 
                           net199648, RN => n112, Q => predict_PC_2_2_port, QN 
                           => net244998);
   predict_PC_reg_2_1_inst : DFFR_X1 port map( D => target_PC_i(1), CK => 
                           net199648, RN => n97, Q => predict_PC_2_1_port, QN 
                           => net244997);
   predict_PC_reg_2_0_inst : DFFR_X1 port map( D => target_PC_i(0), CK => 
                           net199648, RN => n102, Q => predict_PC_2_0_port, QN 
                           => net244996);
   predict_PC_reg_3_31_inst : DFFR_X1 port map( D => target_PC_i(31), CK => 
                           net199653, RN => n102, Q => predict_PC_3_31_port, QN
                           => net244995);
   predict_PC_reg_3_30_inst : DFFR_X1 port map( D => target_PC_i(30), CK => 
                           net199653, RN => n106, Q => predict_PC_3_30_port, QN
                           => net244994);
   predict_PC_reg_3_29_inst : DFFR_X1 port map( D => target_PC_i(29), CK => 
                           net199653, RN => n101, Q => predict_PC_3_29_port, QN
                           => net244993);
   predict_PC_reg_3_28_inst : DFFR_X1 port map( D => target_PC_i(28), CK => 
                           net199653, RN => n99, Q => predict_PC_3_28_port, QN 
                           => net244992);
   predict_PC_reg_3_27_inst : DFFR_X1 port map( D => target_PC_i(27), CK => 
                           net199653, RN => n112, Q => predict_PC_3_27_port, QN
                           => net244991);
   predict_PC_reg_3_26_inst : DFFR_X1 port map( D => target_PC_i(26), CK => 
                           net199653, RN => n110, Q => predict_PC_3_26_port, QN
                           => net244990);
   predict_PC_reg_3_25_inst : DFFR_X1 port map( D => target_PC_i(25), CK => 
                           net199653, RN => n107, Q => predict_PC_3_25_port, QN
                           => net244989);
   predict_PC_reg_3_24_inst : DFFR_X1 port map( D => target_PC_i(24), CK => 
                           net199653, RN => n97, Q => predict_PC_3_24_port, QN 
                           => net244988);
   predict_PC_reg_3_23_inst : DFFR_X1 port map( D => target_PC_i(23), CK => 
                           net199653, RN => n108, Q => predict_PC_3_23_port, QN
                           => net244987);
   predict_PC_reg_3_22_inst : DFFR_X1 port map( D => target_PC_i(22), CK => 
                           net199653, RN => n109, Q => predict_PC_3_22_port, QN
                           => net244986);
   predict_PC_reg_3_21_inst : DFFR_X1 port map( D => target_PC_i(21), CK => 
                           net199653, RN => n105, Q => predict_PC_3_21_port, QN
                           => net244985);
   predict_PC_reg_3_20_inst : DFFR_X1 port map( D => target_PC_i(20), CK => 
                           net199653, RN => n111, Q => predict_PC_3_20_port, QN
                           => net244984);
   predict_PC_reg_3_19_inst : DFFR_X1 port map( D => target_PC_i(19), CK => 
                           net199653, RN => n111, Q => predict_PC_3_19_port, QN
                           => net244983);
   predict_PC_reg_3_18_inst : DFFR_X1 port map( D => target_PC_i(18), CK => 
                           net199653, RN => n96, Q => predict_PC_3_18_port, QN 
                           => net244982);
   predict_PC_reg_3_17_inst : DFFR_X1 port map( D => target_PC_i(17), CK => 
                           net199653, RN => n112, Q => predict_PC_3_17_port, QN
                           => net244981);
   predict_PC_reg_3_16_inst : DFFR_X1 port map( D => target_PC_i(16), CK => 
                           net199653, RN => n103, Q => predict_PC_3_16_port, QN
                           => net244980);
   predict_PC_reg_3_15_inst : DFFR_X1 port map( D => target_PC_i(15), CK => 
                           net199653, RN => n98, Q => predict_PC_3_15_port, QN 
                           => net244979);
   predict_PC_reg_3_14_inst : DFFR_X1 port map( D => target_PC_i(14), CK => 
                           net199653, RN => n113, Q => predict_PC_3_14_port, QN
                           => net244978);
   predict_PC_reg_3_13_inst : DFFR_X1 port map( D => target_PC_i(13), CK => 
                           net199653, RN => n112, Q => predict_PC_3_13_port, QN
                           => net244977);
   predict_PC_reg_3_12_inst : DFFR_X1 port map( D => target_PC_i(12), CK => 
                           net199653, RN => n110, Q => predict_PC_3_12_port, QN
                           => net244976);
   predict_PC_reg_3_11_inst : DFFR_X1 port map( D => target_PC_i(11), CK => 
                           net199653, RN => n104, Q => predict_PC_3_11_port, QN
                           => net244975);
   predict_PC_reg_3_10_inst : DFFR_X1 port map( D => target_PC_i(10), CK => 
                           net199653, RN => n101, Q => predict_PC_3_10_port, QN
                           => net244974);
   predict_PC_reg_3_9_inst : DFFR_X1 port map( D => target_PC_i(9), CK => 
                           net199653, RN => n99, Q => predict_PC_3_9_port, QN 
                           => net244973);
   predict_PC_reg_3_8_inst : DFFR_X1 port map( D => target_PC_i(8), CK => 
                           net199653, RN => n113, Q => predict_PC_3_8_port, QN 
                           => net244972);
   predict_PC_reg_3_7_inst : DFFR_X1 port map( D => target_PC_i(7), CK => 
                           net199653, RN => n113, Q => predict_PC_3_7_port, QN 
                           => net244971);
   predict_PC_reg_3_6_inst : DFFR_X1 port map( D => target_PC_i(6), CK => 
                           net199653, RN => n110, Q => predict_PC_3_6_port, QN 
                           => net244970);
   predict_PC_reg_3_5_inst : DFFR_X1 port map( D => target_PC_i(5), CK => 
                           net199653, RN => n109, Q => predict_PC_3_5_port, QN 
                           => net244969);
   predict_PC_reg_3_4_inst : DFFR_X1 port map( D => target_PC_i(4), CK => 
                           net199653, RN => n107, Q => predict_PC_3_4_port, QN 
                           => net244968);
   predict_PC_reg_3_3_inst : DFFR_X1 port map( D => target_PC_i(3), CK => 
                           net199653, RN => n108, Q => predict_PC_3_3_port, QN 
                           => net244967);
   predict_PC_reg_3_2_inst : DFFR_X1 port map( D => target_PC_i(2), CK => 
                           net199653, RN => n93, Q => predict_PC_3_2_port, QN 
                           => net244966);
   predict_PC_reg_3_1_inst : DFFR_X1 port map( D => target_PC_i(1), CK => 
                           net199653, RN => n90, Q => predict_PC_3_1_port, QN 
                           => net244965);
   predict_PC_reg_3_0_inst : DFFR_X1 port map( D => target_PC_i(0), CK => 
                           net199653, RN => n91, Q => predict_PC_3_0_port, QN 
                           => net244964);
   predict_PC_reg_4_31_inst : DFFR_X1 port map( D => target_PC_i(31), CK => 
                           net199658, RN => n91, Q => predict_PC_4_31_port, QN 
                           => net244963);
   predict_PC_reg_4_30_inst : DFFR_X1 port map( D => target_PC_i(30), CK => 
                           net199658, RN => n92, Q => predict_PC_4_30_port, QN 
                           => net244962);
   predict_PC_reg_4_29_inst : DFFR_X1 port map( D => target_PC_i(29), CK => 
                           net199658, RN => n90, Q => predict_PC_4_29_port, QN 
                           => net244961);
   predict_PC_reg_4_28_inst : DFFR_X1 port map( D => target_PC_i(28), CK => 
                           net199658, RN => n92, Q => predict_PC_4_28_port, QN 
                           => net244960);
   predict_PC_reg_4_27_inst : DFFR_X1 port map( D => target_PC_i(27), CK => 
                           net199658, RN => n91, Q => predict_PC_4_27_port, QN 
                           => net244959);
   predict_PC_reg_4_26_inst : DFFR_X1 port map( D => target_PC_i(26), CK => 
                           net199658, RN => n92, Q => predict_PC_4_26_port, QN 
                           => net244958);
   predict_PC_reg_4_25_inst : DFFR_X1 port map( D => target_PC_i(25), CK => 
                           net199658, RN => n90, Q => predict_PC_4_25_port, QN 
                           => net244957);
   predict_PC_reg_4_24_inst : DFFR_X1 port map( D => target_PC_i(24), CK => 
                           net199658, RN => n90, Q => predict_PC_4_24_port, QN 
                           => net244956);
   predict_PC_reg_4_23_inst : DFFR_X1 port map( D => target_PC_i(23), CK => 
                           net199658, RN => n91, Q => predict_PC_4_23_port, QN 
                           => net244955);
   predict_PC_reg_4_22_inst : DFFR_X1 port map( D => target_PC_i(22), CK => 
                           net199658, RN => n91, Q => predict_PC_4_22_port, QN 
                           => net244954);
   predict_PC_reg_4_21_inst : DFFR_X1 port map( D => target_PC_i(21), CK => 
                           net199658, RN => n90, Q => predict_PC_4_21_port, QN 
                           => net244953);
   predict_PC_reg_4_20_inst : DFFR_X1 port map( D => target_PC_i(20), CK => 
                           net199658, RN => n91, Q => predict_PC_4_20_port, QN 
                           => net244952);
   predict_PC_reg_4_19_inst : DFFR_X1 port map( D => target_PC_i(19), CK => 
                           net199658, RN => n92, Q => predict_PC_4_19_port, QN 
                           => net244951);
   predict_PC_reg_4_18_inst : DFFR_X1 port map( D => target_PC_i(18), CK => 
                           net199658, RN => n90, Q => predict_PC_4_18_port, QN 
                           => net244950);
   predict_PC_reg_4_17_inst : DFFR_X1 port map( D => target_PC_i(17), CK => 
                           net199658, RN => n91, Q => predict_PC_4_17_port, QN 
                           => net244949);
   predict_PC_reg_4_16_inst : DFFR_X1 port map( D => target_PC_i(16), CK => 
                           net199658, RN => n92, Q => predict_PC_4_16_port, QN 
                           => net244948);
   predict_PC_reg_4_15_inst : DFFR_X1 port map( D => target_PC_i(15), CK => 
                           net199658, RN => n90, Q => predict_PC_4_15_port, QN 
                           => net244947);
   predict_PC_reg_4_14_inst : DFFR_X1 port map( D => target_PC_i(14), CK => 
                           net199658, RN => n91, Q => predict_PC_4_14_port, QN 
                           => net244946);
   predict_PC_reg_4_13_inst : DFFR_X1 port map( D => target_PC_i(13), CK => 
                           net199658, RN => n92, Q => predict_PC_4_13_port, QN 
                           => net244945);
   predict_PC_reg_4_12_inst : DFFR_X1 port map( D => target_PC_i(12), CK => 
                           net199658, RN => n90, Q => predict_PC_4_12_port, QN 
                           => net244944);
   predict_PC_reg_4_11_inst : DFFR_X1 port map( D => target_PC_i(11), CK => 
                           net199658, RN => n91, Q => predict_PC_4_11_port, QN 
                           => net244943);
   predict_PC_reg_4_10_inst : DFFR_X1 port map( D => target_PC_i(10), CK => 
                           net199658, RN => n90, Q => predict_PC_4_10_port, QN 
                           => net244942);
   predict_PC_reg_4_9_inst : DFFR_X1 port map( D => target_PC_i(9), CK => 
                           net199658, RN => n90, Q => predict_PC_4_9_port, QN 
                           => net244941);
   predict_PC_reg_4_8_inst : DFFR_X1 port map( D => target_PC_i(8), CK => 
                           net199658, RN => n90, Q => predict_PC_4_8_port, QN 
                           => net244940);
   predict_PC_reg_4_7_inst : DFFR_X1 port map( D => target_PC_i(7), CK => 
                           net199658, RN => n90, Q => predict_PC_4_7_port, QN 
                           => net244939);
   predict_PC_reg_4_6_inst : DFFR_X1 port map( D => target_PC_i(6), CK => 
                           net199658, RN => n90, Q => predict_PC_4_6_port, QN 
                           => net244938);
   predict_PC_reg_4_5_inst : DFFR_X1 port map( D => target_PC_i(5), CK => 
                           net199658, RN => n90, Q => predict_PC_4_5_port, QN 
                           => net244937);
   predict_PC_reg_4_4_inst : DFFR_X1 port map( D => target_PC_i(4), CK => 
                           net199658, RN => n90, Q => predict_PC_4_4_port, QN 
                           => net244936);
   predict_PC_reg_4_3_inst : DFFR_X1 port map( D => target_PC_i(3), CK => 
                           net199658, RN => n90, Q => predict_PC_4_3_port, QN 
                           => net244935);
   predict_PC_reg_4_2_inst : DFFR_X1 port map( D => target_PC_i(2), CK => 
                           net199658, RN => n90, Q => predict_PC_4_2_port, QN 
                           => net244934);
   predict_PC_reg_4_1_inst : DFFR_X1 port map( D => target_PC_i(1), CK => 
                           net199658, RN => n90, Q => predict_PC_4_1_port, QN 
                           => net244933);
   predict_PC_reg_4_0_inst : DFFR_X1 port map( D => target_PC_i(0), CK => 
                           net199658, RN => n90, Q => predict_PC_4_0_port, QN 
                           => net244932);
   predict_PC_reg_5_31_inst : DFFR_X1 port map( D => target_PC_i(31), CK => 
                           net199663, RN => n90, Q => predict_PC_5_31_port, QN 
                           => net244931);
   predict_PC_reg_5_30_inst : DFFR_X1 port map( D => target_PC_i(30), CK => 
                           net199663, RN => n91, Q => predict_PC_5_30_port, QN 
                           => net244930);
   predict_PC_reg_5_29_inst : DFFR_X1 port map( D => target_PC_i(29), CK => 
                           net199663, RN => n91, Q => predict_PC_5_29_port, QN 
                           => net244929);
   predict_PC_reg_5_28_inst : DFFR_X1 port map( D => target_PC_i(28), CK => 
                           net199663, RN => n91, Q => predict_PC_5_28_port, QN 
                           => net244928);
   predict_PC_reg_5_27_inst : DFFR_X1 port map( D => target_PC_i(27), CK => 
                           net199663, RN => n91, Q => predict_PC_5_27_port, QN 
                           => net244927);
   predict_PC_reg_5_26_inst : DFFR_X1 port map( D => target_PC_i(26), CK => 
                           net199663, RN => n91, Q => predict_PC_5_26_port, QN 
                           => net244926);
   predict_PC_reg_5_25_inst : DFFR_X1 port map( D => target_PC_i(25), CK => 
                           net199663, RN => n91, Q => predict_PC_5_25_port, QN 
                           => net244925);
   predict_PC_reg_5_24_inst : DFFR_X1 port map( D => target_PC_i(24), CK => 
                           net199663, RN => n91, Q => predict_PC_5_24_port, QN 
                           => net244924);
   predict_PC_reg_5_23_inst : DFFR_X1 port map( D => target_PC_i(23), CK => 
                           net199663, RN => n91, Q => predict_PC_5_23_port, QN 
                           => net244923);
   predict_PC_reg_5_22_inst : DFFR_X1 port map( D => target_PC_i(22), CK => 
                           net199663, RN => n91, Q => predict_PC_5_22_port, QN 
                           => net244922);
   predict_PC_reg_5_21_inst : DFFR_X1 port map( D => target_PC_i(21), CK => 
                           net199663, RN => n91, Q => predict_PC_5_21_port, QN 
                           => net244921);
   predict_PC_reg_5_20_inst : DFFR_X1 port map( D => target_PC_i(20), CK => 
                           net199663, RN => n91, Q => predict_PC_5_20_port, QN 
                           => net244920);
   predict_PC_reg_5_19_inst : DFFR_X1 port map( D => target_PC_i(19), CK => 
                           net199663, RN => n91, Q => predict_PC_5_19_port, QN 
                           => net244919);
   predict_PC_reg_5_18_inst : DFFR_X1 port map( D => target_PC_i(18), CK => 
                           net199663, RN => n92, Q => predict_PC_5_18_port, QN 
                           => net244918);
   predict_PC_reg_5_17_inst : DFFR_X1 port map( D => target_PC_i(17), CK => 
                           net199663, RN => n92, Q => predict_PC_5_17_port, QN 
                           => net244917);
   predict_PC_reg_5_16_inst : DFFR_X1 port map( D => target_PC_i(16), CK => 
                           net199663, RN => n92, Q => predict_PC_5_16_port, QN 
                           => net244916);
   predict_PC_reg_5_15_inst : DFFR_X1 port map( D => target_PC_i(15), CK => 
                           net199663, RN => n92, Q => predict_PC_5_15_port, QN 
                           => net244915);
   predict_PC_reg_5_14_inst : DFFR_X1 port map( D => target_PC_i(14), CK => 
                           net199663, RN => n92, Q => predict_PC_5_14_port, QN 
                           => net244914);
   predict_PC_reg_5_13_inst : DFFR_X1 port map( D => target_PC_i(13), CK => 
                           net199663, RN => n92, Q => predict_PC_5_13_port, QN 
                           => net244913);
   predict_PC_reg_5_12_inst : DFFR_X1 port map( D => target_PC_i(12), CK => 
                           net199663, RN => n92, Q => predict_PC_5_12_port, QN 
                           => net244912);
   predict_PC_reg_5_11_inst : DFFR_X1 port map( D => target_PC_i(11), CK => 
                           net199663, RN => n92, Q => predict_PC_5_11_port, QN 
                           => net244911);
   predict_PC_reg_5_10_inst : DFFR_X1 port map( D => target_PC_i(10), CK => 
                           net199663, RN => n92, Q => predict_PC_5_10_port, QN 
                           => net244910);
   predict_PC_reg_5_9_inst : DFFR_X1 port map( D => target_PC_i(9), CK => 
                           net199663, RN => n92, Q => predict_PC_5_9_port, QN 
                           => net244909);
   predict_PC_reg_5_8_inst : DFFR_X1 port map( D => target_PC_i(8), CK => 
                           net199663, RN => n92, Q => predict_PC_5_8_port, QN 
                           => net244908);
   predict_PC_reg_5_7_inst : DFFR_X1 port map( D => target_PC_i(7), CK => 
                           net199663, RN => n92, Q => predict_PC_5_7_port, QN 
                           => net244907);
   predict_PC_reg_5_6_inst : DFFR_X1 port map( D => target_PC_i(6), CK => 
                           net199663, RN => n93, Q => predict_PC_5_6_port, QN 
                           => net244906);
   predict_PC_reg_5_5_inst : DFFR_X1 port map( D => target_PC_i(5), CK => 
                           net199663, RN => n94, Q => predict_PC_5_5_port, QN 
                           => net244905);
   predict_PC_reg_5_4_inst : DFFR_X1 port map( D => target_PC_i(4), CK => 
                           net199663, RN => n95, Q => predict_PC_5_4_port, QN 
                           => net244904);
   predict_PC_reg_5_3_inst : DFFR_X1 port map( D => target_PC_i(3), CK => 
                           net199663, RN => n96, Q => predict_PC_5_3_port, QN 
                           => net244903);
   predict_PC_reg_5_2_inst : DFFR_X1 port map( D => target_PC_i(2), CK => 
                           net199663, RN => n96, Q => predict_PC_5_2_port, QN 
                           => net244902);
   predict_PC_reg_5_1_inst : DFFR_X1 port map( D => target_PC_i(1), CK => 
                           net199663, RN => n93, Q => predict_PC_5_1_port, QN 
                           => net244901);
   predict_PC_reg_5_0_inst : DFFR_X1 port map( D => target_PC_i(0), CK => 
                           net199663, RN => n94, Q => predict_PC_5_0_port, QN 
                           => net244900);
   predict_PC_reg_6_31_inst : DFFR_X1 port map( D => target_PC_i(31), CK => 
                           net199668, RN => n95, Q => predict_PC_6_31_port, QN 
                           => net244899);
   predict_PC_reg_6_30_inst : DFFR_X1 port map( D => target_PC_i(30), CK => 
                           net199668, RN => n96, Q => predict_PC_6_30_port, QN 
                           => net244898);
   predict_PC_reg_6_29_inst : DFFR_X1 port map( D => target_PC_i(29), CK => 
                           net199668, RN => n96, Q => predict_PC_6_29_port, QN 
                           => net244897);
   predict_PC_reg_6_28_inst : DFFR_X1 port map( D => target_PC_i(28), CK => 
                           net199668, RN => n94, Q => predict_PC_6_28_port, QN 
                           => net244896);
   predict_PC_reg_6_27_inst : DFFR_X1 port map( D => target_PC_i(27), CK => 
                           net199668, RN => n94, Q => predict_PC_6_27_port, QN 
                           => net244895);
   predict_PC_reg_6_26_inst : DFFR_X1 port map( D => target_PC_i(26), CK => 
                           net199668, RN => n95, Q => predict_PC_6_26_port, QN 
                           => net244894);
   predict_PC_reg_6_25_inst : DFFR_X1 port map( D => target_PC_i(25), CK => 
                           net199668, RN => n96, Q => predict_PC_6_25_port, QN 
                           => net244893);
   predict_PC_reg_6_24_inst : DFFR_X1 port map( D => target_PC_i(24), CK => 
                           net199668, RN => n93, Q => predict_PC_6_24_port, QN 
                           => net244892);
   predict_PC_reg_6_23_inst : DFFR_X1 port map( D => target_PC_i(23), CK => 
                           net199668, RN => n94, Q => predict_PC_6_23_port, QN 
                           => net244891);
   predict_PC_reg_6_22_inst : DFFR_X1 port map( D => target_PC_i(22), CK => 
                           net199668, RN => n95, Q => predict_PC_6_22_port, QN 
                           => net244890);
   predict_PC_reg_6_21_inst : DFFR_X1 port map( D => target_PC_i(21), CK => 
                           net199668, RN => n96, Q => predict_PC_6_21_port, QN 
                           => net244889);
   predict_PC_reg_6_20_inst : DFFR_X1 port map( D => target_PC_i(20), CK => 
                           net199668, RN => n93, Q => predict_PC_6_20_port, QN 
                           => net244888);
   predict_PC_reg_6_19_inst : DFFR_X1 port map( D => target_PC_i(19), CK => 
                           net199668, RN => n94, Q => predict_PC_6_19_port, QN 
                           => net244887);
   predict_PC_reg_6_18_inst : DFFR_X1 port map( D => target_PC_i(18), CK => 
                           net199668, RN => n95, Q => predict_PC_6_18_port, QN 
                           => net244886);
   predict_PC_reg_6_17_inst : DFFR_X1 port map( D => target_PC_i(17), CK => 
                           net199668, RN => n96, Q => predict_PC_6_17_port, QN 
                           => net244885);
   predict_PC_reg_6_16_inst : DFFR_X1 port map( D => target_PC_i(16), CK => 
                           net199668, RN => n93, Q => predict_PC_6_16_port, QN 
                           => net244884);
   predict_PC_reg_6_15_inst : DFFR_X1 port map( D => target_PC_i(15), CK => 
                           net199668, RN => n93, Q => predict_PC_6_15_port, QN 
                           => net244883);
   predict_PC_reg_6_14_inst : DFFR_X1 port map( D => target_PC_i(14), CK => 
                           net199668, RN => n93, Q => predict_PC_6_14_port, QN 
                           => net244882);
   predict_PC_reg_6_13_inst : DFFR_X1 port map( D => target_PC_i(13), CK => 
                           net199668, RN => n93, Q => predict_PC_6_13_port, QN 
                           => net244881);
   predict_PC_reg_6_12_inst : DFFR_X1 port map( D => target_PC_i(12), CK => 
                           net199668, RN => n93, Q => predict_PC_6_12_port, QN 
                           => net244880);
   predict_PC_reg_6_11_inst : DFFR_X1 port map( D => target_PC_i(11), CK => 
                           net199668, RN => n93, Q => predict_PC_6_11_port, QN 
                           => net244879);
   predict_PC_reg_6_10_inst : DFFR_X1 port map( D => target_PC_i(10), CK => 
                           net199668, RN => n93, Q => predict_PC_6_10_port, QN 
                           => net244878);
   predict_PC_reg_6_9_inst : DFFR_X1 port map( D => target_PC_i(9), CK => 
                           net199668, RN => n93, Q => predict_PC_6_9_port, QN 
                           => net244877);
   predict_PC_reg_6_8_inst : DFFR_X1 port map( D => target_PC_i(8), CK => 
                           net199668, RN => n93, Q => predict_PC_6_8_port, QN 
                           => net244876);
   predict_PC_reg_6_7_inst : DFFR_X1 port map( D => target_PC_i(7), CK => 
                           net199668, RN => n93, Q => predict_PC_6_7_port, QN 
                           => net244875);
   predict_PC_reg_6_6_inst : DFFR_X1 port map( D => target_PC_i(6), CK => 
                           net199668, RN => n93, Q => predict_PC_6_6_port, QN 
                           => net244874);
   predict_PC_reg_6_5_inst : DFFR_X1 port map( D => target_PC_i(5), CK => 
                           net199668, RN => n93, Q => predict_PC_6_5_port, QN 
                           => net244873);
   predict_PC_reg_6_4_inst : DFFR_X1 port map( D => target_PC_i(4), CK => 
                           net199668, RN => n93, Q => predict_PC_6_4_port, QN 
                           => net244872);
   predict_PC_reg_6_3_inst : DFFR_X1 port map( D => target_PC_i(3), CK => 
                           net199668, RN => n94, Q => predict_PC_6_3_port, QN 
                           => net244871);
   predict_PC_reg_6_2_inst : DFFR_X1 port map( D => target_PC_i(2), CK => 
                           net199668, RN => n94, Q => predict_PC_6_2_port, QN 
                           => net244870);
   predict_PC_reg_6_1_inst : DFFR_X1 port map( D => target_PC_i(1), CK => 
                           net199668, RN => n94, Q => predict_PC_6_1_port, QN 
                           => net244869);
   predict_PC_reg_6_0_inst : DFFR_X1 port map( D => target_PC_i(0), CK => 
                           net199668, RN => n94, Q => predict_PC_6_0_port, QN 
                           => net244868);
   predict_PC_reg_7_31_inst : DFFR_X1 port map( D => target_PC_i(31), CK => 
                           net199673, RN => n94, Q => predict_PC_7_31_port, QN 
                           => net244867);
   predict_PC_reg_7_30_inst : DFFR_X1 port map( D => target_PC_i(30), CK => 
                           net199673, RN => n94, Q => predict_PC_7_30_port, QN 
                           => net244866);
   predict_PC_reg_7_29_inst : DFFR_X1 port map( D => target_PC_i(29), CK => 
                           net199673, RN => n94, Q => predict_PC_7_29_port, QN 
                           => net244865);
   predict_PC_reg_7_28_inst : DFFR_X1 port map( D => target_PC_i(28), CK => 
                           net199673, RN => n94, Q => predict_PC_7_28_port, QN 
                           => net244864);
   predict_PC_reg_7_27_inst : DFFR_X1 port map( D => target_PC_i(27), CK => 
                           net199673, RN => n94, Q => predict_PC_7_27_port, QN 
                           => net244863);
   predict_PC_reg_7_26_inst : DFFR_X1 port map( D => target_PC_i(26), CK => 
                           net199673, RN => n94, Q => predict_PC_7_26_port, QN 
                           => net244862);
   predict_PC_reg_7_25_inst : DFFR_X1 port map( D => target_PC_i(25), CK => 
                           net199673, RN => n94, Q => predict_PC_7_25_port, QN 
                           => net244861);
   predict_PC_reg_7_24_inst : DFFR_X1 port map( D => target_PC_i(24), CK => 
                           net199673, RN => n94, Q => predict_PC_7_24_port, QN 
                           => net244860);
   predict_PC_reg_7_23_inst : DFFR_X1 port map( D => target_PC_i(23), CK => 
                           net199673, RN => n95, Q => predict_PC_7_23_port, QN 
                           => net244859);
   predict_PC_reg_7_22_inst : DFFR_X1 port map( D => target_PC_i(22), CK => 
                           net199673, RN => n95, Q => predict_PC_7_22_port, QN 
                           => net244858);
   predict_PC_reg_7_21_inst : DFFR_X1 port map( D => target_PC_i(21), CK => 
                           net199673, RN => n95, Q => predict_PC_7_21_port, QN 
                           => net244857);
   predict_PC_reg_7_20_inst : DFFR_X1 port map( D => target_PC_i(20), CK => 
                           net199673, RN => n95, Q => predict_PC_7_20_port, QN 
                           => net244856);
   predict_PC_reg_7_19_inst : DFFR_X1 port map( D => target_PC_i(19), CK => 
                           net199673, RN => n95, Q => predict_PC_7_19_port, QN 
                           => net244855);
   predict_PC_reg_7_18_inst : DFFR_X1 port map( D => target_PC_i(18), CK => 
                           net199673, RN => n95, Q => predict_PC_7_18_port, QN 
                           => net244854);
   predict_PC_reg_7_17_inst : DFFR_X1 port map( D => target_PC_i(17), CK => 
                           net199673, RN => n95, Q => predict_PC_7_17_port, QN 
                           => net244853);
   predict_PC_reg_7_16_inst : DFFR_X1 port map( D => target_PC_i(16), CK => 
                           net199673, RN => n95, Q => predict_PC_7_16_port, QN 
                           => net244852);
   predict_PC_reg_7_15_inst : DFFR_X1 port map( D => target_PC_i(15), CK => 
                           net199673, RN => n95, Q => predict_PC_7_15_port, QN 
                           => net244851);
   predict_PC_reg_7_14_inst : DFFR_X1 port map( D => target_PC_i(14), CK => 
                           net199673, RN => n95, Q => predict_PC_7_14_port, QN 
                           => net244850);
   predict_PC_reg_7_13_inst : DFFR_X1 port map( D => target_PC_i(13), CK => 
                           net199673, RN => n95, Q => predict_PC_7_13_port, QN 
                           => net244849);
   predict_PC_reg_7_12_inst : DFFR_X1 port map( D => target_PC_i(12), CK => 
                           net199673, RN => n95, Q => predict_PC_7_12_port, QN 
                           => net244848);
   predict_PC_reg_7_11_inst : DFFR_X1 port map( D => target_PC_i(11), CK => 
                           net199673, RN => n96, Q => predict_PC_7_11_port, QN 
                           => net244847);
   predict_PC_reg_7_10_inst : DFFR_X1 port map( D => target_PC_i(10), CK => 
                           net199673, RN => n96, Q => predict_PC_7_10_port, QN 
                           => net244846);
   predict_PC_reg_7_9_inst : DFFR_X1 port map( D => target_PC_i(9), CK => 
                           net199673, RN => n96, Q => predict_PC_7_9_port, QN 
                           => net244845);
   predict_PC_reg_7_8_inst : DFFR_X1 port map( D => target_PC_i(8), CK => 
                           net199673, RN => n96, Q => predict_PC_7_8_port, QN 
                           => net244844);
   predict_PC_reg_7_7_inst : DFFR_X1 port map( D => target_PC_i(7), CK => 
                           net199673, RN => n96, Q => predict_PC_7_7_port, QN 
                           => net244843);
   predict_PC_reg_7_6_inst : DFFR_X1 port map( D => target_PC_i(6), CK => 
                           net199673, RN => n96, Q => predict_PC_7_6_port, QN 
                           => net244842);
   predict_PC_reg_7_5_inst : DFFR_X1 port map( D => target_PC_i(5), CK => 
                           net199673, RN => n96, Q => predict_PC_7_5_port, QN 
                           => net244841);
   predict_PC_reg_7_4_inst : DFFR_X1 port map( D => target_PC_i(4), CK => 
                           net199673, RN => n96, Q => predict_PC_7_4_port, QN 
                           => net244840);
   predict_PC_reg_7_3_inst : DFFR_X1 port map( D => target_PC_i(3), CK => 
                           net199673, RN => n96, Q => predict_PC_7_3_port, QN 
                           => net244839);
   predict_PC_reg_7_2_inst : DFFR_X1 port map( D => target_PC_i(2), CK => 
                           net199673, RN => n96, Q => predict_PC_7_2_port, QN 
                           => net244838);
   predict_PC_reg_7_1_inst : DFFR_X1 port map( D => target_PC_i(1), CK => 
                           net199673, RN => n96, Q => predict_PC_7_1_port, QN 
                           => net244837);
   predict_PC_reg_7_0_inst : DFFR_X1 port map( D => target_PC_i(0), CK => 
                           net199673, RN => n96, Q => predict_PC_7_0_port, QN 
                           => net244836);
   predict_PC_reg_8_31_inst : DFFR_X1 port map( D => target_PC_i(31), CK => 
                           net199678, RN => n95, Q => predict_PC_8_31_port, QN 
                           => net244835);
   predict_PC_reg_8_30_inst : DFFR_X1 port map( D => target_PC_i(30), CK => 
                           net199678, RN => n94, Q => predict_PC_8_30_port, QN 
                           => net244834);
   predict_PC_reg_8_29_inst : DFFR_X1 port map( D => target_PC_i(29), CK => 
                           net199678, RN => n93, Q => predict_PC_8_29_port, QN 
                           => net244833);
   predict_PC_reg_8_28_inst : DFFR_X1 port map( D => target_PC_i(28), CK => 
                           net199678, RN => n94, Q => predict_PC_8_28_port, QN 
                           => net244832);
   predict_PC_reg_8_27_inst : DFFR_X1 port map( D => target_PC_i(27), CK => 
                           net199678, RN => n95, Q => predict_PC_8_27_port, QN 
                           => net244831);
   predict_PC_reg_8_26_inst : DFFR_X1 port map( D => target_PC_i(26), CK => 
                           net199678, RN => n96, Q => predict_PC_8_26_port, QN 
                           => net244830);
   predict_PC_reg_8_25_inst : DFFR_X1 port map( D => target_PC_i(25), CK => 
                           net199678, RN => n93, Q => predict_PC_8_25_port, QN 
                           => net244829);
   predict_PC_reg_8_24_inst : DFFR_X1 port map( D => target_PC_i(24), CK => 
                           net199678, RN => n95, Q => predict_PC_8_24_port, QN 
                           => net244828);
   predict_PC_reg_8_23_inst : DFFR_X1 port map( D => target_PC_i(23), CK => 
                           net199678, RN => n93, Q => predict_PC_8_23_port, QN 
                           => net244827);
   predict_PC_reg_8_22_inst : DFFR_X1 port map( D => target_PC_i(22), CK => 
                           net199678, RN => n102, Q => predict_PC_8_22_port, QN
                           => net244826);
   predict_PC_reg_8_21_inst : DFFR_X1 port map( D => target_PC_i(21), CK => 
                           net199678, RN => n97, Q => predict_PC_8_21_port, QN 
                           => net244825);
   predict_PC_reg_8_20_inst : DFFR_X1 port map( D => target_PC_i(20), CK => 
                           net199678, RN => n97, Q => predict_PC_8_20_port, QN 
                           => net244824);
   predict_PC_reg_8_19_inst : DFFR_X1 port map( D => target_PC_i(19), CK => 
                           net199678, RN => n103, Q => predict_PC_8_19_port, QN
                           => net244823);
   predict_PC_reg_8_18_inst : DFFR_X1 port map( D => target_PC_i(18), CK => 
                           net199678, RN => n103, Q => predict_PC_8_18_port, QN
                           => net244822);
   predict_PC_reg_8_17_inst : DFFR_X1 port map( D => target_PC_i(17), CK => 
                           net199678, RN => n113, Q => predict_PC_8_17_port, QN
                           => net244821);
   predict_PC_reg_8_16_inst : DFFR_X1 port map( D => target_PC_i(16), CK => 
                           net199678, RN => n112, Q => predict_PC_8_16_port, QN
                           => net244820);
   predict_PC_reg_8_15_inst : DFFR_X1 port map( D => target_PC_i(15), CK => 
                           net199678, RN => n106, Q => predict_PC_8_15_port, QN
                           => net244819);
   predict_PC_reg_8_14_inst : DFFR_X1 port map( D => target_PC_i(14), CK => 
                           net199678, RN => n96, Q => predict_PC_8_14_port, QN 
                           => net244818);
   predict_PC_reg_8_13_inst : DFFR_X1 port map( D => target_PC_i(13), CK => 
                           net199678, RN => n106, Q => predict_PC_8_13_port, QN
                           => net244817);
   predict_PC_reg_8_12_inst : DFFR_X1 port map( D => target_PC_i(12), CK => 
                           net199678, RN => n101, Q => predict_PC_8_12_port, QN
                           => net244816);
   predict_PC_reg_8_11_inst : DFFR_X1 port map( D => target_PC_i(11), CK => 
                           net199678, RN => n110, Q => predict_PC_8_11_port, QN
                           => net244815);
   predict_PC_reg_8_10_inst : DFFR_X1 port map( D => target_PC_i(10), CK => 
                           net199678, RN => n109, Q => predict_PC_8_10_port, QN
                           => net244814);
   predict_PC_reg_8_9_inst : DFFR_X1 port map( D => target_PC_i(9), CK => 
                           net199678, RN => n105, Q => predict_PC_8_9_port, QN 
                           => net244813);
   predict_PC_reg_8_8_inst : DFFR_X1 port map( D => target_PC_i(8), CK => 
                           net199678, RN => n104, Q => predict_PC_8_8_port, QN 
                           => net244812);
   predict_PC_reg_8_7_inst : DFFR_X1 port map( D => target_PC_i(7), CK => 
                           net199678, RN => n102, Q => predict_PC_8_7_port, QN 
                           => net244811);
   predict_PC_reg_8_6_inst : DFFR_X1 port map( D => target_PC_i(6), CK => 
                           net199678, RN => n111, Q => predict_PC_8_6_port, QN 
                           => net244810);
   predict_PC_reg_8_5_inst : DFFR_X1 port map( D => target_PC_i(5), CK => 
                           net199678, RN => n103, Q => predict_PC_8_5_port, QN 
                           => net244809);
   predict_PC_reg_8_4_inst : DFFR_X1 port map( D => target_PC_i(4), CK => 
                           net199678, RN => n103, Q => predict_PC_8_4_port, QN 
                           => net244808);
   predict_PC_reg_8_3_inst : DFFR_X1 port map( D => target_PC_i(3), CK => 
                           net199678, RN => n103, Q => predict_PC_8_3_port, QN 
                           => net244807);
   predict_PC_reg_8_2_inst : DFFR_X1 port map( D => target_PC_i(2), CK => 
                           net199678, RN => n113, Q => predict_PC_8_2_port, QN 
                           => net244806);
   predict_PC_reg_8_1_inst : DFFR_X1 port map( D => target_PC_i(1), CK => 
                           net199678, RN => n113, Q => predict_PC_8_1_port, QN 
                           => net244805);
   predict_PC_reg_8_0_inst : DFFR_X1 port map( D => target_PC_i(0), CK => 
                           net199678, RN => n112, Q => predict_PC_8_0_port, QN 
                           => net244804);
   predict_PC_reg_9_31_inst : DFFR_X1 port map( D => target_PC_i(31), CK => 
                           net199683, RN => n101, Q => predict_PC_9_31_port, QN
                           => net244803);
   predict_PC_reg_9_30_inst : DFFR_X1 port map( D => target_PC_i(30), CK => 
                           net199683, RN => n107, Q => predict_PC_9_30_port, QN
                           => net244802);
   predict_PC_reg_9_29_inst : DFFR_X1 port map( D => target_PC_i(29), CK => 
                           net199683, RN => n108, Q => predict_PC_9_29_port, QN
                           => net244801);
   predict_PC_reg_9_28_inst : DFFR_X1 port map( D => target_PC_i(28), CK => 
                           net199683, RN => n109, Q => predict_PC_9_28_port, QN
                           => net244800);
   predict_PC_reg_9_27_inst : DFFR_X1 port map( D => target_PC_i(27), CK => 
                           net199683, RN => n105, Q => predict_PC_9_27_port, QN
                           => net244799);
   predict_PC_reg_9_26_inst : DFFR_X1 port map( D => target_PC_i(26), CK => 
                           net199683, RN => n104, Q => predict_PC_9_26_port, QN
                           => net244798);
   predict_PC_reg_9_25_inst : DFFR_X1 port map( D => target_PC_i(25), CK => 
                           net199683, RN => n102, Q => predict_PC_9_25_port, QN
                           => net244797);
   predict_PC_reg_9_24_inst : DFFR_X1 port map( D => target_PC_i(24), CK => 
                           net199683, RN => n111, Q => predict_PC_9_24_port, QN
                           => net244796);
   predict_PC_reg_9_23_inst : DFFR_X1 port map( D => target_PC_i(23), CK => 
                           net199683, RN => n113, Q => predict_PC_9_23_port, QN
                           => net244795);
   predict_PC_reg_9_22_inst : DFFR_X1 port map( D => target_PC_i(22), CK => 
                           net199683, RN => n113, Q => predict_PC_9_22_port, QN
                           => net244794);
   predict_PC_reg_9_21_inst : DFFR_X1 port map( D => target_PC_i(21), CK => 
                           net199683, RN => n98, Q => predict_PC_9_21_port, QN 
                           => net244793);
   predict_PC_reg_9_20_inst : DFFR_X1 port map( D => target_PC_i(20), CK => 
                           net199683, RN => n97, Q => predict_PC_9_20_port, QN 
                           => net244792);
   predict_PC_reg_9_19_inst : DFFR_X1 port map( D => target_PC_i(19), CK => 
                           net199683, RN => n103, Q => predict_PC_9_19_port, QN
                           => net244791);
   predict_PC_reg_9_18_inst : DFFR_X1 port map( D => target_PC_i(18), CK => 
                           net199683, RN => n103, Q => predict_PC_9_18_port, QN
                           => net244790);
   predict_PC_reg_9_17_inst : DFFR_X1 port map( D => target_PC_i(17), CK => 
                           net199683, RN => n110, Q => predict_PC_9_17_port, QN
                           => net244789);
   predict_PC_reg_9_16_inst : DFFR_X1 port map( D => target_PC_i(16), CK => 
                           net199683, RN => n107, Q => predict_PC_9_16_port, QN
                           => net244788);
   predict_PC_reg_9_15_inst : DFFR_X1 port map( D => target_PC_i(15), CK => 
                           net199683, RN => n108, Q => predict_PC_9_15_port, QN
                           => net244787);
   predict_PC_reg_9_14_inst : DFFR_X1 port map( D => target_PC_i(14), CK => 
                           net199683, RN => n109, Q => predict_PC_9_14_port, QN
                           => net244786);
   predict_PC_reg_9_13_inst : DFFR_X1 port map( D => target_PC_i(13), CK => 
                           net199683, RN => n105, Q => predict_PC_9_13_port, QN
                           => net244785);
   predict_PC_reg_9_12_inst : DFFR_X1 port map( D => target_PC_i(12), CK => 
                           net199683, RN => n100, Q => predict_PC_9_12_port, QN
                           => net244784);
   predict_PC_reg_9_11_inst : DFFR_X1 port map( D => target_PC_i(11), CK => 
                           net199683, RN => n104, Q => predict_PC_9_11_port, QN
                           => net244783);
   predict_PC_reg_9_10_inst : DFFR_X1 port map( D => target_PC_i(10), CK => 
                           net199683, RN => n102, Q => predict_PC_9_10_port, QN
                           => net244782);
   predict_PC_reg_9_9_inst : DFFR_X1 port map( D => target_PC_i(9), CK => 
                           net199683, RN => n99, Q => predict_PC_9_9_port, QN 
                           => net244781);
   predict_PC_reg_9_8_inst : DFFR_X1 port map( D => target_PC_i(8), CK => 
                           net199683, RN => n111, Q => predict_PC_9_8_port, QN 
                           => net244780);
   predict_PC_reg_9_7_inst : DFFR_X1 port map( D => target_PC_i(7), CK => 
                           net199683, RN => n113, Q => predict_PC_9_7_port, QN 
                           => net244779);
   predict_PC_reg_9_6_inst : DFFR_X1 port map( D => target_PC_i(6), CK => 
                           net199683, RN => n106, Q => predict_PC_9_6_port, QN 
                           => net244778);
   predict_PC_reg_9_5_inst : DFFR_X1 port map( D => target_PC_i(5), CK => 
                           net199683, RN => n101, Q => predict_PC_9_5_port, QN 
                           => net244777);
   predict_PC_reg_9_4_inst : DFFR_X1 port map( D => target_PC_i(4), CK => 
                           net199683, RN => n113, Q => predict_PC_9_4_port, QN 
                           => net244776);
   predict_PC_reg_9_3_inst : DFFR_X1 port map( D => target_PC_i(3), CK => 
                           net199683, RN => n110, Q => predict_PC_9_3_port, QN 
                           => net244775);
   predict_PC_reg_9_2_inst : DFFR_X1 port map( D => target_PC_i(2), CK => 
                           net199683, RN => n107, Q => predict_PC_9_2_port, QN 
                           => net244774);
   predict_PC_reg_9_1_inst : DFFR_X1 port map( D => target_PC_i(1), CK => 
                           net199683, RN => n108, Q => predict_PC_9_1_port, QN 
                           => net244773);
   predict_PC_reg_9_0_inst : DFFR_X1 port map( D => target_PC_i(0), CK => 
                           net199683, RN => n109, Q => predict_PC_9_0_port, QN 
                           => net244772);
   predict_PC_reg_10_31_inst : DFFR_X1 port map( D => target_PC_i(31), CK => 
                           net199688, RN => n105, Q => predict_PC_10_31_port, 
                           QN => net244771);
   predict_PC_reg_10_30_inst : DFFR_X1 port map( D => target_PC_i(30), CK => 
                           net199688, RN => n100, Q => predict_PC_10_30_port, 
                           QN => net244770);
   predict_PC_reg_10_29_inst : DFFR_X1 port map( D => target_PC_i(29), CK => 
                           net199688, RN => n104, Q => predict_PC_10_29_port, 
                           QN => net244769);
   predict_PC_reg_10_28_inst : DFFR_X1 port map( D => target_PC_i(28), CK => 
                           net199688, RN => n102, Q => predict_PC_10_28_port, 
                           QN => net244768);
   predict_PC_reg_10_27_inst : DFFR_X1 port map( D => target_PC_i(27), CK => 
                           net199688, RN => n106, Q => predict_PC_10_27_port, 
                           QN => net244767);
   predict_PC_reg_10_26_inst : DFFR_X1 port map( D => target_PC_i(26), CK => 
                           net199688, RN => n106, Q => predict_PC_10_26_port, 
                           QN => net244766);
   predict_PC_reg_10_25_inst : DFFR_X1 port map( D => target_PC_i(25), CK => 
                           net199688, RN => n101, Q => predict_PC_10_25_port, 
                           QN => net244765);
   predict_PC_reg_10_24_inst : DFFR_X1 port map( D => target_PC_i(24), CK => 
                           net199688, RN => n112, Q => predict_PC_10_24_port, 
                           QN => net244764);
   predict_PC_reg_10_23_inst : DFFR_X1 port map( D => target_PC_i(23), CK => 
                           net199688, RN => n110, Q => predict_PC_10_23_port, 
                           QN => net244763);
   predict_PC_reg_10_22_inst : DFFR_X1 port map( D => target_PC_i(22), CK => 
                           net199688, RN => n107, Q => predict_PC_10_22_port, 
                           QN => net244762);
   predict_PC_reg_10_21_inst : DFFR_X1 port map( D => target_PC_i(21), CK => 
                           net199688, RN => n108, Q => predict_PC_10_21_port, 
                           QN => net244761);
   predict_PC_reg_10_20_inst : DFFR_X1 port map( D => target_PC_i(20), CK => 
                           net199688, RN => n109, Q => predict_PC_10_20_port, 
                           QN => net244760);
   predict_PC_reg_10_19_inst : DFFR_X1 port map( D => target_PC_i(19), CK => 
                           net199688, RN => n105, Q => predict_PC_10_19_port, 
                           QN => net244759);
   predict_PC_reg_10_18_inst : DFFR_X1 port map( D => target_PC_i(18), CK => 
                           net199688, RN => n100, Q => predict_PC_10_18_port, 
                           QN => net244758);
   predict_PC_reg_10_17_inst : DFFR_X1 port map( D => target_PC_i(17), CK => 
                           net199688, RN => n104, Q => predict_PC_10_17_port, 
                           QN => net244757);
   predict_PC_reg_10_16_inst : DFFR_X1 port map( D => target_PC_i(16), CK => 
                           net199688, RN => n102, Q => predict_PC_10_16_port, 
                           QN => net244756);
   predict_PC_reg_10_15_inst : DFFR_X1 port map( D => target_PC_i(15), CK => 
                           net199688, RN => n112, Q => predict_PC_10_15_port, 
                           QN => net244755);
   predict_PC_reg_10_14_inst : DFFR_X1 port map( D => target_PC_i(14), CK => 
                           net199688, RN => n97, Q => predict_PC_10_14_port, QN
                           => net244754);
   predict_PC_reg_10_13_inst : DFFR_X1 port map( D => target_PC_i(13), CK => 
                           net199688, RN => n111, Q => predict_PC_10_13_port, 
                           QN => net244753);
   predict_PC_reg_10_12_inst : DFFR_X1 port map( D => target_PC_i(12), CK => 
                           net199688, RN => n106, Q => predict_PC_10_12_port, 
                           QN => net244752);
   predict_PC_reg_10_11_inst : DFFR_X1 port map( D => target_PC_i(11), CK => 
                           net199688, RN => n101, Q => predict_PC_10_11_port, 
                           QN => net244751);
   predict_PC_reg_10_10_inst : DFFR_X1 port map( D => target_PC_i(10), CK => 
                           net199688, RN => n96, Q => predict_PC_10_10_port, QN
                           => net244750);
   predict_PC_reg_10_9_inst : DFFR_X1 port map( D => target_PC_i(9), CK => 
                           net199688, RN => n112, Q => predict_PC_10_9_port, QN
                           => net244749);
   predict_PC_reg_10_8_inst : DFFR_X1 port map( D => target_PC_i(8), CK => 
                           net199688, RN => n110, Q => predict_PC_10_8_port, QN
                           => net244748);
   predict_PC_reg_10_7_inst : DFFR_X1 port map( D => target_PC_i(7), CK => 
                           net199688, RN => n107, Q => predict_PC_10_7_port, QN
                           => net244747);
   predict_PC_reg_10_6_inst : DFFR_X1 port map( D => target_PC_i(6), CK => 
                           net199688, RN => n108, Q => predict_PC_10_6_port, QN
                           => net244746);
   predict_PC_reg_10_5_inst : DFFR_X1 port map( D => target_PC_i(5), CK => 
                           net199688, RN => n106, Q => predict_PC_10_5_port, QN
                           => net244745);
   predict_PC_reg_10_4_inst : DFFR_X1 port map( D => target_PC_i(4), CK => 
                           net199688, RN => n101, Q => predict_PC_10_4_port, QN
                           => net244744);
   predict_PC_reg_10_3_inst : DFFR_X1 port map( D => target_PC_i(3), CK => 
                           net199688, RN => n110, Q => predict_PC_10_3_port, QN
                           => net244743);
   predict_PC_reg_10_2_inst : DFFR_X1 port map( D => target_PC_i(2), CK => 
                           net199688, RN => n107, Q => predict_PC_10_2_port, QN
                           => net244742);
   predict_PC_reg_10_1_inst : DFFR_X1 port map( D => target_PC_i(1), CK => 
                           net199688, RN => n107, Q => predict_PC_10_1_port, QN
                           => net244741);
   predict_PC_reg_10_0_inst : DFFR_X1 port map( D => target_PC_i(0), CK => 
                           net199688, RN => n108, Q => predict_PC_10_0_port, QN
                           => net244740);
   predict_PC_reg_11_31_inst : DFFR_X1 port map( D => target_PC_i(31), CK => 
                           net199693, RN => n109, Q => predict_PC_11_31_port, 
                           QN => net244739);
   predict_PC_reg_11_30_inst : DFFR_X1 port map( D => target_PC_i(30), CK => 
                           net199693, RN => n105, Q => predict_PC_11_30_port, 
                           QN => net244738);
   predict_PC_reg_11_29_inst : DFFR_X1 port map( D => target_PC_i(29), CK => 
                           net199693, RN => n100, Q => predict_PC_11_29_port, 
                           QN => net244737);
   predict_PC_reg_11_28_inst : DFFR_X1 port map( D => target_PC_i(28), CK => 
                           net199693, RN => n94, Q => predict_PC_11_28_port, QN
                           => net244736);
   predict_PC_reg_11_27_inst : DFFR_X1 port map( D => target_PC_i(27), CK => 
                           net199693, RN => n104, Q => predict_PC_11_27_port, 
                           QN => net244735);
   predict_PC_reg_11_26_inst : DFFR_X1 port map( D => target_PC_i(26), CK => 
                           net199693, RN => n95, Q => predict_PC_11_26_port, QN
                           => net244734);
   predict_PC_reg_11_25_inst : DFFR_X1 port map( D => target_PC_i(25), CK => 
                           net199693, RN => n101, Q => predict_PC_11_25_port, 
                           QN => net244733);
   predict_PC_reg_11_24_inst : DFFR_X1 port map( D => target_PC_i(24), CK => 
                           net199693, RN => n106, Q => predict_PC_11_24_port, 
                           QN => net244732);
   predict_PC_reg_11_23_inst : DFFR_X1 port map( D => target_PC_i(23), CK => 
                           net199693, RN => n101, Q => predict_PC_11_23_port, 
                           QN => net244731);
   predict_PC_reg_11_22_inst : DFFR_X1 port map( D => target_PC_i(22), CK => 
                           net199693, RN => n110, Q => predict_PC_11_22_port, 
                           QN => net244730);
   predict_PC_reg_11_21_inst : DFFR_X1 port map( D => target_PC_i(21), CK => 
                           net199693, RN => n107, Q => predict_PC_11_21_port, 
                           QN => net244729);
   predict_PC_reg_11_20_inst : DFFR_X1 port map( D => target_PC_i(20), CK => 
                           net199693, RN => n93, Q => predict_PC_11_20_port, QN
                           => net244728);
   predict_PC_reg_11_19_inst : DFFR_X1 port map( D => target_PC_i(19), CK => 
                           net199693, RN => n93, Q => predict_PC_11_19_port, QN
                           => net244727);
   predict_PC_reg_11_18_inst : DFFR_X1 port map( D => target_PC_i(18), CK => 
                           net199693, RN => n109, Q => predict_PC_11_18_port, 
                           QN => net244726);
   predict_PC_reg_11_17_inst : DFFR_X1 port map( D => target_PC_i(17), CK => 
                           net199693, RN => n105, Q => predict_PC_11_17_port, 
                           QN => net244725);
   predict_PC_reg_11_16_inst : DFFR_X1 port map( D => target_PC_i(16), CK => 
                           net199693, RN => n100, Q => predict_PC_11_16_port, 
                           QN => net244724);
   predict_PC_reg_11_15_inst : DFFR_X1 port map( D => target_PC_i(15), CK => 
                           net199693, RN => n94, Q => predict_PC_11_15_port, QN
                           => net244723);
   predict_PC_reg_11_14_inst : DFFR_X1 port map( D => target_PC_i(14), CK => 
                           net199693, RN => n104, Q => predict_PC_11_14_port, 
                           QN => net244722);
   predict_PC_reg_11_13_inst : DFFR_X1 port map( D => target_PC_i(13), CK => 
                           net199693, RN => n112, Q => predict_PC_11_13_port, 
                           QN => net244721);
   predict_PC_reg_11_12_inst : DFFR_X1 port map( D => target_PC_i(12), CK => 
                           net199693, RN => n112, Q => predict_PC_11_12_port, 
                           QN => net244720);
   predict_PC_reg_11_11_inst : DFFR_X1 port map( D => target_PC_i(11), CK => 
                           net199693, RN => n112, Q => predict_PC_11_11_port, 
                           QN => net244719);
   predict_PC_reg_11_10_inst : DFFR_X1 port map( D => target_PC_i(10), CK => 
                           net199693, RN => n112, Q => predict_PC_11_10_port, 
                           QN => net244718);
   predict_PC_reg_11_9_inst : DFFR_X1 port map( D => target_PC_i(9), CK => 
                           net199693, RN => n112, Q => predict_PC_11_9_port, QN
                           => net244717);
   predict_PC_reg_11_8_inst : DFFR_X1 port map( D => target_PC_i(8), CK => 
                           net199693, RN => n112, Q => predict_PC_11_8_port, QN
                           => net244716);
   predict_PC_reg_11_7_inst : DFFR_X1 port map( D => target_PC_i(7), CK => 
                           net199693, RN => n112, Q => predict_PC_11_7_port, QN
                           => net244715);
   predict_PC_reg_11_6_inst : DFFR_X1 port map( D => target_PC_i(6), CK => 
                           net199693, RN => n112, Q => predict_PC_11_6_port, QN
                           => net244714);
   predict_PC_reg_11_5_inst : DFFR_X1 port map( D => target_PC_i(5), CK => 
                           net199693, RN => n108, Q => predict_PC_11_5_port, QN
                           => net244713);
   predict_PC_reg_11_4_inst : DFFR_X1 port map( D => target_PC_i(4), CK => 
                           net199693, RN => n112, Q => predict_PC_11_4_port, QN
                           => net244712);
   predict_PC_reg_11_3_inst : DFFR_X1 port map( D => target_PC_i(3), CK => 
                           net199693, RN => n112, Q => predict_PC_11_3_port, QN
                           => net244711);
   predict_PC_reg_11_2_inst : DFFR_X1 port map( D => target_PC_i(2), CK => 
                           net199693, RN => n112, Q => predict_PC_11_2_port, QN
                           => net244710);
   predict_PC_reg_11_1_inst : DFFR_X1 port map( D => target_PC_i(1), CK => 
                           net199693, RN => n113, Q => predict_PC_11_1_port, QN
                           => net244709);
   predict_PC_reg_11_0_inst : DFFR_X1 port map( D => target_PC_i(0), CK => 
                           net199693, RN => n113, Q => predict_PC_11_0_port, QN
                           => net244708);
   predict_PC_reg_12_31_inst : DFFR_X1 port map( D => target_PC_i(31), CK => 
                           net199698, RN => n113, Q => predict_PC_12_31_port, 
                           QN => net244707);
   predict_PC_reg_12_30_inst : DFFR_X1 port map( D => target_PC_i(30), CK => 
                           net199698, RN => n113, Q => predict_PC_12_30_port, 
                           QN => net244706);
   predict_PC_reg_12_29_inst : DFFR_X1 port map( D => target_PC_i(29), CK => 
                           net199698, RN => n113, Q => predict_PC_12_29_port, 
                           QN => net244705);
   predict_PC_reg_12_28_inst : DFFR_X1 port map( D => target_PC_i(28), CK => 
                           net199698, RN => n113, Q => predict_PC_12_28_port, 
                           QN => net244704);
   predict_PC_reg_12_27_inst : DFFR_X1 port map( D => target_PC_i(27), CK => 
                           net199698, RN => n113, Q => predict_PC_12_27_port, 
                           QN => net244703);
   predict_PC_reg_12_26_inst : DFFR_X1 port map( D => target_PC_i(26), CK => 
                           net199698, RN => n113, Q => predict_PC_12_26_port, 
                           QN => net244702);
   predict_PC_reg_12_25_inst : DFFR_X1 port map( D => target_PC_i(25), CK => 
                           net199698, RN => n113, Q => predict_PC_12_25_port, 
                           QN => net244701);
   predict_PC_reg_12_24_inst : DFFR_X1 port map( D => target_PC_i(24), CK => 
                           net199698, RN => n113, Q => predict_PC_12_24_port, 
                           QN => net244700);
   predict_PC_reg_12_23_inst : DFFR_X1 port map( D => target_PC_i(23), CK => 
                           net199698, RN => n112, Q => predict_PC_12_23_port, 
                           QN => net244699);
   predict_PC_reg_12_22_inst : DFFR_X1 port map( D => target_PC_i(22), CK => 
                           net199698, RN => n113, Q => predict_PC_12_22_port, 
                           QN => net244698);
   predict_PC_reg_12_21_inst : DFFR_X1 port map( D => target_PC_i(21), CK => 
                           net199698, RN => n92, Q => predict_PC_12_21_port, QN
                           => net244697);
   predict_PC_reg_12_20_inst : DFFR_X1 port map( D => target_PC_i(20), CK => 
                           net199698, RN => n92, Q => predict_PC_12_20_port, QN
                           => net244696);
   predict_PC_reg_12_19_inst : DFFR_X1 port map( D => target_PC_i(19), CK => 
                           net199698, RN => n91, Q => predict_PC_12_19_port, QN
                           => net244695);
   predict_PC_reg_12_18_inst : DFFR_X1 port map( D => target_PC_i(18), CK => 
                           net199698, RN => n91, Q => predict_PC_12_18_port, QN
                           => net244694);
   predict_PC_reg_12_17_inst : DFFR_X1 port map( D => target_PC_i(17), CK => 
                           net199698, RN => n92, Q => predict_PC_12_17_port, QN
                           => net244693);
   predict_PC_reg_12_16_inst : DFFR_X1 port map( D => target_PC_i(16), CK => 
                           net199698, RN => n90, Q => predict_PC_12_16_port, QN
                           => net244692);
   predict_PC_reg_12_15_inst : DFFR_X1 port map( D => target_PC_i(15), CK => 
                           net199698, RN => n90, Q => predict_PC_12_15_port, QN
                           => net244691);
   predict_PC_reg_12_14_inst : DFFR_X1 port map( D => target_PC_i(14), CK => 
                           net199698, RN => n90, Q => predict_PC_12_14_port, QN
                           => net244690);
   predict_PC_reg_12_13_inst : DFFR_X1 port map( D => target_PC_i(13), CK => 
                           net199698, RN => n91, Q => predict_PC_12_13_port, QN
                           => net244689);
   predict_PC_reg_12_12_inst : DFFR_X1 port map( D => target_PC_i(12), CK => 
                           net199698, RN => n92, Q => predict_PC_12_12_port, QN
                           => net244688);
   predict_PC_reg_12_11_inst : DFFR_X1 port map( D => target_PC_i(11), CK => 
                           net199698, RN => n113, Q => predict_PC_12_11_port, 
                           QN => net244687);
   predict_PC_reg_12_10_inst : DFFR_X1 port map( D => target_PC_i(10), CK => 
                           net199698, RN => n106, Q => predict_PC_12_10_port, 
                           QN => net244686);
   predict_PC_reg_12_9_inst : DFFR_X1 port map( D => target_PC_i(9), CK => 
                           net199698, RN => n105, Q => predict_PC_12_9_port, QN
                           => net244685);
   predict_PC_reg_12_8_inst : DFFR_X1 port map( D => target_PC_i(8), CK => 
                           net199698, RN => n104, Q => predict_PC_12_8_port, QN
                           => net244684);
   predict_PC_reg_12_7_inst : DFFR_X1 port map( D => target_PC_i(7), CK => 
                           net199698, RN => n102, Q => predict_PC_12_7_port, QN
                           => net244683);
   predict_PC_reg_12_6_inst : DFFR_X1 port map( D => target_PC_i(6), CK => 
                           net199698, RN => n111, Q => predict_PC_12_6_port, QN
                           => net244682);
   predict_PC_reg_12_5_inst : DFFR_X1 port map( D => target_PC_i(5), CK => 
                           net199698, RN => n98, Q => predict_PC_12_5_port, QN 
                           => net244681);
   predict_PC_reg_12_4_inst : DFFR_X1 port map( D => target_PC_i(4), CK => 
                           net199698, RN => n98, Q => predict_PC_12_4_port, QN 
                           => net244680);
   predict_PC_reg_12_3_inst : DFFR_X1 port map( D => target_PC_i(3), CK => 
                           net199698, RN => n101, Q => predict_PC_12_3_port, QN
                           => net244679);
   predict_PC_reg_12_2_inst : DFFR_X1 port map( D => target_PC_i(2), CK => 
                           net199698, RN => n101, Q => predict_PC_12_2_port, QN
                           => net244678);
   predict_PC_reg_12_1_inst : DFFR_X1 port map( D => target_PC_i(1), CK => 
                           net199698, RN => n101, Q => predict_PC_12_1_port, QN
                           => net244677);
   predict_PC_reg_12_0_inst : DFFR_X1 port map( D => target_PC_i(0), CK => 
                           net199698, RN => n101, Q => predict_PC_12_0_port, QN
                           => net244676);
   predict_PC_reg_13_31_inst : DFFR_X1 port map( D => target_PC_i(31), CK => 
                           net199703, RN => n101, Q => predict_PC_13_31_port, 
                           QN => net244675);
   predict_PC_reg_13_30_inst : DFFR_X1 port map( D => target_PC_i(30), CK => 
                           net199703, RN => n101, Q => predict_PC_13_30_port, 
                           QN => net244674);
   predict_PC_reg_13_29_inst : DFFR_X1 port map( D => target_PC_i(29), CK => 
                           net199703, RN => n101, Q => predict_PC_13_29_port, 
                           QN => net244673);
   predict_PC_reg_13_28_inst : DFFR_X1 port map( D => target_PC_i(28), CK => 
                           net199703, RN => n101, Q => predict_PC_13_28_port, 
                           QN => net244672);
   predict_PC_reg_13_27_inst : DFFR_X1 port map( D => target_PC_i(27), CK => 
                           net199703, RN => n101, Q => predict_PC_13_27_port, 
                           QN => net244671);
   predict_PC_reg_13_26_inst : DFFR_X1 port map( D => target_PC_i(26), CK => 
                           net199703, RN => n101, Q => predict_PC_13_26_port, 
                           QN => net244670);
   predict_PC_reg_13_25_inst : DFFR_X1 port map( D => target_PC_i(25), CK => 
                           net199703, RN => n101, Q => predict_PC_13_25_port, 
                           QN => net244669);
   predict_PC_reg_13_24_inst : DFFR_X1 port map( D => target_PC_i(24), CK => 
                           net199703, RN => n101, Q => predict_PC_13_24_port, 
                           QN => net244668);
   predict_PC_reg_13_23_inst : DFFR_X1 port map( D => target_PC_i(23), CK => 
                           net199703, RN => n102, Q => predict_PC_13_23_port, 
                           QN => net244667);
   predict_PC_reg_13_22_inst : DFFR_X1 port map( D => target_PC_i(22), CK => 
                           net199703, RN => n102, Q => predict_PC_13_22_port, 
                           QN => net244666);
   predict_PC_reg_13_21_inst : DFFR_X1 port map( D => target_PC_i(21), CK => 
                           net199703, RN => n102, Q => predict_PC_13_21_port, 
                           QN => net244665);
   predict_PC_reg_13_20_inst : DFFR_X1 port map( D => target_PC_i(20), CK => 
                           net199703, RN => n102, Q => predict_PC_13_20_port, 
                           QN => net244664);
   predict_PC_reg_13_19_inst : DFFR_X1 port map( D => target_PC_i(19), CK => 
                           net199703, RN => n102, Q => predict_PC_13_19_port, 
                           QN => net244663);
   predict_PC_reg_13_18_inst : DFFR_X1 port map( D => target_PC_i(18), CK => 
                           net199703, RN => n102, Q => predict_PC_13_18_port, 
                           QN => net244662);
   predict_PC_reg_13_17_inst : DFFR_X1 port map( D => target_PC_i(17), CK => 
                           net199703, RN => n102, Q => predict_PC_13_17_port, 
                           QN => net244661);
   predict_PC_reg_13_16_inst : DFFR_X1 port map( D => target_PC_i(16), CK => 
                           net199703, RN => n102, Q => predict_PC_13_16_port, 
                           QN => net244660);
   predict_PC_reg_13_15_inst : DFFR_X1 port map( D => target_PC_i(15), CK => 
                           net199703, RN => n102, Q => predict_PC_13_15_port, 
                           QN => net244659);
   predict_PC_reg_13_14_inst : DFFR_X1 port map( D => target_PC_i(14), CK => 
                           net199703, RN => n102, Q => predict_PC_13_14_port, 
                           QN => net244658);
   predict_PC_reg_13_13_inst : DFFR_X1 port map( D => target_PC_i(13), CK => 
                           net199703, RN => n102, Q => predict_PC_13_13_port, 
                           QN => net244657);
   predict_PC_reg_13_12_inst : DFFR_X1 port map( D => target_PC_i(12), CK => 
                           net199703, RN => n102, Q => predict_PC_13_12_port, 
                           QN => net244656);
   predict_PC_reg_13_11_inst : DFFR_X1 port map( D => target_PC_i(11), CK => 
                           net199703, RN => n103, Q => predict_PC_13_11_port, 
                           QN => net244655);
   predict_PC_reg_13_10_inst : DFFR_X1 port map( D => target_PC_i(10), CK => 
                           net199703, RN => n103, Q => predict_PC_13_10_port, 
                           QN => net244654);
   predict_PC_reg_13_9_inst : DFFR_X1 port map( D => target_PC_i(9), CK => 
                           net199703, RN => n103, Q => predict_PC_13_9_port, QN
                           => net244653);
   predict_PC_reg_13_8_inst : DFFR_X1 port map( D => target_PC_i(8), CK => 
                           net199703, RN => n103, Q => predict_PC_13_8_port, QN
                           => net244652);
   predict_PC_reg_13_7_inst : DFFR_X1 port map( D => target_PC_i(7), CK => 
                           net199703, RN => n103, Q => predict_PC_13_7_port, QN
                           => net244651);
   predict_PC_reg_13_6_inst : DFFR_X1 port map( D => target_PC_i(6), CK => 
                           net199703, RN => n103, Q => predict_PC_13_6_port, QN
                           => net244650);
   predict_PC_reg_13_5_inst : DFFR_X1 port map( D => target_PC_i(5), CK => 
                           net199703, RN => n103, Q => predict_PC_13_5_port, QN
                           => net244649);
   predict_PC_reg_13_4_inst : DFFR_X1 port map( D => target_PC_i(4), CK => 
                           net199703, RN => n103, Q => predict_PC_13_4_port, QN
                           => net244648);
   predict_PC_reg_13_3_inst : DFFR_X1 port map( D => target_PC_i(3), CK => 
                           net199703, RN => n103, Q => predict_PC_13_3_port, QN
                           => net244647);
   predict_PC_reg_13_2_inst : DFFR_X1 port map( D => target_PC_i(2), CK => 
                           net199703, RN => n103, Q => predict_PC_13_2_port, QN
                           => net244646);
   predict_PC_reg_13_1_inst : DFFR_X1 port map( D => target_PC_i(1), CK => 
                           net199703, RN => n103, Q => predict_PC_13_1_port, QN
                           => net244645);
   predict_PC_reg_13_0_inst : DFFR_X1 port map( D => target_PC_i(0), CK => 
                           net199703, RN => n103, Q => predict_PC_13_0_port, QN
                           => net244644);
   predict_PC_reg_14_31_inst : DFFR_X1 port map( D => target_PC_i(31), CK => 
                           net199708, RN => n104, Q => predict_PC_14_31_port, 
                           QN => net244643);
   predict_PC_reg_14_30_inst : DFFR_X1 port map( D => target_PC_i(30), CK => 
                           net199708, RN => n104, Q => predict_PC_14_30_port, 
                           QN => net244642);
   predict_PC_reg_14_29_inst : DFFR_X1 port map( D => target_PC_i(29), CK => 
                           net199708, RN => n104, Q => predict_PC_14_29_port, 
                           QN => net244641);
   predict_PC_reg_14_28_inst : DFFR_X1 port map( D => target_PC_i(28), CK => 
                           net199708, RN => n104, Q => predict_PC_14_28_port, 
                           QN => net244640);
   predict_PC_reg_14_27_inst : DFFR_X1 port map( D => target_PC_i(27), CK => 
                           net199708, RN => n104, Q => predict_PC_14_27_port, 
                           QN => net244639);
   predict_PC_reg_14_26_inst : DFFR_X1 port map( D => target_PC_i(26), CK => 
                           net199708, RN => n104, Q => predict_PC_14_26_port, 
                           QN => net244638);
   predict_PC_reg_14_25_inst : DFFR_X1 port map( D => target_PC_i(25), CK => 
                           net199708, RN => n104, Q => predict_PC_14_25_port, 
                           QN => net244637);
   predict_PC_reg_14_24_inst : DFFR_X1 port map( D => target_PC_i(24), CK => 
                           net199708, RN => n104, Q => predict_PC_14_24_port, 
                           QN => net244636);
   predict_PC_reg_14_23_inst : DFFR_X1 port map( D => target_PC_i(23), CK => 
                           net199708, RN => n104, Q => predict_PC_14_23_port, 
                           QN => net244635);
   predict_PC_reg_14_22_inst : DFFR_X1 port map( D => target_PC_i(22), CK => 
                           net199708, RN => n104, Q => predict_PC_14_22_port, 
                           QN => net244634);
   predict_PC_reg_14_21_inst : DFFR_X1 port map( D => target_PC_i(21), CK => 
                           net199708, RN => n104, Q => predict_PC_14_21_port, 
                           QN => net244633);
   predict_PC_reg_14_20_inst : DFFR_X1 port map( D => target_PC_i(20), CK => 
                           net199708, RN => n104, Q => predict_PC_14_20_port, 
                           QN => net244632);
   predict_PC_reg_14_19_inst : DFFR_X1 port map( D => target_PC_i(19), CK => 
                           net199708, RN => n105, Q => predict_PC_14_19_port, 
                           QN => net244631);
   predict_PC_reg_14_18_inst : DFFR_X1 port map( D => target_PC_i(18), CK => 
                           net199708, RN => n105, Q => predict_PC_14_18_port, 
                           QN => net244630);
   predict_PC_reg_14_17_inst : DFFR_X1 port map( D => target_PC_i(17), CK => 
                           net199708, RN => n105, Q => predict_PC_14_17_port, 
                           QN => net244629);
   predict_PC_reg_14_16_inst : DFFR_X1 port map( D => target_PC_i(16), CK => 
                           net199708, RN => n105, Q => predict_PC_14_16_port, 
                           QN => net244628);
   predict_PC_reg_14_15_inst : DFFR_X1 port map( D => target_PC_i(15), CK => 
                           net199708, RN => n105, Q => predict_PC_14_15_port, 
                           QN => net244627);
   predict_PC_reg_14_14_inst : DFFR_X1 port map( D => target_PC_i(14), CK => 
                           net199708, RN => n105, Q => predict_PC_14_14_port, 
                           QN => net244626);
   predict_PC_reg_14_13_inst : DFFR_X1 port map( D => target_PC_i(13), CK => 
                           net199708, RN => n105, Q => predict_PC_14_13_port, 
                           QN => net244625);
   predict_PC_reg_14_12_inst : DFFR_X1 port map( D => target_PC_i(12), CK => 
                           net199708, RN => n105, Q => predict_PC_14_12_port, 
                           QN => net244624);
   predict_PC_reg_14_11_inst : DFFR_X1 port map( D => target_PC_i(11), CK => 
                           net199708, RN => n105, Q => predict_PC_14_11_port, 
                           QN => net244623);
   predict_PC_reg_14_10_inst : DFFR_X1 port map( D => target_PC_i(10), CK => 
                           net199708, RN => n105, Q => predict_PC_14_10_port, 
                           QN => net244622);
   predict_PC_reg_14_9_inst : DFFR_X1 port map( D => target_PC_i(9), CK => 
                           net199708, RN => n105, Q => predict_PC_14_9_port, QN
                           => net244621);
   predict_PC_reg_14_8_inst : DFFR_X1 port map( D => target_PC_i(8), CK => 
                           net199708, RN => n105, Q => predict_PC_14_8_port, QN
                           => net244620);
   predict_PC_reg_14_7_inst : DFFR_X1 port map( D => target_PC_i(7), CK => 
                           net199708, RN => n106, Q => predict_PC_14_7_port, QN
                           => net244619);
   predict_PC_reg_14_6_inst : DFFR_X1 port map( D => target_PC_i(6), CK => 
                           net199708, RN => n106, Q => predict_PC_14_6_port, QN
                           => net244618);
   predict_PC_reg_14_5_inst : DFFR_X1 port map( D => target_PC_i(5), CK => 
                           net199708, RN => n106, Q => predict_PC_14_5_port, QN
                           => net244617);
   predict_PC_reg_14_4_inst : DFFR_X1 port map( D => target_PC_i(4), CK => 
                           net199708, RN => n106, Q => predict_PC_14_4_port, QN
                           => net244616);
   predict_PC_reg_14_3_inst : DFFR_X1 port map( D => target_PC_i(3), CK => 
                           net199708, RN => n111, Q => predict_PC_14_3_port, QN
                           => net244615);
   predict_PC_reg_14_2_inst : DFFR_X1 port map( D => target_PC_i(2), CK => 
                           net199708, RN => n106, Q => predict_PC_14_2_port, QN
                           => net244614);
   predict_PC_reg_14_1_inst : DFFR_X1 port map( D => target_PC_i(1), CK => 
                           net199708, RN => n106, Q => predict_PC_14_1_port, QN
                           => net244613);
   predict_PC_reg_14_0_inst : DFFR_X1 port map( D => target_PC_i(0), CK => 
                           net199708, RN => n106, Q => predict_PC_14_0_port, QN
                           => net244612);
   predict_PC_reg_15_31_inst : DFFR_X1 port map( D => target_PC_i(31), CK => 
                           net199713, RN => n106, Q => predict_PC_15_31_port, 
                           QN => net244611);
   last_PC_reg_31_inst : DFFR_X1 port map( D => predicted_next_PC_o_31_port, CK
                           => net199633, RN => n106, Q => net244610, QN => n483
                           );
   predict_PC_reg_15_30_inst : DFFR_X1 port map( D => target_PC_i(30), CK => 
                           net199713, RN => n106, Q => predict_PC_15_30_port, 
                           QN => net244609);
   last_PC_reg_30_inst : DFFR_X1 port map( D => predicted_next_PC_o_30_port, CK
                           => net199633, RN => n106, Q => net244608, QN => n485
                           );
   predict_PC_reg_15_29_inst : DFFR_X1 port map( D => target_PC_i(29), CK => 
                           net199713, RN => n107, Q => predict_PC_15_29_port, 
                           QN => net244607);
   last_PC_reg_29_inst : DFFR_X1 port map( D => predicted_next_PC_o_29_port, CK
                           => net199633, RN => n107, Q => net244606, QN => n487
                           );
   predict_PC_reg_15_28_inst : DFFR_X1 port map( D => target_PC_i(28), CK => 
                           net199713, RN => n107, Q => predict_PC_15_28_port, 
                           QN => net244605);
   last_PC_reg_28_inst : DFFR_X1 port map( D => predicted_next_PC_o_28_port, CK
                           => net199633, RN => n107, Q => net244604, QN => n489
                           );
   predict_PC_reg_15_27_inst : DFFR_X1 port map( D => target_PC_i(27), CK => 
                           net199713, RN => n107, Q => predict_PC_15_27_port, 
                           QN => net244603);
   last_PC_reg_27_inst : DFFR_X1 port map( D => predicted_next_PC_o_27_port, CK
                           => net199633, RN => n107, Q => net244602, QN => n491
                           );
   predict_PC_reg_15_26_inst : DFFR_X1 port map( D => target_PC_i(26), CK => 
                           net199713, RN => n107, Q => predict_PC_15_26_port, 
                           QN => net244601);
   last_PC_reg_26_inst : DFFR_X1 port map( D => predicted_next_PC_o_26_port, CK
                           => net199633, RN => n107, Q => net244600, QN => n493
                           );
   predict_PC_reg_15_25_inst : DFFR_X1 port map( D => target_PC_i(25), CK => 
                           net199713, RN => n107, Q => predict_PC_15_25_port, 
                           QN => net244599);
   last_PC_reg_25_inst : DFFR_X1 port map( D => predicted_next_PC_o_25_port, CK
                           => net199633, RN => n107, Q => net244598, QN => n495
                           );
   predict_PC_reg_15_24_inst : DFFR_X1 port map( D => target_PC_i(24), CK => 
                           net199713, RN => n107, Q => predict_PC_15_24_port, 
                           QN => net244597);
   last_PC_reg_24_inst : DFFR_X1 port map( D => predicted_next_PC_o_24_port, CK
                           => net199633, RN => n107, Q => net244596, QN => n497
                           );
   predict_PC_reg_15_23_inst : DFFR_X1 port map( D => target_PC_i(23), CK => 
                           net199713, RN => n108, Q => predict_PC_15_23_port, 
                           QN => net244595);
   last_PC_reg_23_inst : DFFR_X1 port map( D => predicted_next_PC_o_23_port, CK
                           => net199633, RN => n108, Q => net244594, QN => n499
                           );
   predict_PC_reg_15_22_inst : DFFR_X1 port map( D => target_PC_i(22), CK => 
                           net199713, RN => n108, Q => predict_PC_15_22_port, 
                           QN => net244593);
   last_PC_reg_22_inst : DFFR_X1 port map( D => predicted_next_PC_o_22_port, CK
                           => net199633, RN => n108, Q => net244592, QN => n501
                           );
   predict_PC_reg_15_21_inst : DFFR_X1 port map( D => target_PC_i(21), CK => 
                           net199713, RN => n108, Q => predict_PC_15_21_port, 
                           QN => net244591);
   last_PC_reg_21_inst : DFFR_X1 port map( D => predicted_next_PC_o_21_port, CK
                           => net199633, RN => n108, Q => net244590, QN => n503
                           );
   predict_PC_reg_15_20_inst : DFFR_X1 port map( D => target_PC_i(20), CK => 
                           net199713, RN => n108, Q => predict_PC_15_20_port, 
                           QN => net244589);
   last_PC_reg_20_inst : DFFR_X1 port map( D => predicted_next_PC_o_20_port, CK
                           => net199633, RN => n108, Q => net244588, QN => n505
                           );
   predict_PC_reg_15_19_inst : DFFR_X1 port map( D => target_PC_i(19), CK => 
                           net199713, RN => n108, Q => predict_PC_15_19_port, 
                           QN => net244587);
   last_PC_reg_19_inst : DFFR_X1 port map( D => predicted_next_PC_o_19_port, CK
                           => net199633, RN => n108, Q => net244586, QN => n507
                           );
   predict_PC_reg_15_18_inst : DFFR_X1 port map( D => target_PC_i(18), CK => 
                           net199713, RN => n108, Q => predict_PC_15_18_port, 
                           QN => net244585);
   last_PC_reg_18_inst : DFFR_X1 port map( D => predicted_next_PC_o_18_port, CK
                           => net199633, RN => n108, Q => net244584, QN => n509
                           );
   predict_PC_reg_15_17_inst : DFFR_X1 port map( D => target_PC_i(17), CK => 
                           net199713, RN => n109, Q => predict_PC_15_17_port, 
                           QN => net244583);
   last_PC_reg_17_inst : DFFR_X1 port map( D => predicted_next_PC_o_17_port, CK
                           => net199633, RN => n109, Q => net244582, QN => n511
                           );
   predict_PC_reg_15_16_inst : DFFR_X1 port map( D => target_PC_i(16), CK => 
                           net199713, RN => n109, Q => predict_PC_15_16_port, 
                           QN => net244581);
   last_PC_reg_16_inst : DFFR_X1 port map( D => predicted_next_PC_o_16_port, CK
                           => net199633, RN => n109, Q => net244580, QN => n513
                           );
   predict_PC_reg_15_15_inst : DFFR_X1 port map( D => target_PC_i(15), CK => 
                           net199713, RN => n109, Q => predict_PC_15_15_port, 
                           QN => net244579);
   last_PC_reg_15_inst : DFFR_X1 port map( D => predicted_next_PC_o_15_port, CK
                           => net199633, RN => n109, Q => net244578, QN => n515
                           );
   predict_PC_reg_15_14_inst : DFFR_X1 port map( D => target_PC_i(14), CK => 
                           net199713, RN => n109, Q => predict_PC_15_14_port, 
                           QN => net244577);
   last_PC_reg_14_inst : DFFR_X1 port map( D => predicted_next_PC_o_14_port, CK
                           => net199633, RN => n109, Q => net244576, QN => n517
                           );
   predict_PC_reg_15_13_inst : DFFR_X1 port map( D => target_PC_i(13), CK => 
                           net199713, RN => n109, Q => predict_PC_15_13_port, 
                           QN => net244575);
   last_PC_reg_13_inst : DFFR_X1 port map( D => predicted_next_PC_o_13_port, CK
                           => net199633, RN => n109, Q => net244574, QN => n519
                           );
   predict_PC_reg_15_12_inst : DFFR_X1 port map( D => target_PC_i(12), CK => 
                           net199713, RN => n109, Q => predict_PC_15_12_port, 
                           QN => net244573);
   last_PC_reg_12_inst : DFFR_X1 port map( D => predicted_next_PC_o_12_port, CK
                           => net199633, RN => n109, Q => net244572, QN => n521
                           );
   predict_PC_reg_15_11_inst : DFFR_X1 port map( D => target_PC_i(11), CK => 
                           net199713, RN => n110, Q => predict_PC_15_11_port, 
                           QN => net244571);
   last_PC_reg_11_inst : DFFR_X1 port map( D => predicted_next_PC_o_11_port, CK
                           => net199633, RN => n110, Q => net244570, QN => n523
                           );
   predict_PC_reg_15_10_inst : DFFR_X1 port map( D => target_PC_i(10), CK => 
                           net199713, RN => n110, Q => predict_PC_15_10_port, 
                           QN => net244569);
   last_PC_reg_10_inst : DFFR_X1 port map( D => predicted_next_PC_o_10_port, CK
                           => net199633, RN => n110, Q => net244568, QN => n525
                           );
   predict_PC_reg_15_9_inst : DFFR_X1 port map( D => target_PC_i(9), CK => 
                           net199713, RN => n110, Q => predict_PC_15_9_port, QN
                           => net244567);
   last_PC_reg_9_inst : DFFR_X1 port map( D => predicted_next_PC_o_9_port, CK 
                           => net199633, RN => n110, Q => net244566, QN => n527
                           );
   predict_PC_reg_15_8_inst : DFFR_X1 port map( D => target_PC_i(8), CK => 
                           net199713, RN => n110, Q => predict_PC_15_8_port, QN
                           => net244565);
   last_PC_reg_8_inst : DFFR_X1 port map( D => predicted_next_PC_o_8_port, CK 
                           => net199633, RN => n110, Q => net244564, QN => n529
                           );
   predict_PC_reg_15_7_inst : DFFR_X1 port map( D => target_PC_i(7), CK => 
                           net199713, RN => n110, Q => predict_PC_15_7_port, QN
                           => net244563);
   last_PC_reg_7_inst : DFFR_X1 port map( D => predicted_next_PC_o_7_port, CK 
                           => net199633, RN => n110, Q => net244562, QN => n531
                           );
   predict_PC_reg_15_6_inst : DFFR_X1 port map( D => target_PC_i(6), CK => 
                           net199713, RN => n110, Q => predict_PC_15_6_port, QN
                           => net244561);
   last_PC_reg_6_inst : DFFR_X1 port map( D => predicted_next_PC_o_6_port, CK 
                           => net199633, RN => n110, Q => net244560, QN => n533
                           );
   predict_PC_reg_15_5_inst : DFFR_X1 port map( D => target_PC_i(5), CK => 
                           net199713, RN => n111, Q => predict_PC_15_5_port, QN
                           => net244559);
   last_PC_reg_5_inst : DFFR_X1 port map( D => predicted_next_PC_o_5_port, CK 
                           => net199633, RN => n111, Q => net244558, QN => n535
                           );
   predict_PC_reg_15_4_inst : DFFR_X1 port map( D => target_PC_i(4), CK => 
                           net199713, RN => n111, Q => predict_PC_15_4_port, QN
                           => net244557);
   last_PC_reg_4_inst : DFFR_X1 port map( D => predicted_next_PC_o_4_port, CK 
                           => net199633, RN => n111, Q => net244556, QN => n537
                           );
   predict_PC_reg_15_3_inst : DFFR_X1 port map( D => target_PC_i(3), CK => 
                           net199713, RN => n111, Q => predict_PC_15_3_port, QN
                           => net244555);
   last_PC_reg_3_inst : DFFR_X1 port map( D => predicted_next_PC_o_3_port, CK 
                           => net199633, RN => n111, Q => net244554, QN => n539
                           );
   predict_PC_reg_15_2_inst : DFFR_X1 port map( D => target_PC_i(2), CK => 
                           net199713, RN => n111, Q => predict_PC_15_2_port, QN
                           => net244553);
   last_PC_reg_2_inst : DFFR_X1 port map( D => predicted_next_PC_o_2_port, CK 
                           => net199633, RN => n111, Q => net244552, QN => n541
                           );
   predict_PC_reg_15_1_inst : DFFR_X1 port map( D => target_PC_i(1), CK => 
                           net199713, RN => n111, Q => predict_PC_15_1_port, QN
                           => net244551);
   last_PC_reg_1_inst : DFFR_X1 port map( D => predicted_next_PC_o_1_port, CK 
                           => net199633, RN => n111, Q => net244550, QN => n543
                           );
   predict_PC_reg_15_0_inst : DFFR_X1 port map( D => target_PC_i(0), CK => 
                           net199713, RN => n111, Q => predict_PC_15_0_port, QN
                           => net244549);
   last_PC_reg_0_inst : DFFR_X1 port map( D => predicted_next_PC_o_0_port, CK 
                           => net199633, RN => n111, Q => net244548, QN => n545
                           );
   last_mispredict_reg : DFFR_X1 port map( D => mispredict_o_port, CK => 
                           net199633, RN => n108, Q => net244547, QN => n546);
   pred_x_0 : predictor_2_0 port map( clock => clock, reset => reset, enable =>
                           write_enable_0_port, taken_i => was_taken_i, 
                           prediction_o => taken_0_port);
   pred_x_1 : predictor_2_15 port map( clock => clock, reset => reset, enable 
                           => write_enable_1_port, taken_i => was_taken_i, 
                           prediction_o => taken_1_port);
   pred_x_2 : predictor_2_14 port map( clock => clock, reset => reset, enable 
                           => write_enable_2_port, taken_i => was_taken_i, 
                           prediction_o => taken_2_port);
   pred_x_3 : predictor_2_13 port map( clock => clock, reset => reset, enable 
                           => write_enable_3_port, taken_i => was_taken_i, 
                           prediction_o => taken_3_port);
   pred_x_4 : predictor_2_12 port map( clock => clock, reset => reset, enable 
                           => write_enable_4_port, taken_i => was_taken_i, 
                           prediction_o => taken_4_port);
   pred_x_5 : predictor_2_11 port map( clock => clock, reset => reset, enable 
                           => write_enable_5_port, taken_i => was_taken_i, 
                           prediction_o => taken_5_port);
   pred_x_6 : predictor_2_10 port map( clock => clock, reset => reset, enable 
                           => write_enable_6_port, taken_i => was_taken_i, 
                           prediction_o => taken_6_port);
   pred_x_7 : predictor_2_9 port map( clock => clock, reset => reset, enable =>
                           write_enable_7_port, taken_i => was_taken_i, 
                           prediction_o => taken_7_port);
   pred_x_8 : predictor_2_8 port map( clock => clock, reset => reset, enable =>
                           write_enable_8_port, taken_i => was_taken_i, 
                           prediction_o => taken_8_port);
   pred_x_9 : predictor_2_7 port map( clock => clock, reset => reset, enable =>
                           write_enable_9_port, taken_i => was_taken_i, 
                           prediction_o => taken_9_port);
   pred_x_10 : predictor_2_6 port map( clock => clock, reset => reset, enable 
                           => write_enable_10_port, taken_i => was_taken_i, 
                           prediction_o => taken_10_port);
   pred_x_11 : predictor_2_5 port map( clock => clock, reset => reset, enable 
                           => write_enable_11_port, taken_i => was_taken_i, 
                           prediction_o => taken_11_port);
   pred_x_12 : predictor_2_4 port map( clock => clock, reset => reset, enable 
                           => write_enable_12_port, taken_i => was_taken_i, 
                           prediction_o => taken_12_port);
   pred_x_13 : predictor_2_3 port map( clock => clock, reset => reset, enable 
                           => write_enable_13_port, taken_i => was_taken_i, 
                           prediction_o => taken_13_port);
   pred_x_14 : predictor_2_2 port map( clock => clock, reset => reset, enable 
                           => write_enable_14_port, taken_i => was_taken_i, 
                           prediction_o => taken_14_port);
   pred_x_15 : predictor_2_1 port map( clock => clock, reset => reset, enable 
                           => write_enable_15_port, taken_i => was_taken_i, 
                           prediction_o => taken_15_port);
   clk_gate_last_TAG_reg : SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_0 port map(
                           CLK => clock, EN => N567, ENCLK => net199633);
   clk_gate_predict_PC_reg_0_inst : SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_16
                           port map( CLK => clock, EN => N566, ENCLK => 
                           net199638);
   clk_gate_predict_PC_reg_1_inst : SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_15
                           port map( CLK => clock, EN => N534, ENCLK => 
                           net199643);
   clk_gate_predict_PC_reg_2_inst : SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_14
                           port map( CLK => clock, EN => N502, ENCLK => 
                           net199648);
   clk_gate_predict_PC_reg_3_inst : SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_13
                           port map( CLK => clock, EN => N470, ENCLK => 
                           net199653);
   clk_gate_predict_PC_reg_4_inst : SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_12
                           port map( CLK => clock, EN => N438, ENCLK => 
                           net199658);
   clk_gate_predict_PC_reg_5_inst : SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_11
                           port map( CLK => clock, EN => N406, ENCLK => 
                           net199663);
   clk_gate_predict_PC_reg_6_inst : SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_10
                           port map( CLK => clock, EN => N374, ENCLK => 
                           net199668);
   clk_gate_predict_PC_reg_7_inst : SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_9 
                           port map( CLK => clock, EN => N342, ENCLK => 
                           net199673);
   clk_gate_predict_PC_reg_8_inst : SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_8 
                           port map( CLK => clock, EN => N310, ENCLK => 
                           net199678);
   clk_gate_predict_PC_reg_9_inst : SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_7 
                           port map( CLK => clock, EN => N278, ENCLK => 
                           net199683);
   clk_gate_predict_PC_reg_10_inst : SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_6
                           port map( CLK => clock, EN => N246, ENCLK => 
                           net199688);
   clk_gate_predict_PC_reg_11_inst : SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_5
                           port map( CLK => clock, EN => N214, ENCLK => 
                           net199693);
   clk_gate_predict_PC_reg_12_inst : SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_4
                           port map( CLK => clock, EN => N182, ENCLK => 
                           net199698);
   clk_gate_predict_PC_reg_13_inst : SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_3
                           port map( CLK => clock, EN => N150, ENCLK => 
                           net199703);
   clk_gate_predict_PC_reg_14_inst : SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_2
                           port map( CLK => clock, EN => N118, ENCLK => 
                           net199708);
   clk_gate_predict_PC_reg_15_inst : SNPS_CLOCK_GATE_HIGH_btb_N_LINES4_SIZE32_1
                           port map( CLK => clock, EN => N86, ENCLK => 
                           net199713);
   U391 : NAND2_X1 port map( A1 => TAG_i(1), A2 => n903, ZN => n895);
   U388 : NAND2_X1 port map( A1 => TAG_i(0), A2 => TAG_i(1), ZN => n894);
   U386 : AOI22_X1 port map( A1 => n557, A2 => taken_10_port, B1 => n558, B2 =>
                           taken_11_port, ZN => n897);
   U383 : NAND2_X1 port map( A1 => TAG_i(0), A2 => n974, ZN => n891);
   U381 : AOI22_X1 port map( A1 => n83, A2 => taken_8_port, B1 => n82, B2 => 
                           taken_9_port, ZN => n898);
   U377 : AOI22_X1 port map( A1 => n553, A2 => taken_14_port, B1 => n554, B2 =>
                           taken_15_port, ZN => n899);
   U374 : AOI22_X1 port map( A1 => n87, A2 => taken_12_port, B1 => n86_port, B2
                           => taken_13_port, ZN => n900);
   U369 : AOI22_X1 port map( A1 => n569, A2 => taken_2_port, B1 => n570, B2 => 
                           taken_3_port, ZN => n887);
   U366 : AOI22_X1 port map( A1 => n75, A2 => taken_0_port, B1 => n74, B2 => 
                           taken_1_port, ZN => n888);
   U365 : NAND2_X1 port map( A1 => TAG_i(2), A2 => n972, ZN => n892);
   U362 : AOI22_X1 port map( A1 => n565, A2 => taken_6_port, B1 => n566_port, 
                           B2 => taken_7_port, ZN => n889);
   U359 : AOI22_X1 port map( A1 => n79, A2 => taken_4_port, B1 => n78, B2 => 
                           taken_5_port, ZN => n890);
   U254 : AOI22_X1 port map( A1 => n75, A2 => predict_PC_0_18_port, B1 => n572,
                           B2 => predict_PC_1_18_port, ZN => n789);
   U253 : AOI22_X1 port map( A1 => n77, A2 => predict_PC_2_18_port, B1 => n76, 
                           B2 => predict_PC_3_18_port, ZN => n790);
   U252 : AOI22_X1 port map( A1 => n567_port, A2 => predict_PC_4_18_port, B1 =>
                           n568, B2 => predict_PC_5_18_port, ZN => n791);
   U251 : AOI22_X1 port map( A1 => n81, A2 => predict_PC_6_18_port, B1 => n80, 
                           B2 => predict_PC_7_18_port, ZN => n792);
   U250 : NAND4_X1 port map( A1 => n789, A2 => n790, A3 => n791, A4 => n792, ZN
                           => n783);
   U249 : AOI22_X1 port map( A1 => n559, A2 => predict_PC_8_18_port, B1 => n560
                           , B2 => predict_PC_9_18_port, ZN => n785);
   U248 : AOI22_X1 port map( A1 => n85, A2 => predict_PC_10_18_port, B1 => n84,
                           B2 => predict_PC_11_18_port, ZN => n786);
   U247 : AOI22_X1 port map( A1 => n555, A2 => predict_PC_12_18_port, B1 => 
                           n556, B2 => predict_PC_13_18_port, ZN => n787);
   U246 : AOI22_X1 port map( A1 => n89, A2 => predict_PC_14_18_port, B1 => n88,
                           B2 => predict_PC_15_18_port, ZN => n788);
   U245 : NAND4_X1 port map( A1 => n785, A2 => n786, A3 => n787, A4 => n788, ZN
                           => n784);
   U243 : AOI22_X1 port map( A1 => n75, A2 => predict_PC_0_19_port, B1 => n74, 
                           B2 => predict_PC_1_19_port, ZN => n779);
   U242 : AOI22_X1 port map( A1 => n77, A2 => predict_PC_2_19_port, B1 => n76, 
                           B2 => predict_PC_3_19_port, ZN => n780);
   U241 : AOI22_X1 port map( A1 => n79, A2 => predict_PC_4_19_port, B1 => n568,
                           B2 => predict_PC_5_19_port, ZN => n781);
   U240 : AOI22_X1 port map( A1 => n81, A2 => predict_PC_6_19_port, B1 => n80, 
                           B2 => predict_PC_7_19_port, ZN => n782);
   U239 : NAND4_X1 port map( A1 => n779, A2 => n780, A3 => n781, A4 => n782, ZN
                           => n773);
   U238 : AOI22_X1 port map( A1 => n83, A2 => predict_PC_8_19_port, B1 => n560,
                           B2 => predict_PC_9_19_port, ZN => n775);
   U237 : AOI22_X1 port map( A1 => n85, A2 => predict_PC_10_19_port, B1 => n84,
                           B2 => predict_PC_11_19_port, ZN => n776);
   U236 : AOI22_X1 port map( A1 => n87, A2 => predict_PC_12_19_port, B1 => n556
                           , B2 => predict_PC_13_19_port, ZN => n777);
   U235 : AOI22_X1 port map( A1 => n89, A2 => predict_PC_14_19_port, B1 => n88,
                           B2 => predict_PC_15_19_port, ZN => n778);
   U234 : NAND4_X1 port map( A1 => n775, A2 => n776, A3 => n777, A4 => n778, ZN
                           => n774);
   U45 : AOI22_X1 port map( A1 => n571, A2 => predict_PC_0_6_port, B1 => n572, 
                           B2 => predict_PC_1_6_port, ZN => n599);
   U44 : AOI22_X1 port map( A1 => n77, A2 => predict_PC_2_6_port, B1 => n76, B2
                           => predict_PC_3_6_port, ZN => n600);
   U43 : AOI22_X1 port map( A1 => n567_port, A2 => predict_PC_4_6_port, B1 => 
                           n568, B2 => predict_PC_5_6_port, ZN => n601);
   U42 : AOI22_X1 port map( A1 => n81, A2 => predict_PC_6_6_port, B1 => n80, B2
                           => predict_PC_7_6_port, ZN => n602);
   U41 : NAND4_X1 port map( A1 => n599, A2 => n600, A3 => n601, A4 => n602, ZN 
                           => n593);
   U40 : AOI22_X1 port map( A1 => n559, A2 => predict_PC_8_6_port, B1 => n560, 
                           B2 => predict_PC_9_6_port, ZN => n595);
   U39 : AOI22_X1 port map( A1 => n85, A2 => predict_PC_10_6_port, B1 => n84, 
                           B2 => predict_PC_11_6_port, ZN => n596);
   U38 : AOI22_X1 port map( A1 => n555, A2 => predict_PC_12_6_port, B1 => n556,
                           B2 => predict_PC_13_6_port, ZN => n597);
   U37 : AOI22_X1 port map( A1 => n89, A2 => predict_PC_14_6_port, B1 => n88, 
                           B2 => predict_PC_15_6_port, ZN => n598);
   U36 : NAND4_X1 port map( A1 => n595, A2 => n596, A3 => n597, A4 => n598, ZN 
                           => n594);
   U232 : AOI22_X1 port map( A1 => n571, A2 => predict_PC_0_1_port, B1 => n74, 
                           B2 => predict_PC_1_1_port, ZN => n769);
   U231 : AOI22_X1 port map( A1 => n77, A2 => predict_PC_2_1_port, B1 => n76, 
                           B2 => predict_PC_3_1_port, ZN => n770);
   U230 : AOI22_X1 port map( A1 => n79, A2 => predict_PC_4_1_port, B1 => n568, 
                           B2 => predict_PC_5_1_port, ZN => n771);
   U229 : AOI22_X1 port map( A1 => n81, A2 => predict_PC_6_1_port, B1 => n80, 
                           B2 => predict_PC_7_1_port, ZN => n772);
   U228 : NAND4_X1 port map( A1 => n769, A2 => n770, A3 => n771, A4 => n772, ZN
                           => n763);
   U227 : AOI22_X1 port map( A1 => n83, A2 => predict_PC_8_1_port, B1 => n560, 
                           B2 => predict_PC_9_1_port, ZN => n765);
   U226 : AOI22_X1 port map( A1 => n85, A2 => predict_PC_10_1_port, B1 => n84, 
                           B2 => predict_PC_11_1_port, ZN => n766);
   U225 : AOI22_X1 port map( A1 => n87, A2 => predict_PC_12_1_port, B1 => n556,
                           B2 => predict_PC_13_1_port, ZN => n767);
   U224 : AOI22_X1 port map( A1 => n89, A2 => predict_PC_14_1_port, B1 => n88, 
                           B2 => predict_PC_15_1_port, ZN => n768);
   U223 : NAND4_X1 port map( A1 => n765, A2 => n766, A3 => n767, A4 => n768, ZN
                           => n764);
   U111 : AOI22_X1 port map( A1 => n571, A2 => predict_PC_0_2_port, B1 => n74, 
                           B2 => predict_PC_1_2_port, ZN => n659);
   U110 : AOI22_X1 port map( A1 => n77, A2 => predict_PC_2_2_port, B1 => n76, 
                           B2 => predict_PC_3_2_port, ZN => n660);
   U109 : AOI22_X1 port map( A1 => n79, A2 => predict_PC_4_2_port, B1 => n78, 
                           B2 => predict_PC_5_2_port, ZN => n661);
   U108 : AOI22_X1 port map( A1 => n81, A2 => predict_PC_6_2_port, B1 => n80, 
                           B2 => predict_PC_7_2_port, ZN => n662);
   U107 : NAND4_X1 port map( A1 => n659, A2 => n660, A3 => n661, A4 => n662, ZN
                           => n653);
   U106 : AOI22_X1 port map( A1 => n83, A2 => predict_PC_8_2_port, B1 => n82, 
                           B2 => predict_PC_9_2_port, ZN => n655);
   U105 : AOI22_X1 port map( A1 => n85, A2 => predict_PC_10_2_port, B1 => n84, 
                           B2 => predict_PC_11_2_port, ZN => n656);
   U104 : AOI22_X1 port map( A1 => n87, A2 => predict_PC_12_2_port, B1 => 
                           n86_port, B2 => predict_PC_13_2_port, ZN => n657);
   U103 : AOI22_X1 port map( A1 => n89, A2 => predict_PC_14_2_port, B1 => n88, 
                           B2 => predict_PC_15_2_port, ZN => n658);
   U102 : NAND4_X1 port map( A1 => n655, A2 => n656, A3 => n657, A4 => n658, ZN
                           => n654);
   U23 : AOI22_X1 port map( A1 => n75, A2 => predict_PC_0_8_port, B1 => n572, 
                           B2 => predict_PC_1_8_port, ZN => n579);
   U22 : AOI22_X1 port map( A1 => n77, A2 => predict_PC_2_8_port, B1 => n76, B2
                           => predict_PC_3_8_port, ZN => n580);
   U21 : AOI22_X1 port map( A1 => n567_port, A2 => predict_PC_4_8_port, B1 => 
                           n568, B2 => predict_PC_5_8_port, ZN => n581);
   U20 : AOI22_X1 port map( A1 => n81, A2 => predict_PC_6_8_port, B1 => n80, B2
                           => predict_PC_7_8_port, ZN => n582);
   U19 : NAND4_X1 port map( A1 => n579, A2 => n580, A3 => n581, A4 => n582, ZN 
                           => n573);
   U18 : AOI22_X1 port map( A1 => n559, A2 => predict_PC_8_8_port, B1 => n560, 
                           B2 => predict_PC_9_8_port, ZN => n575);
   U17 : AOI22_X1 port map( A1 => n85, A2 => predict_PC_10_8_port, B1 => n84, 
                           B2 => predict_PC_11_8_port, ZN => n576);
   U16 : AOI22_X1 port map( A1 => n555, A2 => predict_PC_12_8_port, B1 => n556,
                           B2 => predict_PC_13_8_port, ZN => n577);
   U15 : AOI22_X1 port map( A1 => n89, A2 => predict_PC_14_8_port, B1 => n88, 
                           B2 => predict_PC_15_8_port, ZN => n578);
   U14 : NAND4_X1 port map( A1 => n575, A2 => n576, A3 => n577, A4 => n578, ZN 
                           => n574);
   U276 : AOI22_X1 port map( A1 => n75, A2 => predict_PC_0_16_port, B1 => n74, 
                           B2 => predict_PC_1_16_port, ZN => n809);
   U275 : AOI22_X1 port map( A1 => n569, A2 => predict_PC_2_16_port, B1 => n570
                           , B2 => predict_PC_3_16_port, ZN => n810);
   U274 : AOI22_X1 port map( A1 => n79, A2 => predict_PC_4_16_port, B1 => n78, 
                           B2 => predict_PC_5_16_port, ZN => n811);
   U273 : AOI22_X1 port map( A1 => n565, A2 => predict_PC_6_16_port, B1 => 
                           n566_port, B2 => predict_PC_7_16_port, ZN => n812);
   U272 : NAND4_X1 port map( A1 => n809, A2 => n810, A3 => n811, A4 => n812, ZN
                           => n803);
   U271 : AOI22_X1 port map( A1 => n83, A2 => predict_PC_8_16_port, B1 => n82, 
                           B2 => predict_PC_9_16_port, ZN => n805);
   U270 : AOI22_X1 port map( A1 => n557, A2 => predict_PC_10_16_port, B1 => n84
                           , B2 => predict_PC_11_16_port, ZN => n806);
   U269 : AOI22_X1 port map( A1 => n87, A2 => predict_PC_12_16_port, B1 => 
                           n86_port, B2 => predict_PC_13_16_port, ZN => n807);
   U268 : AOI22_X1 port map( A1 => n553, A2 => predict_PC_14_16_port, B1 => 
                           n554, B2 => predict_PC_15_16_port, ZN => n808);
   U267 : NAND4_X1 port map( A1 => n805, A2 => n806, A3 => n807, A4 => n808, ZN
                           => n804);
   U210 : AOI22_X1 port map( A1 => n75, A2 => predict_PC_0_21_port, B1 => n74, 
                           B2 => predict_PC_1_21_port, ZN => n749);
   U209 : AOI22_X1 port map( A1 => n77, A2 => predict_PC_2_21_port, B1 => n76, 
                           B2 => predict_PC_3_21_port, ZN => n750);
   U208 : AOI22_X1 port map( A1 => n79, A2 => predict_PC_4_21_port, B1 => n568,
                           B2 => predict_PC_5_21_port, ZN => n751);
   U207 : AOI22_X1 port map( A1 => n81, A2 => predict_PC_6_21_port, B1 => n80, 
                           B2 => predict_PC_7_21_port, ZN => n752);
   U206 : NAND4_X1 port map( A1 => n749, A2 => n750, A3 => n751, A4 => n752, ZN
                           => n743);
   U205 : AOI22_X1 port map( A1 => n83, A2 => predict_PC_8_21_port, B1 => n560,
                           B2 => predict_PC_9_21_port, ZN => n745);
   U204 : AOI22_X1 port map( A1 => n85, A2 => predict_PC_10_21_port, B1 => n84,
                           B2 => predict_PC_11_21_port, ZN => n746);
   U203 : AOI22_X1 port map( A1 => n87, A2 => predict_PC_12_21_port, B1 => n556
                           , B2 => predict_PC_13_21_port, ZN => n747);
   U202 : AOI22_X1 port map( A1 => n89, A2 => predict_PC_14_21_port, B1 => n88,
                           B2 => predict_PC_15_21_port, ZN => n748);
   U201 : NAND4_X1 port map( A1 => n745, A2 => n746, A3 => n747, A4 => n748, ZN
                           => n744);
   U342 : AOI22_X1 port map( A1 => n75, A2 => predict_PC_0_10_port, B1 => n74, 
                           B2 => predict_PC_1_10_port, ZN => n869);
   U341 : AOI22_X1 port map( A1 => n569, A2 => predict_PC_2_10_port, B1 => n570
                           , B2 => predict_PC_3_10_port, ZN => n870);
   U340 : AOI22_X1 port map( A1 => n79, A2 => predict_PC_4_10_port, B1 => n78, 
                           B2 => predict_PC_5_10_port, ZN => n871);
   U339 : AOI22_X1 port map( A1 => n565, A2 => predict_PC_6_10_port, B1 => 
                           n566_port, B2 => predict_PC_7_10_port, ZN => n872);
   U338 : NAND4_X1 port map( A1 => n869, A2 => n870, A3 => n871, A4 => n872, ZN
                           => n863);
   U337 : AOI22_X1 port map( A1 => n83, A2 => predict_PC_8_10_port, B1 => n82, 
                           B2 => predict_PC_9_10_port, ZN => n865);
   U336 : AOI22_X1 port map( A1 => n557, A2 => predict_PC_10_10_port, B1 => n84
                           , B2 => predict_PC_11_10_port, ZN => n866);
   U335 : AOI22_X1 port map( A1 => n87, A2 => predict_PC_12_10_port, B1 => 
                           n86_port, B2 => predict_PC_13_10_port, ZN => n867);
   U334 : AOI22_X1 port map( A1 => n553, A2 => predict_PC_14_10_port, B1 => 
                           n554, B2 => predict_PC_15_10_port, ZN => n868);
   U333 : NAND4_X1 port map( A1 => n865, A2 => n866, A3 => n867, A4 => n868, ZN
                           => n864);
   U12 : AOI22_X1 port map( A1 => n75, A2 => predict_PC_0_9_port, B1 => n74, B2
                           => predict_PC_1_9_port, ZN => n561);
   U11 : AOI22_X1 port map( A1 => n77, A2 => predict_PC_2_9_port, B1 => n76, B2
                           => predict_PC_3_9_port, ZN => n562);
   U10 : AOI22_X1 port map( A1 => n79, A2 => predict_PC_4_9_port, B1 => n78, B2
                           => predict_PC_5_9_port, ZN => n563);
   U9 : AOI22_X1 port map( A1 => n81, A2 => predict_PC_6_9_port, B1 => n80, B2 
                           => predict_PC_7_9_port, ZN => n564);
   U8 : NAND4_X1 port map( A1 => n561, A2 => n562, A3 => n563, A4 => n564, ZN 
                           => n547);
   U7 : AOI22_X1 port map( A1 => n83, A2 => predict_PC_8_9_port, B1 => n82, B2 
                           => predict_PC_9_9_port, ZN => n549);
   U6 : AOI22_X1 port map( A1 => n85, A2 => predict_PC_10_9_port, B1 => n84, B2
                           => predict_PC_11_9_port, ZN => n550);
   U5 : AOI22_X1 port map( A1 => n87, A2 => predict_PC_12_9_port, B1 => 
                           n86_port, B2 => predict_PC_13_9_port, ZN => n551);
   U4 : AOI22_X1 port map( A1 => n89, A2 => predict_PC_14_9_port, B1 => n88, B2
                           => predict_PC_15_9_port, ZN => n552);
   U3 : NAND4_X1 port map( A1 => n549, A2 => n550, A3 => n551, A4 => n552, ZN 
                           => n548);
   U309 : AOI22_X1 port map( A1 => n75, A2 => predict_PC_0_13_port, B1 => n74, 
                           B2 => predict_PC_1_13_port, ZN => n839);
   U308 : AOI22_X1 port map( A1 => n569, A2 => predict_PC_2_13_port, B1 => n570
                           , B2 => predict_PC_3_13_port, ZN => n840);
   U307 : AOI22_X1 port map( A1 => n79, A2 => predict_PC_4_13_port, B1 => n78, 
                           B2 => predict_PC_5_13_port, ZN => n841);
   U306 : AOI22_X1 port map( A1 => n565, A2 => predict_PC_6_13_port, B1 => 
                           n566_port, B2 => predict_PC_7_13_port, ZN => n842);
   U305 : NAND4_X1 port map( A1 => n839, A2 => n840, A3 => n841, A4 => n842, ZN
                           => n833);
   U304 : AOI22_X1 port map( A1 => n83, A2 => predict_PC_8_13_port, B1 => n82, 
                           B2 => predict_PC_9_13_port, ZN => n835);
   U303 : AOI22_X1 port map( A1 => n557, A2 => predict_PC_10_13_port, B1 => n84
                           , B2 => predict_PC_11_13_port, ZN => n836);
   U302 : AOI22_X1 port map( A1 => n87, A2 => predict_PC_12_13_port, B1 => 
                           n86_port, B2 => predict_PC_13_13_port, ZN => n837);
   U301 : AOI22_X1 port map( A1 => n553, A2 => predict_PC_14_13_port, B1 => 
                           n554, B2 => predict_PC_15_13_port, ZN => n838);
   U300 : NAND4_X1 port map( A1 => n835, A2 => n836, A3 => n837, A4 => n838, ZN
                           => n834);
   U67 : AOI22_X1 port map( A1 => n571, A2 => predict_PC_0_4_port, B1 => n572, 
                           B2 => predict_PC_1_4_port, ZN => n619);
   U66 : AOI22_X1 port map( A1 => n77, A2 => predict_PC_2_4_port, B1 => n76, B2
                           => predict_PC_3_4_port, ZN => n620);
   U65 : AOI22_X1 port map( A1 => n567_port, A2 => predict_PC_4_4_port, B1 => 
                           n78, B2 => predict_PC_5_4_port, ZN => n621);
   U64 : AOI22_X1 port map( A1 => n81, A2 => predict_PC_6_4_port, B1 => n80, B2
                           => predict_PC_7_4_port, ZN => n622);
   U63 : NAND4_X1 port map( A1 => n619, A2 => n620, A3 => n621, A4 => n622, ZN 
                           => n613);
   U62 : AOI22_X1 port map( A1 => n559, A2 => predict_PC_8_4_port, B1 => n82, 
                           B2 => predict_PC_9_4_port, ZN => n615);
   U61 : AOI22_X1 port map( A1 => n85, A2 => predict_PC_10_4_port, B1 => n84, 
                           B2 => predict_PC_11_4_port, ZN => n616);
   U60 : AOI22_X1 port map( A1 => n555, A2 => predict_PC_12_4_port, B1 => 
                           n86_port, B2 => predict_PC_13_4_port, ZN => n617);
   U59 : AOI22_X1 port map( A1 => n89, A2 => predict_PC_14_4_port, B1 => n88, 
                           B2 => predict_PC_15_4_port, ZN => n618);
   U58 : NAND4_X1 port map( A1 => n615, A2 => n616, A3 => n617, A4 => n618, ZN 
                           => n614);
   U78 : AOI22_X1 port map( A1 => n571, A2 => predict_PC_0_3_port, B1 => n74, 
                           B2 => predict_PC_1_3_port, ZN => n629);
   U77 : AOI22_X1 port map( A1 => n77, A2 => predict_PC_2_3_port, B1 => n76, B2
                           => predict_PC_3_3_port, ZN => n630);
   U76 : AOI22_X1 port map( A1 => n79, A2 => predict_PC_4_3_port, B1 => n78, B2
                           => predict_PC_5_3_port, ZN => n631);
   U75 : AOI22_X1 port map( A1 => n81, A2 => predict_PC_6_3_port, B1 => n80, B2
                           => predict_PC_7_3_port, ZN => n632);
   U74 : NAND4_X1 port map( A1 => n629, A2 => n630, A3 => n631, A4 => n632, ZN 
                           => n623);
   U73 : AOI22_X1 port map( A1 => n83, A2 => predict_PC_8_3_port, B1 => n82, B2
                           => predict_PC_9_3_port, ZN => n625);
   U72 : AOI22_X1 port map( A1 => n85, A2 => predict_PC_10_3_port, B1 => n84, 
                           B2 => predict_PC_11_3_port, ZN => n626);
   U71 : AOI22_X1 port map( A1 => n87, A2 => predict_PC_12_3_port, B1 => 
                           n86_port, B2 => predict_PC_13_3_port, ZN => n627);
   U70 : AOI22_X1 port map( A1 => n89, A2 => predict_PC_14_3_port, B1 => n88, 
                           B2 => predict_PC_15_3_port, ZN => n628);
   U69 : NAND4_X1 port map( A1 => n625, A2 => n626, A3 => n627, A4 => n628, ZN 
                           => n624);
   U56 : AOI22_X1 port map( A1 => n75, A2 => predict_PC_0_5_port, B1 => n74, B2
                           => predict_PC_1_5_port, ZN => n609);
   U55 : AOI22_X1 port map( A1 => n77, A2 => predict_PC_2_5_port, B1 => n76, B2
                           => predict_PC_3_5_port, ZN => n610);
   U54 : AOI22_X1 port map( A1 => n79, A2 => predict_PC_4_5_port, B1 => n78, B2
                           => predict_PC_5_5_port, ZN => n611);
   U53 : AOI22_X1 port map( A1 => n81, A2 => predict_PC_6_5_port, B1 => n80, B2
                           => predict_PC_7_5_port, ZN => n612);
   U52 : NAND4_X1 port map( A1 => n609, A2 => n610, A3 => n611, A4 => n612, ZN 
                           => n603);
   U51 : AOI22_X1 port map( A1 => n83, A2 => predict_PC_8_5_port, B1 => n82, B2
                           => predict_PC_9_5_port, ZN => n605);
   U50 : AOI22_X1 port map( A1 => n85, A2 => predict_PC_10_5_port, B1 => n84, 
                           B2 => predict_PC_11_5_port, ZN => n606);
   U49 : AOI22_X1 port map( A1 => n87, A2 => predict_PC_12_5_port, B1 => 
                           n86_port, B2 => predict_PC_13_5_port, ZN => n607);
   U48 : AOI22_X1 port map( A1 => n89, A2 => predict_PC_14_5_port, B1 => n88, 
                           B2 => predict_PC_15_5_port, ZN => n608);
   U47 : NAND4_X1 port map( A1 => n605, A2 => n606, A3 => n607, A4 => n608, ZN 
                           => n604);
   U133 : AOI22_X1 port map( A1 => n75, A2 => predict_PC_0_28_port, B1 => n74, 
                           B2 => predict_PC_1_28_port, ZN => n679);
   U132 : AOI22_X1 port map( A1 => n77, A2 => predict_PC_2_28_port, B1 => n76, 
                           B2 => predict_PC_3_28_port, ZN => n680);
   U131 : AOI22_X1 port map( A1 => n79, A2 => predict_PC_4_28_port, B1 => n78, 
                           B2 => predict_PC_5_28_port, ZN => n681);
   U130 : AOI22_X1 port map( A1 => n81, A2 => predict_PC_6_28_port, B1 => n80, 
                           B2 => predict_PC_7_28_port, ZN => n682);
   U129 : NAND4_X1 port map( A1 => n679, A2 => n680, A3 => n681, A4 => n682, ZN
                           => n673);
   U128 : AOI22_X1 port map( A1 => n83, A2 => predict_PC_8_28_port, B1 => n82, 
                           B2 => predict_PC_9_28_port, ZN => n675);
   U127 : AOI22_X1 port map( A1 => n85, A2 => predict_PC_10_28_port, B1 => n84,
                           B2 => predict_PC_11_28_port, ZN => n676);
   U126 : AOI22_X1 port map( A1 => n87, A2 => predict_PC_12_28_port, B1 => 
                           n86_port, B2 => predict_PC_13_28_port, ZN => n677);
   U125 : AOI22_X1 port map( A1 => n89, A2 => predict_PC_14_28_port, B1 => n88,
                           B2 => predict_PC_15_28_port, ZN => n678);
   U124 : NAND4_X1 port map( A1 => n675, A2 => n676, A3 => n677, A4 => n678, ZN
                           => n674);
   U122 : AOI22_X1 port map( A1 => n571, A2 => predict_PC_0_29_port, B1 => n74,
                           B2 => predict_PC_1_29_port, ZN => n669);
   U121 : AOI22_X1 port map( A1 => n77, A2 => predict_PC_2_29_port, B1 => n76, 
                           B2 => predict_PC_3_29_port, ZN => n670);
   U120 : AOI22_X1 port map( A1 => n79, A2 => predict_PC_4_29_port, B1 => n78, 
                           B2 => predict_PC_5_29_port, ZN => n671);
   U119 : AOI22_X1 port map( A1 => n81, A2 => predict_PC_6_29_port, B1 => n80, 
                           B2 => predict_PC_7_29_port, ZN => n672);
   U118 : NAND4_X1 port map( A1 => n669, A2 => n670, A3 => n671, A4 => n672, ZN
                           => n663);
   U117 : AOI22_X1 port map( A1 => n83, A2 => predict_PC_8_29_port, B1 => n82, 
                           B2 => predict_PC_9_29_port, ZN => n665);
   U116 : AOI22_X1 port map( A1 => n85, A2 => predict_PC_10_29_port, B1 => n84,
                           B2 => predict_PC_11_29_port, ZN => n666);
   U115 : AOI22_X1 port map( A1 => n87, A2 => predict_PC_12_29_port, B1 => 
                           n86_port, B2 => predict_PC_13_29_port, ZN => n667);
   U114 : AOI22_X1 port map( A1 => n89, A2 => predict_PC_14_29_port, B1 => n88,
                           B2 => predict_PC_15_29_port, ZN => n668);
   U113 : NAND4_X1 port map( A1 => n665, A2 => n666, A3 => n667, A4 => n668, ZN
                           => n664);
   U353 : AOI22_X1 port map( A1 => n75, A2 => predict_PC_0_0_port, B1 => n74, 
                           B2 => predict_PC_1_0_port, ZN => n879);
   U352 : AOI22_X1 port map( A1 => n569, A2 => predict_PC_2_0_port, B1 => n570,
                           B2 => predict_PC_3_0_port, ZN => n880);
   U351 : AOI22_X1 port map( A1 => n79, A2 => predict_PC_4_0_port, B1 => n78, 
                           B2 => predict_PC_5_0_port, ZN => n881);
   U350 : AOI22_X1 port map( A1 => n565, A2 => predict_PC_6_0_port, B1 => 
                           n566_port, B2 => predict_PC_7_0_port, ZN => n882);
   U349 : NAND4_X1 port map( A1 => n879, A2 => n880, A3 => n881, A4 => n882, ZN
                           => n873);
   U348 : AOI22_X1 port map( A1 => n83, A2 => predict_PC_8_0_port, B1 => n82, 
                           B2 => predict_PC_9_0_port, ZN => n875);
   U347 : AOI22_X1 port map( A1 => n557, A2 => predict_PC_10_0_port, B1 => n84,
                           B2 => predict_PC_11_0_port, ZN => n876);
   U346 : AOI22_X1 port map( A1 => n87, A2 => predict_PC_12_0_port, B1 => 
                           n86_port, B2 => predict_PC_13_0_port, ZN => n877);
   U345 : AOI22_X1 port map( A1 => n553, A2 => predict_PC_14_0_port, B1 => n554
                           , B2 => predict_PC_15_0_port, ZN => n878);
   U344 : NAND4_X1 port map( A1 => n875, A2 => n876, A3 => n877, A4 => n878, ZN
                           => n874);
   U298 : AOI22_X1 port map( A1 => n75, A2 => predict_PC_0_14_port, B1 => n74, 
                           B2 => predict_PC_1_14_port, ZN => n829);
   U297 : AOI22_X1 port map( A1 => n569, A2 => predict_PC_2_14_port, B1 => n570
                           , B2 => predict_PC_3_14_port, ZN => n830);
   U296 : AOI22_X1 port map( A1 => n79, A2 => predict_PC_4_14_port, B1 => n78, 
                           B2 => predict_PC_5_14_port, ZN => n831);
   U295 : AOI22_X1 port map( A1 => n565, A2 => predict_PC_6_14_port, B1 => 
                           n566_port, B2 => predict_PC_7_14_port, ZN => n832);
   U294 : NAND4_X1 port map( A1 => n829, A2 => n830, A3 => n831, A4 => n832, ZN
                           => n823);
   U293 : AOI22_X1 port map( A1 => n83, A2 => predict_PC_8_14_port, B1 => n82, 
                           B2 => predict_PC_9_14_port, ZN => n825);
   U292 : AOI22_X1 port map( A1 => n557, A2 => predict_PC_10_14_port, B1 => n84
                           , B2 => predict_PC_11_14_port, ZN => n826);
   U291 : AOI22_X1 port map( A1 => n87, A2 => predict_PC_12_14_port, B1 => 
                           n86_port, B2 => predict_PC_13_14_port, ZN => n827);
   U290 : AOI22_X1 port map( A1 => n553, A2 => predict_PC_14_14_port, B1 => 
                           n554, B2 => predict_PC_15_14_port, ZN => n828);
   U289 : NAND4_X1 port map( A1 => n825, A2 => n826, A3 => n827, A4 => n828, ZN
                           => n824);
   U265 : AOI22_X1 port map( A1 => n75, A2 => predict_PC_0_17_port, B1 => n572,
                           B2 => predict_PC_1_17_port, ZN => n799);
   U264 : AOI22_X1 port map( A1 => n77, A2 => predict_PC_2_17_port, B1 => n76, 
                           B2 => predict_PC_3_17_port, ZN => n800);
   U263 : AOI22_X1 port map( A1 => n567_port, A2 => predict_PC_4_17_port, B1 =>
                           n568, B2 => predict_PC_5_17_port, ZN => n801);
   U262 : AOI22_X1 port map( A1 => n81, A2 => predict_PC_6_17_port, B1 => n80, 
                           B2 => predict_PC_7_17_port, ZN => n802);
   U261 : NAND4_X1 port map( A1 => n799, A2 => n800, A3 => n801, A4 => n802, ZN
                           => n793);
   U260 : AOI22_X1 port map( A1 => n559, A2 => predict_PC_8_17_port, B1 => n560
                           , B2 => predict_PC_9_17_port, ZN => n795);
   U259 : AOI22_X1 port map( A1 => n85, A2 => predict_PC_10_17_port, B1 => n84,
                           B2 => predict_PC_11_17_port, ZN => n796);
   U258 : AOI22_X1 port map( A1 => n555, A2 => predict_PC_12_17_port, B1 => 
                           n556, B2 => predict_PC_13_17_port, ZN => n797);
   U257 : AOI22_X1 port map( A1 => n89, A2 => predict_PC_14_17_port, B1 => n88,
                           B2 => predict_PC_15_17_port, ZN => n798);
   U256 : NAND4_X1 port map( A1 => n795, A2 => n796, A3 => n797, A4 => n798, ZN
                           => n794);
   U221 : AOI22_X1 port map( A1 => n75, A2 => predict_PC_0_20_port, B1 => n572,
                           B2 => predict_PC_1_20_port, ZN => n759);
   U220 : AOI22_X1 port map( A1 => n77, A2 => predict_PC_2_20_port, B1 => n76, 
                           B2 => predict_PC_3_20_port, ZN => n760);
   U219 : AOI22_X1 port map( A1 => n79, A2 => predict_PC_4_20_port, B1 => n78, 
                           B2 => predict_PC_5_20_port, ZN => n761);
   U218 : AOI22_X1 port map( A1 => n81, A2 => predict_PC_6_20_port, B1 => n80, 
                           B2 => predict_PC_7_20_port, ZN => n762);
   U217 : NAND4_X1 port map( A1 => n759, A2 => n760, A3 => n761, A4 => n762, ZN
                           => n753);
   U216 : AOI22_X1 port map( A1 => n83, A2 => predict_PC_8_20_port, B1 => n82, 
                           B2 => predict_PC_9_20_port, ZN => n755);
   U215 : AOI22_X1 port map( A1 => n85, A2 => predict_PC_10_20_port, B1 => n84,
                           B2 => predict_PC_11_20_port, ZN => n756);
   U214 : AOI22_X1 port map( A1 => n87, A2 => predict_PC_12_20_port, B1 => 
                           n86_port, B2 => predict_PC_13_20_port, ZN => n757);
   U213 : AOI22_X1 port map( A1 => n89, A2 => predict_PC_14_20_port, B1 => n88,
                           B2 => predict_PC_15_20_port, ZN => n758);
   U212 : NAND4_X1 port map( A1 => n755, A2 => n756, A3 => n757, A4 => n758, ZN
                           => n754);
   U320 : AOI22_X1 port map( A1 => n75, A2 => predict_PC_0_12_port, B1 => n74, 
                           B2 => predict_PC_1_12_port, ZN => n849);
   U319 : AOI22_X1 port map( A1 => n569, A2 => predict_PC_2_12_port, B1 => n570
                           , B2 => predict_PC_3_12_port, ZN => n850);
   U318 : AOI22_X1 port map( A1 => n79, A2 => predict_PC_4_12_port, B1 => n78, 
                           B2 => predict_PC_5_12_port, ZN => n851);
   U317 : AOI22_X1 port map( A1 => n565, A2 => predict_PC_6_12_port, B1 => 
                           n566_port, B2 => predict_PC_7_12_port, ZN => n852);
   U316 : NAND4_X1 port map( A1 => n849, A2 => n850, A3 => n851, A4 => n852, ZN
                           => n843);
   U315 : AOI22_X1 port map( A1 => n83, A2 => predict_PC_8_12_port, B1 => n82, 
                           B2 => predict_PC_9_12_port, ZN => n845);
   U314 : AOI22_X1 port map( A1 => n557, A2 => predict_PC_10_12_port, B1 => n84
                           , B2 => predict_PC_11_12_port, ZN => n846);
   U313 : AOI22_X1 port map( A1 => n87, A2 => predict_PC_12_12_port, B1 => 
                           n86_port, B2 => predict_PC_13_12_port, ZN => n847);
   U312 : AOI22_X1 port map( A1 => n553, A2 => predict_PC_14_12_port, B1 => 
                           n554, B2 => predict_PC_15_12_port, ZN => n848);
   U311 : NAND4_X1 port map( A1 => n845, A2 => n846, A3 => n847, A4 => n848, ZN
                           => n844);
   U34 : AOI22_X1 port map( A1 => n75, A2 => predict_PC_0_7_port, B1 => n572, 
                           B2 => predict_PC_1_7_port, ZN => n589);
   U33 : AOI22_X1 port map( A1 => n77, A2 => predict_PC_2_7_port, B1 => n76, B2
                           => predict_PC_3_7_port, ZN => n590);
   U32 : AOI22_X1 port map( A1 => n567_port, A2 => predict_PC_4_7_port, B1 => 
                           n78, B2 => predict_PC_5_7_port, ZN => n591);
   U31 : AOI22_X1 port map( A1 => n81, A2 => predict_PC_6_7_port, B1 => n80, B2
                           => predict_PC_7_7_port, ZN => n592);
   U30 : NAND4_X1 port map( A1 => n589, A2 => n590, A3 => n591, A4 => n592, ZN 
                           => n583);
   U29 : AOI22_X1 port map( A1 => n559, A2 => predict_PC_8_7_port, B1 => n82, 
                           B2 => predict_PC_9_7_port, ZN => n585);
   U28 : AOI22_X1 port map( A1 => n85, A2 => predict_PC_10_7_port, B1 => n84, 
                           B2 => predict_PC_11_7_port, ZN => n586);
   U27 : AOI22_X1 port map( A1 => n555, A2 => predict_PC_12_7_port, B1 => 
                           n86_port, B2 => predict_PC_13_7_port, ZN => n587);
   U26 : AOI22_X1 port map( A1 => n89, A2 => predict_PC_14_7_port, B1 => n88, 
                           B2 => predict_PC_15_7_port, ZN => n588);
   U25 : NAND4_X1 port map( A1 => n585, A2 => n586, A3 => n587, A4 => n588, ZN 
                           => n584);
   U100 : AOI22_X1 port map( A1 => n75, A2 => predict_PC_0_30_port, B1 => n74, 
                           B2 => predict_PC_1_30_port, ZN => n649);
   U99 : AOI22_X1 port map( A1 => n77, A2 => predict_PC_2_30_port, B1 => n76, 
                           B2 => predict_PC_3_30_port, ZN => n650);
   U98 : AOI22_X1 port map( A1 => n79, A2 => predict_PC_4_30_port, B1 => n78, 
                           B2 => predict_PC_5_30_port, ZN => n651);
   U97 : AOI22_X1 port map( A1 => n81, A2 => predict_PC_6_30_port, B1 => n80, 
                           B2 => predict_PC_7_30_port, ZN => n652);
   U96 : NAND4_X1 port map( A1 => n649, A2 => n650, A3 => n651, A4 => n652, ZN 
                           => n643);
   U95 : AOI22_X1 port map( A1 => n83, A2 => predict_PC_8_30_port, B1 => n82, 
                           B2 => predict_PC_9_30_port, ZN => n645);
   U94 : AOI22_X1 port map( A1 => n85, A2 => predict_PC_10_30_port, B1 => n84, 
                           B2 => predict_PC_11_30_port, ZN => n646);
   U93 : AOI22_X1 port map( A1 => n87, A2 => predict_PC_12_30_port, B1 => 
                           n86_port, B2 => predict_PC_13_30_port, ZN => n647);
   U92 : AOI22_X1 port map( A1 => n89, A2 => predict_PC_14_30_port, B1 => n88, 
                           B2 => predict_PC_15_30_port, ZN => n648);
   U91 : NAND4_X1 port map( A1 => n645, A2 => n646, A3 => n647, A4 => n648, ZN 
                           => n644);
   U89 : AOI22_X1 port map( A1 => n75, A2 => predict_PC_0_31_port, B1 => n74, 
                           B2 => predict_PC_1_31_port, ZN => n639);
   U88 : AOI22_X1 port map( A1 => n77, A2 => predict_PC_2_31_port, B1 => n76, 
                           B2 => predict_PC_3_31_port, ZN => n640);
   U87 : AOI22_X1 port map( A1 => n79, A2 => predict_PC_4_31_port, B1 => n78, 
                           B2 => predict_PC_5_31_port, ZN => n641);
   U86 : AOI22_X1 port map( A1 => n81, A2 => predict_PC_6_31_port, B1 => n80, 
                           B2 => predict_PC_7_31_port, ZN => n642);
   U85 : NAND4_X1 port map( A1 => n639, A2 => n640, A3 => n641, A4 => n642, ZN 
                           => n633);
   U84 : AOI22_X1 port map( A1 => n83, A2 => predict_PC_8_31_port, B1 => n82, 
                           B2 => predict_PC_9_31_port, ZN => n635);
   U83 : AOI22_X1 port map( A1 => n85, A2 => predict_PC_10_31_port, B1 => n84, 
                           B2 => predict_PC_11_31_port, ZN => n636);
   U82 : AOI22_X1 port map( A1 => n87, A2 => predict_PC_12_31_port, B1 => 
                           n86_port, B2 => predict_PC_13_31_port, ZN => n637);
   U81 : AOI22_X1 port map( A1 => n89, A2 => predict_PC_14_31_port, B1 => n88, 
                           B2 => predict_PC_15_31_port, ZN => n638);
   U80 : NAND4_X1 port map( A1 => n635, A2 => n636, A3 => n637, A4 => n638, ZN 
                           => n634);
   U155 : AOI22_X1 port map( A1 => n75, A2 => predict_PC_0_26_port, B1 => n74, 
                           B2 => predict_PC_1_26_port, ZN => n699);
   U154 : AOI22_X1 port map( A1 => n77, A2 => predict_PC_2_26_port, B1 => n76, 
                           B2 => predict_PC_3_26_port, ZN => n700);
   U153 : AOI22_X1 port map( A1 => n79, A2 => predict_PC_4_26_port, B1 => n78, 
                           B2 => predict_PC_5_26_port, ZN => n701);
   U152 : AOI22_X1 port map( A1 => n81, A2 => predict_PC_6_26_port, B1 => n80, 
                           B2 => predict_PC_7_26_port, ZN => n702);
   U151 : NAND4_X1 port map( A1 => n699, A2 => n700, A3 => n701, A4 => n702, ZN
                           => n693);
   U150 : AOI22_X1 port map( A1 => n83, A2 => predict_PC_8_26_port, B1 => n82, 
                           B2 => predict_PC_9_26_port, ZN => n695);
   U149 : AOI22_X1 port map( A1 => n85, A2 => predict_PC_10_26_port, B1 => n84,
                           B2 => predict_PC_11_26_port, ZN => n696);
   U148 : AOI22_X1 port map( A1 => n87, A2 => predict_PC_12_26_port, B1 => 
                           n86_port, B2 => predict_PC_13_26_port, ZN => n697);
   U147 : AOI22_X1 port map( A1 => n89, A2 => predict_PC_14_26_port, B1 => n88,
                           B2 => predict_PC_15_26_port, ZN => n698);
   U146 : NAND4_X1 port map( A1 => n695, A2 => n696, A3 => n697, A4 => n698, ZN
                           => n694);
   U188 : AOI22_X1 port map( A1 => n75, A2 => predict_PC_0_23_port, B1 => n74, 
                           B2 => predict_PC_1_23_port, ZN => n729);
   U187 : AOI22_X1 port map( A1 => n77, A2 => predict_PC_2_23_port, B1 => n76, 
                           B2 => predict_PC_3_23_port, ZN => n730);
   U186 : AOI22_X1 port map( A1 => n79, A2 => predict_PC_4_23_port, B1 => n78, 
                           B2 => predict_PC_5_23_port, ZN => n731);
   U185 : AOI22_X1 port map( A1 => n81, A2 => predict_PC_6_23_port, B1 => n80, 
                           B2 => predict_PC_7_23_port, ZN => n732);
   U184 : NAND4_X1 port map( A1 => n729, A2 => n730, A3 => n731, A4 => n732, ZN
                           => n723);
   U183 : AOI22_X1 port map( A1 => n83, A2 => predict_PC_8_23_port, B1 => n82, 
                           B2 => predict_PC_9_23_port, ZN => n725);
   U182 : AOI22_X1 port map( A1 => n85, A2 => predict_PC_10_23_port, B1 => n84,
                           B2 => predict_PC_11_23_port, ZN => n726);
   U181 : AOI22_X1 port map( A1 => n87, A2 => predict_PC_12_23_port, B1 => 
                           n86_port, B2 => predict_PC_13_23_port, ZN => n727);
   U180 : AOI22_X1 port map( A1 => n89, A2 => predict_PC_14_23_port, B1 => n88,
                           B2 => predict_PC_15_23_port, ZN => n728);
   U179 : NAND4_X1 port map( A1 => n725, A2 => n726, A3 => n727, A4 => n728, ZN
                           => n724);
   U287 : AOI22_X1 port map( A1 => n75, A2 => predict_PC_0_15_port, B1 => n74, 
                           B2 => predict_PC_1_15_port, ZN => n819);
   U286 : AOI22_X1 port map( A1 => n569, A2 => predict_PC_2_15_port, B1 => n570
                           , B2 => predict_PC_3_15_port, ZN => n820);
   U285 : AOI22_X1 port map( A1 => n79, A2 => predict_PC_4_15_port, B1 => n78, 
                           B2 => predict_PC_5_15_port, ZN => n821);
   U284 : AOI22_X1 port map( A1 => n565, A2 => predict_PC_6_15_port, B1 => 
                           n566_port, B2 => predict_PC_7_15_port, ZN => n822);
   U283 : NAND4_X1 port map( A1 => n819, A2 => n820, A3 => n821, A4 => n822, ZN
                           => n813);
   U282 : AOI22_X1 port map( A1 => n83, A2 => predict_PC_8_15_port, B1 => n82, 
                           B2 => predict_PC_9_15_port, ZN => n815);
   U281 : AOI22_X1 port map( A1 => n557, A2 => predict_PC_10_15_port, B1 => n84
                           , B2 => predict_PC_11_15_port, ZN => n816);
   U280 : AOI22_X1 port map( A1 => n87, A2 => predict_PC_12_15_port, B1 => 
                           n86_port, B2 => predict_PC_13_15_port, ZN => n817);
   U279 : AOI22_X1 port map( A1 => n553, A2 => predict_PC_14_15_port, B1 => 
                           n554, B2 => predict_PC_15_15_port, ZN => n818);
   U278 : NAND4_X1 port map( A1 => n815, A2 => n816, A3 => n817, A4 => n818, ZN
                           => n814);
   U199 : AOI22_X1 port map( A1 => n75, A2 => predict_PC_0_22_port, B1 => n74, 
                           B2 => predict_PC_1_22_port, ZN => n739);
   U198 : AOI22_X1 port map( A1 => n77, A2 => predict_PC_2_22_port, B1 => n76, 
                           B2 => predict_PC_3_22_port, ZN => n740);
   U197 : AOI22_X1 port map( A1 => n79, A2 => predict_PC_4_22_port, B1 => n78, 
                           B2 => predict_PC_5_22_port, ZN => n741);
   U196 : AOI22_X1 port map( A1 => n81, A2 => predict_PC_6_22_port, B1 => n80, 
                           B2 => predict_PC_7_22_port, ZN => n742);
   U195 : NAND4_X1 port map( A1 => n739, A2 => n740, A3 => n741, A4 => n742, ZN
                           => n733);
   U194 : AOI22_X1 port map( A1 => n83, A2 => predict_PC_8_22_port, B1 => n82, 
                           B2 => predict_PC_9_22_port, ZN => n735);
   U193 : AOI22_X1 port map( A1 => n85, A2 => predict_PC_10_22_port, B1 => n84,
                           B2 => predict_PC_11_22_port, ZN => n736);
   U192 : AOI22_X1 port map( A1 => n87, A2 => predict_PC_12_22_port, B1 => 
                           n86_port, B2 => predict_PC_13_22_port, ZN => n737);
   U191 : AOI22_X1 port map( A1 => n89, A2 => predict_PC_14_22_port, B1 => n88,
                           B2 => predict_PC_15_22_port, ZN => n738);
   U190 : NAND4_X1 port map( A1 => n735, A2 => n736, A3 => n737, A4 => n738, ZN
                           => n734);
   U166 : AOI22_X1 port map( A1 => n75, A2 => predict_PC_0_25_port, B1 => n74, 
                           B2 => predict_PC_1_25_port, ZN => n709);
   U165 : AOI22_X1 port map( A1 => n77, A2 => predict_PC_2_25_port, B1 => n76, 
                           B2 => predict_PC_3_25_port, ZN => n710);
   U164 : AOI22_X1 port map( A1 => n79, A2 => predict_PC_4_25_port, B1 => n78, 
                           B2 => predict_PC_5_25_port, ZN => n711);
   U163 : AOI22_X1 port map( A1 => n81, A2 => predict_PC_6_25_port, B1 => n80, 
                           B2 => predict_PC_7_25_port, ZN => n712);
   U162 : NAND4_X1 port map( A1 => n709, A2 => n710, A3 => n711, A4 => n712, ZN
                           => n703);
   U161 : AOI22_X1 port map( A1 => n83, A2 => predict_PC_8_25_port, B1 => n82, 
                           B2 => predict_PC_9_25_port, ZN => n705);
   U160 : AOI22_X1 port map( A1 => n85, A2 => predict_PC_10_25_port, B1 => n84,
                           B2 => predict_PC_11_25_port, ZN => n706);
   U159 : AOI22_X1 port map( A1 => n87, A2 => predict_PC_12_25_port, B1 => 
                           n86_port, B2 => predict_PC_13_25_port, ZN => n707);
   U158 : AOI22_X1 port map( A1 => n89, A2 => predict_PC_14_25_port, B1 => n88,
                           B2 => predict_PC_15_25_port, ZN => n708);
   U157 : NAND4_X1 port map( A1 => n705, A2 => n706, A3 => n707, A4 => n708, ZN
                           => n704);
   U331 : AOI22_X1 port map( A1 => n75, A2 => predict_PC_0_11_port, B1 => n74, 
                           B2 => predict_PC_1_11_port, ZN => n859);
   U330 : AOI22_X1 port map( A1 => n569, A2 => predict_PC_2_11_port, B1 => n570
                           , B2 => predict_PC_3_11_port, ZN => n860);
   U329 : AOI22_X1 port map( A1 => n79, A2 => predict_PC_4_11_port, B1 => n78, 
                           B2 => predict_PC_5_11_port, ZN => n861);
   U328 : AOI22_X1 port map( A1 => n565, A2 => predict_PC_6_11_port, B1 => 
                           n566_port, B2 => predict_PC_7_11_port, ZN => n862);
   U327 : NAND4_X1 port map( A1 => n859, A2 => n860, A3 => n861, A4 => n862, ZN
                           => n853);
   U326 : AOI22_X1 port map( A1 => n83, A2 => predict_PC_8_11_port, B1 => n82, 
                           B2 => predict_PC_9_11_port, ZN => n855);
   U325 : AOI22_X1 port map( A1 => n557, A2 => predict_PC_10_11_port, B1 => n84
                           , B2 => predict_PC_11_11_port, ZN => n856);
   U324 : AOI22_X1 port map( A1 => n87, A2 => predict_PC_12_11_port, B1 => 
                           n86_port, B2 => predict_PC_13_11_port, ZN => n857);
   U323 : AOI22_X1 port map( A1 => n553, A2 => predict_PC_14_11_port, B1 => 
                           n554, B2 => predict_PC_15_11_port, ZN => n858);
   U322 : NAND4_X1 port map( A1 => n855, A2 => n856, A3 => n857, A4 => n858, ZN
                           => n854);
   U144 : AOI22_X1 port map( A1 => n75, A2 => predict_PC_0_27_port, B1 => n74, 
                           B2 => predict_PC_1_27_port, ZN => n689);
   U143 : AOI22_X1 port map( A1 => n77, A2 => predict_PC_2_27_port, B1 => n76, 
                           B2 => predict_PC_3_27_port, ZN => n690);
   U142 : AOI22_X1 port map( A1 => n79, A2 => predict_PC_4_27_port, B1 => n78, 
                           B2 => predict_PC_5_27_port, ZN => n691);
   U141 : AOI22_X1 port map( A1 => n81, A2 => predict_PC_6_27_port, B1 => n80, 
                           B2 => predict_PC_7_27_port, ZN => n692);
   U140 : NAND4_X1 port map( A1 => n689, A2 => n690, A3 => n691, A4 => n692, ZN
                           => n683);
   U139 : AOI22_X1 port map( A1 => n83, A2 => predict_PC_8_27_port, B1 => n82, 
                           B2 => predict_PC_9_27_port, ZN => n685);
   U138 : AOI22_X1 port map( A1 => n85, A2 => predict_PC_10_27_port, B1 => n84,
                           B2 => predict_PC_11_27_port, ZN => n686);
   U137 : AOI22_X1 port map( A1 => n87, A2 => predict_PC_12_27_port, B1 => 
                           n86_port, B2 => predict_PC_13_27_port, ZN => n687);
   U136 : AOI22_X1 port map( A1 => n89, A2 => predict_PC_14_27_port, B1 => n88,
                           B2 => predict_PC_15_27_port, ZN => n688);
   U135 : NAND4_X1 port map( A1 => n685, A2 => n686, A3 => n687, A4 => n688, ZN
                           => n684);
   U177 : AOI22_X1 port map( A1 => n75, A2 => predict_PC_0_24_port, B1 => n74, 
                           B2 => predict_PC_1_24_port, ZN => n719);
   U176 : AOI22_X1 port map( A1 => n77, A2 => predict_PC_2_24_port, B1 => n76, 
                           B2 => predict_PC_3_24_port, ZN => n720);
   U175 : AOI22_X1 port map( A1 => n79, A2 => predict_PC_4_24_port, B1 => n78, 
                           B2 => predict_PC_5_24_port, ZN => n721);
   U174 : AOI22_X1 port map( A1 => n81, A2 => predict_PC_6_24_port, B1 => n80, 
                           B2 => predict_PC_7_24_port, ZN => n722);
   U173 : NAND4_X1 port map( A1 => n719, A2 => n720, A3 => n721, A4 => n722, ZN
                           => n713);
   U172 : AOI22_X1 port map( A1 => n83, A2 => predict_PC_8_24_port, B1 => n82, 
                           B2 => predict_PC_9_24_port, ZN => n715);
   U171 : AOI22_X1 port map( A1 => n85, A2 => predict_PC_10_24_port, B1 => n84,
                           B2 => predict_PC_11_24_port, ZN => n716);
   U170 : AOI22_X1 port map( A1 => n87, A2 => predict_PC_12_24_port, B1 => 
                           n86_port, B2 => predict_PC_13_24_port, ZN => n717);
   U169 : AOI22_X1 port map( A1 => n89, A2 => predict_PC_14_24_port, B1 => n88,
                           B2 => predict_PC_15_24_port, ZN => n718);
   U168 : NAND4_X1 port map( A1 => n715, A2 => n716, A3 => n717, A4 => n718, ZN
                           => n714);
   U479 : NAND2_X1 port map( A1 => n12, A2 => n10, ZN => n943);
   U469 : NAND2_X1 port map( A1 => n979, A2 => n978, ZN => n945);
   U468 : NOR2_X1 port map( A1 => n943, A2 => n945, ZN => N50);
   U449 : NOR2_X1 port map( A1 => n948, A2 => n947, ZN => N39);
   U466 : NAND2_X1 port map( A1 => n11, A2 => n9, ZN => n944);
   U445 : NOR2_X1 port map( A1 => n944, A2 => n947, ZN => N41);
   U450 : NOR2_X1 port map( A1 => n945, A2 => n947, ZN => N38);
   U465 : NAND2_X1 port map( A1 => n976, A2 => n12, ZN => n951);
   U460 : NOR2_X1 port map( A1 => n948, A2 => n951, ZN => N47);
   U477 : NAND2_X1 port map( A1 => n978, A2 => n11, ZN => n949);
   U462 : NOR2_X1 port map( A1 => n949, A2 => n951, ZN => N48);
   U440 : NOR2_X1 port map( A1 => n943, A2 => n944, ZN => N53);
   U456 : NAND2_X1 port map( A1 => n977, A2 => n10, ZN => n946);
   U455 : NOR2_X1 port map( A1 => n944, A2 => n946, ZN => N45);
   U447 : NOR2_X1 port map( A1 => n948, A2 => n946, ZN => N43);
   U471 : NOR2_X1 port map( A1 => n943, A2 => n948, ZN => N51);
   U453 : NOR2_X1 port map( A1 => n949, A2 => n946, ZN => N44);
   U444 : NOR2_X1 port map( A1 => n945, A2 => n946, ZN => N42);
   U464 : NOR2_X1 port map( A1 => n944, A2 => n951, ZN => N49);
   U458 : NOR2_X1 port map( A1 => n945, A2 => n951, ZN => N46);
   U476 : NOR2_X1 port map( A1 => n943, A2 => n949, ZN => N52);
   U448 : NOR2_X1 port map( A1 => n949, A2 => n947, ZN => N40);
   U355 : NOR2_X1 port map( A1 => stall_i, A2 => reset, ZN => n884);
   U354 : OAI22_X1 port map( A1 => stall_i, A2 => n883, B1 => n884, B2 => n975,
                           ZN => n955);
   U472 : NAND2_X1 port map( A1 => n979, A2 => n9, ZN => n948);
   U451 : NAND2_X1 port map( A1 => n977, A2 => n976, ZN => n947);
   U392 : INV_X1 port map( A => TAG_i(0), ZN => n903);
   U393 : INV_X1 port map( A => TAG_i(1), ZN => n974);
   U394 : INV_X1 port map( A => TAG_i(2), ZN => n973);
   U372 : NAND2_X1 port map( A1 => n973, A2 => n972, ZN => n896);
   U385 : NAND2_X1 port map( A1 => n903, A2 => n974, ZN => n893);
   U384 : NOR2_X1 port map( A1 => n902, A2 => n893, ZN => n559);
   U382 : NOR2_X1 port map( A1 => n902, A2 => n891, ZN => n560);
   U376 : NOR2_X1 port map( A1 => n893, A2 => n901, ZN => n555);
   U375 : NOR2_X1 port map( A1 => n891, A2 => n901, ZN => n556);
   U368 : NOR2_X1 port map( A1 => n893, A2 => n896, ZN => n571);
   U361 : NOR2_X1 port map( A1 => n893, A2 => n892, ZN => n567_port);
   U367 : NOR2_X1 port map( A1 => n891, A2 => n896, ZN => n572);
   U360 : NOR2_X1 port map( A1 => n891, A2 => n892, ZN => n568);
   U358 : AND4_X1 port map( A1 => n887, A2 => n888, A3 => n889, A4 => n890, ZN 
                           => n886);
   U373 : AND4_X1 port map( A1 => n897, A2 => n898, A3 => n899, A4 => n900, ZN 
                           => n885);
   U310 : OR2_X1 port map( A1 => n843, A2 => n844, ZN => 
                           predicted_next_PC_o_12_port);
   U123 : OR2_X1 port map( A1 => n673, A2 => n674, ZN => 
                           predicted_next_PC_o_28_port);
   U134 : OR2_X1 port map( A1 => n683, A2 => n684, ZN => 
                           predicted_next_PC_o_27_port);
   U24 : OR2_X1 port map( A1 => n583, A2 => n584, ZN => 
                           predicted_next_PC_o_7_port);
   U79 : OR2_X1 port map( A1 => n633, A2 => n634, ZN => 
                           predicted_next_PC_o_31_port);
   U90 : OR2_X1 port map( A1 => n643, A2 => n644, ZN => 
                           predicted_next_PC_o_30_port);
   U145 : OR2_X1 port map( A1 => n693, A2 => n694, ZN => 
                           predicted_next_PC_o_26_port);
   U222 : OR2_X1 port map( A1 => n763, A2 => n764, ZN => 
                           predicted_next_PC_o_1_port);
   U112 : OR2_X1 port map( A1 => n663, A2 => n664, ZN => 
                           predicted_next_PC_o_29_port);
   U299 : OR2_X1 port map( A1 => n833, A2 => n834, ZN => 
                           predicted_next_PC_o_13_port);
   U156 : OR2_X1 port map( A1 => n703, A2 => n704, ZN => 
                           predicted_next_PC_o_25_port);
   U211 : OR2_X1 port map( A1 => n753, A2 => n754, ZN => 
                           predicted_next_PC_o_20_port);
   U101 : OR2_X1 port map( A1 => n653, A2 => n654, ZN => 
                           predicted_next_PC_o_2_port);
   U244 : OR2_X1 port map( A1 => n783, A2 => n784, ZN => 
                           predicted_next_PC_o_18_port);
   U321 : OR2_X1 port map( A1 => n853, A2 => n854, ZN => 
                           predicted_next_PC_o_11_port);
   U68 : OR2_X1 port map( A1 => n623, A2 => n624, ZN => 
                           predicted_next_PC_o_3_port);
   U266 : OR2_X1 port map( A1 => n803, A2 => n804, ZN => 
                           predicted_next_PC_o_16_port);
   U167 : OR2_X1 port map( A1 => n713, A2 => n714, ZN => 
                           predicted_next_PC_o_24_port);
   U13 : OR2_X1 port map( A1 => n573, A2 => n574, ZN => 
                           predicted_next_PC_o_8_port);
   U233 : OR2_X1 port map( A1 => n773, A2 => n774, ZN => 
                           predicted_next_PC_o_19_port);
   U255 : OR2_X1 port map( A1 => n793, A2 => n794, ZN => 
                           predicted_next_PC_o_17_port);
   U277 : OR2_X1 port map( A1 => n813, A2 => n814, ZN => 
                           predicted_next_PC_o_15_port);
   U46 : OR2_X1 port map( A1 => n603, A2 => n604, ZN => 
                           predicted_next_PC_o_5_port);
   U178 : OR2_X1 port map( A1 => n723, A2 => n724, ZN => 
                           predicted_next_PC_o_23_port);
   U189 : OR2_X1 port map( A1 => n733, A2 => n734, ZN => 
                           predicted_next_PC_o_22_port);
   U35 : OR2_X1 port map( A1 => n593, A2 => n594, ZN => 
                           predicted_next_PC_o_6_port);
   U288 : OR2_X1 port map( A1 => n823, A2 => n824, ZN => 
                           predicted_next_PC_o_14_port);
   U332 : OR2_X1 port map( A1 => n863, A2 => n864, ZN => 
                           predicted_next_PC_o_10_port);
   U343 : OR2_X1 port map( A1 => n873, A2 => n874, ZN => 
                           predicted_next_PC_o_0_port);
   U57 : OR2_X1 port map( A1 => n613, A2 => n614, ZN => 
                           predicted_next_PC_o_4_port);
   U200 : OR2_X1 port map( A1 => n743, A2 => n744, ZN => 
                           predicted_next_PC_o_21_port);
   U2 : OR2_X1 port map( A1 => n547, A2 => n548, ZN => 
                           predicted_next_PC_o_9_port);
   U356 : INV_X1 port map( A => taken_o_port, ZN => n883);
   U459 : AND2_X1 port map( A1 => N47, A2 => N567, ZN => N278);
   U463 : AND2_X1 port map( A1 => N49, A2 => N567, ZN => N214);
   U457 : AND2_X1 port map( A1 => N46, A2 => N567, ZN => N310);
   U467 : AND2_X1 port map( A1 => N50, A2 => N567, ZN => N182);
   U454 : AND2_X1 port map( A1 => N45, A2 => N567, ZN => N342);
   U446 : AND2_X1 port map( A1 => N43, A2 => N567, ZN => N406);
   U452 : AND2_X1 port map( A1 => N44, A2 => N567, ZN => N374);
   U461 : AND2_X1 port map( A1 => N48, A2 => N567, ZN => N246);
   U442 : AND2_X1 port map( A1 => N41, A2 => N567, ZN => N470);
   U436 : AND2_X1 port map( A1 => N53, A2 => N567, ZN => N86);
   U438 : AND2_X1 port map( A1 => N38, A2 => N567, ZN => N566);
   U443 : AND2_X1 port map( A1 => N42, A2 => N567, ZN => N438);
   U441 : AND2_X1 port map( A1 => N40, A2 => N567, ZN => N502);
   U474 : AND2_X1 port map( A1 => N52, A2 => N567, ZN => N118);
   U439 : AND2_X1 port map( A1 => N39, A2 => N567, ZN => N534);
   U470 : AND2_X1 port map( A1 => N51, A2 => N567, ZN => N150);
   U475 : INV_X1 port map( A => stall_i, ZN => N567);
   U357 : AOI22_X1 port map( A1 => target_PC_i(3), A2 => n539, B1 => 
                           target_PC_i(2), B2 => n541, ZN => n1);
   U363 : NOR3_X1 port map( A1 => n53_port, A2 => n51_port, A3 => n52_port, ZN 
                           => n2);
   U364 : NAND3_X1 port map( A1 => n50_port, A2 => n1, A3 => n2, ZN => n49_port
                           );
   U370 : AOI22_X1 port map( A1 => n491, A2 => target_PC_i(27), B1 => n493, B2 
                           => target_PC_i(26), ZN => n3);
   U371 : INV_X1 port map( A => n3, ZN => n33);
   U378 : AOI22_X1 port map( A1 => target_PC_i(17), A2 => n511, B1 => 
                           target_PC_i(16), B2 => n513, ZN => n4);
   U379 : OAI221_X1 port map( B1 => target_PC_i(17), B2 => n511, C1 => 
                           target_PC_i(16), C2 => n513, A => n4, ZN => n63);
   U380 : OAI22_X1 port map( A1 => target_PC_i(5), A2 => n535, B1 => 
                           target_PC_i(4), B2 => n537, ZN => n5);
   U387 : INV_X1 port map( A => n5, ZN => n29);
   U389 : OAI22_X1 port map( A1 => target_PC_i(21), A2 => n503, B1 => 
                           target_PC_i(20), B2 => n505, ZN => n6);
   U390 : INV_X1 port map( A => n6, ZN => n36);
   U395 : OAI22_X1 port map( A1 => target_PC_i(7), A2 => n531, B1 => 
                           target_PC_i(6), B2 => n533, ZN => n7);
   U396 : INV_X1 port map( A => n7, ZN => n23);
   U397 : AOI22_X1 port map( A1 => n525, A2 => target_PC_i(10), B1 => n523, B2 
                           => target_PC_i(11), ZN => n8);
   U398 : OAI221_X1 port map( B1 => n525, B2 => target_PC_i(10), C1 => n523, C2
                           => target_PC_i(11), A => n8, ZN => n64);
   U399 : AND4_X1 port map( A1 => n35, A2 => n36, A3 => n37, A4 => n38_port, ZN
                           => n73);
   U400 : INV_X1 port map( A => n32, ZN => n28);
   U401 : INV_X1 port map( A => n39_port, ZN => n35);
   U402 : INV_X1 port map( A => n27, ZN => n24);
   U403 : BUF_X2 port map( A => n558, Z => n84);
   U404 : BUF_X2 port map( A => n555, Z => n87);
   U405 : BUF_X2 port map( A => n567_port, Z => n79);
   U406 : BUF_X2 port map( A => n571, Z => n75);
   U407 : BUF_X2 port map( A => n559, Z => n83);
   U408 : INV_X1 port map( A => reset, ZN => n95);
   U409 : INV_X1 port map( A => reset, ZN => n104);
   U410 : INV_X1 port map( A => reset, ZN => n99);
   U411 : INV_X1 port map( A => reset, ZN => n90);
   U412 : INV_X1 port map( A => reset, ZN => n94);
   U413 : INV_X1 port map( A => reset, ZN => n92);
   U414 : INV_X1 port map( A => reset, ZN => n100);
   U415 : INV_X1 port map( A => reset, ZN => n105);
   U416 : INV_X1 port map( A => reset, ZN => n109);
   U417 : INV_X1 port map( A => reset, ZN => n91);
   U418 : INV_X1 port map( A => reset, ZN => n108);
   U419 : INV_X1 port map( A => reset, ZN => n93);
   U420 : INV_X1 port map( A => reset, ZN => n107);
   U421 : INV_X1 port map( A => reset, ZN => n110);
   U422 : INV_X1 port map( A => reset, ZN => n101);
   U423 : INV_X1 port map( A => reset, ZN => n106);
   U424 : INV_X1 port map( A => reset, ZN => n112);
   U425 : INV_X1 port map( A => reset, ZN => n113);
   U426 : INV_X1 port map( A => reset, ZN => n103);
   U427 : INV_X1 port map( A => reset, ZN => n97);
   U428 : INV_X1 port map( A => reset, ZN => n98);
   U429 : INV_X1 port map( A => reset, ZN => n96);
   U430 : INV_X1 port map( A => reset, ZN => n111);
   U431 : INV_X1 port map( A => reset, ZN => n102);
   U432 : AOI21_X1 port map( B1 => n14, B2 => n13, A => n15, ZN => 
                           mispredict_o_port);
   U433 : NOR2_X1 port map( A1 => n16, A2 => n17, ZN => n14);
   U434 : OAI21_X1 port map( B1 => was_taken_i, B2 => n13, A => n546, ZN => n15
                           );
   U435 : AOI21_X1 port map( B1 => n885, B2 => n886, A => reset, ZN => 
                           taken_o_port);
   U437 : INV_X1 port map( A => TAG_i(3), ZN => n972);
   U473 : BUF_X1 port map( A => n568, Z => n78);
   U478 : BUF_X1 port map( A => n572, Z => n74);
   U480 : BUF_X1 port map( A => n556, Z => n86_port);
   U481 : BUF_X1 port map( A => n560, Z => n82);
   U482 : BUF_X1 port map( A => n554, Z => n88);
   U483 : BUF_X1 port map( A => n553, Z => n89);
   U484 : BUF_X1 port map( A => n557, Z => n85);
   U485 : BUF_X1 port map( A => n566_port, Z => n80);
   U486 : BUF_X1 port map( A => n565, Z => n81);
   U487 : BUF_X1 port map( A => n570, Z => n76);
   U488 : BUF_X1 port map( A => n569, Z => n77);
   U489 : NOR2_X1 port map( A1 => n33, A2 => n34, ZN => n19);
   U490 : OAI22_X1 port map( A1 => target_PC_i(26), A2 => n493, B1 => 
                           target_PC_i(27), B2 => n491, ZN => n34);
   U491 : NOR2_X1 port map( A1 => n65, A2 => n66, ZN => n45_port);
   U492 : OAI22_X1 port map( A1 => target_PC_i(19), A2 => n507, B1 => n509, B2 
                           => target_PC_i(18), ZN => n66);
   U493 : NAND2_X1 port map( A1 => target_PC_i(18), A2 => n509, ZN => n68);
   U494 : NOR2_X1 port map( A1 => target_PC_i(13), A2 => n519, ZN => n52_port);
   U495 : NOR2_X1 port map( A1 => target_PC_i(9), A2 => n527, ZN => n58);
   U496 : NOR2_X1 port map( A1 => n895, A2 => n896, ZN => n569);
   U497 : NOR2_X1 port map( A1 => n895, A2 => n892, ZN => n565);
   U498 : NOR2_X1 port map( A1 => n895, A2 => n902, ZN => n557);
   U499 : NOR2_X1 port map( A1 => n895, A2 => n901, ZN => n553);
   U500 : NOR2_X1 port map( A1 => n894, A2 => n896, ZN => n570);
   U501 : NOR2_X1 port map( A1 => n894, A2 => n892, ZN => n566_port);
   U502 : NOR2_X1 port map( A1 => n894, A2 => n901, ZN => n554);
   U503 : NOR2_X1 port map( A1 => n902, A2 => n894, ZN => n558);
   U504 : NAND3_X1 port map( A1 => n54, A2 => n55, A3 => n56, ZN => n48_port);
   U505 : NAND2_X1 port map( A1 => target_PC_i(14), A2 => n517, ZN => n61);
   U506 : NAND2_X1 port map( A1 => n61, A2 => n62, ZN => n59);
   U507 : NAND2_X1 port map( A1 => target_PC_i(15), A2 => n515, ZN => n62);
   U508 : NAND4_X1 port map( A1 => n28, A2 => n29, A3 => n31, A4 => n30, ZN => 
                           n21);
   U509 : NOR2_X1 port map( A1 => n21, A2 => n22, ZN => n20);
   U510 : NAND2_X1 port map( A1 => target_PC_i(29), A2 => n487, ZN => n72);
   U511 : NAND2_X1 port map( A1 => n71, A2 => n72, ZN => n69);
   U512 : OAI22_X1 port map( A1 => n517, A2 => target_PC_i(14), B1 => 
                           target_PC_i(15), B2 => n515, ZN => n60);
   U513 : NOR2_X1 port map( A1 => n59, A2 => n60, ZN => n54);
   U514 : AOI22_X1 port map( A1 => n533, A2 => target_PC_i(6), B1 => 
                           target_PC_i(7), B2 => n531, ZN => n25);
   U515 : NAND4_X1 port map( A1 => n23, A2 => n24, A3 => n25, A4 => n26, ZN => 
                           n22);
   U516 : NAND2_X1 port map( A1 => target_PC_i(28), A2 => n489, ZN => n71);
   U517 : NAND2_X1 port map( A1 => target_PC_i(19), A2 => n507, ZN => n67);
   U518 : NAND2_X1 port map( A1 => n67, A2 => n68, ZN => n65);
   U519 : AOI22_X1 port map( A1 => n529, A2 => target_PC_i(8), B1 => 
                           target_PC_i(9), B2 => n527, ZN => n56);
   U520 : AOI22_X1 port map( A1 => n521, A2 => target_PC_i(12), B1 => 
                           target_PC_i(13), B2 => n519, ZN => n50_port);
   U521 : NAND4_X1 port map( A1 => n47_port, A2 => n44_port, A3 => n46_port, A4
                           => n45_port, ZN => n16);
   U522 : NAND2_X1 port map( A1 => target_PC_i(31), A2 => n483, ZN => n42_port)
                           ;
   U523 : NAND2_X1 port map( A1 => n42_port, A2 => n43_port, ZN => n40_port);
   U524 : NAND2_X1 port map( A1 => target_PC_i(30), A2 => n485, ZN => n43_port)
                           ;
   U525 : AOI22_X1 port map( A1 => target_PC_i(24), A2 => n497, B1 => 
                           target_PC_i(25), B2 => n495, ZN => n37);
   U526 : AOI22_X1 port map( A1 => n505, A2 => target_PC_i(20), B1 => 
                           target_PC_i(21), B2 => n503, ZN => n38_port);
   U527 : AOI22_X1 port map( A1 => target_PC_i(1), A2 => n543, B1 => 
                           target_PC_i(0), B2 => n545, ZN => n26);
   U528 : NAND4_X1 port map( A1 => n20, A2 => n73, A3 => n19, A4 => n18, ZN => 
                           n17);
   U529 : OAI22_X1 port map( A1 => target_PC_i(28), A2 => n489, B1 => 
                           target_PC_i(29), B2 => n487, ZN => n70);
   U530 : NOR2_X1 port map( A1 => n69, A2 => n70, ZN => n44_port);
   U531 : NOR2_X1 port map( A1 => target_PC_i(8), A2 => n529, ZN => n57);
   U532 : NOR2_X1 port map( A1 => n57, A2 => n58, ZN => n55);
   U533 : OAI22_X1 port map( A1 => target_PC_i(3), A2 => n539, B1 => 
                           target_PC_i(2), B2 => n541, ZN => n53_port);
   U534 : NOR2_X1 port map( A1 => target_PC_i(12), A2 => n521, ZN => n51_port);
   U535 : OAI22_X1 port map( A1 => target_PC_i(31), A2 => n483, B1 => 
                           target_PC_i(30), B2 => n485, ZN => n41_port);
   U536 : NOR2_X1 port map( A1 => n40_port, A2 => n41_port, ZN => n18);
   U537 : OAI22_X1 port map( A1 => target_PC_i(24), A2 => n497, B1 => 
                           target_PC_i(25), B2 => n495, ZN => n39_port);
   U538 : OAI22_X1 port map( A1 => target_PC_i(23), A2 => n499, B1 => 
                           target_PC_i(22), B2 => n501, ZN => n32);
   U539 : OAI22_X1 port map( A1 => target_PC_i(1), A2 => n543, B1 => 
                           target_PC_i(0), B2 => n545, ZN => n27);
   U540 : NOR2_X1 port map( A1 => n48_port, A2 => n49_port, ZN => n47_port);
   U541 : AOI22_X1 port map( A1 => n537, A2 => target_PC_i(4), B1 => 
                           target_PC_i(5), B2 => n535, ZN => n31);
   U542 : AOI22_X1 port map( A1 => target_PC_i(23), A2 => n499, B1 => 
                           target_PC_i(22), B2 => n501, ZN => n30);
   U543 : NOR2_X1 port map( A1 => n63, A2 => n64, ZN => n46_port);
   U544 : NAND2_X1 port map( A1 => TAG_i(3), A2 => n973, ZN => n902);
   U545 : NAND2_X1 port map( A1 => TAG_i(2), A2 => TAG_i(3), ZN => n901);

end SYN_bhe;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity fetch_block is

   port( branch_target_i, sum_addr_i, A_i, NPC4_i : in std_logic_vector (31 
         downto 0);  S_MUX_PC_BUS_i : in std_logic_vector (1 downto 0);  PC_o, 
         PC4_o, PC_BUS_pre_BTB : out std_logic_vector (31 downto 0);  stall_i, 
         take_prediction_i, mispredict_i : in std_logic;  predicted_PC : in 
         std_logic_vector (31 downto 0);  clk, rst : in std_logic);

end fetch_block;

architecture SYN_Struct of fetch_block is

   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component mux41_1
      port( IN0, IN1, IN2, IN3 : in std_logic_vector (31 downto 0);  CTRL : in 
            std_logic_vector (1 downto 0);  OUT1 : out std_logic_vector (31 
            downto 0));
   end component;
   
   component mux41_0
      port( IN0, IN1, IN2, IN3 : in std_logic_vector (31 downto 0);  CTRL : in 
            std_logic_vector (1 downto 0);  OUT1 : out std_logic_vector (31 
            downto 0));
   end component;
   
   component add4
      port( IN1 : in std_logic_vector (31 downto 0);  OUT1 : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component ff32_en_0
      port( D : in std_logic_vector (31 downto 0);  en, clk, rst : in std_logic
            ;  Q : out std_logic_vector (31 downto 0));
   end component;
   
   signal PC_o_31_port, PC_o_30_port, PC_o_29_port, PC_o_28_port, PC_o_27_port,
      PC_o_26_port, PC_o_25_port, PC_o_24_port, PC_o_23_port, PC_o_22_port, 
      PC_o_21_port, PC_o_20_port, PC_o_19_port, PC_o_18_port, PC_o_17_port, 
      PC_o_16_port, PC_o_15_port, PC_o_14_port, PC_o_13_port, PC_o_12_port, 
      PC_o_11_port, PC_o_10_port, PC_o_9_port, PC_o_8_port, PC_o_7_port, 
      PC_o_6_port, PC_o_5_port, PC_o_4_port, PC_o_3_port, PC_o_2_port, 
      PC_o_1_port, PC_o_0_port, PC4_o_31_port, PC4_o_30_port, PC4_o_29_port, 
      PC4_o_28_port, PC4_o_27_port, PC4_o_26_port, PC4_o_25_port, PC4_o_24_port
      , PC4_o_23_port, PC4_o_22_port, PC4_o_21_port, PC4_o_20_port, 
      PC4_o_19_port, PC4_o_18_port, PC4_o_17_port, PC4_o_16_port, PC4_o_15_port
      , PC4_o_14_port, PC4_o_13_port, PC4_o_12_port, PC4_o_11_port, 
      PC4_o_10_port, PC4_o_9_port, PC4_o_8_port, PC4_o_7_port, PC4_o_6_port, 
      PC4_o_5_port, PC4_o_4_port, PC4_o_3_port, PC4_o_2_port, PC4_o_1_port, 
      PC4_o_0_port, PC_BUS_pre_BTB_31_port, PC_BUS_pre_BTB_30_port, n4, n5, 
      PC_BUS_pre_BTB_27_port, PC_BUS_pre_BTB_26_port, PC_BUS_pre_BTB_25_port, 
      PC_BUS_pre_BTB_24_port, PC_BUS_pre_BTB_23_port, PC_BUS_pre_BTB_22_port, 
      PC_BUS_pre_BTB_21_port, PC_BUS_pre_BTB_20_port, PC_BUS_pre_BTB_19_port, 
      PC_BUS_pre_BTB_18_port, PC_BUS_pre_BTB_17_port, PC_BUS_pre_BTB_16_port, 
      PC_BUS_pre_BTB_15_port, PC_BUS_pre_BTB_14_port, PC_BUS_pre_BTB_13_port, 
      PC_BUS_pre_BTB_12_port, PC_BUS_pre_BTB_11_port, PC_BUS_pre_BTB_10_port, 
      PC_BUS_pre_BTB_9_port, PC_BUS_pre_BTB_8_port, PC_BUS_pre_BTB_7_port, 
      PC_BUS_pre_BTB_6_port, PC_BUS_pre_BTB_5_port, PC_BUS_pre_BTB_4_port, 
      PC_BUS_pre_BTB_3_port, PC_BUS_pre_BTB_2_port, PC_BUS_pre_BTB_1_port, 
      PC_BUS_pre_BTB_0_port, en_IR, PC_BUS_31_port, PC_BUS_30_port, 
      PC_BUS_29_port, PC_BUS_28_port, PC_BUS_27_port, PC_BUS_26_port, 
      PC_BUS_25_port, PC_BUS_24_port, PC_BUS_23_port, PC_BUS_22_port, 
      PC_BUS_21_port, PC_BUS_20_port, PC_BUS_19_port, PC_BUS_18_port, 
      PC_BUS_17_port, PC_BUS_16_port, PC_BUS_15_port, PC_BUS_14_port, 
      PC_BUS_13_port, PC_BUS_12_port, PC_BUS_11_port, PC_BUS_10_port, 
      PC_BUS_9_port, PC_BUS_8_port, PC_BUS_7_port, PC_BUS_6_port, PC_BUS_5_port
      , PC_BUS_4_port, PC_BUS_3_port, PC_BUS_2_port, PC_BUS_1_port, 
      PC_BUS_0_port, PC_BUS_pre_BTB_29_port, PC_BUS_pre_BTB_28_port : std_logic
      ;

begin
   PC_o <= ( PC_o_31_port, PC_o_30_port, PC_o_29_port, PC_o_28_port, 
      PC_o_27_port, PC_o_26_port, PC_o_25_port, PC_o_24_port, PC_o_23_port, 
      PC_o_22_port, PC_o_21_port, PC_o_20_port, PC_o_19_port, PC_o_18_port, 
      PC_o_17_port, PC_o_16_port, PC_o_15_port, PC_o_14_port, PC_o_13_port, 
      PC_o_12_port, PC_o_11_port, PC_o_10_port, PC_o_9_port, PC_o_8_port, 
      PC_o_7_port, PC_o_6_port, PC_o_5_port, PC_o_4_port, PC_o_3_port, 
      PC_o_2_port, PC_o_1_port, PC_o_0_port );
   PC4_o <= ( PC4_o_31_port, PC4_o_30_port, PC4_o_29_port, PC4_o_28_port, 
      PC4_o_27_port, PC4_o_26_port, PC4_o_25_port, PC4_o_24_port, PC4_o_23_port
      , PC4_o_22_port, PC4_o_21_port, PC4_o_20_port, PC4_o_19_port, 
      PC4_o_18_port, PC4_o_17_port, PC4_o_16_port, PC4_o_15_port, PC4_o_14_port
      , PC4_o_13_port, PC4_o_12_port, PC4_o_11_port, PC4_o_10_port, 
      PC4_o_9_port, PC4_o_8_port, PC4_o_7_port, PC4_o_6_port, PC4_o_5_port, 
      PC4_o_4_port, PC4_o_3_port, PC4_o_2_port, PC4_o_1_port, PC4_o_0_port );
   PC_BUS_pre_BTB <= ( PC_BUS_pre_BTB_31_port, PC_BUS_pre_BTB_30_port, 
      PC_BUS_pre_BTB_29_port, PC_BUS_pre_BTB_28_port, PC_BUS_pre_BTB_27_port, 
      PC_BUS_pre_BTB_26_port, PC_BUS_pre_BTB_25_port, PC_BUS_pre_BTB_24_port, 
      PC_BUS_pre_BTB_23_port, PC_BUS_pre_BTB_22_port, PC_BUS_pre_BTB_21_port, 
      PC_BUS_pre_BTB_20_port, PC_BUS_pre_BTB_19_port, PC_BUS_pre_BTB_18_port, 
      PC_BUS_pre_BTB_17_port, PC_BUS_pre_BTB_16_port, PC_BUS_pre_BTB_15_port, 
      PC_BUS_pre_BTB_14_port, PC_BUS_pre_BTB_13_port, PC_BUS_pre_BTB_12_port, 
      PC_BUS_pre_BTB_11_port, PC_BUS_pre_BTB_10_port, PC_BUS_pre_BTB_9_port, 
      PC_BUS_pre_BTB_8_port, PC_BUS_pre_BTB_7_port, PC_BUS_pre_BTB_6_port, 
      PC_BUS_pre_BTB_5_port, PC_BUS_pre_BTB_4_port, PC_BUS_pre_BTB_3_port, 
      PC_BUS_pre_BTB_2_port, PC_BUS_pre_BTB_1_port, PC_BUS_pre_BTB_0_port );
   
   PC : ff32_en_0 port map( D(31) => PC_BUS_31_port, D(30) => PC_BUS_30_port, 
                           D(29) => PC_BUS_29_port, D(28) => PC_BUS_28_port, 
                           D(27) => PC_BUS_27_port, D(26) => PC_BUS_26_port, 
                           D(25) => PC_BUS_25_port, D(24) => PC_BUS_24_port, 
                           D(23) => PC_BUS_23_port, D(22) => PC_BUS_22_port, 
                           D(21) => PC_BUS_21_port, D(20) => PC_BUS_20_port, 
                           D(19) => PC_BUS_19_port, D(18) => PC_BUS_18_port, 
                           D(17) => PC_BUS_17_port, D(16) => PC_BUS_16_port, 
                           D(15) => PC_BUS_15_port, D(14) => PC_BUS_14_port, 
                           D(13) => PC_BUS_13_port, D(12) => PC_BUS_12_port, 
                           D(11) => PC_BUS_11_port, D(10) => PC_BUS_10_port, 
                           D(9) => PC_BUS_9_port, D(8) => PC_BUS_8_port, D(7) 
                           => PC_BUS_7_port, D(6) => PC_BUS_6_port, D(5) => 
                           PC_BUS_5_port, D(4) => PC_BUS_4_port, D(3) => 
                           PC_BUS_3_port, D(2) => PC_BUS_2_port, D(1) => 
                           PC_BUS_1_port, D(0) => PC_BUS_0_port, en => en_IR, 
                           clk => clk, rst => rst, Q(31) => PC_o_31_port, Q(30)
                           => PC_o_30_port, Q(29) => PC_o_29_port, Q(28) => 
                           PC_o_28_port, Q(27) => PC_o_27_port, Q(26) => 
                           PC_o_26_port, Q(25) => PC_o_25_port, Q(24) => 
                           PC_o_24_port, Q(23) => PC_o_23_port, Q(22) => 
                           PC_o_22_port, Q(21) => PC_o_21_port, Q(20) => 
                           PC_o_20_port, Q(19) => PC_o_19_port, Q(18) => 
                           PC_o_18_port, Q(17) => PC_o_17_port, Q(16) => 
                           PC_o_16_port, Q(15) => PC_o_15_port, Q(14) => 
                           PC_o_14_port, Q(13) => PC_o_13_port, Q(12) => 
                           PC_o_12_port, Q(11) => PC_o_11_port, Q(10) => 
                           PC_o_10_port, Q(9) => PC_o_9_port, Q(8) => 
                           PC_o_8_port, Q(7) => PC_o_7_port, Q(6) => 
                           PC_o_6_port, Q(5) => PC_o_5_port, Q(4) => 
                           PC_o_4_port, Q(3) => PC_o_3_port, Q(2) => 
                           PC_o_2_port, Q(1) => PC_o_1_port, Q(0) => 
                           PC_o_0_port);
   PCADD : add4 port map( IN1(31) => PC_o_31_port, IN1(30) => PC_o_30_port, 
                           IN1(29) => PC_o_29_port, IN1(28) => PC_o_28_port, 
                           IN1(27) => PC_o_27_port, IN1(26) => PC_o_26_port, 
                           IN1(25) => PC_o_25_port, IN1(24) => PC_o_24_port, 
                           IN1(23) => PC_o_23_port, IN1(22) => PC_o_22_port, 
                           IN1(21) => PC_o_21_port, IN1(20) => PC_o_20_port, 
                           IN1(19) => PC_o_19_port, IN1(18) => PC_o_18_port, 
                           IN1(17) => PC_o_17_port, IN1(16) => PC_o_16_port, 
                           IN1(15) => PC_o_15_port, IN1(14) => PC_o_14_port, 
                           IN1(13) => PC_o_13_port, IN1(12) => PC_o_12_port, 
                           IN1(11) => PC_o_11_port, IN1(10) => PC_o_10_port, 
                           IN1(9) => PC_o_9_port, IN1(8) => PC_o_8_port, IN1(7)
                           => PC_o_7_port, IN1(6) => PC_o_6_port, IN1(5) => 
                           PC_o_5_port, IN1(4) => PC_o_4_port, IN1(3) => 
                           PC_o_3_port, IN1(2) => PC_o_2_port, IN1(1) => 
                           PC_o_1_port, IN1(0) => PC_o_0_port, OUT1(31) => 
                           PC4_o_31_port, OUT1(30) => PC4_o_30_port, OUT1(29) 
                           => PC4_o_29_port, OUT1(28) => PC4_o_28_port, 
                           OUT1(27) => PC4_o_27_port, OUT1(26) => PC4_o_26_port
                           , OUT1(25) => PC4_o_25_port, OUT1(24) => 
                           PC4_o_24_port, OUT1(23) => PC4_o_23_port, OUT1(22) 
                           => PC4_o_22_port, OUT1(21) => PC4_o_21_port, 
                           OUT1(20) => PC4_o_20_port, OUT1(19) => PC4_o_19_port
                           , OUT1(18) => PC4_o_18_port, OUT1(17) => 
                           PC4_o_17_port, OUT1(16) => PC4_o_16_port, OUT1(15) 
                           => PC4_o_15_port, OUT1(14) => PC4_o_14_port, 
                           OUT1(13) => PC4_o_13_port, OUT1(12) => PC4_o_12_port
                           , OUT1(11) => PC4_o_11_port, OUT1(10) => 
                           PC4_o_10_port, OUT1(9) => PC4_o_9_port, OUT1(8) => 
                           PC4_o_8_port, OUT1(7) => PC4_o_7_port, OUT1(6) => 
                           PC4_o_6_port, OUT1(5) => PC4_o_5_port, OUT1(4) => 
                           PC4_o_4_port, OUT1(3) => PC4_o_3_port, OUT1(2) => 
                           PC4_o_2_port, OUT1(1) => PC4_o_1_port, OUT1(0) => 
                           PC4_o_0_port);
   MUXTARGET : mux41_0 port map( IN0(31) => NPC4_i(31), IN0(30) => NPC4_i(30), 
                           IN0(29) => NPC4_i(29), IN0(28) => NPC4_i(28), 
                           IN0(27) => NPC4_i(27), IN0(26) => NPC4_i(26), 
                           IN0(25) => NPC4_i(25), IN0(24) => NPC4_i(24), 
                           IN0(23) => NPC4_i(23), IN0(22) => NPC4_i(22), 
                           IN0(21) => NPC4_i(21), IN0(20) => NPC4_i(20), 
                           IN0(19) => NPC4_i(19), IN0(18) => NPC4_i(18), 
                           IN0(17) => NPC4_i(17), IN0(16) => NPC4_i(16), 
                           IN0(15) => NPC4_i(15), IN0(14) => NPC4_i(14), 
                           IN0(13) => NPC4_i(13), IN0(12) => NPC4_i(12), 
                           IN0(11) => NPC4_i(11), IN0(10) => NPC4_i(10), IN0(9)
                           => NPC4_i(9), IN0(8) => NPC4_i(8), IN0(7) => 
                           NPC4_i(7), IN0(6) => NPC4_i(6), IN0(5) => NPC4_i(5),
                           IN0(4) => NPC4_i(4), IN0(3) => NPC4_i(3), IN0(2) => 
                           NPC4_i(2), IN0(1) => NPC4_i(1), IN0(0) => NPC4_i(0),
                           IN1(31) => A_i(31), IN1(30) => A_i(30), IN1(29) => 
                           A_i(29), IN1(28) => A_i(28), IN1(27) => A_i(27), 
                           IN1(26) => A_i(26), IN1(25) => A_i(25), IN1(24) => 
                           A_i(24), IN1(23) => A_i(23), IN1(22) => A_i(22), 
                           IN1(21) => A_i(21), IN1(20) => A_i(20), IN1(19) => 
                           A_i(19), IN1(18) => A_i(18), IN1(17) => A_i(17), 
                           IN1(16) => A_i(16), IN1(15) => A_i(15), IN1(14) => 
                           A_i(14), IN1(13) => A_i(13), IN1(12) => A_i(12), 
                           IN1(11) => A_i(11), IN1(10) => A_i(10), IN1(9) => 
                           A_i(9), IN1(8) => A_i(8), IN1(7) => A_i(7), IN1(6) 
                           => A_i(6), IN1(5) => A_i(5), IN1(4) => A_i(4), 
                           IN1(3) => A_i(3), IN1(2) => A_i(2), IN1(1) => A_i(1)
                           , IN1(0) => A_i(0), IN2(31) => sum_addr_i(31), 
                           IN2(30) => sum_addr_i(30), IN2(29) => sum_addr_i(29)
                           , IN2(28) => sum_addr_i(28), IN2(27) => 
                           sum_addr_i(27), IN2(26) => sum_addr_i(26), IN2(25) 
                           => sum_addr_i(25), IN2(24) => sum_addr_i(24), 
                           IN2(23) => sum_addr_i(23), IN2(22) => sum_addr_i(22)
                           , IN2(21) => sum_addr_i(21), IN2(20) => 
                           sum_addr_i(20), IN2(19) => sum_addr_i(19), IN2(18) 
                           => sum_addr_i(18), IN2(17) => sum_addr_i(17), 
                           IN2(16) => sum_addr_i(16), IN2(15) => sum_addr_i(15)
                           , IN2(14) => sum_addr_i(14), IN2(13) => 
                           sum_addr_i(13), IN2(12) => sum_addr_i(12), IN2(11) 
                           => sum_addr_i(11), IN2(10) => sum_addr_i(10), IN2(9)
                           => sum_addr_i(9), IN2(8) => sum_addr_i(8), IN2(7) =>
                           sum_addr_i(7), IN2(6) => sum_addr_i(6), IN2(5) => 
                           sum_addr_i(5), IN2(4) => sum_addr_i(4), IN2(3) => 
                           sum_addr_i(3), IN2(2) => sum_addr_i(2), IN2(1) => 
                           sum_addr_i(1), IN2(0) => sum_addr_i(0), IN3(31) => 
                           branch_target_i(31), IN3(30) => branch_target_i(30),
                           IN3(29) => branch_target_i(29), IN3(28) => 
                           branch_target_i(28), IN3(27) => branch_target_i(27),
                           IN3(26) => branch_target_i(26), IN3(25) => 
                           branch_target_i(25), IN3(24) => branch_target_i(24),
                           IN3(23) => branch_target_i(23), IN3(22) => 
                           branch_target_i(22), IN3(21) => branch_target_i(21),
                           IN3(20) => branch_target_i(20), IN3(19) => 
                           branch_target_i(19), IN3(18) => branch_target_i(18),
                           IN3(17) => branch_target_i(17), IN3(16) => 
                           branch_target_i(16), IN3(15) => branch_target_i(15),
                           IN3(14) => branch_target_i(14), IN3(13) => 
                           branch_target_i(13), IN3(12) => branch_target_i(12),
                           IN3(11) => branch_target_i(11), IN3(10) => 
                           branch_target_i(10), IN3(9) => branch_target_i(9), 
                           IN3(8) => branch_target_i(8), IN3(7) => 
                           branch_target_i(7), IN3(6) => branch_target_i(6), 
                           IN3(5) => branch_target_i(5), IN3(4) => 
                           branch_target_i(4), IN3(3) => branch_target_i(3), 
                           IN3(2) => branch_target_i(2), IN3(1) => 
                           branch_target_i(1), IN3(0) => branch_target_i(0), 
                           CTRL(1) => S_MUX_PC_BUS_i(1), CTRL(0) => 
                           S_MUX_PC_BUS_i(0), OUT1(31) => 
                           PC_BUS_pre_BTB_31_port, OUT1(30) => 
                           PC_BUS_pre_BTB_30_port, OUT1(29) => n4, OUT1(28) => 
                           n5, OUT1(27) => PC_BUS_pre_BTB_27_port, OUT1(26) => 
                           PC_BUS_pre_BTB_26_port, OUT1(25) => 
                           PC_BUS_pre_BTB_25_port, OUT1(24) => 
                           PC_BUS_pre_BTB_24_port, OUT1(23) => 
                           PC_BUS_pre_BTB_23_port, OUT1(22) => 
                           PC_BUS_pre_BTB_22_port, OUT1(21) => 
                           PC_BUS_pre_BTB_21_port, OUT1(20) => 
                           PC_BUS_pre_BTB_20_port, OUT1(19) => 
                           PC_BUS_pre_BTB_19_port, OUT1(18) => 
                           PC_BUS_pre_BTB_18_port, OUT1(17) => 
                           PC_BUS_pre_BTB_17_port, OUT1(16) => 
                           PC_BUS_pre_BTB_16_port, OUT1(15) => 
                           PC_BUS_pre_BTB_15_port, OUT1(14) => 
                           PC_BUS_pre_BTB_14_port, OUT1(13) => 
                           PC_BUS_pre_BTB_13_port, OUT1(12) => 
                           PC_BUS_pre_BTB_12_port, OUT1(11) => 
                           PC_BUS_pre_BTB_11_port, OUT1(10) => 
                           PC_BUS_pre_BTB_10_port, OUT1(9) => 
                           PC_BUS_pre_BTB_9_port, OUT1(8) => 
                           PC_BUS_pre_BTB_8_port, OUT1(7) => 
                           PC_BUS_pre_BTB_7_port, OUT1(6) => 
                           PC_BUS_pre_BTB_6_port, OUT1(5) => 
                           PC_BUS_pre_BTB_5_port, OUT1(4) => 
                           PC_BUS_pre_BTB_4_port, OUT1(3) => 
                           PC_BUS_pre_BTB_3_port, OUT1(2) => 
                           PC_BUS_pre_BTB_2_port, OUT1(1) => 
                           PC_BUS_pre_BTB_1_port, OUT1(0) => 
                           PC_BUS_pre_BTB_0_port);
   MUXPREDICTION : mux41_1 port map( IN0(31) => PC4_o_31_port, IN0(30) => 
                           PC4_o_30_port, IN0(29) => PC4_o_29_port, IN0(28) => 
                           PC4_o_28_port, IN0(27) => PC4_o_27_port, IN0(26) => 
                           PC4_o_26_port, IN0(25) => PC4_o_25_port, IN0(24) => 
                           PC4_o_24_port, IN0(23) => PC4_o_23_port, IN0(22) => 
                           PC4_o_22_port, IN0(21) => PC4_o_21_port, IN0(20) => 
                           PC4_o_20_port, IN0(19) => PC4_o_19_port, IN0(18) => 
                           PC4_o_18_port, IN0(17) => PC4_o_17_port, IN0(16) => 
                           PC4_o_16_port, IN0(15) => PC4_o_15_port, IN0(14) => 
                           PC4_o_14_port, IN0(13) => PC4_o_13_port, IN0(12) => 
                           PC4_o_12_port, IN0(11) => PC4_o_11_port, IN0(10) => 
                           PC4_o_10_port, IN0(9) => PC4_o_9_port, IN0(8) => 
                           PC4_o_8_port, IN0(7) => PC4_o_7_port, IN0(6) => 
                           PC4_o_6_port, IN0(5) => PC4_o_5_port, IN0(4) => 
                           PC4_o_4_port, IN0(3) => PC4_o_3_port, IN0(2) => 
                           PC4_o_2_port, IN0(1) => PC4_o_1_port, IN0(0) => 
                           PC4_o_0_port, IN1(31) => predicted_PC(31), IN1(30) 
                           => predicted_PC(30), IN1(29) => predicted_PC(29), 
                           IN1(28) => predicted_PC(28), IN1(27) => 
                           predicted_PC(27), IN1(26) => predicted_PC(26), 
                           IN1(25) => predicted_PC(25), IN1(24) => 
                           predicted_PC(24), IN1(23) => predicted_PC(23), 
                           IN1(22) => predicted_PC(22), IN1(21) => 
                           predicted_PC(21), IN1(20) => predicted_PC(20), 
                           IN1(19) => predicted_PC(19), IN1(18) => 
                           predicted_PC(18), IN1(17) => predicted_PC(17), 
                           IN1(16) => predicted_PC(16), IN1(15) => 
                           predicted_PC(15), IN1(14) => predicted_PC(14), 
                           IN1(13) => predicted_PC(13), IN1(12) => 
                           predicted_PC(12), IN1(11) => predicted_PC(11), 
                           IN1(10) => predicted_PC(10), IN1(9) => 
                           predicted_PC(9), IN1(8) => predicted_PC(8), IN1(7) 
                           => predicted_PC(7), IN1(6) => predicted_PC(6), 
                           IN1(5) => predicted_PC(5), IN1(4) => predicted_PC(4)
                           , IN1(3) => predicted_PC(3), IN1(2) => 
                           predicted_PC(2), IN1(1) => predicted_PC(1), IN1(0) 
                           => predicted_PC(0), IN2(31) => 
                           PC_BUS_pre_BTB_31_port, IN2(30) => 
                           PC_BUS_pre_BTB_30_port, IN2(29) => 
                           PC_BUS_pre_BTB_29_port, IN2(28) => 
                           PC_BUS_pre_BTB_28_port, IN2(27) => 
                           PC_BUS_pre_BTB_27_port, IN2(26) => 
                           PC_BUS_pre_BTB_26_port, IN2(25) => 
                           PC_BUS_pre_BTB_25_port, IN2(24) => 
                           PC_BUS_pre_BTB_24_port, IN2(23) => 
                           PC_BUS_pre_BTB_23_port, IN2(22) => 
                           PC_BUS_pre_BTB_22_port, IN2(21) => 
                           PC_BUS_pre_BTB_21_port, IN2(20) => 
                           PC_BUS_pre_BTB_20_port, IN2(19) => 
                           PC_BUS_pre_BTB_19_port, IN2(18) => 
                           PC_BUS_pre_BTB_18_port, IN2(17) => 
                           PC_BUS_pre_BTB_17_port, IN2(16) => 
                           PC_BUS_pre_BTB_16_port, IN2(15) => 
                           PC_BUS_pre_BTB_15_port, IN2(14) => 
                           PC_BUS_pre_BTB_14_port, IN2(13) => 
                           PC_BUS_pre_BTB_13_port, IN2(12) => 
                           PC_BUS_pre_BTB_12_port, IN2(11) => 
                           PC_BUS_pre_BTB_11_port, IN2(10) => 
                           PC_BUS_pre_BTB_10_port, IN2(9) => 
                           PC_BUS_pre_BTB_9_port, IN2(8) => 
                           PC_BUS_pre_BTB_8_port, IN2(7) => 
                           PC_BUS_pre_BTB_7_port, IN2(6) => 
                           PC_BUS_pre_BTB_6_port, IN2(5) => 
                           PC_BUS_pre_BTB_5_port, IN2(4) => 
                           PC_BUS_pre_BTB_4_port, IN2(3) => 
                           PC_BUS_pre_BTB_3_port, IN2(2) => 
                           PC_BUS_pre_BTB_2_port, IN2(1) => 
                           PC_BUS_pre_BTB_1_port, IN2(0) => 
                           PC_BUS_pre_BTB_0_port, IN3(31) => 
                           PC_BUS_pre_BTB_31_port, IN3(30) => 
                           PC_BUS_pre_BTB_30_port, IN3(29) => 
                           PC_BUS_pre_BTB_29_port, IN3(28) => 
                           PC_BUS_pre_BTB_28_port, IN3(27) => 
                           PC_BUS_pre_BTB_27_port, IN3(26) => 
                           PC_BUS_pre_BTB_26_port, IN3(25) => 
                           PC_BUS_pre_BTB_25_port, IN3(24) => 
                           PC_BUS_pre_BTB_24_port, IN3(23) => 
                           PC_BUS_pre_BTB_23_port, IN3(22) => 
                           PC_BUS_pre_BTB_22_port, IN3(21) => 
                           PC_BUS_pre_BTB_21_port, IN3(20) => 
                           PC_BUS_pre_BTB_20_port, IN3(19) => 
                           PC_BUS_pre_BTB_19_port, IN3(18) => 
                           PC_BUS_pre_BTB_18_port, IN3(17) => 
                           PC_BUS_pre_BTB_17_port, IN3(16) => 
                           PC_BUS_pre_BTB_16_port, IN3(15) => 
                           PC_BUS_pre_BTB_15_port, IN3(14) => 
                           PC_BUS_pre_BTB_14_port, IN3(13) => 
                           PC_BUS_pre_BTB_13_port, IN3(12) => 
                           PC_BUS_pre_BTB_12_port, IN3(11) => 
                           PC_BUS_pre_BTB_11_port, IN3(10) => 
                           PC_BUS_pre_BTB_10_port, IN3(9) => 
                           PC_BUS_pre_BTB_9_port, IN3(8) => 
                           PC_BUS_pre_BTB_8_port, IN3(7) => 
                           PC_BUS_pre_BTB_7_port, IN3(6) => 
                           PC_BUS_pre_BTB_6_port, IN3(5) => 
                           PC_BUS_pre_BTB_5_port, IN3(4) => 
                           PC_BUS_pre_BTB_4_port, IN3(3) => 
                           PC_BUS_pre_BTB_3_port, IN3(2) => 
                           PC_BUS_pre_BTB_2_port, IN3(1) => 
                           PC_BUS_pre_BTB_1_port, IN3(0) => 
                           PC_BUS_pre_BTB_0_port, CTRL(1) => mispredict_i, 
                           CTRL(0) => take_prediction_i, OUT1(31) => 
                           PC_BUS_31_port, OUT1(30) => PC_BUS_30_port, OUT1(29)
                           => PC_BUS_29_port, OUT1(28) => PC_BUS_28_port, 
                           OUT1(27) => PC_BUS_27_port, OUT1(26) => 
                           PC_BUS_26_port, OUT1(25) => PC_BUS_25_port, OUT1(24)
                           => PC_BUS_24_port, OUT1(23) => PC_BUS_23_port, 
                           OUT1(22) => PC_BUS_22_port, OUT1(21) => 
                           PC_BUS_21_port, OUT1(20) => PC_BUS_20_port, OUT1(19)
                           => PC_BUS_19_port, OUT1(18) => PC_BUS_18_port, 
                           OUT1(17) => PC_BUS_17_port, OUT1(16) => 
                           PC_BUS_16_port, OUT1(15) => PC_BUS_15_port, OUT1(14)
                           => PC_BUS_14_port, OUT1(13) => PC_BUS_13_port, 
                           OUT1(12) => PC_BUS_12_port, OUT1(11) => 
                           PC_BUS_11_port, OUT1(10) => PC_BUS_10_port, OUT1(9) 
                           => PC_BUS_9_port, OUT1(8) => PC_BUS_8_port, OUT1(7) 
                           => PC_BUS_7_port, OUT1(6) => PC_BUS_6_port, OUT1(5) 
                           => PC_BUS_5_port, OUT1(4) => PC_BUS_4_port, OUT1(3) 
                           => PC_BUS_3_port, OUT1(2) => PC_BUS_2_port, OUT1(1) 
                           => PC_BUS_1_port, OUT1(0) => PC_BUS_0_port);
   U1 : INV_X1 port map( A => stall_i, ZN => en_IR);
   U2 : BUF_X2 port map( A => n4, Z => PC_BUS_pre_BTB_29_port);
   U3 : BUF_X2 port map( A => n5, Z => PC_BUS_pre_BTB_28_port);

end SYN_Struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_level.all;

entity top_level is

   port( clock, rst : in std_logic;  IRAM_Addr_o : out std_logic_vector (31 
         downto 0);  IRAM_Dout_i : in std_logic_vector (31 downto 0);  
         DRAM_Enable_o, DRAM_WR_o : out std_logic;  DRAM_Din_o, DRAM_Addr_o : 
         out std_logic_vector (31 downto 0);  DRAM_Dout_i : in std_logic_vector
         (31 downto 0));

end top_level;

architecture SYN_arch of top_level is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component fw_logic
      port( D1_i, rAdec_i, D2_i, D3_i, rA_i, rB_i : in std_logic_vector (4 
            downto 0);  S_mem_W, S_mem_LOAD, S_wb_W, S_exe_W : in std_logic;  
            S_FWAdec, S_FWA, S_FWB : out std_logic_vector (1 downto 0));
   end component;
   
   component mem_block
      port( X_i, LOAD_i : in std_logic_vector (31 downto 0);  S_MUX_MEM_i : in 
            std_logic;  W_o : out std_logic_vector (31 downto 0));
   end component;
   
   component mem_regs
      port( W_i : in std_logic_vector (31 downto 0);  D3_i : in 
            std_logic_vector (4 downto 0);  W_o : out std_logic_vector (31 
            downto 0);  D3_o : out std_logic_vector (4 downto 0);  clk, rst : 
            in std_logic);
   end component;
   
   component execute_block
      port( IMM_i, A_i : in std_logic_vector (31 downto 0);  rB_i, rC_i : in 
            std_logic_vector (4 downto 0);  MUXED_B_i : in std_logic_vector (31
            downto 0);  S_MUX_ALUIN_i : in std_logic;  FW_X_i, FW_W_i : in 
            std_logic_vector (31 downto 0);  S_FW_A_i, S_FW_B_i : in 
            std_logic_vector (1 downto 0);  muxed_dest : out std_logic_vector 
            (4 downto 0);  muxed_B : out std_logic_vector (31 downto 0);  
            S_MUX_DEST_i : in std_logic_vector (1 downto 0);  OP : in 
            std_logic_vector (0 to 4);  ALUW_i : in std_logic_vector (12 downto
            0);  DOUT : out std_logic_vector (31 downto 0);  stall_o : out 
            std_logic;  Clock, Reset : in std_logic);
   end component;
   
   component execute_regs
      port( X_i, S_i : in std_logic_vector (31 downto 0);  D2_i : in 
            std_logic_vector (4 downto 0);  X_o, S_o : out std_logic_vector (31
            downto 0);  D2_o : out std_logic_vector (4 downto 0);  stall_i, clk
            , rst : in std_logic);
   end component;
   
   component decode_regs
      port( A_i, B_i : in std_logic_vector (31 downto 0);  rA_i, rB_i, rC_i : 
            in std_logic_vector (4 downto 0);  IMM_i : in std_logic_vector (31 
            downto 0);  ALUW_i : in std_logic_vector (12 downto 0);  A_o, B_o :
            out std_logic_vector (31 downto 0);  rA_o, rB_o, rC_o : out 
            std_logic_vector (4 downto 0);  IMM_o : out std_logic_vector (31 
            downto 0);  ALUW_o : out std_logic_vector (12 downto 0);  stall_i, 
            clk, rst : in std_logic);
   end component;
   
   component dlx_regfile
      port( Clk, Rst, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, 
            ADD_RD2 : in std_logic_vector (4 downto 0);  DATAIN : in 
            std_logic_vector (31 downto 0);  OUT1, OUT2 : out std_logic_vector 
            (31 downto 0));
   end component;
   
   component 
      dlx_cu_MICROCODE_MEM_SIZE64_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE13
      port( Clk, Rst : in std_logic;  IR_IN : in std_logic_vector (31 downto 0)
            ;  stall_exe_i, mispredict_i : in std_logic;  D1_i, D2_i : in 
            std_logic_vector (4 downto 0);  S1_LATCH_EN, S2_LATCH_EN, 
            S3_LATCH_EN : out std_logic;  S_MUX_PC_BUS : out std_logic_vector 
            (1 downto 0);  S_EXT, S_EXT_SIGN, S_EQ_NEQ : out std_logic;  
            S_MUX_DEST : out std_logic_vector (1 downto 0);  S_MUX_LINK, 
            S_MUX_MEM, S_MEM_W_R, S_MEM_EN, S_RF_W_wb, S_RF_W_mem, S_RF_W_exe, 
            S_MUX_ALUIN, stall_exe_o, stall_dec_o, stall_fetch_o, stall_btb_o, 
            was_branch_o, was_jmp_o : out std_logic;  ALU_WORD_o : out 
            std_logic_vector (12 downto 0);  ALU_OPCODE : out std_logic_vector 
            (0 to 4));
   end component;
   
   component jump_logic
      port( NPCF_i, IR_i, A_i : in std_logic_vector (31 downto 0);  A_o : out 
            std_logic_vector (31 downto 0);  rA_o, rB_o, rC_o : out 
            std_logic_vector (4 downto 0);  branch_target_o, sum_addr_o, 
            extended_imm : out std_logic_vector (31 downto 0);  taken_o : out 
            std_logic;  FW_X_i, FW_W_i : in std_logic_vector (31 downto 0);  
            S_FW_Adec_i : in std_logic_vector (1 downto 0);  S_EXT_i, 
            S_EXT_SIGN_i, S_MUX_LINK_i, S_EQ_NEQ_i : in std_logic);
   end component;
   
   component fetch_regs
      port( NPCF_i, IR_i : in std_logic_vector (31 downto 0);  NPCF_o, IR_o : 
            out std_logic_vector (31 downto 0);  stall_i, clk, rst : in 
            std_logic);
   end component;
   
   component btb_N_LINES4_SIZE32
      port( clock, reset, stall_i : in std_logic;  TAG_i : in std_logic_vector 
            (3 downto 0);  target_PC_i : in std_logic_vector (31 downto 0);  
            was_taken_i : in std_logic;  predicted_next_PC_o : out 
            std_logic_vector (31 downto 0);  taken_o, mispredict_o : out 
            std_logic);
   end component;
   
   component fetch_block
      port( branch_target_i, sum_addr_i, A_i, NPC4_i : in std_logic_vector (31 
            downto 0);  S_MUX_PC_BUS_i : in std_logic_vector (1 downto 0);  
            PC_o, PC4_o, PC_BUS_pre_BTB : out std_logic_vector (31 downto 0);  
            stall_i, take_prediction_i, mispredict_i : in std_logic;  
            predicted_PC : in std_logic_vector (31 downto 0);  clk, rst : in 
            std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, IRAM_Addr_o_31_port, 
      IRAM_Addr_o_30_port, IRAM_Addr_o_29_port, IRAM_Addr_o_28_port, 
      IRAM_Addr_o_27_port, IRAM_Addr_o_26_port, IRAM_Addr_o_25_port, 
      IRAM_Addr_o_24_port, IRAM_Addr_o_23_port, IRAM_Addr_o_22_port, 
      IRAM_Addr_o_21_port, IRAM_Addr_o_20_port, IRAM_Addr_o_19_port, 
      IRAM_Addr_o_18_port, IRAM_Addr_o_17_port, IRAM_Addr_o_16_port, 
      IRAM_Addr_o_15_port, IRAM_Addr_o_14_port, IRAM_Addr_o_13_port, 
      IRAM_Addr_o_12_port, IRAM_Addr_o_11_port, IRAM_Addr_o_10_port, 
      IRAM_Addr_o_9_port, IRAM_Addr_o_8_port, IRAM_Addr_o_7_port, 
      IRAM_Addr_o_6_port, IRAM_Addr_o_5_port, IRAM_Addr_o_4_port, 
      IRAM_Addr_o_3_port, IRAM_Addr_o_2_port, IRAM_Addr_o_1_port, 
      IRAM_Addr_o_0_port, DRAM_Addr_o_31_port, DRAM_Addr_o_30_port, 
      DRAM_Addr_o_29_port, DRAM_Addr_o_28_port, DRAM_Addr_o_27_port, 
      DRAM_Addr_o_26_port, DRAM_Addr_o_25_port, DRAM_Addr_o_24_port, 
      DRAM_Addr_o_23_port, DRAM_Addr_o_22_port, DRAM_Addr_o_21_port, 
      DRAM_Addr_o_20_port, DRAM_Addr_o_19_port, DRAM_Addr_o_18_port, 
      DRAM_Addr_o_17_port, DRAM_Addr_o_16_port, DRAM_Addr_o_15_port, 
      DRAM_Addr_o_14_port, DRAM_Addr_o_13_port, DRAM_Addr_o_12_port, 
      DRAM_Addr_o_11_port, DRAM_Addr_o_10_port, DRAM_Addr_o_9_port, 
      DRAM_Addr_o_8_port, DRAM_Addr_o_7_port, DRAM_Addr_o_6_port, 
      DRAM_Addr_o_5_port, DRAM_Addr_o_4_port, DRAM_Addr_o_3_port, 
      DRAM_Addr_o_2_port, DRAM_Addr_o_1_port, DRAM_Addr_o_0_port, 
      was_taken_from_jl, was_branch, was_jmp, was_taken, 
      dummy_branch_target_31_port, dummy_branch_target_30_port, 
      dummy_branch_target_29_port, dummy_branch_target_28_port, 
      dummy_branch_target_27_port, dummy_branch_target_26_port, 
      dummy_branch_target_25_port, dummy_branch_target_24_port, 
      dummy_branch_target_23_port, dummy_branch_target_22_port, 
      dummy_branch_target_21_port, dummy_branch_target_20_port, 
      dummy_branch_target_19_port, dummy_branch_target_18_port, 
      dummy_branch_target_17_port, dummy_branch_target_16_port, 
      dummy_branch_target_15_port, dummy_branch_target_14_port, 
      dummy_branch_target_13_port, dummy_branch_target_12_port, 
      dummy_branch_target_11_port, dummy_branch_target_10_port, 
      dummy_branch_target_9_port, dummy_branch_target_8_port, 
      dummy_branch_target_7_port, dummy_branch_target_6_port, 
      dummy_branch_target_5_port, dummy_branch_target_4_port, 
      dummy_branch_target_3_port, dummy_branch_target_2_port, 
      dummy_branch_target_1_port, dummy_branch_target_0_port, 
      dummy_sum_addr_31_port, dummy_sum_addr_30_port, dummy_sum_addr_29_port, 
      dummy_sum_addr_28_port, dummy_sum_addr_27_port, dummy_sum_addr_26_port, 
      dummy_sum_addr_25_port, dummy_sum_addr_24_port, dummy_sum_addr_23_port, 
      dummy_sum_addr_22_port, dummy_sum_addr_21_port, dummy_sum_addr_20_port, 
      dummy_sum_addr_19_port, dummy_sum_addr_18_port, dummy_sum_addr_17_port, 
      dummy_sum_addr_16_port, dummy_sum_addr_15_port, dummy_sum_addr_14_port, 
      dummy_sum_addr_13_port, dummy_sum_addr_12_port, dummy_sum_addr_11_port, 
      dummy_sum_addr_10_port, dummy_sum_addr_9_port, dummy_sum_addr_8_port, 
      dummy_sum_addr_7_port, dummy_sum_addr_6_port, dummy_sum_addr_5_port, 
      dummy_sum_addr_4_port, dummy_sum_addr_3_port, dummy_sum_addr_2_port, 
      dummy_sum_addr_1_port, dummy_sum_addr_0_port, dummy_A_31_port, 
      dummy_A_30_port, dummy_A_29_port, dummy_A_28_port, dummy_A_27_port, 
      dummy_A_26_port, dummy_A_25_port, dummy_A_24_port, dummy_A_23_port, 
      dummy_A_22_port, dummy_A_21_port, dummy_A_20_port, dummy_A_19_port, 
      dummy_A_18_port, dummy_A_17_port, dummy_A_16_port, dummy_A_15_port, 
      dummy_A_14_port, dummy_A_13_port, dummy_A_12_port, dummy_A_11_port, 
      dummy_A_10_port, dummy_A_9_port, dummy_A_8_port, dummy_A_7_port, 
      dummy_A_6_port, dummy_A_5_port, dummy_A_4_port, dummy_A_3_port, 
      dummy_A_2_port, dummy_A_1_port, dummy_A_0_port, NPCF_31_port, 
      NPCF_30_port, NPCF_29_port, NPCF_28_port, NPCF_27_port, NPCF_26_port, 
      NPCF_25_port, NPCF_24_port, NPCF_23_port, NPCF_22_port, NPCF_21_port, 
      NPCF_20_port, NPCF_19_port, NPCF_18_port, NPCF_17_port, NPCF_16_port, 
      NPCF_15_port, NPCF_14_port, NPCF_13_port, NPCF_12_port, NPCF_11_port, 
      NPCF_10_port, NPCF_9_port, NPCF_8_port, NPCF_7_port, NPCF_6_port, 
      NPCF_5_port, NPCF_4_port, NPCF_3_port, NPCF_2_port, NPCF_1_port, 
      NPCF_0_port, dummy_S_MUX_PC_BUS_1_port, dummy_S_MUX_PC_BUS_0_port, 
      PC4_31_port, PC4_30_port, PC4_29_port, PC4_28_port, PC4_27_port, 
      PC4_26_port, PC4_25_port, PC4_24_port, PC4_23_port, PC4_22_port, 
      PC4_21_port, PC4_20_port, PC4_19_port, PC4_18_port, PC4_17_port, 
      PC4_16_port, PC4_15_port, PC4_14_port, PC4_13_port, PC4_12_port, 
      PC4_11_port, PC4_10_port, PC4_9_port, PC4_8_port, PC4_7_port, PC4_6_port,
      PC4_5_port, PC4_4_port, PC4_3_port, PC4_2_port, PC4_1_port, PC4_0_port, 
      TARGET_PC_31_port, TARGET_PC_30_port, TARGET_PC_29_port, 
      TARGET_PC_28_port, TARGET_PC_27_port, TARGET_PC_26_port, 
      TARGET_PC_25_port, TARGET_PC_24_port, TARGET_PC_23_port, 
      TARGET_PC_22_port, TARGET_PC_21_port, TARGET_PC_20_port, 
      TARGET_PC_19_port, TARGET_PC_18_port, TARGET_PC_17_port, 
      TARGET_PC_16_port, TARGET_PC_15_port, TARGET_PC_14_port, 
      TARGET_PC_13_port, TARGET_PC_12_port, TARGET_PC_11_port, 
      TARGET_PC_10_port, TARGET_PC_9_port, TARGET_PC_8_port, TARGET_PC_7_port, 
      TARGET_PC_6_port, TARGET_PC_5_port, TARGET_PC_4_port, TARGET_PC_3_port, 
      TARGET_PC_2_port, TARGET_PC_1_port, TARGET_PC_0_port, stall_fetch, 
      take_prediction, predicted_PC_31_port, predicted_PC_30_port, 
      predicted_PC_29_port, predicted_PC_28_port, predicted_PC_27_port, 
      predicted_PC_26_port, predicted_PC_25_port, predicted_PC_24_port, 
      predicted_PC_23_port, predicted_PC_22_port, predicted_PC_21_port, 
      predicted_PC_20_port, predicted_PC_19_port, predicted_PC_18_port, 
      predicted_PC_17_port, predicted_PC_16_port, predicted_PC_15_port, 
      predicted_PC_14_port, predicted_PC_13_port, predicted_PC_12_port, 
      predicted_PC_11_port, predicted_PC_10_port, predicted_PC_9_port, 
      predicted_PC_8_port, predicted_PC_7_port, predicted_PC_6_port, 
      predicted_PC_5_port, predicted_PC_4_port, predicted_PC_3_port, 
      predicted_PC_2_port, predicted_PC_1_port, predicted_PC_0_port, stall_btb,
      IR_31_port, IR_30_port, IR_29_port, IR_28_port, IR_27_port, IR_26_port, 
      IR_25_port, IR_24_port, IR_23_port, IR_22_port, IR_21_port, IR_20_port, 
      IR_19_port, IR_18_port, IR_17_port, IR_16_port, IR_15_port, IR_14_port, 
      IR_13_port, IR_12_port, IR_11_port, IR_10_port, IR_9_port, IR_8_port, 
      IR_7_port, IR_6_port, IR_5_port, IR_4_port, IR_3_port, IR_2_port, 
      IR_1_port, IR_0_port, stall_decode, AtoComp_31_port, AtoComp_30_port, 
      AtoComp_29_port, AtoComp_28_port, AtoComp_27_port, AtoComp_26_port, 
      AtoComp_25_port, AtoComp_24_port, AtoComp_23_port, AtoComp_22_port, 
      AtoComp_21_port, AtoComp_20_port, AtoComp_19_port, AtoComp_18_port, 
      AtoComp_17_port, AtoComp_16_port, AtoComp_15_port, AtoComp_14_port, 
      AtoComp_13_port, AtoComp_12_port, AtoComp_11_port, AtoComp_10_port, 
      AtoComp_9_port, AtoComp_8_port, AtoComp_7_port, AtoComp_6_port, 
      AtoComp_5_port, AtoComp_4_port, AtoComp_3_port, AtoComp_2_port, 
      AtoComp_1_port, AtoComp_0_port, rA2reg_4_port, rA2reg_3_port, 
      rA2reg_2_port, rA2reg_1_port, rA2reg_0_port, rB2reg_4_port, rB2reg_3_port
      , rB2reg_2_port, rB2reg_1_port, rB2reg_0_port, rC2reg_4_port, 
      rC2reg_3_port, rC2reg_2_port, rC2reg_1_port, rC2reg_0_port, 
      help_IMM_31_port, help_IMM_30_port, help_IMM_29_port, help_IMM_28_port, 
      help_IMM_27_port, help_IMM_26_port, help_IMM_25_port, help_IMM_24_port, 
      help_IMM_23_port, help_IMM_22_port, help_IMM_21_port, help_IMM_20_port, 
      help_IMM_19_port, help_IMM_18_port, help_IMM_17_port, help_IMM_16_port, 
      help_IMM_15_port, help_IMM_14_port, help_IMM_13_port, help_IMM_12_port, 
      help_IMM_11_port, help_IMM_10_port, help_IMM_9_port, help_IMM_8_port, 
      help_IMM_7_port, help_IMM_6_port, help_IMM_5_port, help_IMM_4_port, 
      help_IMM_3_port, help_IMM_2_port, help_IMM_1_port, help_IMM_0_port, 
      wb2reg_31_port, wb2reg_30_port, wb2reg_29_port, wb2reg_28_port, 
      wb2reg_27_port, wb2reg_26_port, wb2reg_25_port, wb2reg_24_port, 
      wb2reg_23_port, wb2reg_22_port, wb2reg_21_port, wb2reg_20_port, 
      wb2reg_19_port, wb2reg_18_port, wb2reg_17_port, wb2reg_16_port, 
      wb2reg_15_port, wb2reg_14_port, wb2reg_13_port, wb2reg_12_port, 
      wb2reg_11_port, wb2reg_10_port, wb2reg_9_port, wb2reg_8_port, 
      wb2reg_7_port, wb2reg_6_port, wb2reg_5_port, wb2reg_4_port, wb2reg_3_port
      , wb2reg_2_port, wb2reg_1_port, wb2reg_0_port, dummy_S_FWAdec_1_port, 
      dummy_S_FWAdec_0_port, dummy_S_EXT, dummy_S_EXT_SIGN, dummy_S_EQ_NEQ, 
      exe_stall_cu, muxed_dest2exe_4_port, muxed_dest2exe_3_port, 
      muxed_dest2exe_2_port, muxed_dest2exe_1_port, muxed_dest2exe_0_port, 
      D22D3_4_port, D22D3_3_port, D22D3_2_port, D22D3_1_port, D22D3_0_port, 
      dummy_S_MUX_DEST_1_port, dummy_S_MUX_DEST_0_port, dummy_S_MUX_MEM, 
      dummy_S_RF_W_wb, dummy_S_RF_W_mem, dummy_S_MUX_ALUIN, stall_exe, 
      ALUW_dec_12_port, ALUW_dec_11_port, ALUW_dec_10_port, ALUW_dec_9_port, 
      ALUW_dec_8_port, ALUW_dec_7_port, ALUW_dec_6_port, ALUW_dec_5_port, 
      ALUW_dec_4_port, ALUW_dec_3_port, ALUW_dec_2_port, ALUW_dec_1_port, 
      ALUW_dec_0_port, enable_regfile, W2wb_31_port, W2wb_30_port, W2wb_29_port
      , W2wb_28_port, W2wb_27_port, W2wb_26_port, W2wb_25_port, W2wb_24_port, 
      W2wb_23_port, W2wb_22_port, W2wb_21_port, W2wb_20_port, W2wb_19_port, 
      W2wb_18_port, W2wb_17_port, W2wb_16_port, W2wb_15_port, W2wb_14_port, 
      W2wb_13_port, W2wb_12_port, W2wb_11_port, W2wb_10_port, W2wb_9_port, 
      W2wb_8_port, W2wb_7_port, W2wb_6_port, W2wb_5_port, W2wb_4_port, 
      W2wb_3_port, W2wb_2_port, W2wb_1_port, W2wb_0_port, dummy_B_31_port, 
      dummy_B_30_port, dummy_B_29_port, dummy_B_28_port, dummy_B_27_port, 
      dummy_B_26_port, dummy_B_25_port, dummy_B_24_port, dummy_B_23_port, 
      dummy_B_22_port, dummy_B_21_port, dummy_B_20_port, dummy_B_19_port, 
      dummy_B_18_port, dummy_B_17_port, dummy_B_16_port, dummy_B_15_port, 
      dummy_B_14_port, dummy_B_13_port, dummy_B_12_port, dummy_B_11_port, 
      dummy_B_10_port, dummy_B_9_port, dummy_B_8_port, dummy_B_7_port, 
      dummy_B_6_port, dummy_B_5_port, dummy_B_4_port, dummy_B_3_port, 
      dummy_B_2_port, dummy_B_1_port, dummy_B_0_port, A2exe_31_port, 
      A2exe_30_port, A2exe_29_port, A2exe_28_port, A2exe_27_port, A2exe_26_port
      , A2exe_25_port, A2exe_24_port, A2exe_23_port, A2exe_22_port, 
      A2exe_21_port, A2exe_20_port, A2exe_19_port, A2exe_18_port, A2exe_17_port
      , A2exe_16_port, A2exe_15_port, A2exe_14_port, A2exe_13_port, 
      A2exe_12_port, A2exe_11_port, A2exe_10_port, A2exe_9_port, A2exe_8_port, 
      A2exe_7_port, A2exe_6_port, A2exe_5_port, A2exe_4_port, A2exe_3_port, 
      A2exe_2_port, A2exe_1_port, A2exe_0_port, B2exe_31_port, B2exe_30_port, 
      B2exe_29_port, B2exe_28_port, B2exe_27_port, B2exe_26_port, B2exe_25_port
      , B2exe_24_port, B2exe_23_port, B2exe_22_port, B2exe_21_port, 
      B2exe_20_port, B2exe_19_port, B2exe_18_port, B2exe_17_port, B2exe_16_port
      , B2exe_15_port, B2exe_14_port, B2exe_13_port, B2exe_12_port, 
      B2exe_11_port, B2exe_10_port, B2exe_9_port, B2exe_8_port, B2exe_7_port, 
      B2exe_6_port, B2exe_5_port, B2exe_4_port, B2exe_3_port, B2exe_2_port, 
      B2exe_1_port, B2exe_0_port, rA2fw_4_port, rA2fw_3_port, rA2fw_2_port, 
      rA2fw_1_port, rA2fw_0_port, rB2mux_4_port, rB2mux_3_port, rB2mux_2_port, 
      rB2mux_1_port, rB2mux_0_port, rC2mux_4_port, rC2mux_3_port, rC2mux_2_port
      , rC2mux_1_port, rC2mux_0_port, IMM2exe_31_port, IMM2exe_30_port, 
      IMM2exe_29_port, IMM2exe_28_port, IMM2exe_27_port, IMM2exe_26_port, 
      IMM2exe_25_port, IMM2exe_24_port, IMM2exe_23_port, IMM2exe_22_port, 
      IMM2exe_21_port, IMM2exe_20_port, IMM2exe_19_port, IMM2exe_18_port, 
      IMM2exe_17_port, IMM2exe_16_port, IMM2exe_15_port, IMM2exe_14_port, 
      IMM2exe_13_port, IMM2exe_12_port, IMM2exe_11_port, IMM2exe_10_port, 
      IMM2exe_9_port, IMM2exe_8_port, IMM2exe_7_port, IMM2exe_6_port, 
      IMM2exe_5_port, IMM2exe_4_port, IMM2exe_3_port, IMM2exe_2_port, 
      IMM2exe_1_port, IMM2exe_0_port, ALUW_12_port, ALUW_11_port, ALUW_10_port,
      ALUW_9_port, ALUW_8_port, ALUW_7_port, ALUW_6_port, ALUW_5_port, 
      ALUW_4_port, ALUW_3_port, ALUW_2_port, ALUW_1_port, ALUW_0_port, 
      X2mem_31_port, X2mem_30_port, X2mem_29_port, X2mem_28_port, X2mem_27_port
      , X2mem_26_port, X2mem_25_port, X2mem_24_port, X2mem_23_port, 
      X2mem_22_port, X2mem_21_port, X2mem_20_port, X2mem_19_port, X2mem_18_port
      , X2mem_17_port, X2mem_16_port, X2mem_15_port, X2mem_14_port, 
      X2mem_13_port, X2mem_12_port, X2mem_11_port, X2mem_10_port, X2mem_9_port,
      X2mem_8_port, X2mem_7_port, X2mem_6_port, X2mem_5_port, X2mem_4_port, 
      X2mem_3_port, X2mem_2_port, X2mem_1_port, X2mem_0_port, S2mem_31_port, 
      S2mem_30_port, S2mem_29_port, S2mem_28_port, S2mem_27_port, S2mem_26_port
      , S2mem_25_port, S2mem_24_port, S2mem_23_port, S2mem_22_port, 
      S2mem_21_port, S2mem_20_port, S2mem_19_port, S2mem_18_port, S2mem_17_port
      , S2mem_16_port, S2mem_15_port, S2mem_14_port, S2mem_13_port, 
      S2mem_12_port, S2mem_11_port, S2mem_10_port, S2mem_9_port, S2mem_8_port, 
      S2mem_7_port, S2mem_6_port, S2mem_5_port, S2mem_4_port, S2mem_2_port, 
      S2mem_1_port, S2mem_0_port, dummy_S_FWA2exe_1_port, 
      dummy_S_FWA2exe_0_port, dummy_S_FWB2exe_1_port, dummy_S_FWB2exe_0_port, 
      D32reg_4_port, D32reg_3_port, D32reg_2_port, D32reg_1_port, D32reg_0_port
      , n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18
      , n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, 
      n33, net244538, net244539, net244540, net244541, net244542, net244543, 
      net244544, net244545, net244546 : std_logic;

begin
   IRAM_Addr_o <= ( IRAM_Addr_o_31_port, IRAM_Addr_o_30_port, 
      IRAM_Addr_o_29_port, IRAM_Addr_o_28_port, IRAM_Addr_o_27_port, 
      IRAM_Addr_o_26_port, IRAM_Addr_o_25_port, IRAM_Addr_o_24_port, 
      IRAM_Addr_o_23_port, IRAM_Addr_o_22_port, IRAM_Addr_o_21_port, 
      IRAM_Addr_o_20_port, IRAM_Addr_o_19_port, IRAM_Addr_o_18_port, 
      IRAM_Addr_o_17_port, IRAM_Addr_o_16_port, IRAM_Addr_o_15_port, 
      IRAM_Addr_o_14_port, IRAM_Addr_o_13_port, IRAM_Addr_o_12_port, 
      IRAM_Addr_o_11_port, IRAM_Addr_o_10_port, IRAM_Addr_o_9_port, 
      IRAM_Addr_o_8_port, IRAM_Addr_o_7_port, IRAM_Addr_o_6_port, 
      IRAM_Addr_o_5_port, IRAM_Addr_o_4_port, IRAM_Addr_o_3_port, 
      IRAM_Addr_o_2_port, IRAM_Addr_o_1_port, IRAM_Addr_o_0_port );
   DRAM_Addr_o <= ( DRAM_Addr_o_31_port, DRAM_Addr_o_30_port, 
      DRAM_Addr_o_29_port, DRAM_Addr_o_28_port, DRAM_Addr_o_27_port, 
      DRAM_Addr_o_26_port, DRAM_Addr_o_25_port, DRAM_Addr_o_24_port, 
      DRAM_Addr_o_23_port, DRAM_Addr_o_22_port, DRAM_Addr_o_21_port, 
      DRAM_Addr_o_20_port, DRAM_Addr_o_19_port, DRAM_Addr_o_18_port, 
      DRAM_Addr_o_17_port, DRAM_Addr_o_16_port, DRAM_Addr_o_15_port, 
      DRAM_Addr_o_14_port, DRAM_Addr_o_13_port, DRAM_Addr_o_12_port, 
      DRAM_Addr_o_11_port, DRAM_Addr_o_10_port, DRAM_Addr_o_9_port, 
      DRAM_Addr_o_8_port, DRAM_Addr_o_7_port, DRAM_Addr_o_6_port, 
      DRAM_Addr_o_5_port, DRAM_Addr_o_4_port, DRAM_Addr_o_3_port, 
      DRAM_Addr_o_2_port, DRAM_Addr_o_1_port, DRAM_Addr_o_0_port );
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   UFETCH_BLOCK : fetch_block port map( branch_target_i(31) => 
                           dummy_branch_target_31_port, branch_target_i(30) => 
                           dummy_branch_target_30_port, branch_target_i(29) => 
                           dummy_branch_target_29_port, branch_target_i(28) => 
                           dummy_branch_target_28_port, branch_target_i(27) => 
                           dummy_branch_target_27_port, branch_target_i(26) => 
                           dummy_branch_target_26_port, branch_target_i(25) => 
                           dummy_branch_target_25_port, branch_target_i(24) => 
                           dummy_branch_target_24_port, branch_target_i(23) => 
                           dummy_branch_target_23_port, branch_target_i(22) => 
                           dummy_branch_target_22_port, branch_target_i(21) => 
                           dummy_branch_target_21_port, branch_target_i(20) => 
                           dummy_branch_target_20_port, branch_target_i(19) => 
                           dummy_branch_target_19_port, branch_target_i(18) => 
                           dummy_branch_target_18_port, branch_target_i(17) => 
                           dummy_branch_target_17_port, branch_target_i(16) => 
                           dummy_branch_target_16_port, branch_target_i(15) => 
                           dummy_branch_target_15_port, branch_target_i(14) => 
                           dummy_branch_target_14_port, branch_target_i(13) => 
                           dummy_branch_target_13_port, branch_target_i(12) => 
                           dummy_branch_target_12_port, branch_target_i(11) => 
                           dummy_branch_target_11_port, branch_target_i(10) => 
                           dummy_branch_target_10_port, branch_target_i(9) => 
                           dummy_branch_target_9_port, branch_target_i(8) => 
                           dummy_branch_target_8_port, branch_target_i(7) => 
                           dummy_branch_target_7_port, branch_target_i(6) => 
                           dummy_branch_target_6_port, branch_target_i(5) => 
                           dummy_branch_target_5_port, branch_target_i(4) => 
                           dummy_branch_target_4_port, branch_target_i(3) => 
                           dummy_branch_target_3_port, branch_target_i(2) => 
                           dummy_branch_target_2_port, branch_target_i(1) => 
                           dummy_branch_target_1_port, branch_target_i(0) => 
                           dummy_branch_target_0_port, sum_addr_i(31) => 
                           dummy_sum_addr_31_port, sum_addr_i(30) => 
                           dummy_sum_addr_30_port, sum_addr_i(29) => 
                           dummy_sum_addr_29_port, sum_addr_i(28) => 
                           dummy_sum_addr_28_port, sum_addr_i(27) => 
                           dummy_sum_addr_27_port, sum_addr_i(26) => 
                           dummy_sum_addr_26_port, sum_addr_i(25) => 
                           dummy_sum_addr_25_port, sum_addr_i(24) => 
                           dummy_sum_addr_24_port, sum_addr_i(23) => 
                           dummy_sum_addr_23_port, sum_addr_i(22) => 
                           dummy_sum_addr_22_port, sum_addr_i(21) => 
                           dummy_sum_addr_21_port, sum_addr_i(20) => 
                           dummy_sum_addr_20_port, sum_addr_i(19) => 
                           dummy_sum_addr_19_port, sum_addr_i(18) => 
                           dummy_sum_addr_18_port, sum_addr_i(17) => 
                           dummy_sum_addr_17_port, sum_addr_i(16) => 
                           dummy_sum_addr_16_port, sum_addr_i(15) => 
                           dummy_sum_addr_15_port, sum_addr_i(14) => 
                           dummy_sum_addr_14_port, sum_addr_i(13) => 
                           dummy_sum_addr_13_port, sum_addr_i(12) => 
                           dummy_sum_addr_12_port, sum_addr_i(11) => 
                           dummy_sum_addr_11_port, sum_addr_i(10) => 
                           dummy_sum_addr_10_port, sum_addr_i(9) => 
                           dummy_sum_addr_9_port, sum_addr_i(8) => 
                           dummy_sum_addr_8_port, sum_addr_i(7) => 
                           dummy_sum_addr_7_port, sum_addr_i(6) => 
                           dummy_sum_addr_6_port, sum_addr_i(5) => 
                           dummy_sum_addr_5_port, sum_addr_i(4) => 
                           dummy_sum_addr_4_port, sum_addr_i(3) => 
                           dummy_sum_addr_3_port, sum_addr_i(2) => 
                           dummy_sum_addr_2_port, sum_addr_i(1) => 
                           dummy_sum_addr_1_port, sum_addr_i(0) => 
                           dummy_sum_addr_0_port, A_i(31) => dummy_A_31_port, 
                           A_i(30) => dummy_A_30_port, A_i(29) => 
                           dummy_A_29_port, A_i(28) => dummy_A_28_port, A_i(27)
                           => dummy_A_27_port, A_i(26) => dummy_A_26_port, 
                           A_i(25) => dummy_A_25_port, A_i(24) => 
                           dummy_A_24_port, A_i(23) => dummy_A_23_port, A_i(22)
                           => dummy_A_22_port, A_i(21) => dummy_A_21_port, 
                           A_i(20) => dummy_A_20_port, A_i(19) => 
                           dummy_A_19_port, A_i(18) => dummy_A_18_port, A_i(17)
                           => dummy_A_17_port, A_i(16) => dummy_A_16_port, 
                           A_i(15) => dummy_A_15_port, A_i(14) => 
                           dummy_A_14_port, A_i(13) => dummy_A_13_port, A_i(12)
                           => dummy_A_12_port, A_i(11) => dummy_A_11_port, 
                           A_i(10) => dummy_A_10_port, A_i(9) => dummy_A_9_port
                           , A_i(8) => dummy_A_8_port, A_i(7) => dummy_A_7_port
                           , A_i(6) => dummy_A_6_port, A_i(5) => dummy_A_5_port
                           , A_i(4) => dummy_A_4_port, A_i(3) => dummy_A_3_port
                           , A_i(2) => dummy_A_2_port, A_i(1) => dummy_A_1_port
                           , A_i(0) => dummy_A_0_port, NPC4_i(31) => 
                           NPCF_31_port, NPC4_i(30) => NPCF_30_port, NPC4_i(29)
                           => NPCF_29_port, NPC4_i(28) => NPCF_28_port, 
                           NPC4_i(27) => NPCF_27_port, NPC4_i(26) => 
                           NPCF_26_port, NPC4_i(25) => NPCF_25_port, NPC4_i(24)
                           => NPCF_24_port, NPC4_i(23) => NPCF_23_port, 
                           NPC4_i(22) => NPCF_22_port, NPC4_i(21) => 
                           NPCF_21_port, NPC4_i(20) => NPCF_20_port, NPC4_i(19)
                           => NPCF_19_port, NPC4_i(18) => NPCF_18_port, 
                           NPC4_i(17) => NPCF_17_port, NPC4_i(16) => 
                           NPCF_16_port, NPC4_i(15) => NPCF_15_port, NPC4_i(14)
                           => NPCF_14_port, NPC4_i(13) => NPCF_13_port, 
                           NPC4_i(12) => NPCF_12_port, NPC4_i(11) => 
                           NPCF_11_port, NPC4_i(10) => NPCF_10_port, NPC4_i(9) 
                           => NPCF_9_port, NPC4_i(8) => NPCF_8_port, NPC4_i(7) 
                           => NPCF_7_port, NPC4_i(6) => NPCF_6_port, NPC4_i(5) 
                           => NPCF_5_port, NPC4_i(4) => NPCF_4_port, NPC4_i(3) 
                           => NPCF_3_port, NPC4_i(2) => NPCF_2_port, NPC4_i(1) 
                           => NPCF_1_port, NPC4_i(0) => NPCF_0_port, 
                           S_MUX_PC_BUS_i(1) => dummy_S_MUX_PC_BUS_1_port, 
                           S_MUX_PC_BUS_i(0) => dummy_S_MUX_PC_BUS_0_port, 
                           PC_o(31) => IRAM_Addr_o_31_port, PC_o(30) => 
                           IRAM_Addr_o_30_port, PC_o(29) => IRAM_Addr_o_29_port
                           , PC_o(28) => IRAM_Addr_o_28_port, PC_o(27) => 
                           IRAM_Addr_o_27_port, PC_o(26) => IRAM_Addr_o_26_port
                           , PC_o(25) => IRAM_Addr_o_25_port, PC_o(24) => 
                           IRAM_Addr_o_24_port, PC_o(23) => IRAM_Addr_o_23_port
                           , PC_o(22) => IRAM_Addr_o_22_port, PC_o(21) => 
                           IRAM_Addr_o_21_port, PC_o(20) => IRAM_Addr_o_20_port
                           , PC_o(19) => IRAM_Addr_o_19_port, PC_o(18) => 
                           IRAM_Addr_o_18_port, PC_o(17) => IRAM_Addr_o_17_port
                           , PC_o(16) => IRAM_Addr_o_16_port, PC_o(15) => 
                           IRAM_Addr_o_15_port, PC_o(14) => IRAM_Addr_o_14_port
                           , PC_o(13) => IRAM_Addr_o_13_port, PC_o(12) => 
                           IRAM_Addr_o_12_port, PC_o(11) => IRAM_Addr_o_11_port
                           , PC_o(10) => IRAM_Addr_o_10_port, PC_o(9) => 
                           IRAM_Addr_o_9_port, PC_o(8) => IRAM_Addr_o_8_port, 
                           PC_o(7) => IRAM_Addr_o_7_port, PC_o(6) => 
                           IRAM_Addr_o_6_port, PC_o(5) => IRAM_Addr_o_5_port, 
                           PC_o(4) => IRAM_Addr_o_4_port, PC_o(3) => 
                           IRAM_Addr_o_3_port, PC_o(2) => IRAM_Addr_o_2_port, 
                           PC_o(1) => IRAM_Addr_o_1_port, PC_o(0) => 
                           IRAM_Addr_o_0_port, PC4_o(31) => PC4_31_port, 
                           PC4_o(30) => PC4_30_port, PC4_o(29) => PC4_29_port, 
                           PC4_o(28) => PC4_28_port, PC4_o(27) => PC4_27_port, 
                           PC4_o(26) => PC4_26_port, PC4_o(25) => PC4_25_port, 
                           PC4_o(24) => PC4_24_port, PC4_o(23) => PC4_23_port, 
                           PC4_o(22) => PC4_22_port, PC4_o(21) => PC4_21_port, 
                           PC4_o(20) => PC4_20_port, PC4_o(19) => PC4_19_port, 
                           PC4_o(18) => PC4_18_port, PC4_o(17) => PC4_17_port, 
                           PC4_o(16) => PC4_16_port, PC4_o(15) => PC4_15_port, 
                           PC4_o(14) => PC4_14_port, PC4_o(13) => PC4_13_port, 
                           PC4_o(12) => PC4_12_port, PC4_o(11) => PC4_11_port, 
                           PC4_o(10) => PC4_10_port, PC4_o(9) => PC4_9_port, 
                           PC4_o(8) => PC4_8_port, PC4_o(7) => PC4_7_port, 
                           PC4_o(6) => PC4_6_port, PC4_o(5) => PC4_5_port, 
                           PC4_o(4) => PC4_4_port, PC4_o(3) => PC4_3_port, 
                           PC4_o(2) => PC4_2_port, PC4_o(1) => PC4_1_port, 
                           PC4_o(0) => PC4_0_port, PC_BUS_pre_BTB(31) => 
                           TARGET_PC_31_port, PC_BUS_pre_BTB(30) => 
                           TARGET_PC_30_port, PC_BUS_pre_BTB(29) => 
                           TARGET_PC_29_port, PC_BUS_pre_BTB(28) => 
                           TARGET_PC_28_port, PC_BUS_pre_BTB(27) => 
                           TARGET_PC_27_port, PC_BUS_pre_BTB(26) => 
                           TARGET_PC_26_port, PC_BUS_pre_BTB(25) => 
                           TARGET_PC_25_port, PC_BUS_pre_BTB(24) => 
                           TARGET_PC_24_port, PC_BUS_pre_BTB(23) => 
                           TARGET_PC_23_port, PC_BUS_pre_BTB(22) => 
                           TARGET_PC_22_port, PC_BUS_pre_BTB(21) => 
                           TARGET_PC_21_port, PC_BUS_pre_BTB(20) => 
                           TARGET_PC_20_port, PC_BUS_pre_BTB(19) => 
                           TARGET_PC_19_port, PC_BUS_pre_BTB(18) => 
                           TARGET_PC_18_port, PC_BUS_pre_BTB(17) => 
                           TARGET_PC_17_port, PC_BUS_pre_BTB(16) => 
                           TARGET_PC_16_port, PC_BUS_pre_BTB(15) => 
                           TARGET_PC_15_port, PC_BUS_pre_BTB(14) => 
                           TARGET_PC_14_port, PC_BUS_pre_BTB(13) => 
                           TARGET_PC_13_port, PC_BUS_pre_BTB(12) => 
                           TARGET_PC_12_port, PC_BUS_pre_BTB(11) => 
                           TARGET_PC_11_port, PC_BUS_pre_BTB(10) => 
                           TARGET_PC_10_port, PC_BUS_pre_BTB(9) => 
                           TARGET_PC_9_port, PC_BUS_pre_BTB(8) => 
                           TARGET_PC_8_port, PC_BUS_pre_BTB(7) => 
                           TARGET_PC_7_port, PC_BUS_pre_BTB(6) => 
                           TARGET_PC_6_port, PC_BUS_pre_BTB(5) => 
                           TARGET_PC_5_port, PC_BUS_pre_BTB(4) => 
                           TARGET_PC_4_port, PC_BUS_pre_BTB(3) => 
                           TARGET_PC_3_port, PC_BUS_pre_BTB(2) => 
                           TARGET_PC_2_port, PC_BUS_pre_BTB(1) => 
                           TARGET_PC_1_port, PC_BUS_pre_BTB(0) => 
                           TARGET_PC_0_port, stall_i => stall_fetch, 
                           take_prediction_i => take_prediction, mispredict_i 
                           => n4, predicted_PC(31) => predicted_PC_31_port, 
                           predicted_PC(30) => predicted_PC_30_port, 
                           predicted_PC(29) => predicted_PC_29_port, 
                           predicted_PC(28) => predicted_PC_28_port, 
                           predicted_PC(27) => predicted_PC_27_port, 
                           predicted_PC(26) => predicted_PC_26_port, 
                           predicted_PC(25) => predicted_PC_25_port, 
                           predicted_PC(24) => predicted_PC_24_port, 
                           predicted_PC(23) => predicted_PC_23_port, 
                           predicted_PC(22) => predicted_PC_22_port, 
                           predicted_PC(21) => predicted_PC_21_port, 
                           predicted_PC(20) => predicted_PC_20_port, 
                           predicted_PC(19) => predicted_PC_19_port, 
                           predicted_PC(18) => predicted_PC_18_port, 
                           predicted_PC(17) => predicted_PC_17_port, 
                           predicted_PC(16) => predicted_PC_16_port, 
                           predicted_PC(15) => predicted_PC_15_port, 
                           predicted_PC(14) => predicted_PC_14_port, 
                           predicted_PC(13) => predicted_PC_13_port, 
                           predicted_PC(12) => predicted_PC_12_port, 
                           predicted_PC(11) => predicted_PC_11_port, 
                           predicted_PC(10) => predicted_PC_10_port, 
                           predicted_PC(9) => predicted_PC_9_port, 
                           predicted_PC(8) => predicted_PC_8_port, 
                           predicted_PC(7) => predicted_PC_7_port, 
                           predicted_PC(6) => predicted_PC_6_port, 
                           predicted_PC(5) => predicted_PC_5_port, 
                           predicted_PC(4) => predicted_PC_4_port, 
                           predicted_PC(3) => predicted_PC_3_port, 
                           predicted_PC(2) => predicted_PC_2_port, 
                           predicted_PC(1) => predicted_PC_1_port, 
                           predicted_PC(0) => predicted_PC_0_port, clk => clock
                           , rst => rst);
   UBTB : btb_N_LINES4_SIZE32 port map( clock => clock, reset => rst, stall_i 
                           => stall_btb, TAG_i(3) => IRAM_Addr_o_5_port, 
                           TAG_i(2) => IRAM_Addr_o_4_port, TAG_i(1) => 
                           IRAM_Addr_o_3_port, TAG_i(0) => IRAM_Addr_o_2_port, 
                           target_PC_i(31) => TARGET_PC_31_port, 
                           target_PC_i(30) => TARGET_PC_30_port, 
                           target_PC_i(29) => TARGET_PC_29_port, 
                           target_PC_i(28) => TARGET_PC_28_port, 
                           target_PC_i(27) => TARGET_PC_27_port, 
                           target_PC_i(26) => TARGET_PC_26_port, 
                           target_PC_i(25) => TARGET_PC_25_port, 
                           target_PC_i(24) => TARGET_PC_24_port, 
                           target_PC_i(23) => TARGET_PC_23_port, 
                           target_PC_i(22) => TARGET_PC_22_port, 
                           target_PC_i(21) => TARGET_PC_21_port, 
                           target_PC_i(20) => TARGET_PC_20_port, 
                           target_PC_i(19) => TARGET_PC_19_port, 
                           target_PC_i(18) => TARGET_PC_18_port, 
                           target_PC_i(17) => TARGET_PC_17_port, 
                           target_PC_i(16) => TARGET_PC_16_port, 
                           target_PC_i(15) => TARGET_PC_15_port, 
                           target_PC_i(14) => TARGET_PC_14_port, 
                           target_PC_i(13) => TARGET_PC_13_port, 
                           target_PC_i(12) => TARGET_PC_12_port, 
                           target_PC_i(11) => TARGET_PC_11_port, 
                           target_PC_i(10) => TARGET_PC_10_port, target_PC_i(9)
                           => TARGET_PC_9_port, target_PC_i(8) => 
                           TARGET_PC_8_port, target_PC_i(7) => TARGET_PC_7_port
                           , target_PC_i(6) => TARGET_PC_6_port, target_PC_i(5)
                           => TARGET_PC_5_port, target_PC_i(4) => 
                           TARGET_PC_4_port, target_PC_i(3) => TARGET_PC_3_port
                           , target_PC_i(2) => TARGET_PC_2_port, target_PC_i(1)
                           => TARGET_PC_1_port, target_PC_i(0) => 
                           TARGET_PC_0_port, was_taken_i => was_taken, 
                           predicted_next_PC_o(31) => predicted_PC_31_port, 
                           predicted_next_PC_o(30) => predicted_PC_30_port, 
                           predicted_next_PC_o(29) => predicted_PC_29_port, 
                           predicted_next_PC_o(28) => predicted_PC_28_port, 
                           predicted_next_PC_o(27) => predicted_PC_27_port, 
                           predicted_next_PC_o(26) => predicted_PC_26_port, 
                           predicted_next_PC_o(25) => predicted_PC_25_port, 
                           predicted_next_PC_o(24) => predicted_PC_24_port, 
                           predicted_next_PC_o(23) => predicted_PC_23_port, 
                           predicted_next_PC_o(22) => predicted_PC_22_port, 
                           predicted_next_PC_o(21) => predicted_PC_21_port, 
                           predicted_next_PC_o(20) => predicted_PC_20_port, 
                           predicted_next_PC_o(19) => predicted_PC_19_port, 
                           predicted_next_PC_o(18) => predicted_PC_18_port, 
                           predicted_next_PC_o(17) => predicted_PC_17_port, 
                           predicted_next_PC_o(16) => predicted_PC_16_port, 
                           predicted_next_PC_o(15) => predicted_PC_15_port, 
                           predicted_next_PC_o(14) => predicted_PC_14_port, 
                           predicted_next_PC_o(13) => predicted_PC_13_port, 
                           predicted_next_PC_o(12) => predicted_PC_12_port, 
                           predicted_next_PC_o(11) => predicted_PC_11_port, 
                           predicted_next_PC_o(10) => predicted_PC_10_port, 
                           predicted_next_PC_o(9) => predicted_PC_9_port, 
                           predicted_next_PC_o(8) => predicted_PC_8_port, 
                           predicted_next_PC_o(7) => predicted_PC_7_port, 
                           predicted_next_PC_o(6) => predicted_PC_6_port, 
                           predicted_next_PC_o(5) => predicted_PC_5_port, 
                           predicted_next_PC_o(4) => predicted_PC_4_port, 
                           predicted_next_PC_o(3) => predicted_PC_3_port, 
                           predicted_next_PC_o(2) => predicted_PC_2_port, 
                           predicted_next_PC_o(1) => predicted_PC_1_port, 
                           predicted_next_PC_o(0) => predicted_PC_0_port, 
                           taken_o => take_prediction, mispredict_o => n4);
   UFEETCH_REGS : fetch_regs port map( NPCF_i(31) => PC4_31_port, NPCF_i(30) =>
                           PC4_30_port, NPCF_i(29) => PC4_29_port, NPCF_i(28) 
                           => PC4_28_port, NPCF_i(27) => PC4_27_port, 
                           NPCF_i(26) => PC4_26_port, NPCF_i(25) => PC4_25_port
                           , NPCF_i(24) => PC4_24_port, NPCF_i(23) => 
                           PC4_23_port, NPCF_i(22) => PC4_22_port, NPCF_i(21) 
                           => PC4_21_port, NPCF_i(20) => PC4_20_port, 
                           NPCF_i(19) => PC4_19_port, NPCF_i(18) => PC4_18_port
                           , NPCF_i(17) => PC4_17_port, NPCF_i(16) => 
                           PC4_16_port, NPCF_i(15) => PC4_15_port, NPCF_i(14) 
                           => PC4_14_port, NPCF_i(13) => PC4_13_port, 
                           NPCF_i(12) => PC4_12_port, NPCF_i(11) => PC4_11_port
                           , NPCF_i(10) => PC4_10_port, NPCF_i(9) => PC4_9_port
                           , NPCF_i(8) => PC4_8_port, NPCF_i(7) => PC4_7_port, 
                           NPCF_i(6) => PC4_6_port, NPCF_i(5) => PC4_5_port, 
                           NPCF_i(4) => PC4_4_port, NPCF_i(3) => PC4_3_port, 
                           NPCF_i(2) => PC4_2_port, NPCF_i(1) => PC4_1_port, 
                           NPCF_i(0) => PC4_0_port, IR_i(31) => IRAM_Dout_i(31)
                           , IR_i(30) => IRAM_Dout_i(30), IR_i(29) => 
                           IRAM_Dout_i(29), IR_i(28) => IRAM_Dout_i(28), 
                           IR_i(27) => IRAM_Dout_i(27), IR_i(26) => 
                           IRAM_Dout_i(26), IR_i(25) => IRAM_Dout_i(25), 
                           IR_i(24) => IRAM_Dout_i(24), IR_i(23) => 
                           IRAM_Dout_i(23), IR_i(22) => IRAM_Dout_i(22), 
                           IR_i(21) => IRAM_Dout_i(21), IR_i(20) => 
                           IRAM_Dout_i(20), IR_i(19) => IRAM_Dout_i(19), 
                           IR_i(18) => IRAM_Dout_i(18), IR_i(17) => 
                           IRAM_Dout_i(17), IR_i(16) => IRAM_Dout_i(16), 
                           IR_i(15) => IRAM_Dout_i(15), IR_i(14) => 
                           IRAM_Dout_i(14), IR_i(13) => IRAM_Dout_i(13), 
                           IR_i(12) => IRAM_Dout_i(12), IR_i(11) => 
                           IRAM_Dout_i(11), IR_i(10) => IRAM_Dout_i(10), 
                           IR_i(9) => IRAM_Dout_i(9), IR_i(8) => IRAM_Dout_i(8)
                           , IR_i(7) => IRAM_Dout_i(7), IR_i(6) => 
                           IRAM_Dout_i(6), IR_i(5) => IRAM_Dout_i(5), IR_i(4) 
                           => IRAM_Dout_i(4), IR_i(3) => IRAM_Dout_i(3), 
                           IR_i(2) => IRAM_Dout_i(2), IR_i(1) => IRAM_Dout_i(1)
                           , IR_i(0) => IRAM_Dout_i(0), NPCF_o(31) => 
                           NPCF_31_port, NPCF_o(30) => NPCF_30_port, NPCF_o(29)
                           => NPCF_29_port, NPCF_o(28) => NPCF_28_port, 
                           NPCF_o(27) => NPCF_27_port, NPCF_o(26) => 
                           NPCF_26_port, NPCF_o(25) => NPCF_25_port, NPCF_o(24)
                           => NPCF_24_port, NPCF_o(23) => NPCF_23_port, 
                           NPCF_o(22) => NPCF_22_port, NPCF_o(21) => 
                           NPCF_21_port, NPCF_o(20) => NPCF_20_port, NPCF_o(19)
                           => NPCF_19_port, NPCF_o(18) => NPCF_18_port, 
                           NPCF_o(17) => NPCF_17_port, NPCF_o(16) => 
                           NPCF_16_port, NPCF_o(15) => NPCF_15_port, NPCF_o(14)
                           => NPCF_14_port, NPCF_o(13) => NPCF_13_port, 
                           NPCF_o(12) => NPCF_12_port, NPCF_o(11) => 
                           NPCF_11_port, NPCF_o(10) => NPCF_10_port, NPCF_o(9) 
                           => NPCF_9_port, NPCF_o(8) => NPCF_8_port, NPCF_o(7) 
                           => NPCF_7_port, NPCF_o(6) => NPCF_6_port, NPCF_o(5) 
                           => NPCF_5_port, NPCF_o(4) => NPCF_4_port, NPCF_o(3) 
                           => NPCF_3_port, NPCF_o(2) => NPCF_2_port, NPCF_o(1) 
                           => NPCF_1_port, NPCF_o(0) => NPCF_0_port, IR_o(31) 
                           => IR_31_port, IR_o(30) => IR_30_port, IR_o(29) => 
                           IR_29_port, IR_o(28) => IR_28_port, IR_o(27) => 
                           IR_27_port, IR_o(26) => IR_26_port, IR_o(25) => 
                           IR_25_port, IR_o(24) => IR_24_port, IR_o(23) => 
                           IR_23_port, IR_o(22) => IR_22_port, IR_o(21) => 
                           IR_21_port, IR_o(20) => IR_20_port, IR_o(19) => 
                           IR_19_port, IR_o(18) => IR_18_port, IR_o(17) => 
                           IR_17_port, IR_o(16) => IR_16_port, IR_o(15) => 
                           IR_15_port, IR_o(14) => IR_14_port, IR_o(13) => 
                           IR_13_port, IR_o(12) => IR_12_port, IR_o(11) => 
                           IR_11_port, IR_o(10) => IR_10_port, IR_o(9) => 
                           IR_9_port, IR_o(8) => IR_8_port, IR_o(7) => 
                           IR_7_port, IR_o(6) => IR_6_port, IR_o(5) => 
                           IR_5_port, IR_o(4) => IR_4_port, IR_o(3) => 
                           IR_3_port, IR_o(2) => IR_2_port, IR_o(1) => 
                           IR_1_port, IR_o(0) => IR_0_port, stall_i => 
                           stall_decode, clk => clock, rst => rst);
   UJUMP_LOGIC : jump_logic port map( NPCF_i(31) => NPCF_31_port, NPCF_i(30) =>
                           NPCF_30_port, NPCF_i(29) => NPCF_29_port, NPCF_i(28)
                           => NPCF_28_port, NPCF_i(27) => NPCF_27_port, 
                           NPCF_i(26) => NPCF_26_port, NPCF_i(25) => 
                           NPCF_25_port, NPCF_i(24) => NPCF_24_port, NPCF_i(23)
                           => NPCF_23_port, NPCF_i(22) => NPCF_22_port, 
                           NPCF_i(21) => NPCF_21_port, NPCF_i(20) => 
                           NPCF_20_port, NPCF_i(19) => NPCF_19_port, NPCF_i(18)
                           => NPCF_18_port, NPCF_i(17) => NPCF_17_port, 
                           NPCF_i(16) => NPCF_16_port, NPCF_i(15) => 
                           NPCF_15_port, NPCF_i(14) => NPCF_14_port, NPCF_i(13)
                           => NPCF_13_port, NPCF_i(12) => NPCF_12_port, 
                           NPCF_i(11) => NPCF_11_port, NPCF_i(10) => 
                           NPCF_10_port, NPCF_i(9) => NPCF_9_port, NPCF_i(8) =>
                           NPCF_8_port, NPCF_i(7) => NPCF_7_port, NPCF_i(6) => 
                           NPCF_6_port, NPCF_i(5) => NPCF_5_port, NPCF_i(4) => 
                           NPCF_4_port, NPCF_i(3) => NPCF_3_port, NPCF_i(2) => 
                           NPCF_2_port, NPCF_i(1) => NPCF_1_port, NPCF_i(0) => 
                           NPCF_0_port, IR_i(31) => n12, IR_i(30) => n13, 
                           IR_i(29) => n14, IR_i(28) => n15, IR_i(27) => n16, 
                           IR_i(26) => n17, IR_i(25) => IR_25_port, IR_i(24) =>
                           IR_24_port, IR_i(23) => IR_23_port, IR_i(22) => 
                           IR_22_port, IR_i(21) => IR_21_port, IR_i(20) => 
                           IR_20_port, IR_i(19) => IR_19_port, IR_i(18) => 
                           IR_18_port, IR_i(17) => IR_17_port, IR_i(16) => 
                           IR_16_port, IR_i(15) => IR_15_port, IR_i(14) => 
                           IR_14_port, IR_i(13) => IR_13_port, IR_i(12) => 
                           IR_12_port, IR_i(11) => IR_11_port, IR_i(10) => 
                           IR_10_port, IR_i(9) => IR_9_port, IR_i(8) => 
                           IR_8_port, IR_i(7) => IR_7_port, IR_i(6) => 
                           IR_6_port, IR_i(5) => IR_5_port, IR_i(4) => 
                           IR_4_port, IR_i(3) => IR_3_port, IR_i(2) => 
                           IR_2_port, IR_i(1) => IR_1_port, IR_i(0) => 
                           IR_0_port, A_i(31) => AtoComp_31_port, A_i(30) => 
                           AtoComp_30_port, A_i(29) => AtoComp_29_port, A_i(28)
                           => AtoComp_28_port, A_i(27) => AtoComp_27_port, 
                           A_i(26) => AtoComp_26_port, A_i(25) => 
                           AtoComp_25_port, A_i(24) => AtoComp_24_port, A_i(23)
                           => AtoComp_23_port, A_i(22) => AtoComp_22_port, 
                           A_i(21) => AtoComp_21_port, A_i(20) => 
                           AtoComp_20_port, A_i(19) => AtoComp_19_port, A_i(18)
                           => AtoComp_18_port, A_i(17) => AtoComp_17_port, 
                           A_i(16) => AtoComp_16_port, A_i(15) => 
                           AtoComp_15_port, A_i(14) => AtoComp_14_port, A_i(13)
                           => AtoComp_13_port, A_i(12) => AtoComp_12_port, 
                           A_i(11) => AtoComp_11_port, A_i(10) => 
                           AtoComp_10_port, A_i(9) => AtoComp_9_port, A_i(8) =>
                           AtoComp_8_port, A_i(7) => AtoComp_7_port, A_i(6) => 
                           AtoComp_6_port, A_i(5) => AtoComp_5_port, A_i(4) => 
                           AtoComp_4_port, A_i(3) => AtoComp_3_port, A_i(2) => 
                           AtoComp_2_port, A_i(1) => AtoComp_1_port, A_i(0) => 
                           AtoComp_0_port, A_o(31) => dummy_A_31_port, A_o(30) 
                           => dummy_A_30_port, A_o(29) => dummy_A_29_port, 
                           A_o(28) => dummy_A_28_port, A_o(27) => 
                           dummy_A_27_port, A_o(26) => dummy_A_26_port, A_o(25)
                           => dummy_A_25_port, A_o(24) => dummy_A_24_port, 
                           A_o(23) => dummy_A_23_port, A_o(22) => 
                           dummy_A_22_port, A_o(21) => dummy_A_21_port, A_o(20)
                           => dummy_A_20_port, A_o(19) => dummy_A_19_port, 
                           A_o(18) => dummy_A_18_port, A_o(17) => 
                           dummy_A_17_port, A_o(16) => dummy_A_16_port, A_o(15)
                           => dummy_A_15_port, A_o(14) => dummy_A_14_port, 
                           A_o(13) => dummy_A_13_port, A_o(12) => 
                           dummy_A_12_port, A_o(11) => dummy_A_11_port, A_o(10)
                           => dummy_A_10_port, A_o(9) => dummy_A_9_port, A_o(8)
                           => dummy_A_8_port, A_o(7) => dummy_A_7_port, A_o(6) 
                           => dummy_A_6_port, A_o(5) => dummy_A_5_port, A_o(4) 
                           => dummy_A_4_port, A_o(3) => dummy_A_3_port, A_o(2) 
                           => dummy_A_2_port, A_o(1) => dummy_A_1_port, A_o(0) 
                           => dummy_A_0_port, rA_o(4) => rA2reg_4_port, rA_o(3)
                           => rA2reg_3_port, rA_o(2) => rA2reg_2_port, rA_o(1) 
                           => rA2reg_1_port, rA_o(0) => rA2reg_0_port, rB_o(4) 
                           => rB2reg_4_port, rB_o(3) => rB2reg_3_port, rB_o(2) 
                           => rB2reg_2_port, rB_o(1) => rB2reg_1_port, rB_o(0) 
                           => rB2reg_0_port, rC_o(4) => rC2reg_4_port, rC_o(3) 
                           => rC2reg_3_port, rC_o(2) => rC2reg_2_port, rC_o(1) 
                           => rC2reg_1_port, rC_o(0) => rC2reg_0_port, 
                           branch_target_o(31) => dummy_branch_target_31_port, 
                           branch_target_o(30) => dummy_branch_target_30_port, 
                           branch_target_o(29) => dummy_branch_target_29_port, 
                           branch_target_o(28) => dummy_branch_target_28_port, 
                           branch_target_o(27) => dummy_branch_target_27_port, 
                           branch_target_o(26) => dummy_branch_target_26_port, 
                           branch_target_o(25) => dummy_branch_target_25_port, 
                           branch_target_o(24) => dummy_branch_target_24_port, 
                           branch_target_o(23) => dummy_branch_target_23_port, 
                           branch_target_o(22) => dummy_branch_target_22_port, 
                           branch_target_o(21) => dummy_branch_target_21_port, 
                           branch_target_o(20) => dummy_branch_target_20_port, 
                           branch_target_o(19) => dummy_branch_target_19_port, 
                           branch_target_o(18) => dummy_branch_target_18_port, 
                           branch_target_o(17) => dummy_branch_target_17_port, 
                           branch_target_o(16) => dummy_branch_target_16_port, 
                           branch_target_o(15) => dummy_branch_target_15_port, 
                           branch_target_o(14) => dummy_branch_target_14_port, 
                           branch_target_o(13) => dummy_branch_target_13_port, 
                           branch_target_o(12) => dummy_branch_target_12_port, 
                           branch_target_o(11) => dummy_branch_target_11_port, 
                           branch_target_o(10) => dummy_branch_target_10_port, 
                           branch_target_o(9) => dummy_branch_target_9_port, 
                           branch_target_o(8) => dummy_branch_target_8_port, 
                           branch_target_o(7) => dummy_branch_target_7_port, 
                           branch_target_o(6) => dummy_branch_target_6_port, 
                           branch_target_o(5) => dummy_branch_target_5_port, 
                           branch_target_o(4) => dummy_branch_target_4_port, 
                           branch_target_o(3) => dummy_branch_target_3_port, 
                           branch_target_o(2) => dummy_branch_target_2_port, 
                           branch_target_o(1) => dummy_branch_target_1_port, 
                           branch_target_o(0) => dummy_branch_target_0_port, 
                           sum_addr_o(31) => dummy_sum_addr_31_port, 
                           sum_addr_o(30) => dummy_sum_addr_30_port, 
                           sum_addr_o(29) => dummy_sum_addr_29_port, 
                           sum_addr_o(28) => dummy_sum_addr_28_port, 
                           sum_addr_o(27) => dummy_sum_addr_27_port, 
                           sum_addr_o(26) => dummy_sum_addr_26_port, 
                           sum_addr_o(25) => dummy_sum_addr_25_port, 
                           sum_addr_o(24) => dummy_sum_addr_24_port, 
                           sum_addr_o(23) => dummy_sum_addr_23_port, 
                           sum_addr_o(22) => dummy_sum_addr_22_port, 
                           sum_addr_o(21) => dummy_sum_addr_21_port, 
                           sum_addr_o(20) => dummy_sum_addr_20_port, 
                           sum_addr_o(19) => dummy_sum_addr_19_port, 
                           sum_addr_o(18) => dummy_sum_addr_18_port, 
                           sum_addr_o(17) => dummy_sum_addr_17_port, 
                           sum_addr_o(16) => dummy_sum_addr_16_port, 
                           sum_addr_o(15) => dummy_sum_addr_15_port, 
                           sum_addr_o(14) => dummy_sum_addr_14_port, 
                           sum_addr_o(13) => dummy_sum_addr_13_port, 
                           sum_addr_o(12) => dummy_sum_addr_12_port, 
                           sum_addr_o(11) => dummy_sum_addr_11_port, 
                           sum_addr_o(10) => dummy_sum_addr_10_port, 
                           sum_addr_o(9) => dummy_sum_addr_9_port, 
                           sum_addr_o(8) => dummy_sum_addr_8_port, 
                           sum_addr_o(7) => dummy_sum_addr_7_port, 
                           sum_addr_o(6) => dummy_sum_addr_6_port, 
                           sum_addr_o(5) => dummy_sum_addr_5_port, 
                           sum_addr_o(4) => dummy_sum_addr_4_port, 
                           sum_addr_o(3) => dummy_sum_addr_3_port, 
                           sum_addr_o(2) => dummy_sum_addr_2_port, 
                           sum_addr_o(1) => dummy_sum_addr_1_port, 
                           sum_addr_o(0) => dummy_sum_addr_0_port, 
                           extended_imm(31) => help_IMM_31_port, 
                           extended_imm(30) => help_IMM_30_port, 
                           extended_imm(29) => help_IMM_29_port, 
                           extended_imm(28) => help_IMM_28_port, 
                           extended_imm(27) => help_IMM_27_port, 
                           extended_imm(26) => help_IMM_26_port, 
                           extended_imm(25) => help_IMM_25_port, 
                           extended_imm(24) => help_IMM_24_port, 
                           extended_imm(23) => help_IMM_23_port, 
                           extended_imm(22) => help_IMM_22_port, 
                           extended_imm(21) => help_IMM_21_port, 
                           extended_imm(20) => help_IMM_20_port, 
                           extended_imm(19) => help_IMM_19_port, 
                           extended_imm(18) => help_IMM_18_port, 
                           extended_imm(17) => help_IMM_17_port, 
                           extended_imm(16) => help_IMM_16_port, 
                           extended_imm(15) => help_IMM_15_port, 
                           extended_imm(14) => help_IMM_14_port, 
                           extended_imm(13) => help_IMM_13_port, 
                           extended_imm(12) => help_IMM_12_port, 
                           extended_imm(11) => help_IMM_11_port, 
                           extended_imm(10) => help_IMM_10_port, 
                           extended_imm(9) => help_IMM_9_port, extended_imm(8) 
                           => help_IMM_8_port, extended_imm(7) => 
                           help_IMM_7_port, extended_imm(6) => help_IMM_6_port,
                           extended_imm(5) => help_IMM_5_port, extended_imm(4) 
                           => help_IMM_4_port, extended_imm(3) => 
                           help_IMM_3_port, extended_imm(2) => help_IMM_2_port,
                           extended_imm(1) => help_IMM_1_port, extended_imm(0) 
                           => help_IMM_0_port, taken_o => was_taken_from_jl, 
                           FW_X_i(31) => DRAM_Addr_o_31_port, FW_X_i(30) => 
                           DRAM_Addr_o_30_port, FW_X_i(29) => 
                           DRAM_Addr_o_29_port, FW_X_i(28) => 
                           DRAM_Addr_o_28_port, FW_X_i(27) => 
                           DRAM_Addr_o_27_port, FW_X_i(26) => 
                           DRAM_Addr_o_26_port, FW_X_i(25) => 
                           DRAM_Addr_o_25_port, FW_X_i(24) => 
                           DRAM_Addr_o_24_port, FW_X_i(23) => 
                           DRAM_Addr_o_23_port, FW_X_i(22) => 
                           DRAM_Addr_o_22_port, FW_X_i(21) => 
                           DRAM_Addr_o_21_port, FW_X_i(20) => 
                           DRAM_Addr_o_20_port, FW_X_i(19) => 
                           DRAM_Addr_o_19_port, FW_X_i(18) => 
                           DRAM_Addr_o_18_port, FW_X_i(17) => 
                           DRAM_Addr_o_17_port, FW_X_i(16) => 
                           DRAM_Addr_o_16_port, FW_X_i(15) => 
                           DRAM_Addr_o_15_port, FW_X_i(14) => 
                           DRAM_Addr_o_14_port, FW_X_i(13) => 
                           DRAM_Addr_o_13_port, FW_X_i(12) => 
                           DRAM_Addr_o_12_port, FW_X_i(11) => 
                           DRAM_Addr_o_11_port, FW_X_i(10) => 
                           DRAM_Addr_o_10_port, FW_X_i(9) => DRAM_Addr_o_9_port
                           , FW_X_i(8) => DRAM_Addr_o_8_port, FW_X_i(7) => 
                           DRAM_Addr_o_7_port, FW_X_i(6) => DRAM_Addr_o_6_port,
                           FW_X_i(5) => DRAM_Addr_o_5_port, FW_X_i(4) => 
                           DRAM_Addr_o_4_port, FW_X_i(3) => DRAM_Addr_o_3_port,
                           FW_X_i(2) => DRAM_Addr_o_2_port, FW_X_i(1) => 
                           DRAM_Addr_o_1_port, FW_X_i(0) => DRAM_Addr_o_0_port,
                           FW_W_i(31) => wb2reg_31_port, FW_W_i(30) => 
                           wb2reg_30_port, FW_W_i(29) => wb2reg_29_port, 
                           FW_W_i(28) => wb2reg_28_port, FW_W_i(27) => 
                           wb2reg_27_port, FW_W_i(26) => wb2reg_26_port, 
                           FW_W_i(25) => wb2reg_25_port, FW_W_i(24) => 
                           wb2reg_24_port, FW_W_i(23) => wb2reg_23_port, 
                           FW_W_i(22) => wb2reg_22_port, FW_W_i(21) => 
                           wb2reg_21_port, FW_W_i(20) => wb2reg_20_port, 
                           FW_W_i(19) => wb2reg_19_port, FW_W_i(18) => 
                           wb2reg_18_port, FW_W_i(17) => wb2reg_17_port, 
                           FW_W_i(16) => wb2reg_16_port, FW_W_i(15) => 
                           wb2reg_15_port, FW_W_i(14) => wb2reg_14_port, 
                           FW_W_i(13) => wb2reg_13_port, FW_W_i(12) => 
                           wb2reg_12_port, FW_W_i(11) => wb2reg_11_port, 
                           FW_W_i(10) => wb2reg_10_port, FW_W_i(9) => 
                           wb2reg_9_port, FW_W_i(8) => wb2reg_8_port, FW_W_i(7)
                           => wb2reg_7_port, FW_W_i(6) => wb2reg_6_port, 
                           FW_W_i(5) => wb2reg_5_port, FW_W_i(4) => 
                           wb2reg_4_port, FW_W_i(3) => wb2reg_3_port, FW_W_i(2)
                           => wb2reg_2_port, FW_W_i(1) => wb2reg_1_port, 
                           FW_W_i(0) => wb2reg_0_port, S_FW_Adec_i(1) => 
                           dummy_S_FWAdec_1_port, S_FW_Adec_i(0) => 
                           dummy_S_FWAdec_0_port, S_EXT_i => dummy_S_EXT, 
                           S_EXT_SIGN_i => dummy_S_EXT_SIGN, S_MUX_LINK_i => n6
                           , S_EQ_NEQ_i => dummy_S_EQ_NEQ);
   UCU : 
                           dlx_cu_MICROCODE_MEM_SIZE64_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE13 
                           port map( Clk => clock, Rst => rst, IR_IN(31) => 
                           IR_31_port, IR_IN(30) => IR_30_port, IR_IN(29) => 
                           IR_29_port, IR_IN(28) => IR_28_port, IR_IN(27) => 
                           IR_27_port, IR_IN(26) => IR_26_port, IR_IN(25) => 
                           IR_25_port, IR_IN(24) => IR_24_port, IR_IN(23) => 
                           IR_23_port, IR_IN(22) => IR_22_port, IR_IN(21) => 
                           IR_21_port, IR_IN(20) => IR_20_port, IR_IN(19) => 
                           IR_19_port, IR_IN(18) => IR_18_port, IR_IN(17) => 
                           IR_17_port, IR_IN(16) => IR_16_port, IR_IN(15) => 
                           n18, IR_IN(14) => n19, IR_IN(13) => n20, IR_IN(12) 
                           => n21, IR_IN(11) => n22, IR_IN(10) => IR_10_port, 
                           IR_IN(9) => IR_9_port, IR_IN(8) => IR_8_port, 
                           IR_IN(7) => IR_7_port, IR_IN(6) => IR_6_port, 
                           IR_IN(5) => IR_5_port, IR_IN(4) => IR_4_port, 
                           IR_IN(3) => IR_3_port, IR_IN(2) => IR_2_port, 
                           IR_IN(1) => IR_1_port, IR_IN(0) => IR_0_port, 
                           stall_exe_i => exe_stall_cu, mispredict_i => n4, 
                           D1_i(4) => muxed_dest2exe_4_port, D1_i(3) => 
                           muxed_dest2exe_3_port, D1_i(2) => 
                           muxed_dest2exe_2_port, D1_i(1) => 
                           muxed_dest2exe_1_port, D1_i(0) => 
                           muxed_dest2exe_0_port, D2_i(4) => n7, D2_i(3) => n8,
                           D2_i(2) => n9, D2_i(1) => n11, D2_i(0) => n10, 
                           S1_LATCH_EN => net244538, S2_LATCH_EN => net244539, 
                           S3_LATCH_EN => net244540, S_MUX_PC_BUS(1) => 
                           dummy_S_MUX_PC_BUS_1_port, S_MUX_PC_BUS(0) => 
                           dummy_S_MUX_PC_BUS_0_port, S_EXT => dummy_S_EXT, 
                           S_EXT_SIGN => dummy_S_EXT_SIGN, S_EQ_NEQ => 
                           dummy_S_EQ_NEQ, S_MUX_DEST(1) => 
                           dummy_S_MUX_DEST_1_port, S_MUX_DEST(0) => 
                           dummy_S_MUX_DEST_0_port, S_MUX_LINK => n6, S_MUX_MEM
                           => dummy_S_MUX_MEM, S_MEM_W_R => DRAM_WR_o, S_MEM_EN
                           => DRAM_Enable_o, S_RF_W_wb => dummy_S_RF_W_wb, 
                           S_RF_W_mem => dummy_S_RF_W_mem, S_RF_W_exe => 
                           net244541, S_MUX_ALUIN => dummy_S_MUX_ALUIN, 
                           stall_exe_o => stall_exe, stall_dec_o => 
                           stall_decode, stall_fetch_o => stall_fetch, 
                           stall_btb_o => stall_btb, was_branch_o => was_branch
                           , was_jmp_o => was_jmp, ALU_WORD_o(12) => 
                           ALUW_dec_12_port, ALU_WORD_o(11) => ALUW_dec_11_port
                           , ALU_WORD_o(10) => ALUW_dec_10_port, ALU_WORD_o(9) 
                           => ALUW_dec_9_port, ALU_WORD_o(8) => ALUW_dec_8_port
                           , ALU_WORD_o(7) => ALUW_dec_7_port, ALU_WORD_o(6) =>
                           ALUW_dec_6_port, ALU_WORD_o(5) => ALUW_dec_5_port, 
                           ALU_WORD_o(4) => ALUW_dec_4_port, ALU_WORD_o(3) => 
                           ALUW_dec_3_port, ALU_WORD_o(2) => ALUW_dec_2_port, 
                           ALU_WORD_o(1) => ALUW_dec_1_port, ALU_WORD_o(0) => 
                           ALUW_dec_0_port, ALU_OPCODE(0) => net244542, 
                           ALU_OPCODE(1) => net244543, ALU_OPCODE(2) => 
                           net244544, ALU_OPCODE(3) => net244545, ALU_OPCODE(4)
                           => net244546);
   RF : dlx_regfile port map( Clk => clock, Rst => rst, ENABLE => 
                           enable_regfile, RD1 => X_Logic1_port, RD2 => 
                           X_Logic1_port, WR => dummy_S_RF_W_mem, ADD_WR(4) => 
                           n7, ADD_WR(3) => n8, ADD_WR(2) => n9, ADD_WR(1) => 
                           n11, ADD_WR(0) => n10, ADD_RD1(4) => IRAM_Dout_i(25)
                           , ADD_RD1(3) => IRAM_Dout_i(24), ADD_RD1(2) => 
                           IRAM_Dout_i(23), ADD_RD1(1) => IRAM_Dout_i(22), 
                           ADD_RD1(0) => IRAM_Dout_i(21), ADD_RD2(4) => 
                           IRAM_Dout_i(20), ADD_RD2(3) => IRAM_Dout_i(19), 
                           ADD_RD2(2) => IRAM_Dout_i(18), ADD_RD2(1) => 
                           IRAM_Dout_i(17), ADD_RD2(0) => IRAM_Dout_i(16), 
                           DATAIN(31) => W2wb_31_port, DATAIN(30) => 
                           W2wb_30_port, DATAIN(29) => W2wb_29_port, DATAIN(28)
                           => W2wb_28_port, DATAIN(27) => W2wb_27_port, 
                           DATAIN(26) => W2wb_26_port, DATAIN(25) => 
                           W2wb_25_port, DATAIN(24) => W2wb_24_port, DATAIN(23)
                           => W2wb_23_port, DATAIN(22) => W2wb_22_port, 
                           DATAIN(21) => W2wb_21_port, DATAIN(20) => 
                           W2wb_20_port, DATAIN(19) => W2wb_19_port, DATAIN(18)
                           => W2wb_18_port, DATAIN(17) => W2wb_17_port, 
                           DATAIN(16) => W2wb_16_port, DATAIN(15) => 
                           W2wb_15_port, DATAIN(14) => W2wb_14_port, DATAIN(13)
                           => W2wb_13_port, DATAIN(12) => W2wb_12_port, 
                           DATAIN(11) => W2wb_11_port, DATAIN(10) => 
                           W2wb_10_port, DATAIN(9) => W2wb_9_port, DATAIN(8) =>
                           W2wb_8_port, DATAIN(7) => W2wb_7_port, DATAIN(6) => 
                           W2wb_6_port, DATAIN(5) => W2wb_5_port, DATAIN(4) => 
                           W2wb_4_port, DATAIN(3) => W2wb_3_port, DATAIN(2) => 
                           W2wb_2_port, DATAIN(1) => W2wb_1_port, DATAIN(0) => 
                           W2wb_0_port, OUT1(31) => AtoComp_31_port, OUT1(30) 
                           => AtoComp_30_port, OUT1(29) => AtoComp_29_port, 
                           OUT1(28) => AtoComp_28_port, OUT1(27) => 
                           AtoComp_27_port, OUT1(26) => AtoComp_26_port, 
                           OUT1(25) => AtoComp_25_port, OUT1(24) => 
                           AtoComp_24_port, OUT1(23) => AtoComp_23_port, 
                           OUT1(22) => AtoComp_22_port, OUT1(21) => 
                           AtoComp_21_port, OUT1(20) => AtoComp_20_port, 
                           OUT1(19) => AtoComp_19_port, OUT1(18) => 
                           AtoComp_18_port, OUT1(17) => AtoComp_17_port, 
                           OUT1(16) => AtoComp_16_port, OUT1(15) => 
                           AtoComp_15_port, OUT1(14) => AtoComp_14_port, 
                           OUT1(13) => AtoComp_13_port, OUT1(12) => 
                           AtoComp_12_port, OUT1(11) => AtoComp_11_port, 
                           OUT1(10) => AtoComp_10_port, OUT1(9) => 
                           AtoComp_9_port, OUT1(8) => AtoComp_8_port, OUT1(7) 
                           => AtoComp_7_port, OUT1(6) => AtoComp_6_port, 
                           OUT1(5) => AtoComp_5_port, OUT1(4) => AtoComp_4_port
                           , OUT1(3) => AtoComp_3_port, OUT1(2) => 
                           AtoComp_2_port, OUT1(1) => AtoComp_1_port, OUT1(0) 
                           => AtoComp_0_port, OUT2(31) => dummy_B_31_port, 
                           OUT2(30) => dummy_B_30_port, OUT2(29) => 
                           dummy_B_29_port, OUT2(28) => dummy_B_28_port, 
                           OUT2(27) => dummy_B_27_port, OUT2(26) => 
                           dummy_B_26_port, OUT2(25) => dummy_B_25_port, 
                           OUT2(24) => dummy_B_24_port, OUT2(23) => 
                           dummy_B_23_port, OUT2(22) => dummy_B_22_port, 
                           OUT2(21) => dummy_B_21_port, OUT2(20) => 
                           dummy_B_20_port, OUT2(19) => dummy_B_19_port, 
                           OUT2(18) => dummy_B_18_port, OUT2(17) => 
                           dummy_B_17_port, OUT2(16) => dummy_B_16_port, 
                           OUT2(15) => dummy_B_15_port, OUT2(14) => 
                           dummy_B_14_port, OUT2(13) => dummy_B_13_port, 
                           OUT2(12) => dummy_B_12_port, OUT2(11) => 
                           dummy_B_11_port, OUT2(10) => dummy_B_10_port, 
                           OUT2(9) => dummy_B_9_port, OUT2(8) => dummy_B_8_port
                           , OUT2(7) => dummy_B_7_port, OUT2(6) => 
                           dummy_B_6_port, OUT2(5) => dummy_B_5_port, OUT2(4) 
                           => dummy_B_4_port, OUT2(3) => dummy_B_3_port, 
                           OUT2(2) => dummy_B_2_port, OUT2(1) => dummy_B_1_port
                           , OUT2(0) => dummy_B_0_port);
   UDECODE_REGS : decode_regs port map( A_i(31) => AtoComp_31_port, A_i(30) => 
                           AtoComp_30_port, A_i(29) => AtoComp_29_port, A_i(28)
                           => AtoComp_28_port, A_i(27) => AtoComp_27_port, 
                           A_i(26) => AtoComp_26_port, A_i(25) => 
                           AtoComp_25_port, A_i(24) => AtoComp_24_port, A_i(23)
                           => AtoComp_23_port, A_i(22) => AtoComp_22_port, 
                           A_i(21) => AtoComp_21_port, A_i(20) => 
                           AtoComp_20_port, A_i(19) => AtoComp_19_port, A_i(18)
                           => AtoComp_18_port, A_i(17) => AtoComp_17_port, 
                           A_i(16) => AtoComp_16_port, A_i(15) => 
                           AtoComp_15_port, A_i(14) => AtoComp_14_port, A_i(13)
                           => AtoComp_13_port, A_i(12) => AtoComp_12_port, 
                           A_i(11) => AtoComp_11_port, A_i(10) => 
                           AtoComp_10_port, A_i(9) => AtoComp_9_port, A_i(8) =>
                           AtoComp_8_port, A_i(7) => AtoComp_7_port, A_i(6) => 
                           AtoComp_6_port, A_i(5) => AtoComp_5_port, A_i(4) => 
                           AtoComp_4_port, A_i(3) => AtoComp_3_port, A_i(2) => 
                           AtoComp_2_port, A_i(1) => AtoComp_1_port, A_i(0) => 
                           AtoComp_0_port, B_i(31) => dummy_B_31_port, B_i(30) 
                           => dummy_B_30_port, B_i(29) => dummy_B_29_port, 
                           B_i(28) => dummy_B_28_port, B_i(27) => 
                           dummy_B_27_port, B_i(26) => dummy_B_26_port, B_i(25)
                           => dummy_B_25_port, B_i(24) => dummy_B_24_port, 
                           B_i(23) => dummy_B_23_port, B_i(22) => 
                           dummy_B_22_port, B_i(21) => dummy_B_21_port, B_i(20)
                           => dummy_B_20_port, B_i(19) => dummy_B_19_port, 
                           B_i(18) => dummy_B_18_port, B_i(17) => 
                           dummy_B_17_port, B_i(16) => dummy_B_16_port, B_i(15)
                           => dummy_B_15_port, B_i(14) => dummy_B_14_port, 
                           B_i(13) => dummy_B_13_port, B_i(12) => 
                           dummy_B_12_port, B_i(11) => dummy_B_11_port, B_i(10)
                           => dummy_B_10_port, B_i(9) => dummy_B_9_port, B_i(8)
                           => dummy_B_8_port, B_i(7) => dummy_B_7_port, B_i(6) 
                           => dummy_B_6_port, B_i(5) => dummy_B_5_port, B_i(4) 
                           => dummy_B_4_port, B_i(3) => dummy_B_3_port, B_i(2) 
                           => dummy_B_2_port, B_i(1) => dummy_B_1_port, B_i(0) 
                           => dummy_B_0_port, rA_i(4) => rA2reg_4_port, rA_i(3)
                           => rA2reg_3_port, rA_i(2) => rA2reg_2_port, rA_i(1) 
                           => rA2reg_1_port, rA_i(0) => rA2reg_0_port, rB_i(4) 
                           => rB2reg_4_port, rB_i(3) => rB2reg_3_port, rB_i(2) 
                           => rB2reg_2_port, rB_i(1) => rB2reg_1_port, rB_i(0) 
                           => rB2reg_0_port, rC_i(4) => rC2reg_4_port, rC_i(3) 
                           => rC2reg_3_port, rC_i(2) => rC2reg_2_port, rC_i(1) 
                           => rC2reg_1_port, rC_i(0) => rC2reg_0_port, 
                           IMM_i(31) => help_IMM_31_port, IMM_i(30) => 
                           help_IMM_30_port, IMM_i(29) => help_IMM_29_port, 
                           IMM_i(28) => help_IMM_28_port, IMM_i(27) => 
                           help_IMM_27_port, IMM_i(26) => help_IMM_26_port, 
                           IMM_i(25) => help_IMM_25_port, IMM_i(24) => 
                           help_IMM_24_port, IMM_i(23) => help_IMM_23_port, 
                           IMM_i(22) => help_IMM_22_port, IMM_i(21) => 
                           help_IMM_21_port, IMM_i(20) => help_IMM_20_port, 
                           IMM_i(19) => help_IMM_19_port, IMM_i(18) => 
                           help_IMM_18_port, IMM_i(17) => help_IMM_17_port, 
                           IMM_i(16) => help_IMM_16_port, IMM_i(15) => 
                           help_IMM_15_port, IMM_i(14) => help_IMM_14_port, 
                           IMM_i(13) => help_IMM_13_port, IMM_i(12) => 
                           help_IMM_12_port, IMM_i(11) => help_IMM_11_port, 
                           IMM_i(10) => help_IMM_10_port, IMM_i(9) => 
                           help_IMM_9_port, IMM_i(8) => help_IMM_8_port, 
                           IMM_i(7) => help_IMM_7_port, IMM_i(6) => 
                           help_IMM_6_port, IMM_i(5) => help_IMM_5_port, 
                           IMM_i(4) => help_IMM_4_port, IMM_i(3) => 
                           help_IMM_3_port, IMM_i(2) => help_IMM_2_port, 
                           IMM_i(1) => help_IMM_1_port, IMM_i(0) => 
                           help_IMM_0_port, ALUW_i(12) => ALUW_dec_12_port, 
                           ALUW_i(11) => ALUW_dec_11_port, ALUW_i(10) => 
                           ALUW_dec_10_port, ALUW_i(9) => ALUW_dec_9_port, 
                           ALUW_i(8) => ALUW_dec_8_port, ALUW_i(7) => 
                           ALUW_dec_7_port, ALUW_i(6) => ALUW_dec_6_port, 
                           ALUW_i(5) => ALUW_dec_5_port, ALUW_i(4) => 
                           ALUW_dec_4_port, ALUW_i(3) => ALUW_dec_3_port, 
                           ALUW_i(2) => ALUW_dec_2_port, ALUW_i(1) => 
                           ALUW_dec_1_port, ALUW_i(0) => ALUW_dec_0_port, 
                           A_o(31) => A2exe_31_port, A_o(30) => A2exe_30_port, 
                           A_o(29) => A2exe_29_port, A_o(28) => A2exe_28_port, 
                           A_o(27) => A2exe_27_port, A_o(26) => A2exe_26_port, 
                           A_o(25) => A2exe_25_port, A_o(24) => A2exe_24_port, 
                           A_o(23) => A2exe_23_port, A_o(22) => A2exe_22_port, 
                           A_o(21) => A2exe_21_port, A_o(20) => A2exe_20_port, 
                           A_o(19) => A2exe_19_port, A_o(18) => A2exe_18_port, 
                           A_o(17) => A2exe_17_port, A_o(16) => A2exe_16_port, 
                           A_o(15) => A2exe_15_port, A_o(14) => A2exe_14_port, 
                           A_o(13) => A2exe_13_port, A_o(12) => A2exe_12_port, 
                           A_o(11) => A2exe_11_port, A_o(10) => A2exe_10_port, 
                           A_o(9) => A2exe_9_port, A_o(8) => A2exe_8_port, 
                           A_o(7) => A2exe_7_port, A_o(6) => A2exe_6_port, 
                           A_o(5) => A2exe_5_port, A_o(4) => A2exe_4_port, 
                           A_o(3) => A2exe_3_port, A_o(2) => A2exe_2_port, 
                           A_o(1) => A2exe_1_port, A_o(0) => A2exe_0_port, 
                           B_o(31) => B2exe_31_port, B_o(30) => B2exe_30_port, 
                           B_o(29) => B2exe_29_port, B_o(28) => B2exe_28_port, 
                           B_o(27) => B2exe_27_port, B_o(26) => B2exe_26_port, 
                           B_o(25) => B2exe_25_port, B_o(24) => B2exe_24_port, 
                           B_o(23) => B2exe_23_port, B_o(22) => B2exe_22_port, 
                           B_o(21) => B2exe_21_port, B_o(20) => B2exe_20_port, 
                           B_o(19) => B2exe_19_port, B_o(18) => B2exe_18_port, 
                           B_o(17) => B2exe_17_port, B_o(16) => B2exe_16_port, 
                           B_o(15) => B2exe_15_port, B_o(14) => B2exe_14_port, 
                           B_o(13) => B2exe_13_port, B_o(12) => B2exe_12_port, 
                           B_o(11) => B2exe_11_port, B_o(10) => B2exe_10_port, 
                           B_o(9) => B2exe_9_port, B_o(8) => B2exe_8_port, 
                           B_o(7) => B2exe_7_port, B_o(6) => B2exe_6_port, 
                           B_o(5) => B2exe_5_port, B_o(4) => B2exe_4_port, 
                           B_o(3) => B2exe_3_port, B_o(2) => B2exe_2_port, 
                           B_o(1) => B2exe_1_port, B_o(0) => B2exe_0_port, 
                           rA_o(4) => rA2fw_4_port, rA_o(3) => rA2fw_3_port, 
                           rA_o(2) => rA2fw_2_port, rA_o(1) => rA2fw_1_port, 
                           rA_o(0) => rA2fw_0_port, rB_o(4) => rB2mux_4_port, 
                           rB_o(3) => rB2mux_3_port, rB_o(2) => rB2mux_2_port, 
                           rB_o(1) => rB2mux_1_port, rB_o(0) => rB2mux_0_port, 
                           rC_o(4) => rC2mux_4_port, rC_o(3) => rC2mux_3_port, 
                           rC_o(2) => rC2mux_2_port, rC_o(1) => rC2mux_1_port, 
                           rC_o(0) => rC2mux_0_port, IMM_o(31) => 
                           IMM2exe_31_port, IMM_o(30) => IMM2exe_30_port, 
                           IMM_o(29) => IMM2exe_29_port, IMM_o(28) => 
                           IMM2exe_28_port, IMM_o(27) => IMM2exe_27_port, 
                           IMM_o(26) => IMM2exe_26_port, IMM_o(25) => 
                           IMM2exe_25_port, IMM_o(24) => IMM2exe_24_port, 
                           IMM_o(23) => IMM2exe_23_port, IMM_o(22) => 
                           IMM2exe_22_port, IMM_o(21) => IMM2exe_21_port, 
                           IMM_o(20) => IMM2exe_20_port, IMM_o(19) => 
                           IMM2exe_19_port, IMM_o(18) => IMM2exe_18_port, 
                           IMM_o(17) => IMM2exe_17_port, IMM_o(16) => 
                           IMM2exe_16_port, IMM_o(15) => IMM2exe_15_port, 
                           IMM_o(14) => IMM2exe_14_port, IMM_o(13) => 
                           IMM2exe_13_port, IMM_o(12) => IMM2exe_12_port, 
                           IMM_o(11) => IMM2exe_11_port, IMM_o(10) => 
                           IMM2exe_10_port, IMM_o(9) => IMM2exe_9_port, 
                           IMM_o(8) => IMM2exe_8_port, IMM_o(7) => 
                           IMM2exe_7_port, IMM_o(6) => IMM2exe_6_port, IMM_o(5)
                           => IMM2exe_5_port, IMM_o(4) => IMM2exe_4_port, 
                           IMM_o(3) => IMM2exe_3_port, IMM_o(2) => 
                           IMM2exe_2_port, IMM_o(1) => IMM2exe_1_port, IMM_o(0)
                           => IMM2exe_0_port, ALUW_o(12) => ALUW_12_port, 
                           ALUW_o(11) => ALUW_11_port, ALUW_o(10) => 
                           ALUW_10_port, ALUW_o(9) => ALUW_9_port, ALUW_o(8) =>
                           ALUW_8_port, ALUW_o(7) => ALUW_7_port, ALUW_o(6) => 
                           ALUW_6_port, ALUW_o(5) => ALUW_5_port, ALUW_o(4) => 
                           ALUW_4_port, ALUW_o(3) => ALUW_3_port, ALUW_o(2) => 
                           ALUW_2_port, ALUW_o(1) => ALUW_1_port, ALUW_o(0) => 
                           ALUW_0_port, stall_i => stall_exe, clk => clock, rst
                           => rst);
   UEXECUTE_REGS : execute_regs port map( X_i(31) => X2mem_31_port, X_i(30) => 
                           X2mem_30_port, X_i(29) => X2mem_29_port, X_i(28) => 
                           X2mem_28_port, X_i(27) => X2mem_27_port, X_i(26) => 
                           X2mem_26_port, X_i(25) => X2mem_25_port, X_i(24) => 
                           X2mem_24_port, X_i(23) => X2mem_23_port, X_i(22) => 
                           X2mem_22_port, X_i(21) => X2mem_21_port, X_i(20) => 
                           X2mem_20_port, X_i(19) => X2mem_19_port, X_i(18) => 
                           X2mem_18_port, X_i(17) => X2mem_17_port, X_i(16) => 
                           X2mem_16_port, X_i(15) => X2mem_15_port, X_i(14) => 
                           X2mem_14_port, X_i(13) => X2mem_13_port, X_i(12) => 
                           X2mem_12_port, X_i(11) => X2mem_11_port, X_i(10) => 
                           X2mem_10_port, X_i(9) => X2mem_9_port, X_i(8) => 
                           X2mem_8_port, X_i(7) => X2mem_7_port, X_i(6) => 
                           X2mem_6_port, X_i(5) => X2mem_5_port, X_i(4) => 
                           X2mem_4_port, X_i(3) => X2mem_3_port, X_i(2) => 
                           X2mem_2_port, X_i(1) => X2mem_1_port, X_i(0) => 
                           X2mem_0_port, S_i(31) => S2mem_31_port, S_i(30) => 
                           S2mem_30_port, S_i(29) => S2mem_29_port, S_i(28) => 
                           S2mem_28_port, S_i(27) => S2mem_27_port, S_i(26) => 
                           S2mem_26_port, S_i(25) => S2mem_25_port, S_i(24) => 
                           S2mem_24_port, S_i(23) => S2mem_23_port, S_i(22) => 
                           S2mem_22_port, S_i(21) => S2mem_21_port, S_i(20) => 
                           S2mem_20_port, S_i(19) => S2mem_19_port, S_i(18) => 
                           S2mem_18_port, S_i(17) => S2mem_17_port, S_i(16) => 
                           S2mem_16_port, S_i(15) => S2mem_15_port, S_i(14) => 
                           S2mem_14_port, S_i(13) => S2mem_13_port, S_i(12) => 
                           S2mem_12_port, S_i(11) => S2mem_11_port, S_i(10) => 
                           S2mem_10_port, S_i(9) => S2mem_9_port, S_i(8) => 
                           S2mem_8_port, S_i(7) => S2mem_7_port, S_i(6) => 
                           S2mem_6_port, S_i(5) => S2mem_5_port, S_i(4) => 
                           S2mem_4_port, S_i(3) => n5, S_i(2) => S2mem_2_port, 
                           S_i(1) => S2mem_1_port, S_i(0) => S2mem_0_port, 
                           D2_i(4) => muxed_dest2exe_4_port, D2_i(3) => 
                           muxed_dest2exe_3_port, D2_i(2) => 
                           muxed_dest2exe_2_port, D2_i(1) => 
                           muxed_dest2exe_1_port, D2_i(0) => 
                           muxed_dest2exe_0_port, X_o(31) => 
                           DRAM_Addr_o_31_port, X_o(30) => DRAM_Addr_o_30_port,
                           X_o(29) => DRAM_Addr_o_29_port, X_o(28) => 
                           DRAM_Addr_o_28_port, X_o(27) => DRAM_Addr_o_27_port,
                           X_o(26) => DRAM_Addr_o_26_port, X_o(25) => 
                           DRAM_Addr_o_25_port, X_o(24) => DRAM_Addr_o_24_port,
                           X_o(23) => DRAM_Addr_o_23_port, X_o(22) => 
                           DRAM_Addr_o_22_port, X_o(21) => DRAM_Addr_o_21_port,
                           X_o(20) => DRAM_Addr_o_20_port, X_o(19) => 
                           DRAM_Addr_o_19_port, X_o(18) => DRAM_Addr_o_18_port,
                           X_o(17) => DRAM_Addr_o_17_port, X_o(16) => 
                           DRAM_Addr_o_16_port, X_o(15) => DRAM_Addr_o_15_port,
                           X_o(14) => DRAM_Addr_o_14_port, X_o(13) => 
                           DRAM_Addr_o_13_port, X_o(12) => DRAM_Addr_o_12_port,
                           X_o(11) => DRAM_Addr_o_11_port, X_o(10) => 
                           DRAM_Addr_o_10_port, X_o(9) => DRAM_Addr_o_9_port, 
                           X_o(8) => DRAM_Addr_o_8_port, X_o(7) => 
                           DRAM_Addr_o_7_port, X_o(6) => DRAM_Addr_o_6_port, 
                           X_o(5) => DRAM_Addr_o_5_port, X_o(4) => 
                           DRAM_Addr_o_4_port, X_o(3) => DRAM_Addr_o_3_port, 
                           X_o(2) => DRAM_Addr_o_2_port, X_o(1) => 
                           DRAM_Addr_o_1_port, X_o(0) => DRAM_Addr_o_0_port, 
                           S_o(31) => DRAM_Din_o(31), S_o(30) => DRAM_Din_o(30)
                           , S_o(29) => DRAM_Din_o(29), S_o(28) => 
                           DRAM_Din_o(28), S_o(27) => DRAM_Din_o(27), S_o(26) 
                           => DRAM_Din_o(26), S_o(25) => DRAM_Din_o(25), 
                           S_o(24) => DRAM_Din_o(24), S_o(23) => DRAM_Din_o(23)
                           , S_o(22) => DRAM_Din_o(22), S_o(21) => 
                           DRAM_Din_o(21), S_o(20) => DRAM_Din_o(20), S_o(19) 
                           => DRAM_Din_o(19), S_o(18) => DRAM_Din_o(18), 
                           S_o(17) => DRAM_Din_o(17), S_o(16) => DRAM_Din_o(16)
                           , S_o(15) => DRAM_Din_o(15), S_o(14) => 
                           DRAM_Din_o(14), S_o(13) => DRAM_Din_o(13), S_o(12) 
                           => DRAM_Din_o(12), S_o(11) => DRAM_Din_o(11), 
                           S_o(10) => DRAM_Din_o(10), S_o(9) => DRAM_Din_o(9), 
                           S_o(8) => DRAM_Din_o(8), S_o(7) => DRAM_Din_o(7), 
                           S_o(6) => DRAM_Din_o(6), S_o(5) => DRAM_Din_o(5), 
                           S_o(4) => DRAM_Din_o(4), S_o(3) => DRAM_Din_o(3), 
                           S_o(2) => DRAM_Din_o(2), S_o(1) => DRAM_Din_o(1), 
                           S_o(0) => DRAM_Din_o(0), D2_o(4) => D22D3_4_port, 
                           D2_o(3) => D22D3_3_port, D2_o(2) => D22D3_2_port, 
                           D2_o(1) => D22D3_1_port, D2_o(0) => D22D3_0_port, 
                           stall_i => X_Logic0_port, clk => clock, rst => rst);
   UEXECUTE_BLOCK : execute_block port map( IMM_i(31) => IMM2exe_31_port, 
                           IMM_i(30) => IMM2exe_30_port, IMM_i(29) => 
                           IMM2exe_29_port, IMM_i(28) => IMM2exe_28_port, 
                           IMM_i(27) => IMM2exe_27_port, IMM_i(26) => 
                           IMM2exe_26_port, IMM_i(25) => IMM2exe_25_port, 
                           IMM_i(24) => IMM2exe_24_port, IMM_i(23) => 
                           IMM2exe_23_port, IMM_i(22) => IMM2exe_22_port, 
                           IMM_i(21) => IMM2exe_21_port, IMM_i(20) => 
                           IMM2exe_20_port, IMM_i(19) => IMM2exe_19_port, 
                           IMM_i(18) => IMM2exe_18_port, IMM_i(17) => 
                           IMM2exe_17_port, IMM_i(16) => IMM2exe_16_port, 
                           IMM_i(15) => IMM2exe_15_port, IMM_i(14) => 
                           IMM2exe_14_port, IMM_i(13) => IMM2exe_13_port, 
                           IMM_i(12) => IMM2exe_12_port, IMM_i(11) => 
                           IMM2exe_11_port, IMM_i(10) => IMM2exe_10_port, 
                           IMM_i(9) => IMM2exe_9_port, IMM_i(8) => 
                           IMM2exe_8_port, IMM_i(7) => IMM2exe_7_port, IMM_i(6)
                           => IMM2exe_6_port, IMM_i(5) => IMM2exe_5_port, 
                           IMM_i(4) => IMM2exe_4_port, IMM_i(3) => 
                           IMM2exe_3_port, IMM_i(2) => IMM2exe_2_port, IMM_i(1)
                           => IMM2exe_1_port, IMM_i(0) => IMM2exe_0_port, 
                           A_i(31) => A2exe_31_port, A_i(30) => A2exe_30_port, 
                           A_i(29) => A2exe_29_port, A_i(28) => A2exe_28_port, 
                           A_i(27) => A2exe_27_port, A_i(26) => A2exe_26_port, 
                           A_i(25) => A2exe_25_port, A_i(24) => A2exe_24_port, 
                           A_i(23) => A2exe_23_port, A_i(22) => A2exe_22_port, 
                           A_i(21) => A2exe_21_port, A_i(20) => A2exe_20_port, 
                           A_i(19) => A2exe_19_port, A_i(18) => A2exe_18_port, 
                           A_i(17) => A2exe_17_port, A_i(16) => A2exe_16_port, 
                           A_i(15) => A2exe_15_port, A_i(14) => A2exe_14_port, 
                           A_i(13) => A2exe_13_port, A_i(12) => A2exe_12_port, 
                           A_i(11) => A2exe_11_port, A_i(10) => A2exe_10_port, 
                           A_i(9) => A2exe_9_port, A_i(8) => A2exe_8_port, 
                           A_i(7) => A2exe_7_port, A_i(6) => A2exe_6_port, 
                           A_i(5) => A2exe_5_port, A_i(4) => A2exe_4_port, 
                           A_i(3) => A2exe_3_port, A_i(2) => A2exe_2_port, 
                           A_i(1) => A2exe_1_port, A_i(0) => A2exe_0_port, 
                           rB_i(4) => rB2mux_4_port, rB_i(3) => rB2mux_3_port, 
                           rB_i(2) => rB2mux_2_port, rB_i(1) => rB2mux_1_port, 
                           rB_i(0) => rB2mux_0_port, rC_i(4) => rC2mux_4_port, 
                           rC_i(3) => rC2mux_3_port, rC_i(2) => rC2mux_2_port, 
                           rC_i(1) => rC2mux_1_port, rC_i(0) => rC2mux_0_port, 
                           MUXED_B_i(31) => B2exe_31_port, MUXED_B_i(30) => 
                           B2exe_30_port, MUXED_B_i(29) => B2exe_29_port, 
                           MUXED_B_i(28) => B2exe_28_port, MUXED_B_i(27) => 
                           B2exe_27_port, MUXED_B_i(26) => B2exe_26_port, 
                           MUXED_B_i(25) => B2exe_25_port, MUXED_B_i(24) => 
                           B2exe_24_port, MUXED_B_i(23) => B2exe_23_port, 
                           MUXED_B_i(22) => B2exe_22_port, MUXED_B_i(21) => 
                           B2exe_21_port, MUXED_B_i(20) => B2exe_20_port, 
                           MUXED_B_i(19) => B2exe_19_port, MUXED_B_i(18) => 
                           B2exe_18_port, MUXED_B_i(17) => B2exe_17_port, 
                           MUXED_B_i(16) => B2exe_16_port, MUXED_B_i(15) => 
                           B2exe_15_port, MUXED_B_i(14) => B2exe_14_port, 
                           MUXED_B_i(13) => B2exe_13_port, MUXED_B_i(12) => 
                           B2exe_12_port, MUXED_B_i(11) => B2exe_11_port, 
                           MUXED_B_i(10) => B2exe_10_port, MUXED_B_i(9) => 
                           B2exe_9_port, MUXED_B_i(8) => B2exe_8_port, 
                           MUXED_B_i(7) => B2exe_7_port, MUXED_B_i(6) => 
                           B2exe_6_port, MUXED_B_i(5) => B2exe_5_port, 
                           MUXED_B_i(4) => B2exe_4_port, MUXED_B_i(3) => 
                           B2exe_3_port, MUXED_B_i(2) => B2exe_2_port, 
                           MUXED_B_i(1) => B2exe_1_port, MUXED_B_i(0) => 
                           B2exe_0_port, S_MUX_ALUIN_i => dummy_S_MUX_ALUIN, 
                           FW_X_i(31) => DRAM_Addr_o_31_port, FW_X_i(30) => 
                           DRAM_Addr_o_30_port, FW_X_i(29) => 
                           DRAM_Addr_o_29_port, FW_X_i(28) => 
                           DRAM_Addr_o_28_port, FW_X_i(27) => 
                           DRAM_Addr_o_27_port, FW_X_i(26) => 
                           DRAM_Addr_o_26_port, FW_X_i(25) => 
                           DRAM_Addr_o_25_port, FW_X_i(24) => 
                           DRAM_Addr_o_24_port, FW_X_i(23) => 
                           DRAM_Addr_o_23_port, FW_X_i(22) => 
                           DRAM_Addr_o_22_port, FW_X_i(21) => 
                           DRAM_Addr_o_21_port, FW_X_i(20) => 
                           DRAM_Addr_o_20_port, FW_X_i(19) => 
                           DRAM_Addr_o_19_port, FW_X_i(18) => 
                           DRAM_Addr_o_18_port, FW_X_i(17) => 
                           DRAM_Addr_o_17_port, FW_X_i(16) => 
                           DRAM_Addr_o_16_port, FW_X_i(15) => 
                           DRAM_Addr_o_15_port, FW_X_i(14) => 
                           DRAM_Addr_o_14_port, FW_X_i(13) => 
                           DRAM_Addr_o_13_port, FW_X_i(12) => 
                           DRAM_Addr_o_12_port, FW_X_i(11) => 
                           DRAM_Addr_o_11_port, FW_X_i(10) => 
                           DRAM_Addr_o_10_port, FW_X_i(9) => DRAM_Addr_o_9_port
                           , FW_X_i(8) => DRAM_Addr_o_8_port, FW_X_i(7) => 
                           DRAM_Addr_o_7_port, FW_X_i(6) => DRAM_Addr_o_6_port,
                           FW_X_i(5) => DRAM_Addr_o_5_port, FW_X_i(4) => 
                           DRAM_Addr_o_4_port, FW_X_i(3) => DRAM_Addr_o_3_port,
                           FW_X_i(2) => DRAM_Addr_o_2_port, FW_X_i(1) => 
                           DRAM_Addr_o_1_port, FW_X_i(0) => DRAM_Addr_o_0_port,
                           FW_W_i(31) => wb2reg_31_port, FW_W_i(30) => 
                           wb2reg_30_port, FW_W_i(29) => wb2reg_29_port, 
                           FW_W_i(28) => wb2reg_28_port, FW_W_i(27) => 
                           wb2reg_27_port, FW_W_i(26) => wb2reg_26_port, 
                           FW_W_i(25) => wb2reg_25_port, FW_W_i(24) => 
                           wb2reg_24_port, FW_W_i(23) => wb2reg_23_port, 
                           FW_W_i(22) => wb2reg_22_port, FW_W_i(21) => 
                           wb2reg_21_port, FW_W_i(20) => wb2reg_20_port, 
                           FW_W_i(19) => wb2reg_19_port, FW_W_i(18) => 
                           wb2reg_18_port, FW_W_i(17) => wb2reg_17_port, 
                           FW_W_i(16) => wb2reg_16_port, FW_W_i(15) => 
                           wb2reg_15_port, FW_W_i(14) => wb2reg_14_port, 
                           FW_W_i(13) => wb2reg_13_port, FW_W_i(12) => 
                           wb2reg_12_port, FW_W_i(11) => wb2reg_11_port, 
                           FW_W_i(10) => wb2reg_10_port, FW_W_i(9) => 
                           wb2reg_9_port, FW_W_i(8) => wb2reg_8_port, FW_W_i(7)
                           => wb2reg_7_port, FW_W_i(6) => wb2reg_6_port, 
                           FW_W_i(5) => wb2reg_5_port, FW_W_i(4) => 
                           wb2reg_4_port, FW_W_i(3) => wb2reg_3_port, FW_W_i(2)
                           => wb2reg_2_port, FW_W_i(1) => wb2reg_1_port, 
                           FW_W_i(0) => wb2reg_0_port, S_FW_A_i(1) => 
                           dummy_S_FWA2exe_1_port, S_FW_A_i(0) => 
                           dummy_S_FWA2exe_0_port, S_FW_B_i(1) => 
                           dummy_S_FWB2exe_1_port, S_FW_B_i(0) => 
                           dummy_S_FWB2exe_0_port, muxed_dest(4) => 
                           muxed_dest2exe_4_port, muxed_dest(3) => 
                           muxed_dest2exe_3_port, muxed_dest(2) => 
                           muxed_dest2exe_2_port, muxed_dest(1) => 
                           muxed_dest2exe_1_port, muxed_dest(0) => 
                           muxed_dest2exe_0_port, muxed_B(31) => S2mem_31_port,
                           muxed_B(30) => S2mem_30_port, muxed_B(29) => 
                           S2mem_29_port, muxed_B(28) => S2mem_28_port, 
                           muxed_B(27) => S2mem_27_port, muxed_B(26) => 
                           S2mem_26_port, muxed_B(25) => S2mem_25_port, 
                           muxed_B(24) => S2mem_24_port, muxed_B(23) => 
                           S2mem_23_port, muxed_B(22) => S2mem_22_port, 
                           muxed_B(21) => S2mem_21_port, muxed_B(20) => 
                           S2mem_20_port, muxed_B(19) => S2mem_19_port, 
                           muxed_B(18) => S2mem_18_port, muxed_B(17) => 
                           S2mem_17_port, muxed_B(16) => S2mem_16_port, 
                           muxed_B(15) => S2mem_15_port, muxed_B(14) => 
                           S2mem_14_port, muxed_B(13) => S2mem_13_port, 
                           muxed_B(12) => S2mem_12_port, muxed_B(11) => 
                           S2mem_11_port, muxed_B(10) => S2mem_10_port, 
                           muxed_B(9) => S2mem_9_port, muxed_B(8) => 
                           S2mem_8_port, muxed_B(7) => S2mem_7_port, muxed_B(6)
                           => S2mem_6_port, muxed_B(5) => S2mem_5_port, 
                           muxed_B(4) => S2mem_4_port, muxed_B(3) => n5, 
                           muxed_B(2) => S2mem_2_port, muxed_B(1) => 
                           S2mem_1_port, muxed_B(0) => S2mem_0_port, 
                           S_MUX_DEST_i(1) => dummy_S_MUX_DEST_1_port, 
                           S_MUX_DEST_i(0) => dummy_S_MUX_DEST_0_port, OP(0) =>
                           n23, OP(1) => n24, OP(2) => n25, OP(3) => n26, OP(4)
                           => n27, ALUW_i(12) => ALUW_12_port, ALUW_i(11) => 
                           ALUW_11_port, ALUW_i(10) => ALUW_10_port, ALUW_i(9) 
                           => ALUW_9_port, ALUW_i(8) => ALUW_8_port, ALUW_i(7) 
                           => ALUW_7_port, ALUW_i(6) => ALUW_6_port, ALUW_i(5) 
                           => ALUW_5_port, ALUW_i(4) => ALUW_4_port, ALUW_i(3) 
                           => ALUW_3_port, ALUW_i(2) => ALUW_2_port, ALUW_i(1) 
                           => ALUW_1_port, ALUW_i(0) => ALUW_0_port, DOUT(31) 
                           => X2mem_31_port, DOUT(30) => X2mem_30_port, 
                           DOUT(29) => X2mem_29_port, DOUT(28) => X2mem_28_port
                           , DOUT(27) => X2mem_27_port, DOUT(26) => 
                           X2mem_26_port, DOUT(25) => X2mem_25_port, DOUT(24) 
                           => X2mem_24_port, DOUT(23) => X2mem_23_port, 
                           DOUT(22) => X2mem_22_port, DOUT(21) => X2mem_21_port
                           , DOUT(20) => X2mem_20_port, DOUT(19) => 
                           X2mem_19_port, DOUT(18) => X2mem_18_port, DOUT(17) 
                           => X2mem_17_port, DOUT(16) => X2mem_16_port, 
                           DOUT(15) => X2mem_15_port, DOUT(14) => X2mem_14_port
                           , DOUT(13) => X2mem_13_port, DOUT(12) => 
                           X2mem_12_port, DOUT(11) => X2mem_11_port, DOUT(10) 
                           => X2mem_10_port, DOUT(9) => X2mem_9_port, DOUT(8) 
                           => X2mem_8_port, DOUT(7) => X2mem_7_port, DOUT(6) =>
                           X2mem_6_port, DOUT(5) => X2mem_5_port, DOUT(4) => 
                           X2mem_4_port, DOUT(3) => X2mem_3_port, DOUT(2) => 
                           X2mem_2_port, DOUT(1) => X2mem_1_port, DOUT(0) => 
                           X2mem_0_port, stall_o => exe_stall_cu, Clock => 
                           clock, Reset => rst);
   UMEM_REGS : mem_regs port map( W_i(31) => W2wb_31_port, W_i(30) => 
                           W2wb_30_port, W_i(29) => W2wb_29_port, W_i(28) => 
                           W2wb_28_port, W_i(27) => W2wb_27_port, W_i(26) => 
                           W2wb_26_port, W_i(25) => W2wb_25_port, W_i(24) => 
                           W2wb_24_port, W_i(23) => W2wb_23_port, W_i(22) => 
                           W2wb_22_port, W_i(21) => W2wb_21_port, W_i(20) => 
                           W2wb_20_port, W_i(19) => W2wb_19_port, W_i(18) => 
                           W2wb_18_port, W_i(17) => W2wb_17_port, W_i(16) => 
                           W2wb_16_port, W_i(15) => W2wb_15_port, W_i(14) => 
                           W2wb_14_port, W_i(13) => W2wb_13_port, W_i(12) => 
                           W2wb_12_port, W_i(11) => W2wb_11_port, W_i(10) => 
                           W2wb_10_port, W_i(9) => W2wb_9_port, W_i(8) => 
                           W2wb_8_port, W_i(7) => W2wb_7_port, W_i(6) => 
                           W2wb_6_port, W_i(5) => W2wb_5_port, W_i(4) => 
                           W2wb_4_port, W_i(3) => W2wb_3_port, W_i(2) => 
                           W2wb_2_port, W_i(1) => W2wb_1_port, W_i(0) => 
                           W2wb_0_port, D3_i(4) => n7, D3_i(3) => n8, D3_i(2) 
                           => n9, D3_i(1) => n11, D3_i(0) => n10, W_o(31) => 
                           wb2reg_31_port, W_o(30) => wb2reg_30_port, W_o(29) 
                           => wb2reg_29_port, W_o(28) => wb2reg_28_port, 
                           W_o(27) => wb2reg_27_port, W_o(26) => wb2reg_26_port
                           , W_o(25) => wb2reg_25_port, W_o(24) => 
                           wb2reg_24_port, W_o(23) => wb2reg_23_port, W_o(22) 
                           => wb2reg_22_port, W_o(21) => wb2reg_21_port, 
                           W_o(20) => wb2reg_20_port, W_o(19) => wb2reg_19_port
                           , W_o(18) => wb2reg_18_port, W_o(17) => 
                           wb2reg_17_port, W_o(16) => wb2reg_16_port, W_o(15) 
                           => wb2reg_15_port, W_o(14) => wb2reg_14_port, 
                           W_o(13) => wb2reg_13_port, W_o(12) => wb2reg_12_port
                           , W_o(11) => wb2reg_11_port, W_o(10) => 
                           wb2reg_10_port, W_o(9) => wb2reg_9_port, W_o(8) => 
                           wb2reg_8_port, W_o(7) => wb2reg_7_port, W_o(6) => 
                           wb2reg_6_port, W_o(5) => wb2reg_5_port, W_o(4) => 
                           wb2reg_4_port, W_o(3) => wb2reg_3_port, W_o(2) => 
                           wb2reg_2_port, W_o(1) => wb2reg_1_port, W_o(0) => 
                           wb2reg_0_port, D3_o(4) => D32reg_4_port, D3_o(3) => 
                           D32reg_3_port, D3_o(2) => D32reg_2_port, D3_o(1) => 
                           D32reg_1_port, D3_o(0) => D32reg_0_port, clk => 
                           clock, rst => rst);
   UMEM_BLOCK : mem_block port map( X_i(31) => DRAM_Addr_o_31_port, X_i(30) => 
                           DRAM_Addr_o_30_port, X_i(29) => DRAM_Addr_o_29_port,
                           X_i(28) => DRAM_Addr_o_28_port, X_i(27) => 
                           DRAM_Addr_o_27_port, X_i(26) => DRAM_Addr_o_26_port,
                           X_i(25) => DRAM_Addr_o_25_port, X_i(24) => 
                           DRAM_Addr_o_24_port, X_i(23) => DRAM_Addr_o_23_port,
                           X_i(22) => DRAM_Addr_o_22_port, X_i(21) => 
                           DRAM_Addr_o_21_port, X_i(20) => DRAM_Addr_o_20_port,
                           X_i(19) => DRAM_Addr_o_19_port, X_i(18) => 
                           DRAM_Addr_o_18_port, X_i(17) => DRAM_Addr_o_17_port,
                           X_i(16) => DRAM_Addr_o_16_port, X_i(15) => 
                           DRAM_Addr_o_15_port, X_i(14) => DRAM_Addr_o_14_port,
                           X_i(13) => DRAM_Addr_o_13_port, X_i(12) => 
                           DRAM_Addr_o_12_port, X_i(11) => DRAM_Addr_o_11_port,
                           X_i(10) => DRAM_Addr_o_10_port, X_i(9) => 
                           DRAM_Addr_o_9_port, X_i(8) => DRAM_Addr_o_8_port, 
                           X_i(7) => DRAM_Addr_o_7_port, X_i(6) => 
                           DRAM_Addr_o_6_port, X_i(5) => DRAM_Addr_o_5_port, 
                           X_i(4) => DRAM_Addr_o_4_port, X_i(3) => 
                           DRAM_Addr_o_3_port, X_i(2) => DRAM_Addr_o_2_port, 
                           X_i(1) => DRAM_Addr_o_1_port, X_i(0) => 
                           DRAM_Addr_o_0_port, LOAD_i(31) => DRAM_Dout_i(31), 
                           LOAD_i(30) => DRAM_Dout_i(30), LOAD_i(29) => 
                           DRAM_Dout_i(29), LOAD_i(28) => DRAM_Dout_i(28), 
                           LOAD_i(27) => DRAM_Dout_i(27), LOAD_i(26) => 
                           DRAM_Dout_i(26), LOAD_i(25) => DRAM_Dout_i(25), 
                           LOAD_i(24) => DRAM_Dout_i(24), LOAD_i(23) => 
                           DRAM_Dout_i(23), LOAD_i(22) => DRAM_Dout_i(22), 
                           LOAD_i(21) => DRAM_Dout_i(21), LOAD_i(20) => 
                           DRAM_Dout_i(20), LOAD_i(19) => DRAM_Dout_i(19), 
                           LOAD_i(18) => DRAM_Dout_i(18), LOAD_i(17) => 
                           DRAM_Dout_i(17), LOAD_i(16) => DRAM_Dout_i(16), 
                           LOAD_i(15) => DRAM_Dout_i(15), LOAD_i(14) => 
                           DRAM_Dout_i(14), LOAD_i(13) => DRAM_Dout_i(13), 
                           LOAD_i(12) => DRAM_Dout_i(12), LOAD_i(11) => 
                           DRAM_Dout_i(11), LOAD_i(10) => DRAM_Dout_i(10), 
                           LOAD_i(9) => DRAM_Dout_i(9), LOAD_i(8) => 
                           DRAM_Dout_i(8), LOAD_i(7) => DRAM_Dout_i(7), 
                           LOAD_i(6) => DRAM_Dout_i(6), LOAD_i(5) => 
                           DRAM_Dout_i(5), LOAD_i(4) => DRAM_Dout_i(4), 
                           LOAD_i(3) => DRAM_Dout_i(3), LOAD_i(2) => 
                           DRAM_Dout_i(2), LOAD_i(1) => DRAM_Dout_i(1), 
                           LOAD_i(0) => DRAM_Dout_i(0), S_MUX_MEM_i => 
                           dummy_S_MUX_MEM, W_o(31) => W2wb_31_port, W_o(30) =>
                           W2wb_30_port, W_o(29) => W2wb_29_port, W_o(28) => 
                           W2wb_28_port, W_o(27) => W2wb_27_port, W_o(26) => 
                           W2wb_26_port, W_o(25) => W2wb_25_port, W_o(24) => 
                           W2wb_24_port, W_o(23) => W2wb_23_port, W_o(22) => 
                           W2wb_22_port, W_o(21) => W2wb_21_port, W_o(20) => 
                           W2wb_20_port, W_o(19) => W2wb_19_port, W_o(18) => 
                           W2wb_18_port, W_o(17) => W2wb_17_port, W_o(16) => 
                           W2wb_16_port, W_o(15) => W2wb_15_port, W_o(14) => 
                           W2wb_14_port, W_o(13) => W2wb_13_port, W_o(12) => 
                           W2wb_12_port, W_o(11) => W2wb_11_port, W_o(10) => 
                           W2wb_10_port, W_o(9) => W2wb_9_port, W_o(8) => 
                           W2wb_8_port, W_o(7) => W2wb_7_port, W_o(6) => 
                           W2wb_6_port, W_o(5) => W2wb_5_port, W_o(4) => 
                           W2wb_4_port, W_o(3) => W2wb_3_port, W_o(2) => 
                           W2wb_2_port, W_o(1) => W2wb_1_port, W_o(0) => 
                           W2wb_0_port);
   UFW_LOGIC : fw_logic port map( D1_i(4) => n28, D1_i(3) => n29, D1_i(2) => 
                           n30, D1_i(1) => n31, D1_i(0) => n32, rAdec_i(4) => 
                           IR_25_port, rAdec_i(3) => IR_24_port, rAdec_i(2) => 
                           IR_23_port, rAdec_i(1) => IR_22_port, rAdec_i(0) => 
                           IR_21_port, D2_i(4) => D22D3_4_port, D2_i(3) => 
                           D22D3_3_port, D2_i(2) => D22D3_2_port, D2_i(1) => 
                           D22D3_1_port, D2_i(0) => D22D3_0_port, D3_i(4) => 
                           D32reg_4_port, D3_i(3) => D32reg_3_port, D3_i(2) => 
                           D32reg_2_port, D3_i(1) => D32reg_1_port, D3_i(0) => 
                           D32reg_0_port, rA_i(4) => rA2fw_4_port, rA_i(3) => 
                           rA2fw_3_port, rA_i(2) => rA2fw_2_port, rA_i(1) => 
                           rA2fw_1_port, rA_i(0) => rA2fw_0_port, rB_i(4) => 
                           rB2mux_4_port, rB_i(3) => rB2mux_3_port, rB_i(2) => 
                           rB2mux_2_port, rB_i(1) => rB2mux_1_port, rB_i(0) => 
                           rB2mux_0_port, S_mem_W => dummy_S_RF_W_mem, 
                           S_mem_LOAD => dummy_S_MUX_MEM, S_wb_W => 
                           dummy_S_RF_W_wb, S_exe_W => n33, S_FWAdec(1) => 
                           dummy_S_FWAdec_1_port, S_FWAdec(0) => 
                           dummy_S_FWAdec_0_port, S_FWA(1) => 
                           dummy_S_FWA2exe_1_port, S_FWA(0) => 
                           dummy_S_FWA2exe_0_port, S_FWB(1) => 
                           dummy_S_FWB2exe_1_port, S_FWB(0) => 
                           dummy_S_FWB2exe_0_port);
   U5 : INV_X1 port map( A => stall_decode, ZN => enable_regfile);
   U4 : AOI21_X1 port map( B1 => was_taken_from_jl, B2 => was_branch, A => 
                           was_jmp, ZN => n3);
   U6 : INV_X2 port map( A => n3, ZN => was_taken);
   U7 : BUF_X1 port map( A => D22D3_4_port, Z => n7);
   U8 : BUF_X1 port map( A => D22D3_1_port, Z => n11);
   U9 : BUF_X1 port map( A => D22D3_2_port, Z => n9);
   U10 : BUF_X1 port map( A => D22D3_0_port, Z => n10);
   U11 : BUF_X1 port map( A => D22D3_3_port, Z => n8);
   n12 <= '0';
   n13 <= '0';
   n14 <= '0';
   n15 <= '0';
   n16 <= '0';
   n17 <= '0';
   n18 <= '0';
   n19 <= '0';
   n20 <= '0';
   n21 <= '0';
   n22 <= '0';
   n23 <= '0';
   n24 <= '0';
   n25 <= '0';
   n26 <= '0';
   n27 <= '0';
   n28 <= '0';
   n29 <= '0';
   n30 <= '0';
   n31 <= '0';
   n32 <= '0';
   n33 <= '0';

end SYN_arch;
