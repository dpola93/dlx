
module mux21_4 ( IN0, IN1, CTRL, OUT1 );
  input [31:0] IN0;
  input [31:0] IN1;
  output [31:0] OUT1;
  input CTRL;


  MUX2_X1 U1 ( .A(IN0[9]), .B(IN1[9]), .S(CTRL), .Z(OUT1[9]) );
  MUX2_X1 U2 ( .A(IN0[8]), .B(IN1[8]), .S(CTRL), .Z(OUT1[8]) );
  MUX2_X1 U3 ( .A(IN0[7]), .B(IN1[7]), .S(CTRL), .Z(OUT1[7]) );
  MUX2_X1 U4 ( .A(IN0[6]), .B(IN1[6]), .S(CTRL), .Z(OUT1[6]) );
  MUX2_X1 U5 ( .A(IN0[5]), .B(IN1[5]), .S(CTRL), .Z(OUT1[5]) );
  MUX2_X1 U6 ( .A(IN0[4]), .B(IN1[4]), .S(CTRL), .Z(OUT1[4]) );
  MUX2_X1 U7 ( .A(IN0[3]), .B(IN1[3]), .S(CTRL), .Z(OUT1[3]) );
  MUX2_X1 U8 ( .A(IN0[31]), .B(IN1[31]), .S(CTRL), .Z(OUT1[31]) );
  MUX2_X1 U9 ( .A(IN0[30]), .B(IN1[30]), .S(CTRL), .Z(OUT1[30]) );
  MUX2_X1 U10 ( .A(IN0[2]), .B(IN1[2]), .S(CTRL), .Z(OUT1[2]) );
  MUX2_X1 U11 ( .A(IN0[29]), .B(IN1[29]), .S(CTRL), .Z(OUT1[29]) );
  MUX2_X1 U12 ( .A(IN0[28]), .B(IN1[28]), .S(CTRL), .Z(OUT1[28]) );
  MUX2_X1 U13 ( .A(IN0[27]), .B(IN1[27]), .S(CTRL), .Z(OUT1[27]) );
  MUX2_X1 U14 ( .A(IN0[26]), .B(IN1[26]), .S(CTRL), .Z(OUT1[26]) );
  MUX2_X1 U15 ( .A(IN0[25]), .B(IN1[25]), .S(CTRL), .Z(OUT1[25]) );
  MUX2_X1 U16 ( .A(IN0[24]), .B(IN1[24]), .S(CTRL), .Z(OUT1[24]) );
  MUX2_X1 U17 ( .A(IN0[23]), .B(IN1[23]), .S(CTRL), .Z(OUT1[23]) );
  MUX2_X1 U18 ( .A(IN0[22]), .B(IN1[22]), .S(CTRL), .Z(OUT1[22]) );
  MUX2_X1 U19 ( .A(IN0[21]), .B(IN1[21]), .S(CTRL), .Z(OUT1[21]) );
  MUX2_X1 U20 ( .A(IN0[20]), .B(IN1[20]), .S(CTRL), .Z(OUT1[20]) );
  MUX2_X1 U21 ( .A(IN0[1]), .B(IN1[1]), .S(CTRL), .Z(OUT1[1]) );
  MUX2_X1 U22 ( .A(IN0[19]), .B(IN1[19]), .S(CTRL), .Z(OUT1[19]) );
  MUX2_X1 U23 ( .A(IN0[18]), .B(IN1[18]), .S(CTRL), .Z(OUT1[18]) );
  MUX2_X1 U24 ( .A(IN0[17]), .B(IN1[17]), .S(CTRL), .Z(OUT1[17]) );
  MUX2_X1 U25 ( .A(IN0[16]), .B(IN1[16]), .S(CTRL), .Z(OUT1[16]) );
  MUX2_X1 U26 ( .A(IN0[15]), .B(IN1[15]), .S(CTRL), .Z(OUT1[15]) );
  MUX2_X1 U27 ( .A(IN0[14]), .B(IN1[14]), .S(CTRL), .Z(OUT1[14]) );
  MUX2_X1 U28 ( .A(IN0[13]), .B(IN1[13]), .S(CTRL), .Z(OUT1[13]) );
  MUX2_X1 U29 ( .A(IN0[12]), .B(IN1[12]), .S(CTRL), .Z(OUT1[12]) );
  MUX2_X1 U30 ( .A(IN0[11]), .B(IN1[11]), .S(CTRL), .Z(OUT1[11]) );
  MUX2_X1 U31 ( .A(IN0[10]), .B(IN1[10]), .S(CTRL), .Z(OUT1[10]) );
  MUX2_X1 U32 ( .A(IN0[0]), .B(IN1[0]), .S(CTRL), .Z(OUT1[0]) );
endmodule


module mux21_3 ( IN0, IN1, OUT1, CTRL_BAR );
  input [31:0] IN0;
  input [31:0] IN1;
  output [31:0] OUT1;
  input CTRL_BAR;
  wire   CTRL, n1, n2, n3;
  assign CTRL = CTRL_BAR;

  MUX2_X1 U32 ( .A(IN0[0]), .B(IN1[0]), .S(n1), .Z(OUT1[0]) );
  MUX2_X1 U9 ( .A(IN0[30]), .B(IN1[30]), .S(n2), .Z(OUT1[30]) );
  MUX2_X1 U11 ( .A(IN0[29]), .B(IN1[29]), .S(n2), .Z(OUT1[29]) );
  MUX2_X1 U12 ( .A(IN0[28]), .B(IN1[28]), .S(n2), .Z(OUT1[28]) );
  MUX2_X1 U8 ( .A(IN0[31]), .B(IN1[31]), .S(n2), .Z(OUT1[31]) );
  MUX2_X1 U15 ( .A(IN0[25]), .B(IN1[25]), .S(n3), .Z(OUT1[25]) );
  MUX2_X1 U26 ( .A(IN0[15]), .B(IN1[15]), .S(n1), .Z(OUT1[15]) );
  MUX2_X1 U27 ( .A(IN0[14]), .B(IN1[14]), .S(n1), .Z(OUT1[14]) );
  MUX2_X1 U1 ( .A(IN0[9]), .B(IN1[9]), .S(n2), .Z(OUT1[9]) );
  MUX2_X1 U28 ( .A(IN0[13]), .B(IN1[13]), .S(n1), .Z(OUT1[13]) );
  MUX2_X1 U24 ( .A(IN0[17]), .B(IN1[17]), .S(n3), .Z(OUT1[17]) );
  MUX2_X1 U10 ( .A(IN0[2]), .B(IN1[2]), .S(n2), .Z(OUT1[2]) );
  MUX2_X1 U29 ( .A(IN0[12]), .B(IN1[12]), .S(n1), .Z(OUT1[12]) );
  MUX2_X1 U31 ( .A(IN0[10]), .B(IN1[10]), .S(n1), .Z(OUT1[10]) );
  MUX2_X1 U30 ( .A(IN0[11]), .B(IN1[11]), .S(n1), .Z(OUT1[11]) );
  MUX2_X1 U7 ( .A(IN0[3]), .B(IN1[3]), .S(n2), .Z(OUT1[3]) );
  MUX2_X1 U22 ( .A(IN0[19]), .B(IN1[19]), .S(n3), .Z(OUT1[19]) );
  MUX2_X1 U20 ( .A(IN0[20]), .B(IN1[20]), .S(n3), .Z(OUT1[20]) );
  MUX2_X1 U23 ( .A(IN0[18]), .B(IN1[18]), .S(n3), .Z(OUT1[18]) );
  MUX2_X1 U16 ( .A(IN0[24]), .B(IN1[24]), .S(n3), .Z(OUT1[24]) );
  MUX2_X1 U19 ( .A(IN0[21]), .B(IN1[21]), .S(n3), .Z(OUT1[21]) );
  MUX2_X1 U25 ( .A(IN0[16]), .B(IN1[16]), .S(n1), .Z(OUT1[16]) );
  MUX2_X1 U2 ( .A(IN0[8]), .B(IN1[8]), .S(n2), .Z(OUT1[8]) );
  MUX2_X1 U4 ( .A(IN0[6]), .B(IN1[6]), .S(n2), .Z(OUT1[6]) );
  MUX2_X1 U18 ( .A(IN0[22]), .B(IN1[22]), .S(n3), .Z(OUT1[22]) );
  MUX2_X1 U13 ( .A(IN0[27]), .B(IN1[27]), .S(n3), .Z(OUT1[27]) );
  MUX2_X1 U17 ( .A(IN0[23]), .B(IN1[23]), .S(n3), .Z(OUT1[23]) );
  MUX2_X1 U5 ( .A(IN0[5]), .B(IN1[5]), .S(n2), .Z(OUT1[5]) );
  MUX2_X1 U21 ( .A(IN0[1]), .B(IN1[1]), .S(n3), .Z(OUT1[1]) );
  MUX2_X1 U6 ( .A(IN0[4]), .B(IN1[4]), .S(n2), .Z(OUT1[4]) );
  MUX2_X1 U3 ( .A(IN0[7]), .B(IN1[7]), .S(n2), .Z(OUT1[7]) );
  MUX2_X1 U14 ( .A(IN0[26]), .B(IN1[26]), .S(n3), .Z(OUT1[26]) );
  INV_X1 U33 ( .A(CTRL), .ZN(n1) );
  INV_X1 U34 ( .A(CTRL), .ZN(n3) );
  INV_X1 U35 ( .A(CTRL), .ZN(n2) );
endmodule


module FA_47 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n10, n11, n12;

  XNOR2_X1 U1 ( .A(Ci), .B(n12), .ZN(S) );
  NAND2_X1 U3 ( .A1(n11), .A2(n10), .ZN(Co) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n12) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n10) );
  OAI21_X1 U5 ( .B1(A), .B2(B), .A(Ci), .ZN(n11) );
endmodule


module FA_96 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n6;

  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n6) );
  XNOR2_X1 U1 ( .A(n6), .B(B), .ZN(S) );
endmodule


module FA_37 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n6;

  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n6) );
  XNOR2_X1 U1 ( .A(n6), .B(B), .ZN(S) );
endmodule


module FA_33 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n6;

  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n6) );
  XNOR2_X1 U1 ( .A(n6), .B(B), .ZN(S) );
endmodule


module FA_111 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(S) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Co) );
endmodule


module FA_103 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(S) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Co) );
endmodule


module FA_95 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(S) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Co) );
endmodule


module FA_87 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(S) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Co) );
endmodule


module FA_79 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(S) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Co) );
endmodule


module FA_71 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(S) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Co) );
endmodule


module FA_56 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(S) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Co) );
endmodule


module FA_48 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(S) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Co) );
endmodule


module FA_40 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(S) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Co) );
endmodule


module FA_32 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(S) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Co) );
endmodule


module FA_24 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(S) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Co) );
endmodule


module FA_16 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(S) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Co) );
endmodule


module FA_8 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(S) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Co) );
endmodule


module FA_115 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(S) );
  OR2_X1 U2 ( .A1(A), .A2(B), .ZN(Co) );
endmodule


module FA_107 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(S) );
  OR2_X1 U2 ( .A1(A), .A2(B), .ZN(Co) );
endmodule


module FA_99 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(S) );
  OR2_X1 U2 ( .A1(A), .A2(B), .ZN(Co) );
endmodule


module FA_91 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(S) );
  OR2_X1 U2 ( .A1(A), .A2(B), .ZN(Co) );
endmodule


module FA_83 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(S) );
  OR2_X1 U2 ( .A1(A), .A2(B), .ZN(Co) );
endmodule


module FA_75 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(S) );
  OR2_X1 U2 ( .A1(A), .A2(B), .ZN(Co) );
endmodule


module FA_67 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(S) );
endmodule


module FA_60 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(S) );
endmodule


module FA_52 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(S) );
  OR2_X1 U2 ( .A1(A), .A2(B), .ZN(Co) );
endmodule


module FA_44 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(S) );
endmodule


module FA_36 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Co) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(S) );
endmodule


module FA_28 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(S) );
  OR2_X1 U2 ( .A1(A), .A2(B), .ZN(Co) );
endmodule


module FA_20 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(S) );
  OR2_X1 U2 ( .A1(A), .A2(B), .ZN(Co) );
endmodule


module FA_12 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(S) );
  OR2_X1 U2 ( .A1(A), .A2(B), .ZN(Co) );
endmodule


module FA_4 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(S) );
  OR2_X1 U2 ( .A1(A), .A2(B), .ZN(Co) );
endmodule


module FA_125 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11;

  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n11) );
  XNOR2_X1 U1 ( .A(Ci), .B(n11), .ZN(S) );
  OAI21_X1 U5 ( .B1(A), .B2(B), .A(Ci), .ZN(n10) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n9) );
  NAND2_X1 U3 ( .A1(n10), .A2(n9), .ZN(Co) );
endmodule


module FA_118 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11;

  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n11) );
  XNOR2_X1 U1 ( .A(Ci), .B(n11), .ZN(S) );
  OAI21_X1 U5 ( .B1(A), .B2(B), .A(Ci), .ZN(n10) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n9) );
  NAND2_X1 U3 ( .A1(n10), .A2(n9), .ZN(Co) );
endmodule


module FA_117 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11;

  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n11) );
  XNOR2_X1 U1 ( .A(Ci), .B(n11), .ZN(S) );
  OAI21_X1 U5 ( .B1(A), .B2(B), .A(Ci), .ZN(n10) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n9) );
  NAND2_X1 U3 ( .A1(n10), .A2(n9), .ZN(Co) );
endmodule


module FA_114 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11;

  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n11) );
  XNOR2_X1 U1 ( .A(Ci), .B(n11), .ZN(S) );
  OAI21_X1 U5 ( .B1(A), .B2(B), .A(Ci), .ZN(n10) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n9) );
  NAND2_X1 U3 ( .A1(n10), .A2(n9), .ZN(Co) );
endmodule


module FA_113 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11;

  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n11) );
  XNOR2_X1 U1 ( .A(Ci), .B(n11), .ZN(S) );
  OAI21_X1 U5 ( .B1(A), .B2(B), .A(Ci), .ZN(n10) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n9) );
  NAND2_X1 U3 ( .A1(n10), .A2(n9), .ZN(Co) );
endmodule


module FA_109 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11;

  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n11) );
  XNOR2_X1 U1 ( .A(Ci), .B(n11), .ZN(S) );
  OAI21_X1 U5 ( .B1(A), .B2(B), .A(Ci), .ZN(n10) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n9) );
  NAND2_X1 U3 ( .A1(n10), .A2(n9), .ZN(Co) );
endmodule


module FA_106 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11;

  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n11) );
  XNOR2_X1 U1 ( .A(Ci), .B(n11), .ZN(S) );
  OAI21_X1 U5 ( .B1(A), .B2(B), .A(Ci), .ZN(n10) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n9) );
  NAND2_X1 U3 ( .A1(n10), .A2(n9), .ZN(Co) );
endmodule


module FA_105 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11;

  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n11) );
  XNOR2_X1 U1 ( .A(Ci), .B(n11), .ZN(S) );
  OAI21_X1 U5 ( .B1(A), .B2(B), .A(Ci), .ZN(n10) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n9) );
  NAND2_X1 U3 ( .A1(n10), .A2(n9), .ZN(Co) );
endmodule


module FA_102 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11;

  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n11) );
  XNOR2_X1 U1 ( .A(Ci), .B(n11), .ZN(S) );
  OAI21_X1 U5 ( .B1(A), .B2(B), .A(Ci), .ZN(n10) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n9) );
  NAND2_X1 U3 ( .A1(n10), .A2(n9), .ZN(Co) );
endmodule


module FA_101 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11;

  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n11) );
  XNOR2_X1 U1 ( .A(Ci), .B(n11), .ZN(S) );
  OAI21_X1 U5 ( .B1(A), .B2(B), .A(Ci), .ZN(n10) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n9) );
  NAND2_X1 U3 ( .A1(n10), .A2(n9), .ZN(Co) );
endmodule


module FA_98 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11;

  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n11) );
  XNOR2_X1 U1 ( .A(Ci), .B(n11), .ZN(S) );
  OAI21_X1 U5 ( .B1(A), .B2(B), .A(Ci), .ZN(n10) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n9) );
  NAND2_X1 U3 ( .A1(n10), .A2(n9), .ZN(Co) );
endmodule


module FA_97 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11;

  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n11) );
  XNOR2_X1 U1 ( .A(Ci), .B(n11), .ZN(S) );
  OAI21_X1 U5 ( .B1(A), .B2(B), .A(Ci), .ZN(n10) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n9) );
  NAND2_X1 U3 ( .A1(n10), .A2(n9), .ZN(Co) );
endmodule


module FA_94 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11;

  NAND2_X1 U3 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U1 ( .A(Ci), .B(n11), .ZN(S) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n11) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n9) );
  OAI21_X1 U5 ( .B1(A), .B2(B), .A(Ci), .ZN(n10) );
endmodule


module FA_93 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11;

  XNOR2_X1 U1 ( .A(Ci), .B(n11), .ZN(S) );
  NAND2_X1 U3 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n11) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n9) );
  OAI21_X1 U5 ( .B1(A), .B2(B), .A(Ci), .ZN(n10) );
endmodule


module FA_90 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11;

  NAND2_X1 U3 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U1 ( .A(Ci), .B(n11), .ZN(S) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n11) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n9) );
  OAI21_X1 U5 ( .B1(A), .B2(B), .A(Ci), .ZN(n10) );
endmodule


module FA_89 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11;

  XNOR2_X1 U1 ( .A(Ci), .B(n11), .ZN(S) );
  NAND2_X1 U3 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n11) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n9) );
  OAI21_X1 U5 ( .B1(A), .B2(B), .A(Ci), .ZN(n10) );
endmodule


module FA_86 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11;

  XNOR2_X1 U1 ( .A(Ci), .B(n11), .ZN(S) );
  NAND2_X1 U3 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n11) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n9) );
  OAI21_X1 U5 ( .B1(A), .B2(B), .A(Ci), .ZN(n10) );
endmodule


module FA_85 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11;

  XNOR2_X1 U1 ( .A(Ci), .B(n11), .ZN(S) );
  NAND2_X1 U3 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n11) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n9) );
  OAI21_X1 U5 ( .B1(A), .B2(B), .A(Ci), .ZN(n10) );
endmodule


module FA_82 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11;

  XNOR2_X1 U1 ( .A(Ci), .B(n11), .ZN(S) );
  NAND2_X1 U3 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n11) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n9) );
  OAI21_X1 U5 ( .B1(A), .B2(B), .A(Ci), .ZN(n10) );
endmodule


module FA_81 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11;

  XNOR2_X1 U1 ( .A(Ci), .B(n11), .ZN(S) );
  NAND2_X1 U3 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n11) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n9) );
  OAI21_X1 U5 ( .B1(A), .B2(B), .A(Ci), .ZN(n10) );
endmodule


module FA_78 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11;

  XNOR2_X1 U1 ( .A(Ci), .B(n11), .ZN(S) );
  NAND2_X1 U3 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n11) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n9) );
  OAI21_X1 U5 ( .B1(A), .B2(B), .A(Ci), .ZN(n10) );
endmodule


module FA_77 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11;

  XNOR2_X1 U1 ( .A(Ci), .B(n11), .ZN(S) );
  NAND2_X1 U3 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n11) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n9) );
  OAI21_X1 U5 ( .B1(A), .B2(B), .A(Ci), .ZN(n10) );
endmodule


module FA_74 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11;

  XNOR2_X1 U1 ( .A(Ci), .B(n11), .ZN(S) );
  NAND2_X1 U3 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n11) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n9) );
  OAI21_X1 U5 ( .B1(A), .B2(B), .A(Ci), .ZN(n10) );
endmodule


module FA_73 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11;

  XNOR2_X1 U1 ( .A(Ci), .B(n11), .ZN(S) );
  NAND2_X1 U3 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n11) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n9) );
  OAI21_X1 U5 ( .B1(A), .B2(B), .A(Ci), .ZN(n10) );
endmodule


module FA_70 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11;

  NAND2_X1 U3 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U1 ( .A(Ci), .B(n11), .ZN(S) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n11) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n9) );
  OAI21_X1 U5 ( .B1(A), .B2(B), .A(Ci), .ZN(n10) );
endmodule


module FA_69 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11;

  NAND2_X1 U3 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U1 ( .A(Ci), .B(n11), .ZN(S) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n11) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n9) );
  OAI21_X1 U5 ( .B1(A), .B2(B), .A(Ci), .ZN(n10) );
endmodule


module FA_66 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11;

  NAND2_X1 U3 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U1 ( .A(Ci), .B(n11), .ZN(S) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n11) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n9) );
  OAI21_X1 U5 ( .B1(A), .B2(B), .A(Ci), .ZN(n10) );
endmodule


module FA_65 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11;

  NAND2_X1 U3 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U1 ( .A(Ci), .B(n11), .ZN(S) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n11) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n9) );
  OAI21_X1 U5 ( .B1(A), .B2(B), .A(Ci), .ZN(n10) );
endmodule


module FA_63 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11;

  NAND2_X1 U3 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U1 ( .A(Ci), .B(n11), .ZN(S) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n11) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n9) );
  OAI21_X1 U5 ( .B1(A), .B2(B), .A(Ci), .ZN(n10) );
endmodule


module FA_62 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11;

  NAND2_X1 U3 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U1 ( .A(Ci), .B(n11), .ZN(S) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n11) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n9) );
  OAI21_X1 U5 ( .B1(A), .B2(B), .A(Ci), .ZN(n10) );
endmodule


module FA_59 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11;

  NAND2_X1 U3 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U1 ( .A(Ci), .B(n11), .ZN(S) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n11) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n9) );
  OAI21_X1 U5 ( .B1(A), .B2(B), .A(Ci), .ZN(n10) );
endmodule


module FA_58 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11;

  NAND2_X1 U3 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U1 ( .A(Ci), .B(n11), .ZN(S) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n11) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n9) );
  OAI21_X1 U5 ( .B1(A), .B2(B), .A(Ci), .ZN(n10) );
endmodule


module FA_55 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11;

  XNOR2_X1 U1 ( .A(Ci), .B(n11), .ZN(S) );
  NAND2_X1 U3 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n11) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n9) );
  OAI21_X1 U5 ( .B1(A), .B2(B), .A(Ci), .ZN(n10) );
endmodule


module FA_54 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11;

  NAND2_X1 U3 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U1 ( .A(Ci), .B(n11), .ZN(S) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n11) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n9) );
  OAI21_X1 U5 ( .B1(A), .B2(B), .A(Ci), .ZN(n10) );
endmodule


module FA_51 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11;

  XNOR2_X1 U1 ( .A(Ci), .B(n11), .ZN(S) );
  NAND2_X1 U3 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n11) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n9) );
  OAI21_X1 U5 ( .B1(A), .B2(B), .A(Ci), .ZN(n10) );
endmodule


module FA_50 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11;

  NAND2_X1 U3 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U1 ( .A(Ci), .B(n11), .ZN(S) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n11) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n9) );
  OAI21_X1 U5 ( .B1(A), .B2(B), .A(Ci), .ZN(n10) );
endmodule


module FA_46 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11;

  NAND2_X1 U3 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U1 ( .A(Ci), .B(n11), .ZN(S) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n11) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n9) );
  OAI21_X1 U5 ( .B1(A), .B2(B), .A(Ci), .ZN(n10) );
endmodule


module FA_43 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11;

  XNOR2_X1 U1 ( .A(Ci), .B(n11), .ZN(S) );
  NAND2_X1 U3 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n11) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n9) );
  OAI21_X1 U5 ( .B1(A), .B2(B), .A(Ci), .ZN(n10) );
endmodule


module FA_42 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11;

  NAND2_X1 U3 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U1 ( .A(Ci), .B(n11), .ZN(S) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n11) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n9) );
  OAI21_X1 U5 ( .B1(A), .B2(B), .A(Ci), .ZN(n10) );
endmodule


module FA_39 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11;

  NAND2_X1 U3 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U1 ( .A(Ci), .B(n11), .ZN(S) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n9) );
  XNOR2_X1 U4 ( .A(B), .B(A), .ZN(n11) );
  OAI21_X1 U5 ( .B1(A), .B2(B), .A(Ci), .ZN(n10) );
endmodule


module FA_38 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11;

  NAND2_X1 U3 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U1 ( .A(Ci), .B(n11), .ZN(S) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n11) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n9) );
  OAI21_X1 U5 ( .B1(A), .B2(B), .A(Ci), .ZN(n10) );
endmodule


module FA_35 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11;

  NAND2_X1 U3 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U1 ( .A(Ci), .B(n11), .ZN(S) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n9) );
  XNOR2_X1 U4 ( .A(B), .B(A), .ZN(n11) );
  OAI21_X1 U5 ( .B1(A), .B2(B), .A(Ci), .ZN(n10) );
endmodule


module FA_34 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11;

  NAND2_X1 U3 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U1 ( .A(Ci), .B(n11), .ZN(S) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n11) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n9) );
  OAI21_X1 U5 ( .B1(A), .B2(B), .A(Ci), .ZN(n10) );
endmodule


module FA_31 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11;

  NAND2_X1 U3 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U1 ( .A(Ci), .B(n11), .ZN(S) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n11) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n9) );
  OAI21_X1 U5 ( .B1(A), .B2(B), .A(Ci), .ZN(n10) );
endmodule


module FA_30 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11;

  OAI21_X1 U5 ( .B1(A), .B2(B), .A(Ci), .ZN(n10) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n9) );
  NAND2_X1 U3 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n11) );
  XNOR2_X1 U1 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_27 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11;

  NAND2_X1 U3 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U1 ( .A(Ci), .B(n11), .ZN(S) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n11) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n9) );
  OAI21_X1 U5 ( .B1(A), .B2(B), .A(Ci), .ZN(n10) );
endmodule


module FA_26 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11;

  OAI21_X1 U5 ( .B1(A), .B2(B), .A(Ci), .ZN(n10) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n9) );
  NAND2_X1 U3 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n11) );
  XNOR2_X1 U1 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_23 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11;

  OAI21_X1 U5 ( .B1(A), .B2(B), .A(Ci), .ZN(n10) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n9) );
  NAND2_X1 U3 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n11) );
  XNOR2_X1 U1 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_22 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11;

  NAND2_X1 U3 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U1 ( .A(Ci), .B(n11), .ZN(S) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n11) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n9) );
  OAI21_X1 U5 ( .B1(A), .B2(B), .A(Ci), .ZN(n10) );
endmodule


module FA_19 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11;

  OAI21_X1 U5 ( .B1(A), .B2(B), .A(Ci), .ZN(n10) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n9) );
  NAND2_X1 U3 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n11) );
  XNOR2_X1 U1 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_18 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11;

  NAND2_X1 U3 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U1 ( .A(Ci), .B(n11), .ZN(S) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n11) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n9) );
  OAI21_X1 U5 ( .B1(A), .B2(B), .A(Ci), .ZN(n10) );
endmodule


module FA_15 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11;

  OAI21_X1 U5 ( .B1(A), .B2(B), .A(Ci), .ZN(n10) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n9) );
  NAND2_X1 U3 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n11) );
  XNOR2_X1 U1 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_14 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11;

  NAND2_X1 U3 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U1 ( .A(Ci), .B(n11), .ZN(S) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n11) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n9) );
  OAI21_X1 U5 ( .B1(A), .B2(B), .A(Ci), .ZN(n10) );
endmodule


module FA_11 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11;

  OAI21_X1 U5 ( .B1(A), .B2(B), .A(Ci), .ZN(n10) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n9) );
  NAND2_X1 U3 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n11) );
  XNOR2_X1 U1 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_10 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11;

  NAND2_X1 U3 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U1 ( .A(Ci), .B(n11), .ZN(S) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n11) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n9) );
  OAI21_X1 U5 ( .B1(A), .B2(B), .A(Ci), .ZN(n10) );
endmodule


module FA_7 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11;

  OAI21_X1 U5 ( .B1(A), .B2(B), .A(Ci), .ZN(n10) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n9) );
  NAND2_X1 U3 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n11) );
  XNOR2_X1 U1 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_6 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11;

  OAI21_X1 U5 ( .B1(A), .B2(B), .A(Ci), .ZN(n10) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n9) );
  NAND2_X1 U3 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n11) );
  XNOR2_X1 U1 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_3 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11;

  OAI21_X1 U5 ( .B1(A), .B2(B), .A(Ci), .ZN(n10) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n9) );
  NAND2_X1 U3 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n11) );
  XNOR2_X1 U1 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_2 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11;

  OAI21_X1 U5 ( .B1(A), .B2(B), .A(Ci), .ZN(n10) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n9) );
  NAND2_X1 U3 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n11) );
  XNOR2_X1 U1 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_116 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5;

  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n5) );
  XNOR2_X1 U1 ( .A(n5), .B(B), .ZN(S) );
endmodule


module FA_112 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5;

  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n5) );
  XNOR2_X1 U1 ( .A(n5), .B(B), .ZN(S) );
endmodule


module FA_108 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5;

  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n5) );
  XNOR2_X1 U1 ( .A(n5), .B(B), .ZN(S) );
endmodule


module FA_104 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5;

  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n5) );
  XNOR2_X1 U1 ( .A(n5), .B(B), .ZN(S) );
endmodule


module FA_92 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n6;

  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n6) );
  XNOR2_X1 U1 ( .A(n6), .B(B), .ZN(S) );
endmodule


module FA_88 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n6;

  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n6) );
  XNOR2_X1 U1 ( .A(n6), .B(B), .ZN(S) );
endmodule


module FA_84 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5;

  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n5) );
  XNOR2_X1 U1 ( .A(n5), .B(B), .ZN(S) );
endmodule


module FA_80 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5;

  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n5) );
  XNOR2_X1 U1 ( .A(n5), .B(B), .ZN(S) );
endmodule


module FA_76 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5;

  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n5) );
  XNOR2_X1 U1 ( .A(n5), .B(B), .ZN(S) );
endmodule


module FA_72 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5;

  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n5) );
  XNOR2_X1 U1 ( .A(n5), .B(B), .ZN(S) );
endmodule


module FA_68 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5;

  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n5) );
  XNOR2_X1 U1 ( .A(n5), .B(B), .ZN(S) );
endmodule


module FA_64 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5;

  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n5) );
  XNOR2_X1 U1 ( .A(n5), .B(B), .ZN(S) );
endmodule


module FA_61 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5;

  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n5) );
  XNOR2_X1 U1 ( .A(n5), .B(B), .ZN(S) );
endmodule


module FA_57 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5;

  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n5) );
  XNOR2_X1 U1 ( .A(n5), .B(B), .ZN(S) );
endmodule


module FA_53 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5;

  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n5) );
  XNOR2_X1 U1 ( .A(n5), .B(B), .ZN(S) );
endmodule


module FA_49 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5;

  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n5) );
  XNOR2_X1 U1 ( .A(n5), .B(B), .ZN(S) );
endmodule


module FA_45 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5;

  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n5) );
  XNOR2_X1 U1 ( .A(n5), .B(B), .ZN(S) );
endmodule


module FA_41 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5;

  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n5) );
  XNOR2_X1 U1 ( .A(n5), .B(B), .ZN(S) );
endmodule


module FA_29 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5;

  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n5) );
  XNOR2_X1 U1 ( .A(n5), .B(B), .ZN(S) );
endmodule


module FA_25 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5;

  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n5) );
  XNOR2_X1 U1 ( .A(n5), .B(B), .ZN(S) );
endmodule


module FA_21 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5;

  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n5) );
  XNOR2_X1 U1 ( .A(n5), .B(B), .ZN(S) );
endmodule


module FA_17 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5;

  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n5) );
  XNOR2_X1 U1 ( .A(n5), .B(B), .ZN(S) );
endmodule


module FA_13 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5;

  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n5) );
  XNOR2_X1 U1 ( .A(n5), .B(B), .ZN(S) );
endmodule


module FA_9 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5;

  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n5) );
  XNOR2_X1 U1 ( .A(n5), .B(B), .ZN(S) );
endmodule


module FA_5 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n5) );
  XNOR2_X1 U2 ( .A(Ci), .B(n5), .ZN(S) );
endmodule


module FA_1 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n5;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n5) );
  XNOR2_X1 U2 ( .A(Ci), .B(n5), .ZN(S) );
endmodule


module mux21_SIZE4_13 ( IN0, IN1, CTRL, OUT1 );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] OUT1;
  input CTRL;


  MUX2_X1 U1 ( .A(IN0[3]), .B(IN1[3]), .S(CTRL), .Z(OUT1[3]) );
  MUX2_X1 U2 ( .A(IN0[2]), .B(IN1[2]), .S(CTRL), .Z(OUT1[2]) );
  MUX2_X1 U3 ( .A(IN0[1]), .B(IN1[1]), .S(CTRL), .Z(OUT1[1]) );
  MUX2_X1 U4 ( .A(IN0[0]), .B(IN1[0]), .S(CTRL), .Z(OUT1[0]) );
endmodule


module mux21_SIZE4_12 ( IN0, IN1, CTRL, OUT1 );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] OUT1;
  input CTRL;


  MUX2_X1 U1 ( .A(IN0[3]), .B(IN1[3]), .S(CTRL), .Z(OUT1[3]) );
  MUX2_X1 U2 ( .A(IN0[2]), .B(IN1[2]), .S(CTRL), .Z(OUT1[2]) );
  MUX2_X1 U3 ( .A(IN0[1]), .B(IN1[1]), .S(CTRL), .Z(OUT1[1]) );
  MUX2_X1 U4 ( .A(IN0[0]), .B(IN1[0]), .S(CTRL), .Z(OUT1[0]) );
endmodule


module mux21_SIZE4_11 ( IN0, IN1, CTRL, OUT1 );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] OUT1;
  input CTRL;


  MUX2_X1 U1 ( .A(IN0[3]), .B(IN1[3]), .S(CTRL), .Z(OUT1[3]) );
  MUX2_X1 U2 ( .A(IN0[2]), .B(IN1[2]), .S(CTRL), .Z(OUT1[2]) );
  MUX2_X1 U3 ( .A(IN0[1]), .B(IN1[1]), .S(CTRL), .Z(OUT1[1]) );
  MUX2_X1 U4 ( .A(IN0[0]), .B(IN1[0]), .S(CTRL), .Z(OUT1[0]) );
endmodule


module mux21_SIZE4_10 ( IN0, IN1, CTRL, OUT1 );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] OUT1;
  input CTRL;


  MUX2_X1 U1 ( .A(IN0[3]), .B(IN1[3]), .S(CTRL), .Z(OUT1[3]) );
  MUX2_X1 U2 ( .A(IN0[2]), .B(IN1[2]), .S(CTRL), .Z(OUT1[2]) );
  MUX2_X1 U3 ( .A(IN0[1]), .B(IN1[1]), .S(CTRL), .Z(OUT1[1]) );
  MUX2_X1 U4 ( .A(IN0[0]), .B(IN1[0]), .S(CTRL), .Z(OUT1[0]) );
endmodule


module mux21_SIZE4_9 ( IN0, IN1, CTRL, OUT1 );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] OUT1;
  input CTRL;


  MUX2_X1 U1 ( .A(IN0[3]), .B(IN1[3]), .S(CTRL), .Z(OUT1[3]) );
  MUX2_X1 U3 ( .A(IN0[1]), .B(IN1[1]), .S(CTRL), .Z(OUT1[1]) );
  MUX2_X1 U4 ( .A(IN0[0]), .B(IN1[0]), .S(CTRL), .Z(OUT1[0]) );
  MUX2_X1 U2 ( .A(IN0[2]), .B(IN1[2]), .S(CTRL), .Z(OUT1[2]) );
endmodule


module mux21_SIZE4_8 ( IN0, IN1, CTRL, OUT1 );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] OUT1;
  input CTRL;


  MUX2_X1 U1 ( .A(IN0[3]), .B(IN1[3]), .S(CTRL), .Z(OUT1[3]) );
  MUX2_X1 U2 ( .A(IN0[2]), .B(IN1[2]), .S(CTRL), .Z(OUT1[2]) );
  MUX2_X1 U3 ( .A(IN0[1]), .B(IN1[1]), .S(CTRL), .Z(OUT1[1]) );
  MUX2_X1 U4 ( .A(IN0[0]), .B(IN1[0]), .S(CTRL), .Z(OUT1[0]) );
endmodule


module mux21_SIZE4_7 ( IN0, IN1, CTRL, OUT1 );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] OUT1;
  input CTRL;


  MUX2_X1 U1 ( .A(IN0[3]), .B(IN1[3]), .S(CTRL), .Z(OUT1[3]) );
  MUX2_X1 U2 ( .A(IN0[2]), .B(IN1[2]), .S(CTRL), .Z(OUT1[2]) );
  MUX2_X1 U3 ( .A(IN0[1]), .B(IN1[1]), .S(CTRL), .Z(OUT1[1]) );
  MUX2_X1 U4 ( .A(IN0[0]), .B(IN1[0]), .S(CTRL), .Z(OUT1[0]) );
endmodule


module mux21_SIZE4_6 ( IN0, IN1, CTRL, OUT1 );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] OUT1;
  input CTRL;


  MUX2_X1 U1 ( .A(IN0[3]), .B(IN1[3]), .S(CTRL), .Z(OUT1[3]) );
  MUX2_X1 U2 ( .A(IN0[2]), .B(IN1[2]), .S(CTRL), .Z(OUT1[2]) );
  MUX2_X1 U3 ( .A(IN0[1]), .B(IN1[1]), .S(CTRL), .Z(OUT1[1]) );
  MUX2_X1 U4 ( .A(IN0[0]), .B(IN1[0]), .S(CTRL), .Z(OUT1[0]) );
endmodule


module mux21_SIZE4_5 ( IN0, IN1, CTRL, OUT1 );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] OUT1;
  input CTRL;


  MUX2_X1 U1 ( .A(IN0[3]), .B(IN1[3]), .S(CTRL), .Z(OUT1[3]) );
  MUX2_X1 U2 ( .A(IN0[2]), .B(IN1[2]), .S(CTRL), .Z(OUT1[2]) );
  MUX2_X1 U3 ( .A(IN0[1]), .B(IN1[1]), .S(CTRL), .Z(OUT1[1]) );
  MUX2_X1 U4 ( .A(IN0[0]), .B(IN1[0]), .S(CTRL), .Z(OUT1[0]) );
endmodule


module mux21_SIZE4_4 ( IN0, IN1, CTRL, OUT1 );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] OUT1;
  input CTRL;


  MUX2_X1 U1 ( .A(IN0[3]), .B(IN1[3]), .S(CTRL), .Z(OUT1[3]) );
  MUX2_X1 U2 ( .A(IN0[2]), .B(IN1[2]), .S(CTRL), .Z(OUT1[2]) );
  MUX2_X1 U3 ( .A(IN0[1]), .B(IN1[1]), .S(CTRL), .Z(OUT1[1]) );
  MUX2_X1 U4 ( .A(IN0[0]), .B(IN1[0]), .S(CTRL), .Z(OUT1[0]) );
endmodule


module mux21_SIZE4_3 ( IN0, IN1, CTRL, OUT1 );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] OUT1;
  input CTRL;


  MUX2_X1 U1 ( .A(IN0[3]), .B(IN1[3]), .S(CTRL), .Z(OUT1[3]) );
  MUX2_X1 U2 ( .A(IN0[2]), .B(IN1[2]), .S(CTRL), .Z(OUT1[2]) );
  MUX2_X1 U3 ( .A(IN0[1]), .B(IN1[1]), .S(CTRL), .Z(OUT1[1]) );
  MUX2_X1 U4 ( .A(IN0[0]), .B(IN1[0]), .S(CTRL), .Z(OUT1[0]) );
endmodule


module mux21_SIZE4_2 ( IN0, IN1, CTRL, OUT1 );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] OUT1;
  input CTRL;


  MUX2_X1 U1 ( .A(IN0[3]), .B(IN1[3]), .S(CTRL), .Z(OUT1[3]) );
  MUX2_X1 U2 ( .A(IN0[2]), .B(IN1[2]), .S(CTRL), .Z(OUT1[2]) );
  MUX2_X1 U3 ( .A(IN0[0]), .B(IN1[0]), .S(CTRL), .Z(OUT1[0]) );
  MUX2_X1 U4 ( .A(IN0[1]), .B(IN1[1]), .S(CTRL), .Z(OUT1[1]) );
endmodule


module mux21_SIZE4_1 ( IN0, IN1, CTRL, OUT1 );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] OUT1;
  input CTRL;


  MUX2_X1 U2 ( .A(IN0[2]), .B(IN1[2]), .S(CTRL), .Z(OUT1[2]) );
  MUX2_X1 U1 ( .A(IN0[0]), .B(IN1[0]), .S(CTRL), .Z(OUT1[0]) );
  MUX2_X1 U3 ( .A(IN0[3]), .B(IN1[3]), .S(CTRL), .Z(OUT1[3]) );
  MUX2_X1 U4 ( .A(IN0[1]), .B(IN1[1]), .S(CTRL), .Z(OUT1[1]) );
endmodule


module RCA_N4_12 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;
  wire   n1;
  wire   [3:1] CTMP;

  FA_48 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(1'b0), .S(S[0]), .Co(n1) );
  FA_47 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(n1), .S(S[1]), .Co(CTMP[2]) );
  FA_46 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_45 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module RCA_N4_10 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_40 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(1'b0), .S(S[0]), .Co(CTMP[1]) );
  FA_39 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_38 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_37 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module RCA_N4_9 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_36 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(1'b1), .S(S[0]), .Co(CTMP[1]) );
  FA_35 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_34 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_33 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module RCA_N4_23 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_95 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(1'b0), .S(S[0]), .Co(CTMP[1]) );
  FA_94 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_93 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_92 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module RCA_N4_21 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_87 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(1'b0), .S(S[0]), .Co(CTMP[1]) );
  FA_86 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_85 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_84 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module RCA_N4_19 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_79 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(1'b0), .S(S[0]), .Co(CTMP[1]) );
  FA_78 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_77 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_76 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module RCA_N4_17 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_71 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(1'b0), .S(S[0]), .Co(CTMP[1]) );
  FA_70 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_69 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_68 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module RCA_N4_14 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_56 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(1'b0), .S(S[0]), .Co(CTMP[1]) );
  FA_55 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_54 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_53 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module RCA_N4_8 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_32 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(1'b0), .S(S[0]), .Co(CTMP[1]) );
  FA_31 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_30 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_29 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module RCA_N4_6 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_24 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(1'b0), .S(S[0]), .Co(CTMP[1]) );
  FA_23 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_22 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_21 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module RCA_N4_4 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_16 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(1'b0), .S(S[0]), .Co(CTMP[1]) );
  FA_15 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_14 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_13 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module RCA_N4_2 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_8 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(1'b0), .S(S[0]), .Co(CTMP[1]) );
  FA_7 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_6 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_5 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module RCA_N4_28 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_115 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(1'b1), .S(S[0]), .Co(CTMP[1]) );
  FA_114 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_113 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_112 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module RCA_N4_26 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_107 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(1'b1), .S(S[0]), .Co(CTMP[1]) );
  FA_106 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_105 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_104 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module RCA_N4_22 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_91 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(1'b1), .S(S[0]), .Co(CTMP[1]) );
  FA_90 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_89 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_88 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module RCA_N4_20 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_83 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(1'b1), .S(S[0]), .Co(CTMP[1]) );
  FA_82 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_81 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_80 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module RCA_N4_18 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_75 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(1'b1), .S(S[0]), .Co(CTMP[1]) );
  FA_74 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_73 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_72 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module RCA_N4_16 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_67 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(1'b1), .S(S[0]), .Co(CTMP[1]) );
  FA_66 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_65 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_64 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module RCA_N4_15 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_60 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(1'b1), .S(S[0]), .Co(CTMP[1]) );
  FA_59 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_58 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_57 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module RCA_N4_13 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_52 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(1'b1), .S(S[0]), .Co(CTMP[1]) );
  FA_51 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_50 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_49 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module RCA_N4_11 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_44 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(1'b1), .S(S[0]), .Co(CTMP[1]) );
  FA_43 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_42 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_41 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module RCA_N4_7 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_28 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(1'b1), .S(S[0]), .Co(CTMP[1]) );
  FA_27 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_26 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_25 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module RCA_N4_5 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_20 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(1'b1), .S(S[0]), .Co(CTMP[1]) );
  FA_19 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_18 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_17 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module RCA_N4_3 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_12 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(1'b1), .S(S[0]), .Co(CTMP[1]) );
  FA_11 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_10 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_9 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module RCA_N4_1 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_4 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(1'b1), .S(S[0]), .Co(CTMP[1]) );
  FA_3 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_2 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module carry_sel_gen_N4_6 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:0] nocarry_sum_to_mux;
  wire   [3:0] carry_sum_to_mux;

  RCA_N4_12 rca_nocarry ( .A(A), .B(B), .Ci(1'b0), .S(nocarry_sum_to_mux) );
  RCA_N4_11 rca_carry ( .A(A), .B(B), .Ci(1'b1), .S(carry_sum_to_mux) );
  mux21_SIZE4_6 outmux ( .IN0(nocarry_sum_to_mux), .IN1(carry_sum_to_mux), 
        .CTRL(Ci), .OUT1(S) );
endmodule


module carry_sel_gen_N4_5 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:0] nocarry_sum_to_mux;
  wire   [3:0] carry_sum_to_mux;

  RCA_N4_10 rca_nocarry ( .A(A), .B(B), .Ci(1'b0), .S(nocarry_sum_to_mux) );
  RCA_N4_9 rca_carry ( .A(A), .B(B), .Ci(1'b1), .S(carry_sum_to_mux) );
  mux21_SIZE4_5 outmux ( .IN0(nocarry_sum_to_mux), .IN1(carry_sum_to_mux), 
        .CTRL(Ci), .OUT1(S) );
endmodule


module carry_sel_gen_N4_4 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:0] nocarry_sum_to_mux;
  wire   [3:0] carry_sum_to_mux;

  RCA_N4_8 rca_nocarry ( .A(A), .B(B), .Ci(1'b0), .S(nocarry_sum_to_mux) );
  RCA_N4_7 rca_carry ( .A(A), .B(B), .Ci(1'b1), .S(carry_sum_to_mux) );
  mux21_SIZE4_4 outmux ( .IN0(nocarry_sum_to_mux), .IN1(carry_sum_to_mux), 
        .CTRL(Ci), .OUT1(S) );
endmodule


module carry_sel_gen_N4_10 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:0] nocarry_sum_to_mux;
  wire   [3:0] carry_sum_to_mux;

  RCA_N4_21 rca_nocarry ( .A(A), .B(B), .Ci(1'b0), .S(nocarry_sum_to_mux) );
  RCA_N4_20 rca_carry ( .A(A), .B(B), .Ci(1'b1), .S(carry_sum_to_mux) );
  mux21_SIZE4_10 outmux ( .IN0(nocarry_sum_to_mux), .IN1(carry_sum_to_mux), 
        .CTRL(Ci), .OUT1(S) );
endmodule


module carry_sel_gen_N4_9 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:0] nocarry_sum_to_mux;
  wire   [3:0] carry_sum_to_mux;

  RCA_N4_19 rca_nocarry ( .A(A), .B(B), .Ci(1'b0), .S(nocarry_sum_to_mux) );
  RCA_N4_18 rca_carry ( .A(A), .B(B), .Ci(1'b1), .S(carry_sum_to_mux) );
  mux21_SIZE4_9 outmux ( .IN0(nocarry_sum_to_mux), .IN1(carry_sum_to_mux), 
        .CTRL(Ci), .OUT1(S) );
endmodule


module carry_sel_gen_N4_8 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:0] nocarry_sum_to_mux;
  wire   [3:0] carry_sum_to_mux;

  RCA_N4_17 rca_nocarry ( .A(A), .B(B), .Ci(1'b0), .S(nocarry_sum_to_mux) );
  RCA_N4_16 rca_carry ( .A(A), .B(B), .Ci(1'b1), .S(carry_sum_to_mux) );
  mux21_SIZE4_8 outmux ( .IN0(nocarry_sum_to_mux), .IN1(carry_sum_to_mux), 
        .CTRL(Ci), .OUT1(S) );
endmodule


module carry_sel_gen_N4_7 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:0] nocarry_sum_to_mux;
  wire   [3:0] carry_sum_to_mux;

  RCA_N4_14 rca_nocarry ( .A(A), .B(B), .Ci(1'b0), .S(nocarry_sum_to_mux) );
  RCA_N4_13 rca_carry ( .A(A), .B(B), .Ci(1'b1), .S(carry_sum_to_mux) );
  mux21_SIZE4_7 outmux ( .IN0(nocarry_sum_to_mux), .IN1(carry_sum_to_mux), 
        .CTRL(Ci), .OUT1(S) );
endmodule


module carry_sel_gen_N4_3 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:0] nocarry_sum_to_mux;
  wire   [3:0] carry_sum_to_mux;

  RCA_N4_6 rca_nocarry ( .A(A), .B(B), .Ci(1'b0), .S(nocarry_sum_to_mux) );
  RCA_N4_5 rca_carry ( .A(A), .B(B), .Ci(1'b1), .S(carry_sum_to_mux) );
  mux21_SIZE4_3 outmux ( .IN0(nocarry_sum_to_mux), .IN1(carry_sum_to_mux), 
        .CTRL(Ci), .OUT1(S) );
endmodule


module carry_sel_gen_N4_2 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:0] nocarry_sum_to_mux;
  wire   [3:0] carry_sum_to_mux;

  RCA_N4_4 rca_nocarry ( .A(A), .B(B), .Ci(1'b0), .S(nocarry_sum_to_mux) );
  RCA_N4_3 rca_carry ( .A(A), .B(B), .Ci(1'b1), .S(carry_sum_to_mux) );
  mux21_SIZE4_2 outmux ( .IN0(nocarry_sum_to_mux), .IN1(carry_sum_to_mux), 
        .CTRL(Ci), .OUT1(S) );
endmodule


module carry_sel_gen_N4_1 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:0] nocarry_sum_to_mux;
  wire   [3:0] carry_sum_to_mux;

  RCA_N4_2 rca_nocarry ( .A(A), .B(B), .Ci(1'b0), .S(nocarry_sum_to_mux) );
  RCA_N4_1 rca_carry ( .A(A), .B(B), .Ci(1'b1), .S(carry_sum_to_mux) );
  mux21_SIZE4_1 outmux ( .IN0(nocarry_sum_to_mux), .IN1(carry_sum_to_mux), 
        .CTRL(Ci), .OUT1(S) );
endmodule


module pg_20 ( g, p, g_prec, p_prec, g_out, p_out );
  input g, p, g_prec, p_prec;
  output g_out, p_out;
  wire   n6, n7;

  INV_X1 U1 ( .A(g), .ZN(n7) );
  AND2_X1 U2 ( .A1(p), .A2(p_prec), .ZN(p_out) );
  NAND2_X1 U3 ( .A1(p), .A2(g_prec), .ZN(n6) );
  NAND2_X1 U4 ( .A1(n6), .A2(n7), .ZN(g_out) );
endmodule


module pg_12 ( p, g_prec, p_prec, g_out, p_out, g_BAR );
  input p, g_prec, p_prec, g_BAR;
  output g_out, p_out;
  wire   g, n5;
  assign g = g_BAR;

  AND2_X1 U1 ( .A1(p), .A2(p_prec), .ZN(p_out) );
  NAND2_X1 U2 ( .A1(p), .A2(g_prec), .ZN(n5) );
  NAND2_X1 U3 ( .A1(n5), .A2(g), .ZN(g_out) );
endmodule


module pg_49 ( g, p, g_prec, p_prec, p_out, g_out_BAR );
  input g, p, g_prec, p_prec;
  output p_out, g_out_BAR;


  AOI21_X1 U2 ( .B1(g_prec), .B2(p), .A(g), .ZN(g_out_BAR) );
  AND2_X1 U1 ( .A1(p), .A2(p_prec), .ZN(p_out) );
endmodule


module pg_47 ( g, p, g_prec, p_prec, p_out, g_out_BAR );
  input g, p, g_prec, p_prec;
  output p_out, g_out_BAR;


  AOI21_X1 U2 ( .B1(g_prec), .B2(p), .A(g), .ZN(g_out_BAR) );
  AND2_X1 U1 ( .A1(p), .A2(p_prec), .ZN(p_out) );
endmodule


module pg_45 ( g, p, g_prec, p_prec, p_out, g_out_BAR );
  input g, p, g_prec, p_prec;
  output p_out, g_out_BAR;


  AOI21_X1 U2 ( .B1(g_prec), .B2(p), .A(g), .ZN(g_out_BAR) );
  AND2_X1 U1 ( .A1(p_prec), .A2(p), .ZN(p_out) );
endmodule


module pg_34 ( g, p, g_prec, p_prec, p_out, g_out_BAR );
  input g, p, g_prec, p_prec;
  output p_out, g_out_BAR;


  AOI21_X1 U2 ( .B1(g_prec), .B2(p), .A(g), .ZN(g_out_BAR) );
  AND2_X1 U1 ( .A1(p_prec), .A2(p), .ZN(p_out) );
endmodule


module pg_25 ( g, p, g_prec, p_prec, p_out, g_out_BAR );
  input g, p, g_prec, p_prec;
  output p_out, g_out_BAR;


  AOI21_X1 U2 ( .B1(p), .B2(g_prec), .A(g), .ZN(g_out_BAR) );
  AND2_X1 U1 ( .A1(p), .A2(p_prec), .ZN(p_out) );
endmodule


module pg_23 ( g, p, g_prec, p_prec, p_out, g_out_BAR );
  input g, p, g_prec, p_prec;
  output p_out, g_out_BAR;


  AOI21_X1 U2 ( .B1(p), .B2(g_prec), .A(g), .ZN(g_out_BAR) );
  AND2_X1 U1 ( .A1(p), .A2(p_prec), .ZN(p_out) );
endmodule


module pg_21 ( g, p, g_prec, p_prec, p_out, g_out_BAR );
  input g, p, g_prec, p_prec;
  output p_out, g_out_BAR;


  AND2_X1 U1 ( .A1(p), .A2(p_prec), .ZN(p_out) );
  AOI21_X1 U2 ( .B1(p), .B2(g_prec), .A(g), .ZN(g_out_BAR) );
endmodule


module pg_19 ( g, p, g_prec, p_prec, p_out, g_out_BAR );
  input g, p, g_prec, p_prec;
  output p_out, g_out_BAR;


  AND2_X1 U1 ( .A1(p_prec), .A2(p), .ZN(p_out) );
  AOI21_X1 U2 ( .B1(g_prec), .B2(p), .A(g), .ZN(g_out_BAR) );
endmodule


module pg_8 ( g, p, g_prec, p_prec, p_out, g_out_BAR );
  input g, p, g_prec, p_prec;
  output p_out, g_out_BAR;


  AND2_X1 U1 ( .A1(p_prec), .A2(p), .ZN(p_out) );
  AOI21_X1 U2 ( .B1(g_prec), .B2(p), .A(g), .ZN(g_out_BAR) );
endmodule


module pg_36 ( p, g_prec, p_prec, g_out, p_out, g_BAR );
  input p, g_prec, p_prec, g_BAR;
  output g_out, p_out;
  wire   g, n4;
  assign g = g_BAR;

  NAND2_X1 U3 ( .A1(p), .A2(g_prec), .ZN(n4) );
  NAND2_X1 U2 ( .A1(g), .A2(n4), .ZN(g_out) );
  AND2_X1 U1 ( .A1(p), .A2(p_prec), .ZN(p_out) );
endmodule


module pg_35 ( p, g_prec, p_prec, g_out, p_out, g_BAR );
  input p, g_prec, p_prec, g_BAR;
  output g_out, p_out;
  wire   g, n4;
  assign g = g_BAR;

  AND2_X1 U1 ( .A1(p), .A2(p_prec), .ZN(p_out) );
  NAND2_X1 U2 ( .A1(g_prec), .A2(p), .ZN(n4) );
  NAND2_X1 U3 ( .A1(n4), .A2(g), .ZN(g_out) );
endmodule


module pg_30 ( p, g_prec, p_prec, g_out, p_out, g_BAR );
  input p, g_prec, p_prec, g_BAR;
  output g_out, p_out;
  wire   g, n4;
  assign g = g_BAR;

  AND2_X1 U1 ( .A1(p), .A2(p_prec), .ZN(p_out) );
  NAND2_X1 U2 ( .A1(g_prec), .A2(p), .ZN(n4) );
  NAND2_X1 U3 ( .A1(n4), .A2(g), .ZN(g_out) );
endmodule


module pg_11 ( p, g_prec, p_prec, g_out, p_out, g_BAR );
  input p, g_prec, p_prec, g_BAR;
  output g_out, p_out;
  wire   g, n4;
  assign g = g_BAR;

  AND2_X1 U1 ( .A1(p), .A2(p_prec), .ZN(p_out) );
  NAND2_X1 U2 ( .A1(g_prec), .A2(p), .ZN(n4) );
  NAND2_X1 U3 ( .A1(n4), .A2(g), .ZN(g_out) );
endmodule


module pg_10 ( p, g_prec, p_prec, g_out, p_out, g_BAR );
  input p, g_prec, p_prec, g_BAR;
  output g_out, p_out;
  wire   g, n4;
  assign g = g_BAR;

  AND2_X1 U1 ( .A1(p), .A2(p_prec), .ZN(p_out) );
  NAND2_X1 U2 ( .A1(p), .A2(g_prec), .ZN(n4) );
  NAND2_X1 U3 ( .A1(n4), .A2(g), .ZN(g_out) );
endmodule


module pg_9 ( p, g_prec, p_prec, g_out, p_out, g_BAR );
  input p, g_prec, p_prec, g_BAR;
  output g_out, p_out;
  wire   g, n4;
  assign g = g_BAR;

  AND2_X1 U1 ( .A1(p), .A2(p_prec), .ZN(p_out) );
  NAND2_X1 U2 ( .A1(g_prec), .A2(p), .ZN(n4) );
  NAND2_X1 U3 ( .A1(n4), .A2(g), .ZN(g_out) );
endmodule


module pg_4 ( p, g_prec, p_prec, g_out, p_out, g_BAR );
  input p, g_prec, p_prec, g_BAR;
  output g_out, p_out;
  wire   g, n4;
  assign g = g_BAR;

  AND2_X1 U1 ( .A1(p), .A2(p_prec), .ZN(p_out) );
  NAND2_X1 U2 ( .A1(p), .A2(g_prec), .ZN(n4) );
  NAND2_X1 U3 ( .A1(n4), .A2(g), .ZN(g_out) );
endmodule


module pg_50 ( g, p, g_prec, p_prec, g_out, p_out );
  input g, p, g_prec, p_prec;
  output g_out, p_out;
  wire   n5;

  AOI21_X1 U3 ( .B1(g_prec), .B2(p), .A(g), .ZN(n5) );
  AND2_X1 U1 ( .A1(p), .A2(p_prec), .ZN(p_out) );
  INV_X1 U2 ( .A(n5), .ZN(g_out) );
endmodule


module pg_48 ( g, p, g_prec, p_prec, g_out, p_out );
  input g, p, g_prec, p_prec;
  output g_out, p_out;
  wire   n5;

  AOI21_X1 U3 ( .B1(g_prec), .B2(p), .A(g), .ZN(n5) );
  AND2_X1 U1 ( .A1(p), .A2(p_prec), .ZN(p_out) );
  INV_X1 U2 ( .A(n5), .ZN(g_out) );
endmodule


module pg_44 ( g, p, g_prec, p_prec, g_out, p_out );
  input g, p, g_prec, p_prec;
  output g_out, p_out;
  wire   n5;

  AOI21_X1 U3 ( .B1(g_prec), .B2(p), .A(g), .ZN(n5) );
  INV_X1 U2 ( .A(n5), .ZN(g_out) );
  AND2_X1 U1 ( .A1(p), .A2(p_prec), .ZN(p_out) );
endmodule


module pg_43 ( g, p, g_prec, p_prec, g_out, p_out );
  input g, p, g_prec, p_prec;
  output g_out, p_out;
  wire   n5;

  AOI21_X1 U3 ( .B1(g_prec), .B2(p), .A(g), .ZN(n5) );
  INV_X1 U2 ( .A(n5), .ZN(g_out) );
  AND2_X1 U1 ( .A1(p_prec), .A2(p), .ZN(p_out) );
endmodule


module pg_42 ( g, p, g_prec, p_prec, g_out, p_out );
  input g, p, g_prec, p_prec;
  output g_out, p_out;
  wire   n5;

  AND2_X1 U1 ( .A1(p), .A2(p_prec), .ZN(p_out) );
  INV_X1 U2 ( .A(n5), .ZN(g_out) );
  AOI21_X1 U3 ( .B1(g_prec), .B2(p), .A(g), .ZN(n5) );
endmodule


module pg_41 ( g, p, g_prec, p_prec, p_out, g_out_BAR );
  input g, p, g_prec, p_prec;
  output p_out, g_out_BAR;


  AND2_X1 U1 ( .A1(p_prec), .A2(p), .ZN(p_out) );
  AOI21_X1 U2 ( .B1(p), .B2(g_prec), .A(g), .ZN(g_out_BAR) );
endmodule


module pg_33 ( p, g_prec, p_prec, g_out, p_out, g_BAR );
  input p, g_prec, p_prec, g_BAR;
  output g_out, p_out;
  wire   g, n5;
  assign g = g_BAR;

  AND2_X1 U1 ( .A1(p), .A2(p_prec), .ZN(p_out) );
  NAND2_X1 U2 ( .A1(g_prec), .A2(p), .ZN(n5) );
  NAND2_X1 U3 ( .A1(n5), .A2(g), .ZN(g_out) );
endmodule


module pg_31 ( g, p, g_prec, p_prec, g_out, p_out );
  input g, p, g_prec, p_prec;
  output g_out, p_out;
  wire   n5;

  AOI21_X1 U3 ( .B1(g_prec), .B2(p), .A(g), .ZN(n5) );
  AND2_X1 U1 ( .A1(p), .A2(p_prec), .ZN(p_out) );
  INV_X1 U2 ( .A(n5), .ZN(g_out) );
endmodule


module pg_28 ( g, p, g_prec, p_prec, g_out, p_out );
  input g, p, g_prec, p_prec;
  output g_out, p_out;
  wire   n5, n6;

  AND2_X1 U1 ( .A1(p_prec), .A2(p), .ZN(p_out) );
  INV_X1 U2 ( .A(g), .ZN(n6) );
  NAND2_X1 U3 ( .A1(g_prec), .A2(p), .ZN(n5) );
  NAND2_X1 U4 ( .A1(n5), .A2(n6), .ZN(g_out) );
endmodule


module pg_26 ( g, p, g_prec, p_prec, g_out, p_out );
  input g, p, g_prec, p_prec;
  output g_out, p_out;
  wire   n5;

  AOI21_X1 U1 ( .B1(g_prec), .B2(p), .A(g), .ZN(n5) );
  INV_X1 U2 ( .A(n5), .ZN(g_out) );
  AND2_X1 U3 ( .A1(p), .A2(p_prec), .ZN(p_out) );
endmodule


module pg_24 ( g, p, g_prec, p_prec, g_out, p_out );
  input g, p, g_prec, p_prec;
  output g_out, p_out;
  wire   n5;

  AOI21_X1 U1 ( .B1(p), .B2(g_prec), .A(g), .ZN(n5) );
  INV_X1 U2 ( .A(n5), .ZN(g_out) );
  AND2_X1 U3 ( .A1(p), .A2(p_prec), .ZN(p_out) );
endmodule


module pg_22 ( g, p, g_prec, p_prec, g_out, p_out );
  input g, p, g_prec, p_prec;
  output g_out, p_out;
  wire   n5, n6;

  INV_X1 U1 ( .A(g), .ZN(n6) );
  AND2_X1 U2 ( .A1(p_prec), .A2(p), .ZN(p_out) );
  NAND2_X1 U3 ( .A1(p), .A2(g_prec), .ZN(n5) );
  NAND2_X1 U4 ( .A1(n5), .A2(n6), .ZN(g_out) );
endmodule


module pg_18 ( g, p, g_prec, p_prec, g_out, p_out );
  input g, p, g_prec, p_prec;
  output g_out, p_out;
  wire   n5;

  AOI21_X1 U3 ( .B1(p), .B2(g_prec), .A(g), .ZN(n5) );
  INV_X1 U1 ( .A(n5), .ZN(g_out) );
  AND2_X1 U2 ( .A1(p), .A2(p_prec), .ZN(p_out) );
endmodule


module pg_17 ( g, p, g_prec, p_prec, g_out, p_out );
  input g, p, g_prec, p_prec;
  output g_out, p_out;
  wire   n5;

  AOI21_X1 U3 ( .B1(p), .B2(g_prec), .A(g), .ZN(n5) );
  INV_X1 U1 ( .A(n5), .ZN(g_out) );
  AND2_X1 U2 ( .A1(p), .A2(p_prec), .ZN(p_out) );
endmodule


module pg_16 ( g, p, g_prec, p_prec, g_out, p_out );
  input g, p, g_prec, p_prec;
  output g_out, p_out;
  wire   n6;

  AOI21_X1 U3 ( .B1(p), .B2(g_prec), .A(g), .ZN(n6) );
  AND2_X1 U1 ( .A1(p), .A2(p_prec), .ZN(p_out) );
  INV_X1 U2 ( .A(n6), .ZN(g_out) );
endmodule


module pg_15 ( g, p, g_prec, p_prec, g_out, p_out );
  input g, p, g_prec, p_prec;
  output g_out, p_out;
  wire   n5;

  AOI21_X1 U3 ( .B1(g_prec), .B2(p), .A(g), .ZN(n5) );
  INV_X1 U1 ( .A(n5), .ZN(g_out) );
  AND2_X1 U2 ( .A1(p_prec), .A2(p), .ZN(p_out) );
endmodule


module pg_14 ( g, p, g_prec, p_prec, g_out, p_out );
  input g, p, g_prec, p_prec;
  output g_out, p_out;
  wire   n5;

  AOI21_X1 U3 ( .B1(g_prec), .B2(p), .A(g), .ZN(n5) );
  AND2_X1 U1 ( .A1(p), .A2(p_prec), .ZN(p_out) );
  INV_X1 U2 ( .A(n5), .ZN(g_out) );
endmodule


module pg_13 ( g, p, g_prec, p_prec, g_out, p_out );
  input g, p, g_prec, p_prec;
  output g_out, p_out;
  wire   n5;

  AOI21_X1 U3 ( .B1(g_prec), .B2(p), .A(g), .ZN(n5) );
  AND2_X1 U1 ( .A1(p), .A2(p_prec), .ZN(p_out) );
  INV_X1 U2 ( .A(n5), .ZN(g_out) );
endmodule


module pg_7 ( g, p, g_prec, p_prec, g_out, p_out );
  input g, p, g_prec, p_prec;
  output g_out, p_out;
  wire   n5;

  AND2_X1 U1 ( .A1(p), .A2(p_prec), .ZN(p_out) );
  INV_X1 U2 ( .A(n5), .ZN(g_out) );
  AOI21_X1 U3 ( .B1(g_prec), .B2(p), .A(g), .ZN(n5) );
endmodule


module pg_6 ( g, p, g_prec, p_prec, g_out, p_out );
  input g, p, g_prec, p_prec;
  output g_out, p_out;
  wire   n5;

  AOI21_X1 U3 ( .B1(g_prec), .B2(p), .A(g), .ZN(n5) );
  AND2_X1 U1 ( .A1(p), .A2(p_prec), .ZN(p_out) );
  INV_X1 U2 ( .A(n5), .ZN(g_out) );
endmodule


module pg_5 ( g, p, g_prec, p_prec, g_out, p_out );
  input g, p, g_prec, p_prec;
  output g_out, p_out;
  wire   n5, n6;

  AND2_X1 U1 ( .A1(p), .A2(p_prec), .ZN(p_out) );
  INV_X1 U2 ( .A(g), .ZN(n6) );
  NAND2_X1 U3 ( .A1(g_prec), .A2(p), .ZN(n5) );
  NAND2_X1 U4 ( .A1(n5), .A2(n6), .ZN(g_out) );
endmodule


module pg_3 ( g, p, g_prec, p_prec, g_out, p_out );
  input g, p, g_prec, p_prec;
  output g_out, p_out;
  wire   n5;

  AOI21_X1 U3 ( .B1(g_prec), .B2(p), .A(g), .ZN(n5) );
  AND2_X1 U1 ( .A1(p), .A2(p_prec), .ZN(p_out) );
  INV_X1 U2 ( .A(n5), .ZN(g_out) );
endmodule


module pg_2 ( g, p, g_prec, p_prec, g_out, p_out );
  input g, p, g_prec, p_prec;
  output g_out, p_out;
  wire   n5, n6;

  AND2_X1 U1 ( .A1(p), .A2(p_prec), .ZN(p_out) );
  INV_X1 U2 ( .A(g), .ZN(n6) );
  NAND2_X1 U3 ( .A1(g_prec), .A2(p), .ZN(n5) );
  NAND2_X1 U4 ( .A1(n5), .A2(n6), .ZN(g_out) );
endmodule


module pg_1 ( g, p, g_prec, p_prec, g_out, p_out );
  input g, p, g_prec, p_prec;
  output g_out, p_out;
  wire   n5;

  AND2_X1 U1 ( .A1(p), .A2(p_prec), .ZN(p_out) );
  INV_X1 U2 ( .A(n5), .ZN(g_out) );
  AOI21_X1 U3 ( .B1(g_prec), .B2(p), .A(g), .ZN(n5) );
endmodule


module g_9 ( g, p, g_prec, g_out );
  input g, p, g_prec;
  output g_out;
  wire   n4;

  AOI21_X1 U1 ( .B1(p), .B2(g_prec), .A(g), .ZN(n4) );
  INV_X1 U2 ( .A(n4), .ZN(g_out) );
endmodule


module g_16 ( g, p, g_prec, g_out );
  input g, p, g_prec;
  output g_out;
  wire   n5;

  AOI21_X1 U2 ( .B1(p), .B2(g_prec), .A(g), .ZN(n5) );
  INV_X1 U1 ( .A(n5), .ZN(g_out) );
endmodule


module g_15 ( g, p, g_prec, g_out );
  input g, p, g_prec;
  output g_out;
  wire   n5;

  AOI21_X1 U2 ( .B1(p), .B2(g_prec), .A(g), .ZN(n5) );
  INV_X1 U1 ( .A(n5), .ZN(g_out) );
endmodule


module g_14 ( g, p, g_prec, g_out );
  input g, p, g_prec;
  output g_out;
  wire   n5;

  AOI21_X1 U2 ( .B1(p), .B2(g_prec), .A(g), .ZN(n5) );
  INV_X1 U1 ( .A(n5), .ZN(g_out) );
endmodule


module g_13 ( g, p, g_prec, g_out );
  input g, p, g_prec;
  output g_out;
  wire   n5;

  INV_X1 U1 ( .A(n5), .ZN(g_out) );
  AOI21_X1 U2 ( .B1(p), .B2(g_prec), .A(g), .ZN(n5) );
endmodule


module g_12 ( g, p, g_prec, g_out );
  input g, p, g_prec;
  output g_out;
  wire   n5;

  AND2_X1 U1 ( .A1(p), .A2(g_prec), .ZN(n5) );
  OR2_X1 U2 ( .A1(g), .A2(n5), .ZN(g_out) );
endmodule


module g_11 ( g, p, g_prec, g_out );
  input g, p, g_prec;
  output g_out;
  wire   n5;

  AND2_X1 U1 ( .A1(p), .A2(g_prec), .ZN(n5) );
  OR2_X2 U2 ( .A1(g), .A2(n5), .ZN(g_out) );
endmodule


module g_8 ( g, p, g_prec, g_out );
  input g, p, g_prec;
  output g_out;
  wire   n5, n6;

  INV_X1 U1 ( .A(g), .ZN(n5) );
  NAND2_X1 U2 ( .A1(n6), .A2(n5), .ZN(g_out) );
  NAND2_X1 U3 ( .A1(g_prec), .A2(p), .ZN(n6) );
endmodule


module g_7 ( g, p, g_prec, g_out );
  input g, p, g_prec;
  output g_out;
  wire   n5, n6;

  NAND2_X1 U1 ( .A1(n6), .A2(n5), .ZN(g_out) );
  INV_X1 U2 ( .A(g), .ZN(n5) );
  NAND2_X1 U3 ( .A1(g_prec), .A2(p), .ZN(n6) );
endmodule


module g_6 ( g, p, g_prec, g_out );
  input g, p, g_prec;
  output g_out;
  wire   n5;

  INV_X1 U1 ( .A(n5), .ZN(g_out) );
  AOI21_X1 U2 ( .B1(p), .B2(g_prec), .A(g), .ZN(n5) );
endmodule


module g_5 ( g, p, g_prec, g_out );
  input g, p, g_prec;
  output g_out;
  wire   n5;

  INV_X1 U1 ( .A(n5), .ZN(g_out) );
  AOI21_X1 U2 ( .B1(g_prec), .B2(p), .A(g), .ZN(n5) );
endmodule


module g_4 ( g, p, g_prec, g_out );
  input g, p, g_prec;
  output g_out;
  wire   n5, n6;

  NAND2_X1 U1 ( .A1(n5), .A2(n6), .ZN(g_out) );
  INV_X1 U2 ( .A(g), .ZN(n6) );
  NAND2_X1 U3 ( .A1(g_prec), .A2(p), .ZN(n5) );
endmodule


module g_3 ( g, p, g_prec, g_out );
  input g, p, g_prec;
  output g_out;
  wire   n5, n6;

  INV_X1 U1 ( .A(g), .ZN(n6) );
  NAND2_X1 U2 ( .A1(n5), .A2(n6), .ZN(g_out) );
  NAND2_X1 U3 ( .A1(g_prec), .A2(p), .ZN(n5) );
endmodule


module g_2 ( g, p, g_prec, g_out );
  input g, p, g_prec;
  output g_out;
  wire   n5;

  INV_X1 U1 ( .A(n5), .ZN(g_out) );
  AOI21_X1 U2 ( .B1(g_prec), .B2(p), .A(g), .ZN(n5) );
endmodule


module g_1 ( g, p, g_prec, g_out );
  input g, p, g_prec;
  output g_out;
  wire   n5;

  INV_X1 U1 ( .A(n5), .ZN(g_out) );
  AOI21_X1 U2 ( .B1(p), .B2(g_prec), .A(g), .ZN(n5) );
endmodule


module pg_net_18 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p_out) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g_out) );
endmodule


module pg_net_61 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p_out) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g_out) );
endmodule


module pg_net_60 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p_out) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g_out) );
endmodule


module pg_net_59 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p_out) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g_out) );
endmodule


module pg_net_58 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p_out) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g_out) );
endmodule


module pg_net_57 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p_out) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g_out) );
endmodule


module pg_net_56 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p_out) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g_out) );
endmodule


module pg_net_55 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p_out) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g_out) );
endmodule


module pg_net_54 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p_out) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g_out) );
endmodule


module pg_net_53 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p_out) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g_out) );
endmodule


module pg_net_52 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p_out) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g_out) );
endmodule


module pg_net_51 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p_out) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g_out) );
endmodule


module pg_net_50 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p_out) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g_out) );
endmodule


module pg_net_48 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p_out) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g_out) );
endmodule


module pg_net_47 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;
  wire   n2;

  INV_X1 U1 ( .A(a), .ZN(n2) );
  AND2_X1 U2 ( .A1(b), .A2(a), .ZN(g_out) );
  XNOR2_X1 U3 ( .A(b), .B(n2), .ZN(p_out) );
endmodule


module pg_net_46 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p_out) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g_out) );
endmodule


module pg_net_45 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p_out) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g_out) );
endmodule


module pg_net_44 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p_out) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g_out) );
endmodule


module pg_net_43 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;
  wire   n2;

  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g_out) );
  INV_X1 U2 ( .A(a), .ZN(n2) );
  XNOR2_X1 U3 ( .A(b), .B(n2), .ZN(p_out) );
endmodule


module pg_net_42 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p_out) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g_out) );
endmodule


module pg_net_41 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;
  wire   n2;

  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g_out) );
  INV_X1 U2 ( .A(a), .ZN(n2) );
  XNOR2_X1 U3 ( .A(b), .B(n2), .ZN(p_out) );
endmodule


module pg_net_40 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p_out) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g_out) );
endmodule


module pg_net_39 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p_out) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g_out) );
endmodule


module pg_net_38 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;


  XOR2_X1 U1 ( .A(a), .B(b), .Z(p_out) );
  AND2_X1 U2 ( .A1(b), .A2(a), .ZN(g_out) );
endmodule


module pg_net_37 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p_out) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g_out) );
endmodule


module pg_net_32 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g_out) );
endmodule


module pg_net_31 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;
  wire   n2;

  INV_X1 U1 ( .A(a), .ZN(n2) );
  AND2_X1 U2 ( .A1(b), .A2(a), .ZN(g_out) );
  XNOR2_X1 U3 ( .A(b), .B(n2), .ZN(p_out) );
endmodule


module pg_net_30 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;


  XOR2_X1 U1 ( .A(a), .B(b), .Z(p_out) );
  AND2_X1 U2 ( .A1(b), .A2(a), .ZN(g_out) );
endmodule


module pg_net_29 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p_out) );
  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g_out) );
endmodule


module pg_net_28 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;
  wire   n2;

  INV_X1 U1 ( .A(a), .ZN(n2) );
  AND2_X1 U2 ( .A1(b), .A2(a), .ZN(g_out) );
  XNOR2_X1 U3 ( .A(b), .B(n2), .ZN(p_out) );
endmodule


module pg_net_27 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;
  wire   n3;

  INV_X1 U1 ( .A(a), .ZN(n3) );
  AND2_X1 U2 ( .A1(b), .A2(a), .ZN(g_out) );
  XNOR2_X1 U3 ( .A(b), .B(n3), .ZN(p_out) );
endmodule


module pg_net_26 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p_out) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g_out) );
endmodule


module pg_net_25 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p_out) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g_out) );
endmodule


module pg_net_24 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p_out) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g_out) );
endmodule


module pg_net_23 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;
  wire   n2;

  INV_X1 U1 ( .A(a), .ZN(n2) );
  AND2_X1 U2 ( .A1(b), .A2(a), .ZN(g_out) );
  XNOR2_X1 U3 ( .A(b), .B(n2), .ZN(p_out) );
endmodule


module pg_net_22 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p_out) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g_out) );
endmodule


module pg_net_21 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p_out) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g_out) );
endmodule


module pg_net_20 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;
  wire   n2;

  INV_X1 U1 ( .A(a), .ZN(n2) );
  AND2_X1 U2 ( .A1(b), .A2(a), .ZN(g_out) );
  XNOR2_X1 U3 ( .A(b), .B(n2), .ZN(p_out) );
endmodule


module pg_net_19 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p_out) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g_out) );
endmodule


module pg_net_17 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p_out) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g_out) );
endmodule


module pg_net_16 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p_out) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g_out) );
endmodule


module pg_net_15 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;


  XOR2_X1 U1 ( .A(a), .B(b), .Z(p_out) );
  AND2_X1 U2 ( .A1(b), .A2(a), .ZN(g_out) );
endmodule


module pg_net_14 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p_out) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g_out) );
endmodule


module pg_net_13 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p_out) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g_out) );
endmodule


module pg_net_12 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;
  wire   n2;

  INV_X1 U1 ( .A(a), .ZN(n2) );
  AND2_X1 U2 ( .A1(b), .A2(a), .ZN(g_out) );
  XNOR2_X1 U3 ( .A(b), .B(n2), .ZN(p_out) );
endmodule


module pg_net_11 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p_out) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g_out) );
endmodule


module pg_net_10 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p_out) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g_out) );
endmodule


module pg_net_9 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p_out) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g_out) );
endmodule


module pg_net_8 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p_out) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g_out) );
endmodule


module pg_net_7 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p_out) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g_out) );
endmodule


module pg_net_6 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p_out) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g_out) );
endmodule


module pg_net_5 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p_out) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g_out) );
endmodule


module pg_net_4 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p_out) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g_out) );
endmodule


module pg_net_3 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p_out) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g_out) );
endmodule


module pg_net_2 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p_out) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g_out) );
endmodule


module pg_net_1 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;
  wire   n2;

  INV_X1 U1 ( .A(a), .ZN(n2) );
  AND2_X1 U2 ( .A1(b), .A2(a), .ZN(g_out) );
  XNOR2_X1 U3 ( .A(b), .B(n2), .ZN(p_out) );
endmodule


module FA_0_1 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(S) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Co) );
endmodule


module mux21_SIZE4_0_1 ( IN0, IN1, CTRL, OUT1 );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] OUT1;
  input CTRL;


  MUX2_X1 U1 ( .A(IN0[3]), .B(IN1[3]), .S(CTRL), .Z(OUT1[3]) );
  MUX2_X1 U2 ( .A(IN0[2]), .B(IN1[2]), .S(CTRL), .Z(OUT1[2]) );
  MUX2_X1 U3 ( .A(IN0[1]), .B(IN1[1]), .S(CTRL), .Z(OUT1[1]) );
  MUX2_X1 U4 ( .A(IN0[0]), .B(IN1[0]), .S(CTRL), .Z(OUT1[0]) );
endmodule


module RCA_N4_0_1 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_0_1 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(1'b0), .S(S[0]), .Co(CTMP[1]) );
  FA_63 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_62 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_61 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module carry_sel_gen_N4_0_1 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:0] nocarry_sum_to_mux;
  wire   [3:0] carry_sum_to_mux;

  RCA_N4_0_1 rca_nocarry ( .A(A), .B(B), .Ci(1'b0), .S(nocarry_sum_to_mux) );
  RCA_N4_15 rca_carry ( .A(A), .B(B), .Ci(1'b1), .S(carry_sum_to_mux) );
  mux21_SIZE4_0_1 outmux ( .IN0(nocarry_sum_to_mux), .IN1(carry_sum_to_mux), 
        .CTRL(Ci), .OUT1(S) );
endmodule


module pg_0_1 ( g, p, g_prec, p_prec, g_out, p_out );
  input g, p, g_prec, p_prec;
  output g_out, p_out;
  wire   n5, n6;

  INV_X1 U1 ( .A(g), .ZN(n6) );
  AND2_X1 U2 ( .A1(p), .A2(p_prec), .ZN(p_out) );
  NAND2_X1 U3 ( .A1(p), .A2(g_prec), .ZN(n5) );
  NAND2_X1 U4 ( .A1(n5), .A2(n6), .ZN(g_out) );
endmodule


module g_0_1 ( g, p, g_prec, g_out );
  input g, p, g_prec;
  output g_out;
  wire   n4;

  AOI21_X1 U1 ( .B1(p), .B2(g_prec), .A(g), .ZN(n4) );
  INV_X1 U2 ( .A(n4), .ZN(g_out) );
endmodule


module pg_net_0_1 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;
  wire   n3;

  INV_X1 U1 ( .A(a), .ZN(n3) );
  AND2_X1 U2 ( .A1(b), .A2(a), .ZN(g_out) );
  XNOR2_X1 U3 ( .A(n3), .B(b), .ZN(p_out) );
endmodule


module sum_gen_N32_1 ( A, B, Cin, S );
  input [31:0] A;
  input [31:0] B;
  input [8:0] Cin;
  output [31:0] S;


  carry_sel_gen_N4_0_1 csel_N_0 ( .A(A[3:0]), .B(B[3:0]), .Ci(Cin[0]), .S(
        S[3:0]) );
  carry_sel_gen_N4_7 csel_N_1 ( .A(A[7:4]), .B(B[7:4]), .Ci(Cin[1]), .S(S[7:4]) );
  carry_sel_gen_N4_6 csel_N_2 ( .A(A[11:8]), .B(B[11:8]), .Ci(Cin[2]), .S(
        S[11:8]) );
  carry_sel_gen_N4_5 csel_N_3 ( .A(A[15:12]), .B(B[15:12]), .Ci(Cin[3]), .S(
        S[15:12]) );
  carry_sel_gen_N4_4 csel_N_4 ( .A(A[19:16]), .B(B[19:16]), .Ci(Cin[4]), .S(
        S[19:16]) );
  carry_sel_gen_N4_3 csel_N_5 ( .A(A[23:20]), .B(B[23:20]), .Ci(Cin[5]), .S(
        S[23:20]) );
  carry_sel_gen_N4_2 csel_N_6 ( .A(A[27:24]), .B(B[27:24]), .Ci(Cin[6]), .S(
        S[27:24]) );
  carry_sel_gen_N4_1 csel_N_7 ( .A(A[31:28]), .B(B[31:28]), .Ci(Cin[7]), .S(
        S[31:28]) );
endmodule


module carry_tree_N32_logN5_1 ( A, B, Cin, Cout );
  input [31:0] A;
  input [31:0] B;
  output [7:0] Cout;
  input Cin;
  wire   \pg_1[15][1] , \pg_1[15][0] , \pg_1[14][1] , \pg_1[14][0] ,
         \pg_1[13][1] , \pg_1[13][0] , \pg_1[12][1] , \pg_1[12][0] ,
         \pg_1[11][1] , \pg_1[11][0] , \pg_1[10][1] , \pg_1[10][0] ,
         \pg_1[9][1] , \pg_1[9][0] , \pg_1[8][1] , \pg_1[8][0] , \pg_1[7][1] ,
         \pg_1[7][0] , \pg_1[6][1] , \pg_1[6][0] , \pg_1[5][1] , \pg_1[5][0] ,
         \pg_1[4][1] , \pg_1[4][0] , \pg_1[3][1] , \pg_1[3][0] , \pg_1[2][1] ,
         \pg_1[2][0] , \pg_1[1][1] , \pg_1[1][0] , \pg_1[0][0] ,
         \pg_n[4][7][1] , \pg_n[4][7][0] , \pg_n[4][6][1] , \pg_n[4][6][0] ,
         \pg_n[3][7][1] , \pg_n[3][7][0] , \pg_n[3][5][1] , \pg_n[3][3][1] ,
         \pg_n[3][3][0] , \pg_n[2][7][1] , \pg_n[2][7][0] , \pg_n[2][6][1] ,
         \pg_n[2][6][0] , \pg_n[2][5][1] , \pg_n[2][5][0] , \pg_n[2][4][1] ,
         \pg_n[2][3][1] , \pg_n[2][3][0] , \pg_n[2][2][1] , \pg_n[2][2][0] ,
         \pg_n[2][1][1] , \pg_n[2][1][0] , n1, n5, n26, n7, n8, n12, n18, n20,
         n22, n23;
  wire   [31:1] p_net;
  wire   [31:0] g_net;
  wire   [1:0] magic_pro;

  pg_net_0_1 pg_net_x_1 ( .a(A[1]), .b(B[1]), .g_out(g_net[1]), .p_out(
        p_net[1]) );
  pg_net_31 pg_net_x_2 ( .a(A[2]), .b(B[2]), .g_out(g_net[2]), .p_out(p_net[2]) );
  pg_net_30 pg_net_x_3 ( .a(A[3]), .b(B[3]), .g_out(g_net[3]), .p_out(p_net[3]) );
  pg_net_29 pg_net_x_4 ( .a(A[4]), .b(B[4]), .g_out(g_net[4]), .p_out(p_net[4]) );
  pg_net_28 pg_net_x_5 ( .a(A[5]), .b(B[5]), .g_out(g_net[5]), .p_out(p_net[5]) );
  pg_net_27 pg_net_x_6 ( .a(A[6]), .b(B[6]), .g_out(g_net[6]), .p_out(p_net[6]) );
  pg_net_26 pg_net_x_7 ( .a(A[7]), .b(B[7]), .g_out(g_net[7]), .p_out(p_net[7]) );
  pg_net_25 pg_net_x_8 ( .a(A[8]), .b(B[8]), .g_out(g_net[8]), .p_out(p_net[8]) );
  pg_net_24 pg_net_x_9 ( .a(A[9]), .b(B[9]), .g_out(g_net[9]), .p_out(p_net[9]) );
  pg_net_23 pg_net_x_10 ( .a(A[10]), .b(B[10]), .g_out(g_net[10]), .p_out(
        p_net[10]) );
  pg_net_22 pg_net_x_11 ( .a(A[11]), .b(B[11]), .g_out(g_net[11]), .p_out(
        p_net[11]) );
  pg_net_21 pg_net_x_12 ( .a(A[12]), .b(B[12]), .g_out(g_net[12]), .p_out(
        p_net[12]) );
  pg_net_20 pg_net_x_13 ( .a(A[13]), .b(B[13]), .g_out(g_net[13]), .p_out(
        p_net[13]) );
  pg_net_19 pg_net_x_14 ( .a(A[14]), .b(B[14]), .g_out(g_net[14]), .p_out(
        p_net[14]) );
  pg_net_18 pg_net_x_15 ( .a(A[15]), .b(B[15]), .g_out(g_net[15]), .p_out(
        p_net[15]) );
  pg_net_17 pg_net_x_16 ( .a(A[16]), .b(B[16]), .g_out(g_net[16]), .p_out(
        p_net[16]) );
  pg_net_16 pg_net_x_17 ( .a(A[17]), .b(B[17]), .g_out(g_net[17]), .p_out(
        p_net[17]) );
  pg_net_15 pg_net_x_18 ( .a(A[18]), .b(B[18]), .g_out(g_net[18]), .p_out(
        p_net[18]) );
  pg_net_14 pg_net_x_19 ( .a(A[19]), .b(B[19]), .g_out(g_net[19]), .p_out(
        p_net[19]) );
  pg_net_13 pg_net_x_20 ( .a(A[20]), .b(B[20]), .g_out(g_net[20]), .p_out(
        p_net[20]) );
  pg_net_12 pg_net_x_21 ( .a(A[21]), .b(B[21]), .g_out(g_net[21]), .p_out(
        p_net[21]) );
  pg_net_11 pg_net_x_22 ( .a(A[22]), .b(B[22]), .g_out(g_net[22]), .p_out(
        p_net[22]) );
  pg_net_10 pg_net_x_23 ( .a(A[23]), .b(B[23]), .g_out(g_net[23]), .p_out(
        p_net[23]) );
  pg_net_9 pg_net_x_24 ( .a(A[24]), .b(B[24]), .g_out(g_net[24]), .p_out(
        p_net[24]) );
  pg_net_8 pg_net_x_25 ( .a(A[25]), .b(B[25]), .g_out(g_net[25]), .p_out(n18)
         );
  pg_net_7 pg_net_x_26 ( .a(A[26]), .b(B[26]), .g_out(g_net[26]), .p_out(
        p_net[26]) );
  pg_net_6 pg_net_x_27 ( .a(A[27]), .b(B[27]), .g_out(g_net[27]), .p_out(
        p_net[27]) );
  pg_net_5 pg_net_x_28 ( .a(A[28]), .b(B[28]), .g_out(g_net[28]), .p_out(
        p_net[28]) );
  pg_net_4 pg_net_x_29 ( .a(A[29]), .b(B[29]), .g_out(g_net[29]), .p_out(
        p_net[29]) );
  pg_net_3 pg_net_x_30 ( .a(A[30]), .b(B[30]), .g_out(g_net[30]), .p_out(
        p_net[30]) );
  pg_net_2 pg_net_x_31 ( .a(A[31]), .b(B[31]), .g_out(g_net[31]), .p_out(
        p_net[31]) );
  pg_net_1 pg_net_0_MAGIC ( .a(A[0]), .b(B[0]), .g_out(magic_pro[0]), .p_out(
        magic_pro[1]) );
  g_0_1 xG_0_0_MAGIC ( .g(magic_pro[0]), .p(magic_pro[1]), .g_prec(Cin), 
        .g_out(g_net[0]) );
  g_9 xG_1_0 ( .g(g_net[1]), .p(p_net[1]), .g_prec(g_net[0]), .g_out(
        \pg_1[0][0] ) );
  pg_0_1 xPG_1_1 ( .g(g_net[3]), .p(p_net[3]), .g_prec(g_net[2]), .p_prec(
        p_net[2]), .g_out(\pg_1[1][0] ), .p_out(\pg_1[1][1] ) );
  pg_26 xPG_1_2 ( .g(g_net[5]), .p(p_net[5]), .g_prec(g_net[4]), .p_prec(
        p_net[4]), .g_out(\pg_1[2][0] ), .p_out(\pg_1[2][1] ) );
  pg_25 xPG_1_3 ( .g(g_net[7]), .p(p_net[7]), .g_prec(g_net[6]), .p_prec(
        p_net[6]), .p_out(\pg_1[3][1] ), .g_out_BAR(\pg_1[3][0] ) );
  pg_24 xPG_1_4 ( .g(g_net[9]), .p(p_net[9]), .g_prec(g_net[8]), .p_prec(
        p_net[8]), .g_out(\pg_1[4][0] ), .p_out(\pg_1[4][1] ) );
  pg_23 xPG_1_5 ( .g(g_net[11]), .p(p_net[11]), .g_prec(g_net[10]), .p_prec(
        p_net[10]), .p_out(\pg_1[5][1] ), .g_out_BAR(\pg_1[5][0] ) );
  pg_22 xPG_1_6 ( .g(g_net[13]), .p(p_net[13]), .g_prec(g_net[12]), .p_prec(
        p_net[12]), .g_out(\pg_1[6][0] ), .p_out(\pg_1[6][1] ) );
  pg_21 xPG_1_7 ( .g(g_net[15]), .p(p_net[15]), .g_prec(g_net[14]), .p_prec(
        p_net[14]), .p_out(\pg_1[7][1] ), .g_out_BAR(\pg_1[7][0] ) );
  pg_20 xPG_1_8 ( .g(g_net[17]), .p(p_net[17]), .g_prec(g_net[16]), .p_prec(
        p_net[16]), .g_out(\pg_1[8][0] ), .p_out(\pg_1[8][1] ) );
  pg_19 xPG_1_9 ( .g(g_net[19]), .p(p_net[19]), .g_prec(g_net[18]), .p_prec(
        p_net[18]), .p_out(\pg_1[9][1] ), .g_out_BAR(\pg_1[9][0] ) );
  pg_18 xPG_1_10 ( .g(g_net[21]), .p(p_net[21]), .g_prec(g_net[20]), .p_prec(
        p_net[20]), .g_out(\pg_1[10][0] ), .p_out(\pg_1[10][1] ) );
  pg_17 xPG_1_11 ( .g(g_net[23]), .p(p_net[23]), .g_prec(g_net[22]), .p_prec(
        p_net[22]), .g_out(\pg_1[11][0] ), .p_out(\pg_1[11][1] ) );
  pg_16 xPG_1_12 ( .g(g_net[25]), .p(n18), .g_prec(g_net[24]), .p_prec(
        p_net[24]), .g_out(\pg_1[12][0] ), .p_out(\pg_1[12][1] ) );
  pg_15 xPG_1_13 ( .g(g_net[27]), .p(p_net[27]), .g_prec(g_net[26]), .p_prec(
        p_net[26]), .g_out(\pg_1[13][0] ), .p_out(\pg_1[13][1] ) );
  pg_14 xPG_1_14 ( .g(g_net[29]), .p(p_net[29]), .g_prec(g_net[28]), .p_prec(
        p_net[28]), .g_out(\pg_1[14][0] ), .p_out(\pg_1[14][1] ) );
  pg_13 xPG_1_15 ( .g(g_net[31]), .p(p_net[31]), .g_prec(g_net[30]), .p_prec(
        p_net[30]), .g_out(\pg_1[15][0] ), .p_out(\pg_1[15][1] ) );
  g_8 xG_2_0 ( .g(\pg_1[1][0] ), .p(\pg_1[1][1] ), .g_prec(\pg_1[0][0] ), 
        .g_out(n26) );
  pg_12 xPG_2_1 ( .p(\pg_1[3][1] ), .g_prec(\pg_1[2][0] ), .p_prec(
        \pg_1[2][1] ), .g_out(\pg_n[2][1][0] ), .p_out(\pg_n[2][1][1] ), 
        .g_BAR(\pg_1[3][0] ) );
  pg_11 xPG_2_2 ( .p(\pg_1[5][1] ), .g_prec(\pg_1[4][0] ), .p_prec(
        \pg_1[4][1] ), .g_out(\pg_n[2][2][0] ), .p_out(\pg_n[2][2][1] ), 
        .g_BAR(\pg_1[5][0] ) );
  pg_10 xPG_2_3 ( .p(\pg_1[7][1] ), .g_prec(\pg_1[6][0] ), .p_prec(
        \pg_1[6][1] ), .g_out(\pg_n[2][3][0] ), .p_out(\pg_n[2][3][1] ), 
        .g_BAR(\pg_1[7][0] ) );
  pg_9 xPG_2_4 ( .p(\pg_1[9][1] ), .g_prec(\pg_1[8][0] ), .p_prec(\pg_1[8][1] ), .g_out(n5), .p_out(\pg_n[2][4][1] ), .g_BAR(\pg_1[9][0] ) );
  pg_8 xPG_2_5 ( .g(\pg_1[11][0] ), .p(\pg_1[11][1] ), .g_prec(\pg_1[10][0] ), 
        .p_prec(\pg_1[10][1] ), .p_out(\pg_n[2][5][1] ), .g_out_BAR(
        \pg_n[2][5][0] ) );
  pg_7 xPG_2_6 ( .g(\pg_1[13][0] ), .p(\pg_1[13][1] ), .g_prec(\pg_1[12][0] ), 
        .p_prec(\pg_1[12][1] ), .g_out(\pg_n[2][6][0] ), .p_out(
        \pg_n[2][6][1] ) );
  pg_6 xPG_2_7 ( .g(\pg_1[15][0] ), .p(\pg_1[15][1] ), .g_prec(\pg_1[14][0] ), 
        .p_prec(\pg_1[14][1] ), .g_out(\pg_n[2][7][0] ), .p_out(
        \pg_n[2][7][1] ) );
  g_7 xG_3_1 ( .g(\pg_n[2][1][0] ), .p(\pg_n[2][1][1] ), .g_prec(n26), .g_out(
        n8) );
  g_6 xG_4_2 ( .g(n20), .p(\pg_n[2][2][1] ), .g_prec(n23), .g_out(Cout[2]) );
  g_5 xG_4_3 ( .g(\pg_n[3][3][0] ), .p(\pg_n[3][3][1] ), .g_prec(n8), .g_out(
        n1) );
  g_4 xG_5_4 ( .g(n12), .p(\pg_n[2][4][1] ), .g_prec(n1), .g_out(Cout[4]) );
  g_3 xG_5_5 ( .g(n22), .p(\pg_n[3][5][1] ), .g_prec(n1), .g_out(Cout[5]) );
  g_2 xG_5_6 ( .g(\pg_n[4][6][0] ), .p(\pg_n[4][6][1] ), .g_prec(n1), .g_out(
        Cout[6]) );
  g_1 xG_5_7 ( .g(\pg_n[4][7][0] ), .p(\pg_n[4][7][1] ), .g_prec(Cout[3]), 
        .g_out(Cout[7]) );
  pg_5 xPG_3_3 ( .g(\pg_n[2][3][0] ), .p(\pg_n[2][3][1] ), .g_prec(
        \pg_n[2][2][0] ), .p_prec(\pg_n[2][2][1] ), .g_out(\pg_n[3][3][0] ), 
        .p_out(\pg_n[3][3][1] ) );
  pg_4 xPG_3_5 ( .p(\pg_n[2][5][1] ), .g_prec(n5), .p_prec(\pg_n[2][4][1] ), 
        .g_out(n7), .p_out(\pg_n[3][5][1] ), .g_BAR(\pg_n[2][5][0] ) );
  pg_3 xPG_3_7 ( .g(\pg_n[2][7][0] ), .p(\pg_n[2][7][1] ), .g_prec(
        \pg_n[2][6][0] ), .p_prec(\pg_n[2][6][1] ), .g_out(\pg_n[3][7][0] ), 
        .p_out(\pg_n[3][7][1] ) );
  pg_2 xPG_4_6 ( .g(\pg_n[2][6][0] ), .p(\pg_n[2][6][1] ), .g_prec(n7), 
        .p_prec(\pg_n[3][5][1] ), .g_out(\pg_n[4][6][0] ), .p_out(
        \pg_n[4][6][1] ) );
  pg_1 xPG_4_7 ( .g(\pg_n[3][7][0] ), .p(\pg_n[3][7][1] ), .g_prec(n22), 
        .p_prec(\pg_n[3][5][1] ), .g_out(\pg_n[4][7][0] ), .p_out(
        \pg_n[4][7][1] ) );
  CLKBUF_X1 U1 ( .A(n5), .Z(n12) );
  CLKBUF_X1 U2 ( .A(n7), .Z(n22) );
  CLKBUF_X1 U3 ( .A(\pg_n[2][2][0] ), .Z(n20) );
  BUF_X1 U4 ( .A(n8), .Z(n23) );
  BUF_X1 U5 ( .A(n1), .Z(Cout[3]) );
  CLKBUF_X1 U6 ( .A(n26), .Z(Cout[0]) );
  BUF_X1 U7 ( .A(n23), .Z(Cout[1]) );
endmodule


module xor_gen_N32_1 ( A, B, S );
  input [31:0] A;
  output [31:0] S;
  input B;
  wire   n15, n16, n17, n19, n20, n21, n22, n23;

  XOR2_X1 U8 ( .A(B), .B(A[31]), .Z(S[31]) );
  XOR2_X1 U9 ( .A(B), .B(A[30]), .Z(S[30]) );
  XOR2_X1 U12 ( .A(B), .B(A[28]), .Z(S[28]) );
  XOR2_X1 U13 ( .A(B), .B(A[27]), .Z(S[27]) );
  XOR2_X1 U14 ( .A(B), .B(A[26]), .Z(S[26]) );
  XOR2_X1 U16 ( .A(B), .B(A[24]), .Z(S[24]) );
  XOR2_X1 U17 ( .A(B), .B(A[23]), .Z(S[23]) );
  XOR2_X1 U20 ( .A(B), .B(A[20]), .Z(S[20]) );
  XOR2_X1 U29 ( .A(B), .B(A[12]), .Z(S[12]) );
  XNOR2_X1 U1 ( .A(A[0]), .B(n19), .ZN(S[0]) );
  XNOR2_X1 U2 ( .A(A[3]), .B(n19), .ZN(S[3]) );
  MUX2_X1 U3 ( .A(B), .B(n19), .S(A[9]), .Z(S[9]) );
  XOR2_X1 U4 ( .A(B), .B(A[14]), .Z(S[14]) );
  XOR2_X1 U5 ( .A(B), .B(A[21]), .Z(S[21]) );
  XOR2_X1 U6 ( .A(B), .B(A[29]), .Z(S[29]) );
  MUX2_X1 U7 ( .A(B), .B(n19), .S(A[5]), .Z(S[5]) );
  XOR2_X2 U10 ( .A(A[18]), .B(B), .Z(S[18]) );
  XOR2_X1 U11 ( .A(A[8]), .B(B), .Z(S[8]) );
  XOR2_X1 U15 ( .A(B), .B(A[16]), .Z(S[16]) );
  INV_X1 U18 ( .A(B), .ZN(n19) );
  INV_X1 U19 ( .A(A[13]), .ZN(n21) );
  XNOR2_X1 U21 ( .A(A[19]), .B(n19), .ZN(S[19]) );
  NAND2_X1 U22 ( .A1(n16), .A2(n17), .ZN(S[10]) );
  XOR2_X1 U23 ( .A(B), .B(A[25]), .Z(S[25]) );
  XOR2_X1 U24 ( .A(B), .B(A[22]), .Z(S[22]) );
  NAND2_X1 U25 ( .A1(n22), .A2(n23), .ZN(S[13]) );
  XOR2_X1 U26 ( .A(B), .B(A[6]), .Z(S[6]) );
  XOR2_X1 U27 ( .A(B), .B(A[17]), .Z(S[17]) );
  XOR2_X1 U28 ( .A(A[2]), .B(B), .Z(S[2]) );
  NAND2_X1 U30 ( .A1(A[10]), .A2(n19), .ZN(n16) );
  NAND2_X1 U31 ( .A1(n15), .A2(B), .ZN(n17) );
  INV_X1 U32 ( .A(A[10]), .ZN(n15) );
  OAI21_X2 U33 ( .B1(A[1]), .B2(n19), .A(n20), .ZN(S[1]) );
  XOR2_X1 U34 ( .A(A[11]), .B(B), .Z(S[11]) );
  XOR2_X1 U35 ( .A(A[15]), .B(B), .Z(S[15]) );
  XOR2_X1 U36 ( .A(A[4]), .B(B), .Z(S[4]) );
  XOR2_X1 U37 ( .A(A[7]), .B(B), .Z(S[7]) );
  NAND2_X1 U38 ( .A1(A[1]), .A2(n19), .ZN(n20) );
  NAND2_X1 U39 ( .A1(n21), .A2(B), .ZN(n22) );
  NAND2_X1 U40 ( .A1(A[13]), .A2(n19), .ZN(n23) );
endmodule


module ff32_en_SIZE5_2 ( D, en, clk, rst, Q );
  input [4:0] D;
  output [4:0] Q;
  input en, clk, rst;
  wire   n1, n3, n4, n5, n6, net645267, net645268, net645269, net645270,
         net645271, n13, n14, n15, n16, n17, n18, n19;

  DFFR_X1 \Q_reg[4]  ( .D(n1), .CK(clk), .RN(n14), .Q(Q[4]), .QN(net645271) );
  DFFR_X1 \Q_reg[3]  ( .D(n3), .CK(clk), .RN(n14), .Q(Q[3]), .QN(net645270) );
  DFFR_X1 \Q_reg[2]  ( .D(n4), .CK(clk), .RN(n14), .Q(Q[2]), .QN(net645269) );
  DFFR_X1 \Q_reg[1]  ( .D(n5), .CK(clk), .RN(n14), .Q(Q[1]), .QN(net645268) );
  DFFR_X1 \Q_reg[0]  ( .D(n6), .CK(clk), .RN(n14), .Q(Q[0]), .QN(net645267) );
  NAND2_X1 U7 ( .A1(n13), .A2(D[2]), .ZN(n17) );
  OAI21_X1 U6 ( .B1(n13), .B2(net645269), .A(n17), .ZN(n4) );
  NAND2_X1 U9 ( .A1(n13), .A2(D[3]), .ZN(n16) );
  OAI21_X1 U8 ( .B1(n13), .B2(net645270), .A(n16), .ZN(n3) );
  NAND2_X1 U12 ( .A1(n13), .A2(D[4]), .ZN(n15) );
  OAI21_X1 U11 ( .B1(n13), .B2(net645271), .A(n15), .ZN(n1) );
  NAND2_X1 U3 ( .A1(n13), .A2(D[0]), .ZN(n19) );
  OAI21_X1 U2 ( .B1(n13), .B2(net645267), .A(n19), .ZN(n6) );
  NAND2_X1 U5 ( .A1(n13), .A2(D[1]), .ZN(n18) );
  OAI21_X1 U4 ( .B1(n13), .B2(net645268), .A(n18), .ZN(n5) );
  INV_X1 U10 ( .A(rst), .ZN(n14) );
  BUF_X1 U13 ( .A(en), .Z(n13) );
endmodule


module ff32_en_SIZE5_1 ( D, en, clk, rst, Q );
  input [4:0] D;
  output [4:0] Q;
  input en, clk, rst;
  wire   n19, n20, n21, n22, n23;

  DFFR_X1 \Q_reg[1]  ( .D(D[1]), .CK(clk), .RN(n19), .Q(Q[1]) );
  DFFS_X1 \Q_reg[0]  ( .D(n23), .CK(clk), .SN(n19), .QN(Q[0]) );
  DFFS_X1 \Q_reg[3]  ( .D(n21), .CK(clk), .SN(n19), .QN(Q[3]) );
  DFFS_X1 \Q_reg[2]  ( .D(n22), .CK(clk), .SN(n19), .QN(Q[2]) );
  DFFS_X2 \Q_reg[4]  ( .D(n20), .CK(clk), .SN(n19), .QN(Q[4]) );
  INV_X1 U2 ( .A(D[0]), .ZN(n23) );
  INV_X1 U3 ( .A(rst), .ZN(n19) );
  INV_X1 U4 ( .A(D[4]), .ZN(n20) );
  INV_X1 U5 ( .A(D[3]), .ZN(n21) );
  INV_X1 U6 ( .A(D[2]), .ZN(n22) );
endmodule


module ff32_en_SIZE32_5 ( D, en, clk, rst, Q );
  input [31:0] D;
  output [31:0] Q;
  input en, clk, rst;
  wire   n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n97, net645107, net645108, net645109, net645110,
         net645111, net645112, net645113, net645114, net645115, net645116,
         net645117, net645118, net645119, net645120, net645121, net645122,
         net645123, net645124, net645125, net645126, net645127, net645128,
         net645129, net645130, net645131, net645132, net645133, net645134,
         net645135, net645136, net645137, net645138, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n96, n98, n99, n100
;

  DFFR_X1 \Q_reg[31]  ( .D(n97), .CK(clk), .RN(n36), .Q(Q[31]), .QN(net645138)
         );
  DFFR_X1 \Q_reg[30]  ( .D(n95), .CK(clk), .RN(n36), .Q(Q[30]), .QN(net645137)
         );
  DFFR_X1 \Q_reg[29]  ( .D(n94), .CK(clk), .RN(n36), .Q(Q[29]), .QN(net645136)
         );
  DFFR_X1 \Q_reg[28]  ( .D(n93), .CK(clk), .RN(n36), .Q(Q[28]), .QN(net645135)
         );
  DFFR_X1 \Q_reg[27]  ( .D(n92), .CK(clk), .RN(n36), .Q(Q[27]), .QN(net645134)
         );
  DFFR_X1 \Q_reg[26]  ( .D(n91), .CK(clk), .RN(n36), .Q(Q[26]), .QN(net645133)
         );
  DFFR_X1 \Q_reg[25]  ( .D(n90), .CK(clk), .RN(n36), .Q(Q[25]), .QN(net645132)
         );
  DFFR_X1 \Q_reg[24]  ( .D(n89), .CK(clk), .RN(n36), .Q(Q[24]), .QN(net645131)
         );
  DFFR_X1 \Q_reg[23]  ( .D(n88), .CK(clk), .RN(n36), .Q(Q[23]), .QN(net645130)
         );
  DFFR_X1 \Q_reg[22]  ( .D(n87), .CK(clk), .RN(n36), .Q(Q[22]), .QN(net645129)
         );
  DFFR_X1 \Q_reg[21]  ( .D(n86), .CK(clk), .RN(n36), .Q(Q[21]), .QN(net645128)
         );
  DFFR_X1 \Q_reg[19]  ( .D(n84), .CK(clk), .RN(n36), .Q(Q[19]), .QN(net645127)
         );
  DFFR_X1 \Q_reg[18]  ( .D(n83), .CK(clk), .RN(n36), .Q(Q[18]), .QN(net645126)
         );
  DFFR_X1 \Q_reg[17]  ( .D(n82), .CK(clk), .RN(n36), .Q(Q[17]), .QN(net645125)
         );
  DFFR_X1 \Q_reg[16]  ( .D(n81), .CK(clk), .RN(n36), .Q(Q[16]), .QN(net645124)
         );
  DFFR_X1 \Q_reg[15]  ( .D(n80), .CK(clk), .RN(n36), .Q(Q[15]), .QN(net645123)
         );
  DFFR_X1 \Q_reg[14]  ( .D(n79), .CK(clk), .RN(n36), .Q(Q[14]), .QN(net645122)
         );
  DFFR_X1 \Q_reg[13]  ( .D(n78), .CK(clk), .RN(n36), .Q(Q[13]), .QN(net645121)
         );
  DFFR_X1 \Q_reg[12]  ( .D(n77), .CK(clk), .RN(n36), .Q(Q[12]), .QN(net645120)
         );
  DFFR_X1 \Q_reg[11]  ( .D(n76), .CK(clk), .RN(n36), .Q(Q[11]), .QN(net645119)
         );
  DFFR_X1 \Q_reg[10]  ( .D(n75), .CK(clk), .RN(n36), .Q(Q[10]), .QN(net645118)
         );
  DFFR_X1 \Q_reg[9]  ( .D(n74), .CK(clk), .RN(n36), .Q(Q[9]), .QN(net645117)
         );
  DFFR_X1 \Q_reg[8]  ( .D(n73), .CK(clk), .RN(n36), .Q(Q[8]), .QN(net645116)
         );
  DFFR_X1 \Q_reg[7]  ( .D(n72), .CK(clk), .RN(n36), .Q(Q[7]), .QN(net645115)
         );
  DFFR_X1 \Q_reg[6]  ( .D(n71), .CK(clk), .RN(n36), .Q(Q[6]), .QN(net645114)
         );
  DFFR_X1 \Q_reg[5]  ( .D(n70), .CK(clk), .RN(n36), .Q(Q[5]), .QN(net645113)
         );
  DFFR_X1 \Q_reg[4]  ( .D(n69), .CK(clk), .RN(n36), .Q(Q[4]), .QN(net645112)
         );
  DFFR_X1 \Q_reg[3]  ( .D(n68), .CK(clk), .RN(n36), .Q(Q[3]), .QN(net645111)
         );
  DFFR_X1 \Q_reg[2]  ( .D(n67), .CK(clk), .RN(n36), .Q(Q[2]), .QN(net645110)
         );
  DFFR_X1 \Q_reg[1]  ( .D(n66), .CK(clk), .RN(n36), .Q(Q[1]), .QN(net645109)
         );
  DFFR_X1 \Q_reg[0]  ( .D(n65), .CK(clk), .RN(n36), .Q(Q[0]), .QN(net645108)
         );
  DFFR_X1 \Q_reg[20]  ( .D(n85), .CK(clk), .RN(n36), .Q(Q[20]), .QN(net645107)
         );
  NAND2_X1 U43 ( .A1(en), .A2(D[11]), .ZN(n48) );
  OAI21_X1 U42 ( .B1(en), .B2(net645119), .A(n48), .ZN(n76) );
  NAND2_X1 U45 ( .A1(en), .A2(D[10]), .ZN(n47) );
  OAI21_X1 U44 ( .B1(en), .B2(net645118), .A(n47), .ZN(n75) );
  NAND2_X1 U37 ( .A1(en), .A2(D[14]), .ZN(n51) );
  OAI21_X1 U36 ( .B1(en), .B2(net645122), .A(n51), .ZN(n79) );
  NAND2_X1 U39 ( .A1(en), .A2(D[13]), .ZN(n50) );
  OAI21_X1 U38 ( .B1(en), .B2(net645121), .A(n50), .ZN(n78) );
  NAND2_X1 U55 ( .A1(en), .A2(D[5]), .ZN(n42) );
  OAI21_X1 U54 ( .B1(en), .B2(net645113), .A(n42), .ZN(n70) );
  NAND2_X1 U57 ( .A1(en), .A2(D[4]), .ZN(n41) );
  OAI21_X1 U56 ( .B1(en), .B2(net645112), .A(n41), .ZN(n69) );
  NAND2_X1 U13 ( .A1(en), .A2(D[26]), .ZN(n63) );
  OAI21_X1 U12 ( .B1(en), .B2(net645133), .A(n63), .ZN(n91) );
  NAND2_X1 U49 ( .A1(en), .A2(D[8]), .ZN(n45) );
  OAI21_X1 U48 ( .B1(en), .B2(net645116), .A(n45), .ZN(n73) );
  NAND2_X1 U23 ( .A1(en), .A2(D[21]), .ZN(n58) );
  OAI21_X1 U22 ( .B1(en), .B2(net645128), .A(n58), .ZN(n86) );
  NAND2_X1 U61 ( .A1(en), .A2(D[2]), .ZN(n39) );
  OAI21_X1 U60 ( .B1(en), .B2(net645110), .A(n39), .ZN(n67) );
  NAND2_X1 U59 ( .A1(en), .A2(D[3]), .ZN(n40) );
  OAI21_X1 U58 ( .B1(en), .B2(net645111), .A(n40), .ZN(n68) );
  NAND2_X1 U53 ( .A1(en), .A2(D[6]), .ZN(n43) );
  OAI21_X1 U52 ( .B1(en), .B2(net645114), .A(n43), .ZN(n71) );
  NAND2_X1 U21 ( .A1(en), .A2(D[22]), .ZN(n59) );
  OAI21_X1 U20 ( .B1(en), .B2(net645129), .A(n59), .ZN(n87) );
  NAND2_X1 U17 ( .A1(en), .A2(D[24]), .ZN(n61) );
  OAI21_X1 U16 ( .B1(en), .B2(net645131), .A(n61), .ZN(n89) );
  NAND2_X1 U25 ( .A1(en), .A2(D[20]), .ZN(n57) );
  OAI21_X1 U24 ( .B1(en), .B2(net645107), .A(n57), .ZN(n85) );
  NAND2_X1 U27 ( .A1(en), .A2(D[19]), .ZN(n56) );
  OAI21_X1 U26 ( .B1(en), .B2(net645127), .A(n56), .ZN(n84) );
  NAND2_X1 U51 ( .A1(en), .A2(D[7]), .ZN(n44) );
  OAI21_X1 U50 ( .B1(en), .B2(net645115), .A(n44), .ZN(n72) );
  NAND2_X1 U7 ( .A1(en), .A2(D[29]), .ZN(n98) );
  OAI21_X1 U6 ( .B1(en), .B2(net645136), .A(n98), .ZN(n94) );
  NAND2_X1 U9 ( .A1(en), .A2(D[28]), .ZN(n96) );
  OAI21_X1 U8 ( .B1(en), .B2(net645135), .A(n96), .ZN(n93) );
  NAND2_X1 U11 ( .A1(en), .A2(D[27]), .ZN(n64) );
  OAI21_X1 U10 ( .B1(en), .B2(net645134), .A(n64), .ZN(n92) );
  NAND2_X1 U19 ( .A1(en), .A2(D[23]), .ZN(n60) );
  OAI21_X1 U18 ( .B1(en), .B2(net645130), .A(n60), .ZN(n88) );
  NAND2_X1 U15 ( .A1(en), .A2(D[25]), .ZN(n62) );
  OAI21_X1 U14 ( .B1(en), .B2(net645132), .A(n62), .ZN(n90) );
  NAND2_X1 U35 ( .A1(en), .A2(D[15]), .ZN(n52) );
  OAI21_X1 U34 ( .B1(en), .B2(net645123), .A(n52), .ZN(n80) );
  NAND2_X1 U33 ( .A1(en), .A2(D[16]), .ZN(n53) );
  OAI21_X1 U32 ( .B1(en), .B2(net645124), .A(n53), .ZN(n81) );
  NAND2_X1 U31 ( .A1(en), .A2(D[17]), .ZN(n54) );
  OAI21_X1 U30 ( .B1(en), .B2(net645125), .A(n54), .ZN(n82) );
  NAND2_X1 U29 ( .A1(en), .A2(D[18]), .ZN(n55) );
  OAI21_X1 U28 ( .B1(en), .B2(net645126), .A(n55), .ZN(n83) );
  NAND2_X1 U47 ( .A1(en), .A2(D[9]), .ZN(n46) );
  OAI21_X1 U46 ( .B1(en), .B2(net645117), .A(n46), .ZN(n74) );
  NAND2_X1 U41 ( .A1(en), .A2(D[12]), .ZN(n49) );
  OAI21_X1 U40 ( .B1(en), .B2(net645120), .A(n49), .ZN(n77) );
  NAND2_X1 U63 ( .A1(en), .A2(D[1]), .ZN(n38) );
  OAI21_X1 U62 ( .B1(en), .B2(net645109), .A(n38), .ZN(n66) );
  NAND2_X1 U65 ( .A1(en), .A2(D[0]), .ZN(n37) );
  OAI21_X1 U64 ( .B1(en), .B2(net645108), .A(n37), .ZN(n65) );
  NAND2_X1 U3 ( .A1(en), .A2(D[31]), .ZN(n100) );
  OAI21_X1 U2 ( .B1(en), .B2(net645138), .A(n100), .ZN(n97) );
  NAND2_X1 U5 ( .A1(en), .A2(D[30]), .ZN(n99) );
  OAI21_X1 U4 ( .B1(en), .B2(net645137), .A(n99), .ZN(n95) );
  INV_X2 U66 ( .A(rst), .ZN(n36) );
endmodule


module ff32_en_SIZE32_4 ( D, en, clk, rst, Q );
  input [31:0] D;
  output [31:0] Q;
  input en, clk, rst;
  wire   n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n97, net645107, net645108, net645109, net645110,
         net645111, net645112, net645113, net645114, net645115, net645116,
         net645117, net645118, net645119, net645120, net645121, net645122,
         net645123, net645124, net645125, net645126, net645127, net645128,
         net645129, net645130, net645131, net645132, net645133, net645134,
         net645135, net645136, net645137, net645138, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n96, n98, n99, n100,
         n101, n102, n103, n104;

  DFFR_X1 \Q_reg[31]  ( .D(n97), .CK(clk), .RN(n40), .Q(Q[31]), .QN(net645138)
         );
  DFFR_X1 \Q_reg[30]  ( .D(n95), .CK(clk), .RN(n40), .Q(Q[30]), .QN(net645137)
         );
  DFFR_X1 \Q_reg[29]  ( .D(n94), .CK(clk), .RN(n40), .Q(Q[29]), .QN(net645136)
         );
  DFFR_X1 \Q_reg[28]  ( .D(n93), .CK(clk), .RN(n40), .Q(Q[28]), .QN(net645135)
         );
  DFFR_X1 \Q_reg[27]  ( .D(n92), .CK(clk), .RN(n40), .Q(Q[27]), .QN(net645134)
         );
  DFFR_X1 \Q_reg[26]  ( .D(n91), .CK(clk), .RN(n40), .Q(Q[26]), .QN(net645133)
         );
  DFFR_X1 \Q_reg[25]  ( .D(n90), .CK(clk), .RN(n40), .Q(Q[25]), .QN(net645132)
         );
  DFFR_X1 \Q_reg[24]  ( .D(n89), .CK(clk), .RN(n40), .Q(Q[24]), .QN(net645131)
         );
  DFFR_X1 \Q_reg[23]  ( .D(n88), .CK(clk), .RN(n40), .Q(Q[23]), .QN(net645130)
         );
  DFFR_X1 \Q_reg[22]  ( .D(n87), .CK(clk), .RN(n40), .Q(Q[22]), .QN(net645129)
         );
  DFFR_X1 \Q_reg[21]  ( .D(n86), .CK(clk), .RN(n40), .Q(Q[21]), .QN(net645128)
         );
  DFFR_X1 \Q_reg[19]  ( .D(n84), .CK(clk), .RN(n40), .Q(Q[19]), .QN(net645127)
         );
  DFFR_X1 \Q_reg[18]  ( .D(n83), .CK(clk), .RN(n40), .Q(Q[18]), .QN(net645126)
         );
  DFFR_X1 \Q_reg[17]  ( .D(n82), .CK(clk), .RN(n40), .Q(Q[17]), .QN(net645125)
         );
  DFFR_X1 \Q_reg[16]  ( .D(n81), .CK(clk), .RN(n40), .Q(Q[16]), .QN(net645124)
         );
  DFFR_X1 \Q_reg[15]  ( .D(n80), .CK(clk), .RN(n40), .Q(Q[15]), .QN(net645123)
         );
  DFFR_X1 \Q_reg[14]  ( .D(n79), .CK(clk), .RN(n40), .Q(Q[14]), .QN(net645122)
         );
  DFFR_X1 \Q_reg[13]  ( .D(n78), .CK(clk), .RN(n40), .Q(Q[13]), .QN(net645121)
         );
  DFFR_X1 \Q_reg[12]  ( .D(n77), .CK(clk), .RN(n40), .Q(Q[12]), .QN(net645120)
         );
  DFFR_X1 \Q_reg[11]  ( .D(n76), .CK(clk), .RN(n40), .Q(Q[11]), .QN(net645119)
         );
  DFFR_X1 \Q_reg[10]  ( .D(n75), .CK(clk), .RN(n40), .Q(Q[10]), .QN(net645118)
         );
  DFFR_X1 \Q_reg[9]  ( .D(n74), .CK(clk), .RN(n40), .Q(Q[9]), .QN(net645117)
         );
  DFFR_X1 \Q_reg[8]  ( .D(n73), .CK(clk), .RN(n40), .Q(Q[8]), .QN(net645116)
         );
  DFFR_X1 \Q_reg[7]  ( .D(n72), .CK(clk), .RN(n40), .Q(Q[7]), .QN(net645115)
         );
  DFFR_X1 \Q_reg[6]  ( .D(n71), .CK(clk), .RN(n40), .Q(Q[6]), .QN(net645114)
         );
  DFFR_X1 \Q_reg[5]  ( .D(n70), .CK(clk), .RN(n40), .Q(Q[5]), .QN(net645113)
         );
  DFFR_X1 \Q_reg[4]  ( .D(n69), .CK(clk), .RN(n40), .Q(Q[4]), .QN(net645112)
         );
  DFFR_X1 \Q_reg[3]  ( .D(n68), .CK(clk), .RN(n40), .Q(Q[3]), .QN(net645111)
         );
  DFFR_X1 \Q_reg[2]  ( .D(n67), .CK(clk), .RN(n40), .Q(Q[2]), .QN(net645110)
         );
  DFFR_X1 \Q_reg[1]  ( .D(n66), .CK(clk), .RN(n40), .Q(Q[1]), .QN(net645109)
         );
  DFFR_X1 \Q_reg[0]  ( .D(n65), .CK(clk), .RN(n40), .Q(Q[0]), .QN(net645108)
         );
  DFFR_X1 \Q_reg[20]  ( .D(n85), .CK(clk), .RN(n40), .Q(Q[20]), .QN(net645107)
         );
  NAND2_X1 U39 ( .A1(n39), .A2(D[13]), .ZN(n54) );
  OAI21_X1 U38 ( .B1(n37), .B2(net645121), .A(n54), .ZN(n78) );
  NAND2_X1 U3 ( .A1(n39), .A2(D[31]), .ZN(n104) );
  OAI21_X1 U2 ( .B1(n37), .B2(net645138), .A(n104), .ZN(n97) );
  NAND2_X1 U43 ( .A1(n39), .A2(D[11]), .ZN(n52) );
  OAI21_X1 U42 ( .B1(n37), .B2(net645119), .A(n52), .ZN(n76) );
  NAND2_X1 U63 ( .A1(n39), .A2(D[1]), .ZN(n42) );
  OAI21_X1 U62 ( .B1(n36), .B2(net645109), .A(n42), .ZN(n66) );
  NAND2_X1 U5 ( .A1(n39), .A2(D[30]), .ZN(n103) );
  OAI21_X1 U4 ( .B1(n36), .B2(net645137), .A(n103), .ZN(n95) );
  NAND2_X1 U45 ( .A1(n39), .A2(D[10]), .ZN(n51) );
  OAI21_X1 U44 ( .B1(n37), .B2(net645118), .A(n51), .ZN(n75) );
  NAND2_X1 U37 ( .A1(n39), .A2(D[14]), .ZN(n55) );
  OAI21_X1 U36 ( .B1(n37), .B2(net645122), .A(n55), .ZN(n79) );
  NAND2_X1 U33 ( .A1(en), .A2(D[16]), .ZN(n57) );
  OAI21_X1 U32 ( .B1(n37), .B2(net645124), .A(n57), .ZN(n81) );
  NAND2_X1 U27 ( .A1(en), .A2(D[19]), .ZN(n60) );
  OAI21_X1 U26 ( .B1(n36), .B2(net645127), .A(n60), .ZN(n84) );
  NAND2_X1 U41 ( .A1(en), .A2(D[12]), .ZN(n53) );
  OAI21_X1 U40 ( .B1(n37), .B2(net645120), .A(n53), .ZN(n77) );
  NAND2_X1 U19 ( .A1(n38), .A2(D[23]), .ZN(n64) );
  OAI21_X1 U18 ( .B1(n36), .B2(net645130), .A(n64), .ZN(n88) );
  NAND2_X1 U9 ( .A1(n38), .A2(D[28]), .ZN(n101) );
  OAI21_X1 U8 ( .B1(n36), .B2(net645135), .A(n101), .ZN(n93) );
  NAND2_X1 U23 ( .A1(n38), .A2(D[21]), .ZN(n62) );
  OAI21_X1 U22 ( .B1(n36), .B2(net645128), .A(n62), .ZN(n86) );
  NAND2_X1 U31 ( .A1(en), .A2(D[17]), .ZN(n58) );
  OAI21_X1 U30 ( .B1(n37), .B2(net645125), .A(n58), .ZN(n82) );
  NAND2_X1 U17 ( .A1(n38), .A2(D[24]), .ZN(n96) );
  OAI21_X1 U16 ( .B1(n36), .B2(net645131), .A(n96), .ZN(n89) );
  NAND2_X1 U29 ( .A1(en), .A2(D[18]), .ZN(n59) );
  OAI21_X1 U28 ( .B1(n37), .B2(net645126), .A(n59), .ZN(n83) );
  NAND2_X1 U21 ( .A1(en), .A2(D[22]), .ZN(n63) );
  OAI21_X1 U20 ( .B1(n36), .B2(net645129), .A(n63), .ZN(n87) );
  NAND2_X1 U61 ( .A1(n38), .A2(D[2]), .ZN(n43) );
  OAI21_X1 U60 ( .B1(n37), .B2(net645110), .A(n43), .ZN(n67) );
  NAND2_X1 U51 ( .A1(en), .A2(D[7]), .ZN(n48) );
  OAI21_X1 U50 ( .B1(n37), .B2(net645115), .A(n48), .ZN(n72) );
  NAND2_X1 U7 ( .A1(n38), .A2(D[29]), .ZN(n102) );
  OAI21_X1 U6 ( .B1(n36), .B2(net645136), .A(n102), .ZN(n94) );
  NAND2_X1 U49 ( .A1(en), .A2(D[8]), .ZN(n49) );
  OAI21_X1 U48 ( .B1(n36), .B2(net645116), .A(n49), .ZN(n73) );
  NAND2_X1 U25 ( .A1(en), .A2(D[20]), .ZN(n61) );
  OAI21_X1 U24 ( .B1(n36), .B2(net645107), .A(n61), .ZN(n85) );
  NAND2_X1 U13 ( .A1(n38), .A2(D[26]), .ZN(n99) );
  OAI21_X1 U12 ( .B1(n36), .B2(net645133), .A(n99), .ZN(n91) );
  NAND2_X1 U15 ( .A1(n38), .A2(D[25]), .ZN(n98) );
  OAI21_X1 U14 ( .B1(n36), .B2(net645132), .A(n98), .ZN(n90) );
  NAND2_X1 U11 ( .A1(n38), .A2(D[27]), .ZN(n100) );
  OAI21_X1 U10 ( .B1(n36), .B2(net645134), .A(n100), .ZN(n92) );
  NAND2_X1 U35 ( .A1(en), .A2(D[15]), .ZN(n56) );
  OAI21_X1 U34 ( .B1(n37), .B2(net645123), .A(n56), .ZN(n80) );
  NAND2_X1 U53 ( .A1(n38), .A2(D[6]), .ZN(n47) );
  OAI21_X1 U52 ( .B1(n37), .B2(net645114), .A(n47), .ZN(n71) );
  NAND2_X1 U47 ( .A1(en), .A2(D[9]), .ZN(n50) );
  OAI21_X1 U46 ( .B1(n37), .B2(net645117), .A(n50), .ZN(n74) );
  NAND2_X1 U65 ( .A1(n39), .A2(D[0]), .ZN(n41) );
  OAI21_X1 U64 ( .B1(n39), .B2(net645108), .A(n41), .ZN(n65) );
  NAND2_X1 U57 ( .A1(n38), .A2(D[4]), .ZN(n45) );
  OAI21_X1 U56 ( .B1(n39), .B2(net645112), .A(n45), .ZN(n69) );
  NAND2_X1 U59 ( .A1(n38), .A2(D[3]), .ZN(n44) );
  OAI21_X1 U58 ( .B1(n39), .B2(net645111), .A(n44), .ZN(n68) );
  NAND2_X1 U55 ( .A1(en), .A2(D[5]), .ZN(n46) );
  OAI21_X1 U54 ( .B1(n39), .B2(net645113), .A(n46), .ZN(n70) );
  INV_X2 U66 ( .A(rst), .ZN(n40) );
  BUF_X1 U67 ( .A(en), .Z(n36) );
  BUF_X1 U68 ( .A(en), .Z(n37) );
  BUF_X1 U69 ( .A(en), .Z(n38) );
  BUF_X1 U70 ( .A(en), .Z(n39) );
endmodule


module ff32_en_SIZE32_3 ( D, en, clk, rst, Q );
  input [31:0] D;
  output [31:0] Q;
  input en, clk, rst;
  wire   n35;

  DFFR_X1 \Q_reg[31]  ( .D(D[31]), .CK(clk), .RN(n35), .Q(Q[31]) );
  DFFR_X1 \Q_reg[30]  ( .D(D[30]), .CK(clk), .RN(n35), .Q(Q[30]) );
  DFFR_X1 \Q_reg[29]  ( .D(D[29]), .CK(clk), .RN(n35), .Q(Q[29]) );
  DFFR_X1 \Q_reg[28]  ( .D(D[28]), .CK(clk), .RN(n35), .Q(Q[28]) );
  DFFR_X1 \Q_reg[27]  ( .D(D[27]), .CK(clk), .RN(n35), .Q(Q[27]) );
  DFFR_X1 \Q_reg[26]  ( .D(D[26]), .CK(clk), .RN(n35), .Q(Q[26]) );
  DFFR_X1 \Q_reg[25]  ( .D(D[25]), .CK(clk), .RN(n35), .Q(Q[25]) );
  DFFR_X1 \Q_reg[24]  ( .D(D[24]), .CK(clk), .RN(n35), .Q(Q[24]) );
  DFFR_X1 \Q_reg[23]  ( .D(D[23]), .CK(clk), .RN(n35), .Q(Q[23]) );
  DFFR_X1 \Q_reg[22]  ( .D(D[22]), .CK(clk), .RN(n35), .Q(Q[22]) );
  DFFR_X1 \Q_reg[21]  ( .D(D[21]), .CK(clk), .RN(n35), .Q(Q[21]) );
  DFFR_X1 \Q_reg[19]  ( .D(D[19]), .CK(clk), .RN(n35), .Q(Q[19]) );
  DFFR_X1 \Q_reg[18]  ( .D(D[18]), .CK(clk), .RN(n35), .Q(Q[18]) );
  DFFR_X1 \Q_reg[17]  ( .D(D[17]), .CK(clk), .RN(n35), .Q(Q[17]) );
  DFFR_X1 \Q_reg[16]  ( .D(D[16]), .CK(clk), .RN(n35), .Q(Q[16]) );
  DFFR_X1 \Q_reg[15]  ( .D(D[15]), .CK(clk), .RN(n35), .Q(Q[15]) );
  DFFR_X1 \Q_reg[14]  ( .D(D[14]), .CK(clk), .RN(n35), .Q(Q[14]) );
  DFFR_X1 \Q_reg[13]  ( .D(D[13]), .CK(clk), .RN(n35), .Q(Q[13]) );
  DFFR_X1 \Q_reg[12]  ( .D(D[12]), .CK(clk), .RN(n35), .Q(Q[12]) );
  DFFR_X1 \Q_reg[11]  ( .D(D[11]), .CK(clk), .RN(n35), .Q(Q[11]) );
  DFFR_X1 \Q_reg[10]  ( .D(D[10]), .CK(clk), .RN(n35), .Q(Q[10]) );
  DFFR_X1 \Q_reg[9]  ( .D(D[9]), .CK(clk), .RN(n35), .Q(Q[9]) );
  DFFR_X1 \Q_reg[8]  ( .D(D[8]), .CK(clk), .RN(n35), .Q(Q[8]) );
  DFFR_X1 \Q_reg[7]  ( .D(D[7]), .CK(clk), .RN(n35), .Q(Q[7]) );
  DFFR_X1 \Q_reg[6]  ( .D(D[6]), .CK(clk), .RN(n35), .Q(Q[6]) );
  DFFR_X1 \Q_reg[5]  ( .D(D[5]), .CK(clk), .RN(n35), .Q(Q[5]) );
  DFFR_X1 \Q_reg[4]  ( .D(D[4]), .CK(clk), .RN(n35), .Q(Q[4]) );
  DFFR_X1 \Q_reg[3]  ( .D(D[3]), .CK(clk), .RN(n35), .Q(Q[3]) );
  DFFR_X1 \Q_reg[2]  ( .D(D[2]), .CK(clk), .RN(n35), .Q(Q[2]) );
  DFFR_X1 \Q_reg[1]  ( .D(D[1]), .CK(clk), .RN(n35), .Q(Q[1]) );
  DFFR_X1 \Q_reg[0]  ( .D(D[0]), .CK(clk), .RN(n35), .Q(Q[0]) );
  DFFR_X1 \Q_reg[20]  ( .D(D[20]), .CK(clk), .RN(n35), .Q(Q[20]) );
  INV_X2 U2 ( .A(rst), .ZN(n35) );
endmodule


module ff32_en_SIZE32_2 ( D, en, clk, rst, Q );
  input [31:0] D;
  output [31:0] Q;
  input en, clk, rst;
  wire   n37;

  DFFR_X1 \Q_reg[31]  ( .D(D[31]), .CK(clk), .RN(n37), .Q(Q[31]) );
  DFFR_X1 \Q_reg[30]  ( .D(D[30]), .CK(clk), .RN(n37), .Q(Q[30]) );
  DFFR_X1 \Q_reg[29]  ( .D(D[29]), .CK(clk), .RN(n37), .Q(Q[29]) );
  DFFR_X1 \Q_reg[28]  ( .D(D[28]), .CK(clk), .RN(n37), .Q(Q[28]) );
  DFFR_X1 \Q_reg[27]  ( .D(D[27]), .CK(clk), .RN(n37), .Q(Q[27]) );
  DFFR_X1 \Q_reg[26]  ( .D(D[26]), .CK(clk), .RN(n37), .Q(Q[26]) );
  DFFR_X1 \Q_reg[25]  ( .D(D[25]), .CK(clk), .RN(n37), .Q(Q[25]) );
  DFFR_X1 \Q_reg[24]  ( .D(D[24]), .CK(clk), .RN(n37), .Q(Q[24]) );
  DFFR_X1 \Q_reg[23]  ( .D(D[23]), .CK(clk), .RN(n37), .Q(Q[23]) );
  DFFR_X1 \Q_reg[22]  ( .D(D[22]), .CK(clk), .RN(n37), .Q(Q[22]) );
  DFFR_X1 \Q_reg[21]  ( .D(D[21]), .CK(clk), .RN(n37), .Q(Q[21]) );
  DFFR_X1 \Q_reg[19]  ( .D(D[19]), .CK(clk), .RN(n37), .Q(Q[19]) );
  DFFR_X1 \Q_reg[18]  ( .D(D[18]), .CK(clk), .RN(n37), .Q(Q[18]) );
  DFFR_X1 \Q_reg[17]  ( .D(D[17]), .CK(clk), .RN(n37), .Q(Q[17]) );
  DFFR_X1 \Q_reg[16]  ( .D(D[16]), .CK(clk), .RN(n37), .Q(Q[16]) );
  DFFR_X1 \Q_reg[15]  ( .D(D[15]), .CK(clk), .RN(n37), .Q(Q[15]) );
  DFFR_X1 \Q_reg[14]  ( .D(D[14]), .CK(clk), .RN(n37), .Q(Q[14]) );
  DFFR_X1 \Q_reg[13]  ( .D(D[13]), .CK(clk), .RN(n37), .Q(Q[13]) );
  DFFR_X1 \Q_reg[12]  ( .D(D[12]), .CK(clk), .RN(n37), .Q(Q[12]) );
  DFFR_X1 \Q_reg[11]  ( .D(D[11]), .CK(clk), .RN(n37), .Q(Q[11]) );
  DFFR_X1 \Q_reg[10]  ( .D(D[10]), .CK(clk), .RN(n37), .Q(Q[10]) );
  DFFR_X1 \Q_reg[9]  ( .D(D[9]), .CK(clk), .RN(n37), .Q(Q[9]) );
  DFFR_X1 \Q_reg[8]  ( .D(D[8]), .CK(clk), .RN(n37), .Q(Q[8]) );
  DFFR_X1 \Q_reg[7]  ( .D(D[7]), .CK(clk), .RN(n37), .Q(Q[7]) );
  DFFR_X1 \Q_reg[6]  ( .D(D[6]), .CK(clk), .RN(n37), .Q(Q[6]) );
  DFFR_X1 \Q_reg[5]  ( .D(D[5]), .CK(clk), .RN(n37), .Q(Q[5]) );
  DFFR_X1 \Q_reg[4]  ( .D(D[4]), .CK(clk), .RN(n37), .Q(Q[4]) );
  DFFR_X1 \Q_reg[3]  ( .D(D[3]), .CK(clk), .RN(n37), .Q(Q[3]) );
  DFFR_X1 \Q_reg[2]  ( .D(D[2]), .CK(clk), .RN(n37), .Q(Q[2]) );
  DFFR_X1 \Q_reg[1]  ( .D(D[1]), .CK(clk), .RN(n37), .Q(Q[1]) );
  DFFR_X1 \Q_reg[0]  ( .D(D[0]), .CK(clk), .RN(n37), .Q(Q[0]) );
  DFFR_X1 \Q_reg[20]  ( .D(D[20]), .CK(clk), .RN(n37), .Q(Q[20]) );
  INV_X2 U2 ( .A(rst), .ZN(n37) );
endmodule


module ff32_en_SIZE32_1 ( D, en, clk, rst, Q );
  input [31:0] D;
  output [31:0] Q;
  input en, clk, rst;
  wire   n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n97, net645107, net645108, net645109, net645110,
         net645111, net645112, net645113, net645114, net645115, net645116,
         net645117, net645118, net645119, net645120, net645121, net645122,
         net645123, net645124, net645125, net645126, net645127, net645128,
         net645129, net645130, net645131, net645132, net645133, net645134,
         net645135, net645136, net645137, net645138, n35, n36, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n96, n98, n99, n100,
         n101;

  DFFR_X1 \Q_reg[31]  ( .D(n97), .CK(clk), .RN(n39), .Q(Q[31]), .QN(net645138)
         );
  DFFR_X1 \Q_reg[30]  ( .D(n95), .CK(clk), .RN(n39), .Q(Q[30]), .QN(net645137)
         );
  DFFR_X1 \Q_reg[29]  ( .D(n94), .CK(clk), .RN(n39), .Q(Q[29]), .QN(net645136)
         );
  DFFR_X1 \Q_reg[28]  ( .D(n93), .CK(clk), .RN(n39), .Q(Q[28]), .QN(net645135)
         );
  DFFR_X1 \Q_reg[27]  ( .D(n92), .CK(clk), .RN(n39), .Q(Q[27]), .QN(net645134)
         );
  DFFR_X1 \Q_reg[26]  ( .D(n91), .CK(clk), .RN(n39), .Q(Q[26]), .QN(net645133)
         );
  DFFR_X1 \Q_reg[25]  ( .D(n90), .CK(clk), .RN(n39), .Q(Q[25]), .QN(net645132)
         );
  DFFR_X1 \Q_reg[24]  ( .D(n89), .CK(clk), .RN(n39), .Q(Q[24]), .QN(net645131)
         );
  DFFR_X1 \Q_reg[23]  ( .D(n88), .CK(clk), .RN(n39), .Q(Q[23]), .QN(net645130)
         );
  DFFR_X1 \Q_reg[22]  ( .D(n87), .CK(clk), .RN(n39), .Q(Q[22]), .QN(net645129)
         );
  DFFR_X1 \Q_reg[21]  ( .D(n86), .CK(clk), .RN(n39), .Q(Q[21]), .QN(net645128)
         );
  DFFR_X1 \Q_reg[19]  ( .D(n84), .CK(clk), .RN(n39), .Q(Q[19]), .QN(net645127)
         );
  DFFR_X1 \Q_reg[18]  ( .D(n83), .CK(clk), .RN(n39), .Q(Q[18]), .QN(net645126)
         );
  DFFR_X1 \Q_reg[17]  ( .D(n82), .CK(clk), .RN(n39), .Q(Q[17]), .QN(net645125)
         );
  DFFR_X1 \Q_reg[16]  ( .D(n81), .CK(clk), .RN(n39), .Q(Q[16]), .QN(net645124)
         );
  DFFR_X1 \Q_reg[15]  ( .D(n80), .CK(clk), .RN(n39), .Q(Q[15]), .QN(net645123)
         );
  DFFR_X1 \Q_reg[14]  ( .D(n79), .CK(clk), .RN(n39), .Q(Q[14]), .QN(net645122)
         );
  DFFR_X1 \Q_reg[13]  ( .D(n78), .CK(clk), .RN(n39), .Q(Q[13]), .QN(net645121)
         );
  DFFR_X1 \Q_reg[12]  ( .D(n77), .CK(clk), .RN(n39), .Q(Q[12]), .QN(net645120)
         );
  DFFR_X1 \Q_reg[11]  ( .D(n76), .CK(clk), .RN(n39), .Q(Q[11]), .QN(net645119)
         );
  DFFR_X1 \Q_reg[10]  ( .D(n75), .CK(clk), .RN(n39), .Q(Q[10]), .QN(net645118)
         );
  DFFR_X1 \Q_reg[9]  ( .D(n74), .CK(clk), .RN(n39), .Q(Q[9]), .QN(net645117)
         );
  DFFR_X1 \Q_reg[8]  ( .D(n73), .CK(clk), .RN(n39), .Q(Q[8]), .QN(net645116)
         );
  DFFR_X1 \Q_reg[7]  ( .D(n72), .CK(clk), .RN(n39), .Q(Q[7]), .QN(net645115)
         );
  DFFR_X1 \Q_reg[6]  ( .D(n71), .CK(clk), .RN(n39), .Q(Q[6]), .QN(net645114)
         );
  DFFR_X1 \Q_reg[5]  ( .D(n70), .CK(clk), .RN(n39), .Q(Q[5]), .QN(net645113)
         );
  DFFR_X1 \Q_reg[4]  ( .D(n69), .CK(clk), .RN(n39), .Q(Q[4]), .QN(net645112)
         );
  DFFR_X1 \Q_reg[3]  ( .D(n68), .CK(clk), .RN(n39), .Q(Q[3]), .QN(net645111)
         );
  DFFR_X1 \Q_reg[2]  ( .D(n67), .CK(clk), .RN(n39), .Q(Q[2]), .QN(net645110)
         );
  DFFR_X1 \Q_reg[1]  ( .D(n66), .CK(clk), .RN(n39), .Q(Q[1]), .QN(net645109)
         );
  DFFR_X1 \Q_reg[0]  ( .D(n65), .CK(clk), .RN(n39), .Q(Q[0]), .QN(net645108)
         );
  DFFR_X1 \Q_reg[20]  ( .D(n85), .CK(clk), .RN(n39), .Q(Q[20]), .QN(net645107)
         );
  NAND2_X1 U3 ( .A1(en), .A2(D[31]), .ZN(n101) );
  OAI21_X1 U2 ( .B1(en), .B2(net645138), .A(n101), .ZN(n97) );
  NAND2_X1 U19 ( .A1(en), .A2(D[23]), .ZN(n62) );
  OAI21_X1 U18 ( .B1(en), .B2(net645130), .A(n62), .ZN(n88) );
  NAND2_X1 U11 ( .A1(en), .A2(D[27]), .ZN(n98) );
  OAI21_X1 U10 ( .B1(en), .B2(net645134), .A(n98), .ZN(n92) );
  NAND2_X1 U21 ( .A1(en), .A2(D[22]), .ZN(n61) );
  OAI21_X1 U20 ( .B1(n38), .B2(net645129), .A(n61), .ZN(n87) );
  NAND2_X1 U13 ( .A1(en), .A2(D[26]), .ZN(n96) );
  OAI21_X1 U12 ( .B1(en), .B2(net645133), .A(n96), .ZN(n91) );
  NAND2_X1 U7 ( .A1(en), .A2(D[29]), .ZN(n100) );
  OAI21_X1 U6 ( .B1(n38), .B2(net645136), .A(n100), .ZN(n94) );
  NAND2_X1 U9 ( .A1(en), .A2(D[28]), .ZN(n99) );
  OAI21_X1 U8 ( .B1(en), .B2(net645135), .A(n99), .ZN(n93) );
  NAND2_X1 U15 ( .A1(en), .A2(D[25]), .ZN(n64) );
  OAI21_X1 U14 ( .B1(en), .B2(net645132), .A(n64), .ZN(n90) );
  NAND2_X1 U23 ( .A1(en), .A2(D[21]), .ZN(n60) );
  OAI21_X1 U22 ( .B1(en), .B2(net645128), .A(n60), .ZN(n86) );
  NAND2_X1 U25 ( .A1(en), .A2(D[20]), .ZN(n59) );
  OAI21_X1 U24 ( .B1(en), .B2(net645107), .A(n59), .ZN(n85) );
  NAND2_X1 U17 ( .A1(en), .A2(D[24]), .ZN(n63) );
  OAI21_X1 U16 ( .B1(en), .B2(net645131), .A(n63), .ZN(n89) );
  NAND2_X1 U27 ( .A1(en), .A2(D[19]), .ZN(n58) );
  OAI21_X1 U26 ( .B1(en), .B2(net645127), .A(n58), .ZN(n84) );
  NAND2_X1 U39 ( .A1(n38), .A2(D[13]), .ZN(n53) );
  OAI21_X1 U38 ( .B1(en), .B2(net645121), .A(n53), .ZN(n78) );
  NAND2_X1 U37 ( .A1(n38), .A2(D[14]), .ZN(n54) );
  OAI21_X1 U36 ( .B1(n38), .B2(net645122), .A(n54), .ZN(n79) );
  NAND2_X1 U41 ( .A1(en), .A2(D[12]), .ZN(n52) );
  OAI21_X1 U40 ( .B1(en), .B2(net645120), .A(n52), .ZN(n77) );
  NAND2_X1 U35 ( .A1(en), .A2(D[15]), .ZN(n55) );
  OAI21_X1 U34 ( .B1(en), .B2(net645123), .A(n55), .ZN(n80) );
  NAND2_X1 U51 ( .A1(en), .A2(D[7]), .ZN(n47) );
  OAI21_X1 U50 ( .B1(en), .B2(net645115), .A(n47), .ZN(n72) );
  NAND2_X1 U43 ( .A1(n38), .A2(D[11]), .ZN(n51) );
  OAI21_X1 U42 ( .B1(en), .B2(net645119), .A(n51), .ZN(n76) );
  NAND2_X1 U49 ( .A1(en), .A2(D[8]), .ZN(n48) );
  OAI21_X1 U48 ( .B1(n38), .B2(net645116), .A(n48), .ZN(n73) );
  NAND2_X1 U47 ( .A1(en), .A2(D[9]), .ZN(n49) );
  OAI21_X1 U46 ( .B1(en), .B2(net645117), .A(n49), .ZN(n74) );
  NAND2_X1 U31 ( .A1(en), .A2(D[17]), .ZN(n56) );
  OAI21_X1 U30 ( .B1(en), .B2(net645125), .A(n56), .ZN(n82) );
  NAND2_X1 U29 ( .A1(en), .A2(D[18]), .ZN(n57) );
  OAI21_X1 U28 ( .B1(en), .B2(net645126), .A(n57), .ZN(n83) );
  NAND2_X1 U45 ( .A1(n38), .A2(D[10]), .ZN(n50) );
  OAI21_X1 U44 ( .B1(en), .B2(net645118), .A(n50), .ZN(n75) );
  NAND2_X1 U59 ( .A1(en), .A2(D[3]), .ZN(n43) );
  OAI21_X1 U58 ( .B1(n38), .B2(net645111), .A(n43), .ZN(n68) );
  NAND2_X1 U53 ( .A1(en), .A2(D[6]), .ZN(n46) );
  OAI21_X1 U52 ( .B1(n38), .B2(net645114), .A(n46), .ZN(n71) );
  NAND2_X1 U55 ( .A1(en), .A2(D[5]), .ZN(n45) );
  OAI21_X1 U54 ( .B1(n38), .B2(net645113), .A(n45), .ZN(n70) );
  NAND2_X1 U57 ( .A1(en), .A2(D[4]), .ZN(n44) );
  OAI21_X1 U56 ( .B1(n38), .B2(net645112), .A(n44), .ZN(n69) );
  NAND2_X1 U61 ( .A1(en), .A2(D[2]), .ZN(n42) );
  OAI21_X1 U60 ( .B1(n38), .B2(net645110), .A(n42), .ZN(n67) );
  NAND2_X1 U63 ( .A1(en), .A2(D[1]), .ZN(n41) );
  OAI21_X1 U62 ( .B1(n38), .B2(net645109), .A(n41), .ZN(n66) );
  NAND2_X1 U65 ( .A1(en), .A2(D[0]), .ZN(n40) );
  OAI21_X1 U64 ( .B1(n38), .B2(net645108), .A(n40), .ZN(n65) );
  NAND2_X1 U4 ( .A1(en), .A2(D[16]), .ZN(n35) );
  OAI21_X1 U5 ( .B1(en), .B2(net645124), .A(n35), .ZN(n81) );
  NAND2_X1 U32 ( .A1(en), .A2(D[30]), .ZN(n36) );
  OAI21_X1 U33 ( .B1(en), .B2(net645137), .A(n36), .ZN(n95) );
  INV_X2 U66 ( .A(rst), .ZN(n39) );
  BUF_X1 U67 ( .A(en), .Z(n38) );
endmodule


module p4add_N32_logN5_1 ( A, B, Cin, sign, S, Cout );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input Cin, sign;
  output Cout;
  wire   n1, n2, n3, n5, n6, n10, n11, n12, n13, n14, n15, n16, n17, n19, n22,
         n23, n24, n27, n28, n29, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47;
  wire   [31:0] new_B;
  wire   [7:0] carry_pro;

  xor_gen_N32_1 xor32 ( .A(B), .B(sign), .S({new_B[31:28], n29, n1, n14, 
        new_B[24:21], n33, n13, n28, n22, new_B[16], n3, n16, n6, new_B[12], 
        n2, n17, n15, n5, n32, n31, n19, n23, n12, n11, n24, n10}) );
  carry_tree_N32_logN5_1 ct ( .A(A), .B({new_B[31:28], n29, n1, n14, 
        new_B[24:21], n33, n13, n28, n22, new_B[16], n3, n16, n6, new_B[12], 
        n2, n17, n15, n5, n32, n31, n19, n23, n12, n11, n24, n10}), .Cin(sign), 
        .Cout({Cout, carry_pro[7:1]}) );
  sum_gen_N32_1 add ( .A(A), .B({new_B[31:28], n29, n1, n40, new_B[24], n47, 
        n41, n34, n33, n38, n28, n45, new_B[16], n3, n42, n36, new_B[12], n37, 
        n39, n27, n5, n32, n43, n19, n23, n35, n46, n24, n44}), .Cin({1'b0, 
        carry_pro[7:1], sign}), .S(S) );
  BUF_X1 U1 ( .A(n15), .Z(n27) );
  BUF_X1 U2 ( .A(n6), .Z(n36) );
  BUF_X1 U3 ( .A(n12), .Z(n35) );
  BUF_X1 U4 ( .A(new_B[22]), .Z(n41) );
  BUF_X1 U5 ( .A(n13), .Z(n38) );
  BUF_X1 U6 ( .A(n10), .Z(n44) );
  BUF_X1 U7 ( .A(n31), .Z(n43) );
  BUF_X1 U8 ( .A(new_B[21]), .Z(n34) );
  BUF_X1 U9 ( .A(n14), .Z(n40) );
  CLKBUF_X1 U10 ( .A(n2), .Z(n37) );
  CLKBUF_X1 U11 ( .A(n17), .Z(n39) );
  CLKBUF_X1 U12 ( .A(new_B[23]), .Z(n47) );
  CLKBUF_X1 U13 ( .A(n16), .Z(n42) );
  CLKBUF_X1 U14 ( .A(n22), .Z(n45) );
  CLKBUF_X1 U15 ( .A(n11), .Z(n46) );
endmodule


module predictor_2_14 ( clock, reset, enable, taken_i, prediction_o );
  input clock, reset, enable, taken_i;
  output prediction_o;
  wire   N11, N12, n5, n6, n8, n10, n12, n13, n14;
  wire   [1:0] next_STATE;

  DLH_X1 \next_STATE_reg[0]  ( .G(enable), .D(N11), .Q(next_STATE[0]) );
  DFFR_X1 \STATE_reg[0]  ( .D(n6), .CK(clock), .RN(n12), .Q(n5), .QN(n10) );
  DLH_X1 \next_STATE_reg[1]  ( .G(enable), .D(N12), .Q(next_STATE[1]) );
  DFFR_X1 \STATE_reg[1]  ( .D(n8), .CK(clock), .RN(n12), .Q(prediction_o) );
  MUX2_X1 U8 ( .A(prediction_o), .B(next_STATE[1]), .S(enable), .Z(n8) );
  MUX2_X1 U9 ( .A(n5), .B(next_STATE[0]), .S(enable), .Z(n6) );
  NOR2_X1 U7 ( .A1(prediction_o), .A2(taken_i), .ZN(n14) );
  NAND2_X1 U6 ( .A1(prediction_o), .A2(taken_i), .ZN(n13) );
  OAI21_X1 U3 ( .B1(n14), .B2(n10), .A(n13), .ZN(N12) );
  OAI21_X1 U5 ( .B1(n5), .B2(n14), .A(n13), .ZN(N11) );
  INV_X1 U2 ( .A(reset), .ZN(n12) );
endmodule


module predictor_2_13 ( clock, reset, enable, taken_i, prediction_o );
  input clock, reset, enable, taken_i;
  output prediction_o;
  wire   N11, N12, n5, n6, n8, n10, n12, n13, n14;
  wire   [1:0] next_STATE;

  DLH_X1 \next_STATE_reg[0]  ( .G(enable), .D(N11), .Q(next_STATE[0]) );
  DFFR_X1 \STATE_reg[0]  ( .D(n6), .CK(clock), .RN(n12), .Q(n5), .QN(n10) );
  DLH_X1 \next_STATE_reg[1]  ( .G(enable), .D(N12), .Q(next_STATE[1]) );
  DFFR_X1 \STATE_reg[1]  ( .D(n8), .CK(clock), .RN(n12), .Q(prediction_o) );
  MUX2_X1 U8 ( .A(prediction_o), .B(next_STATE[1]), .S(enable), .Z(n8) );
  MUX2_X1 U9 ( .A(n5), .B(next_STATE[0]), .S(enable), .Z(n6) );
  NOR2_X1 U7 ( .A1(prediction_o), .A2(taken_i), .ZN(n14) );
  NAND2_X1 U6 ( .A1(prediction_o), .A2(taken_i), .ZN(n13) );
  OAI21_X1 U5 ( .B1(n5), .B2(n14), .A(n13), .ZN(N11) );
  OAI21_X1 U3 ( .B1(n14), .B2(n10), .A(n13), .ZN(N12) );
  INV_X1 U2 ( .A(reset), .ZN(n12) );
endmodule


module predictor_2_12 ( clock, reset, enable, taken_i, prediction_o );
  input clock, reset, enable, taken_i;
  output prediction_o;
  wire   N11, N12, n5, n6, n8, n10, n12, n13, n14;
  wire   [1:0] next_STATE;

  DLH_X1 \next_STATE_reg[0]  ( .G(enable), .D(N11), .Q(next_STATE[0]) );
  DFFR_X1 \STATE_reg[0]  ( .D(n6), .CK(clock), .RN(n12), .Q(n5), .QN(n10) );
  DLH_X1 \next_STATE_reg[1]  ( .G(enable), .D(N12), .Q(next_STATE[1]) );
  DFFR_X1 \STATE_reg[1]  ( .D(n8), .CK(clock), .RN(n12), .Q(prediction_o) );
  MUX2_X1 U8 ( .A(prediction_o), .B(next_STATE[1]), .S(enable), .Z(n8) );
  MUX2_X1 U9 ( .A(n5), .B(next_STATE[0]), .S(enable), .Z(n6) );
  NOR2_X1 U7 ( .A1(prediction_o), .A2(taken_i), .ZN(n14) );
  NAND2_X1 U6 ( .A1(prediction_o), .A2(taken_i), .ZN(n13) );
  OAI21_X1 U5 ( .B1(n5), .B2(n14), .A(n13), .ZN(N11) );
  OAI21_X1 U3 ( .B1(n14), .B2(n10), .A(n13), .ZN(N12) );
  INV_X1 U2 ( .A(reset), .ZN(n12) );
endmodule


module predictor_2_11 ( clock, reset, enable, taken_i, prediction_o );
  input clock, reset, enable, taken_i;
  output prediction_o;
  wire   N11, N12, n5, n6, n8, n10, n12, n13, n14;
  wire   [1:0] next_STATE;

  DLH_X1 \next_STATE_reg[0]  ( .G(enable), .D(N11), .Q(next_STATE[0]) );
  DFFR_X1 \STATE_reg[0]  ( .D(n6), .CK(clock), .RN(n12), .Q(n5), .QN(n10) );
  DLH_X1 \next_STATE_reg[1]  ( .G(enable), .D(N12), .Q(next_STATE[1]) );
  DFFR_X1 \STATE_reg[1]  ( .D(n8), .CK(clock), .RN(n12), .Q(prediction_o) );
  MUX2_X1 U8 ( .A(prediction_o), .B(next_STATE[1]), .S(enable), .Z(n8) );
  MUX2_X1 U9 ( .A(n5), .B(next_STATE[0]), .S(enable), .Z(n6) );
  NOR2_X1 U7 ( .A1(prediction_o), .A2(taken_i), .ZN(n14) );
  NAND2_X1 U6 ( .A1(prediction_o), .A2(taken_i), .ZN(n13) );
  OAI21_X1 U5 ( .B1(n5), .B2(n14), .A(n13), .ZN(N11) );
  OAI21_X1 U3 ( .B1(n14), .B2(n10), .A(n13), .ZN(N12) );
  INV_X1 U2 ( .A(reset), .ZN(n12) );
endmodule


module predictor_2_10 ( clock, reset, enable, taken_i, prediction_o );
  input clock, reset, enable, taken_i;
  output prediction_o;
  wire   N11, N12, n5, n6, n8, n10, n12, n13, n14;
  wire   [1:0] next_STATE;

  DLH_X1 \next_STATE_reg[0]  ( .G(enable), .D(N11), .Q(next_STATE[0]) );
  DFFR_X1 \STATE_reg[0]  ( .D(n6), .CK(clock), .RN(n12), .Q(n5), .QN(n10) );
  DLH_X1 \next_STATE_reg[1]  ( .G(enable), .D(N12), .Q(next_STATE[1]) );
  DFFR_X1 \STATE_reg[1]  ( .D(n8), .CK(clock), .RN(n12), .Q(prediction_o) );
  MUX2_X1 U8 ( .A(prediction_o), .B(next_STATE[1]), .S(enable), .Z(n8) );
  MUX2_X1 U9 ( .A(n5), .B(next_STATE[0]), .S(enable), .Z(n6) );
  NOR2_X1 U7 ( .A1(prediction_o), .A2(taken_i), .ZN(n14) );
  NAND2_X1 U6 ( .A1(prediction_o), .A2(taken_i), .ZN(n13) );
  OAI21_X1 U3 ( .B1(n14), .B2(n10), .A(n13), .ZN(N12) );
  OAI21_X1 U5 ( .B1(n5), .B2(n14), .A(n13), .ZN(N11) );
  INV_X1 U2 ( .A(reset), .ZN(n12) );
endmodule


module predictor_2_9 ( clock, reset, enable, taken_i, prediction_o );
  input clock, reset, enable, taken_i;
  output prediction_o;
  wire   N11, N12, n5, n6, n8, n10, n12, n13, n14;
  wire   [1:0] next_STATE;

  DLH_X1 \next_STATE_reg[0]  ( .G(enable), .D(N11), .Q(next_STATE[0]) );
  DFFR_X1 \STATE_reg[0]  ( .D(n6), .CK(clock), .RN(n12), .Q(n5), .QN(n10) );
  DLH_X1 \next_STATE_reg[1]  ( .G(enable), .D(N12), .Q(next_STATE[1]) );
  DFFR_X1 \STATE_reg[1]  ( .D(n8), .CK(clock), .RN(n12), .Q(prediction_o) );
  MUX2_X1 U8 ( .A(prediction_o), .B(next_STATE[1]), .S(enable), .Z(n8) );
  MUX2_X1 U9 ( .A(n5), .B(next_STATE[0]), .S(enable), .Z(n6) );
  NOR2_X1 U7 ( .A1(prediction_o), .A2(taken_i), .ZN(n14) );
  NAND2_X1 U6 ( .A1(prediction_o), .A2(taken_i), .ZN(n13) );
  OAI21_X1 U3 ( .B1(n14), .B2(n10), .A(n13), .ZN(N12) );
  OAI21_X1 U5 ( .B1(n5), .B2(n14), .A(n13), .ZN(N11) );
  INV_X1 U2 ( .A(reset), .ZN(n12) );
endmodule


module predictor_2_8 ( clock, reset, enable, taken_i, prediction_o );
  input clock, reset, enable, taken_i;
  output prediction_o;
  wire   N11, N12, n5, n6, n8, n10, n12, n13, n14;
  wire   [1:0] next_STATE;

  DLH_X1 \next_STATE_reg[0]  ( .G(enable), .D(N11), .Q(next_STATE[0]) );
  DFFR_X1 \STATE_reg[0]  ( .D(n6), .CK(clock), .RN(n12), .Q(n5), .QN(n10) );
  DLH_X1 \next_STATE_reg[1]  ( .G(enable), .D(N12), .Q(next_STATE[1]) );
  DFFR_X1 \STATE_reg[1]  ( .D(n8), .CK(clock), .RN(n12), .Q(prediction_o) );
  MUX2_X1 U8 ( .A(prediction_o), .B(next_STATE[1]), .S(enable), .Z(n8) );
  MUX2_X1 U9 ( .A(n5), .B(next_STATE[0]), .S(enable), .Z(n6) );
  NOR2_X1 U7 ( .A1(prediction_o), .A2(taken_i), .ZN(n14) );
  NAND2_X1 U6 ( .A1(prediction_o), .A2(taken_i), .ZN(n13) );
  OAI21_X1 U3 ( .B1(n14), .B2(n10), .A(n13), .ZN(N12) );
  OAI21_X1 U5 ( .B1(n5), .B2(n14), .A(n13), .ZN(N11) );
  INV_X1 U2 ( .A(reset), .ZN(n12) );
endmodule


module predictor_2_7 ( clock, reset, enable, taken_i, prediction_o );
  input clock, reset, enable, taken_i;
  output prediction_o;
  wire   N11, N12, n5, n6, n8, n10, n12, n13, n14;
  wire   [1:0] next_STATE;

  DLH_X1 \next_STATE_reg[0]  ( .G(enable), .D(N11), .Q(next_STATE[0]) );
  DFFR_X1 \STATE_reg[0]  ( .D(n6), .CK(clock), .RN(n12), .Q(n5), .QN(n10) );
  DLH_X1 \next_STATE_reg[1]  ( .G(enable), .D(N12), .Q(next_STATE[1]) );
  DFFR_X1 \STATE_reg[1]  ( .D(n8), .CK(clock), .RN(n12), .Q(prediction_o) );
  MUX2_X1 U8 ( .A(prediction_o), .B(next_STATE[1]), .S(enable), .Z(n8) );
  MUX2_X1 U9 ( .A(n5), .B(next_STATE[0]), .S(enable), .Z(n6) );
  NOR2_X1 U7 ( .A1(prediction_o), .A2(taken_i), .ZN(n14) );
  NAND2_X1 U6 ( .A1(prediction_o), .A2(taken_i), .ZN(n13) );
  OAI21_X1 U3 ( .B1(n14), .B2(n10), .A(n13), .ZN(N12) );
  OAI21_X1 U5 ( .B1(n5), .B2(n14), .A(n13), .ZN(N11) );
  INV_X1 U2 ( .A(reset), .ZN(n12) );
endmodule


module predictor_2_6 ( clock, reset, enable, taken_i, prediction_o );
  input clock, reset, enable, taken_i;
  output prediction_o;
  wire   N11, N12, n5, n6, n8, n10, n12, n13, n14;
  wire   [1:0] next_STATE;

  DLH_X1 \next_STATE_reg[0]  ( .G(enable), .D(N11), .Q(next_STATE[0]) );
  DFFR_X1 \STATE_reg[0]  ( .D(n6), .CK(clock), .RN(n12), .Q(n5), .QN(n10) );
  DLH_X1 \next_STATE_reg[1]  ( .G(enable), .D(N12), .Q(next_STATE[1]) );
  DFFR_X1 \STATE_reg[1]  ( .D(n8), .CK(clock), .RN(n12), .Q(prediction_o) );
  MUX2_X1 U8 ( .A(prediction_o), .B(next_STATE[1]), .S(enable), .Z(n8) );
  MUX2_X1 U9 ( .A(n5), .B(next_STATE[0]), .S(enable), .Z(n6) );
  NOR2_X1 U7 ( .A1(prediction_o), .A2(taken_i), .ZN(n14) );
  NAND2_X1 U6 ( .A1(prediction_o), .A2(taken_i), .ZN(n13) );
  OAI21_X1 U3 ( .B1(n14), .B2(n10), .A(n13), .ZN(N12) );
  OAI21_X1 U5 ( .B1(n5), .B2(n14), .A(n13), .ZN(N11) );
  INV_X1 U2 ( .A(reset), .ZN(n12) );
endmodule


module predictor_2_5 ( clock, reset, enable, taken_i, prediction_o );
  input clock, reset, enable, taken_i;
  output prediction_o;
  wire   N11, N12, n5, n6, n8, n10, n12, n13, n14;
  wire   [1:0] next_STATE;

  DLH_X1 \next_STATE_reg[0]  ( .G(enable), .D(N11), .Q(next_STATE[0]) );
  DFFR_X1 \STATE_reg[0]  ( .D(n6), .CK(clock), .RN(n12), .Q(n5), .QN(n10) );
  DLH_X1 \next_STATE_reg[1]  ( .G(enable), .D(N12), .Q(next_STATE[1]) );
  DFFR_X1 \STATE_reg[1]  ( .D(n8), .CK(clock), .RN(n12), .Q(prediction_o) );
  MUX2_X1 U8 ( .A(prediction_o), .B(next_STATE[1]), .S(enable), .Z(n8) );
  MUX2_X1 U9 ( .A(n5), .B(next_STATE[0]), .S(enable), .Z(n6) );
  NOR2_X1 U7 ( .A1(prediction_o), .A2(taken_i), .ZN(n14) );
  NAND2_X1 U6 ( .A1(prediction_o), .A2(taken_i), .ZN(n13) );
  OAI21_X1 U5 ( .B1(n5), .B2(n14), .A(n13), .ZN(N11) );
  OAI21_X1 U3 ( .B1(n14), .B2(n10), .A(n13), .ZN(N12) );
  INV_X1 U2 ( .A(reset), .ZN(n12) );
endmodule


module predictor_2_4 ( clock, reset, enable, taken_i, prediction_o );
  input clock, reset, enable, taken_i;
  output prediction_o;
  wire   N11, N12, n5, n6, n8, n10, n12, n13, n14;
  wire   [1:0] next_STATE;

  DLH_X1 \next_STATE_reg[0]  ( .G(enable), .D(N11), .Q(next_STATE[0]) );
  DFFR_X1 \STATE_reg[0]  ( .D(n6), .CK(clock), .RN(n12), .Q(n5), .QN(n10) );
  DLH_X1 \next_STATE_reg[1]  ( .G(enable), .D(N12), .Q(next_STATE[1]) );
  DFFR_X1 \STATE_reg[1]  ( .D(n8), .CK(clock), .RN(n12), .Q(prediction_o) );
  MUX2_X1 U8 ( .A(prediction_o), .B(next_STATE[1]), .S(enable), .Z(n8) );
  MUX2_X1 U9 ( .A(n5), .B(next_STATE[0]), .S(enable), .Z(n6) );
  NOR2_X1 U7 ( .A1(prediction_o), .A2(taken_i), .ZN(n14) );
  NAND2_X1 U6 ( .A1(prediction_o), .A2(taken_i), .ZN(n13) );
  OAI21_X1 U3 ( .B1(n14), .B2(n10), .A(n13), .ZN(N12) );
  OAI21_X1 U5 ( .B1(n5), .B2(n14), .A(n13), .ZN(N11) );
  INV_X1 U2 ( .A(reset), .ZN(n12) );
endmodule


module predictor_2_3 ( clock, reset, enable, taken_i, prediction_o );
  input clock, reset, enable, taken_i;
  output prediction_o;
  wire   N11, N12, n5, n6, n8, n10, n12, n13, n14;
  wire   [1:0] next_STATE;

  DLH_X1 \next_STATE_reg[0]  ( .G(enable), .D(N11), .Q(next_STATE[0]) );
  DFFR_X1 \STATE_reg[0]  ( .D(n6), .CK(clock), .RN(n12), .Q(n5), .QN(n10) );
  DLH_X1 \next_STATE_reg[1]  ( .G(enable), .D(N12), .Q(next_STATE[1]) );
  DFFR_X1 \STATE_reg[1]  ( .D(n8), .CK(clock), .RN(n12), .Q(prediction_o) );
  MUX2_X1 U8 ( .A(prediction_o), .B(next_STATE[1]), .S(enable), .Z(n8) );
  MUX2_X1 U9 ( .A(n5), .B(next_STATE[0]), .S(enable), .Z(n6) );
  NOR2_X1 U7 ( .A1(prediction_o), .A2(taken_i), .ZN(n14) );
  NAND2_X1 U6 ( .A1(prediction_o), .A2(taken_i), .ZN(n13) );
  OAI21_X1 U5 ( .B1(n5), .B2(n14), .A(n13), .ZN(N11) );
  OAI21_X1 U3 ( .B1(n14), .B2(n10), .A(n13), .ZN(N12) );
  INV_X1 U2 ( .A(reset), .ZN(n12) );
endmodule


module predictor_2_2 ( clock, reset, enable, taken_i, prediction_o );
  input clock, reset, enable, taken_i;
  output prediction_o;
  wire   N11, N12, n5, n6, n8, n10, n12, n13, n14;
  wire   [1:0] next_STATE;

  DLH_X1 \next_STATE_reg[0]  ( .G(enable), .D(N11), .Q(next_STATE[0]) );
  DFFR_X1 \STATE_reg[0]  ( .D(n6), .CK(clock), .RN(n12), .Q(n5), .QN(n10) );
  DLH_X1 \next_STATE_reg[1]  ( .G(enable), .D(N12), .Q(next_STATE[1]) );
  DFFR_X1 \STATE_reg[1]  ( .D(n8), .CK(clock), .RN(n12), .Q(prediction_o) );
  MUX2_X1 U8 ( .A(prediction_o), .B(next_STATE[1]), .S(enable), .Z(n8) );
  MUX2_X1 U9 ( .A(n5), .B(next_STATE[0]), .S(enable), .Z(n6) );
  NOR2_X1 U7 ( .A1(prediction_o), .A2(taken_i), .ZN(n14) );
  NAND2_X1 U6 ( .A1(prediction_o), .A2(taken_i), .ZN(n13) );
  OAI21_X1 U5 ( .B1(n5), .B2(n14), .A(n13), .ZN(N11) );
  OAI21_X1 U3 ( .B1(n14), .B2(n10), .A(n13), .ZN(N12) );
  INV_X1 U2 ( .A(reset), .ZN(n12) );
endmodule


module predictor_2_1 ( clock, reset, enable, taken_i, prediction_o );
  input clock, reset, enable, taken_i;
  output prediction_o;
  wire   N11, N12, n5, n6, n8, n10, n12, n13, n14;
  wire   [1:0] next_STATE;

  DLH_X1 \next_STATE_reg[0]  ( .G(enable), .D(N11), .Q(next_STATE[0]) );
  DFFR_X1 \STATE_reg[0]  ( .D(n6), .CK(clock), .RN(n12), .Q(n5), .QN(n10) );
  DLH_X1 \next_STATE_reg[1]  ( .G(enable), .D(N12), .Q(next_STATE[1]) );
  DFFR_X1 \STATE_reg[1]  ( .D(n8), .CK(clock), .RN(n12), .Q(prediction_o) );
  MUX2_X1 U8 ( .A(prediction_o), .B(next_STATE[1]), .S(enable), .Z(n8) );
  MUX2_X1 U9 ( .A(n5), .B(next_STATE[0]), .S(enable), .Z(n6) );
  NOR2_X1 U7 ( .A1(prediction_o), .A2(taken_i), .ZN(n14) );
  NAND2_X1 U6 ( .A1(prediction_o), .A2(taken_i), .ZN(n13) );
  OAI21_X1 U3 ( .B1(n14), .B2(n10), .A(n13), .ZN(N12) );
  OAI21_X1 U5 ( .B1(n5), .B2(n14), .A(n13), .ZN(N11) );
  INV_X1 U2 ( .A(reset), .ZN(n12) );
endmodule


module mux41_1 ( IN0, IN1, IN2, IN3, CTRL, OUT1 );
  input [31:0] IN0;
  input [31:0] IN1;
  input [31:0] IN2;
  input [31:0] IN3;
  input [1:0] CTRL;
  output [31:0] OUT1;
  wire   n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n157, n158;

  NAND2_X1 U1 ( .A1(n91), .A2(n90), .ZN(OUT1[11]) );
  CLKBUF_X3 U2 ( .A(n156), .Z(n127) );
  INV_X1 U3 ( .A(CTRL[0]), .ZN(n110) );
  AND2_X1 U4 ( .A1(CTRL[1]), .A2(n110), .ZN(n78) );
  AND2_X1 U5 ( .A1(CTRL[1]), .A2(CTRL[0]), .ZN(n158) );
  CLKBUF_X3 U6 ( .A(n157), .Z(n130) );
  CLKBUF_X3 U7 ( .A(n157), .Z(n129) );
  CLKBUF_X3 U8 ( .A(n157), .Z(n128) );
  CLKBUF_X3 U9 ( .A(n156), .Z(n125) );
  CLKBUF_X3 U10 ( .A(n156), .Z(n126) );
  BUF_X2 U11 ( .A(n78), .Z(n79) );
  BUF_X2 U12 ( .A(n158), .Z(n133) );
  BUF_X2 U13 ( .A(n158), .Z(n132) );
  BUF_X2 U14 ( .A(n78), .Z(n80) );
  BUF_X2 U15 ( .A(n78), .Z(n81) );
  BUF_X2 U16 ( .A(n158), .Z(n131) );
  AOI22_X1 U17 ( .A1(n131), .A2(IN3[15]), .B1(n80), .B2(IN2[15]), .ZN(n83) );
  AOI22_X1 U18 ( .A1(n131), .A2(IN3[18]), .B1(n79), .B2(IN2[18]), .ZN(n103) );
  AOI22_X1 U19 ( .A1(n132), .A2(IN3[29]), .B1(n80), .B2(IN2[29]), .ZN(n105) );
  AOI22_X1 U20 ( .A1(n131), .A2(IN3[16]), .B1(n81), .B2(IN2[16]), .ZN(n112) );
  AOI22_X1 U21 ( .A1(n132), .A2(IN3[22]), .B1(n79), .B2(IN2[22]), .ZN(n116) );
  AOI22_X1 U22 ( .A1(n131), .A2(IN3[19]), .B1(n79), .B2(IN2[19]), .ZN(n118) );
  AOI22_X1 U23 ( .A1(n131), .A2(IN3[12]), .B1(n80), .B2(IN2[12]), .ZN(n120) );
  AOI22_X1 U24 ( .A1(n133), .A2(IN3[4]), .B1(n79), .B2(IN2[4]), .ZN(n124) );
  AOI22_X1 U25 ( .A1(n133), .A2(IN3[6]), .B1(n81), .B2(IN2[6]), .ZN(n152) );
  AOI22_X1 U26 ( .A1(n131), .A2(IN3[1]), .B1(n81), .B2(IN2[1]), .ZN(n138) );
  AOI22_X1 U27 ( .A1(n133), .A2(IN3[31]), .B1(n79), .B2(IN2[31]), .ZN(n85) );
  AOI22_X1 U28 ( .A1(n131), .A2(IN3[10]), .B1(n81), .B2(IN2[10]), .ZN(n93) );
  AOI22_X1 U29 ( .A1(n132), .A2(IN3[23]), .B1(n81), .B2(IN2[23]), .ZN(n97) );
  AOI22_X1 U30 ( .A1(n133), .A2(IN3[3]), .B1(n79), .B2(IN2[3]), .ZN(n107) );
  AOI22_X1 U31 ( .A1(n132), .A2(IN3[2]), .B1(n79), .B2(IN2[2]), .ZN(n109) );
  AOI22_X1 U32 ( .A1(n133), .A2(IN3[5]), .B1(n80), .B2(IN2[5]), .ZN(n114) );
  AOI22_X1 U33 ( .A1(n131), .A2(IN3[17]), .B1(n79), .B2(IN2[17]), .ZN(n122) );
  AOI22_X1 U34 ( .A1(n131), .A2(IN3[13]), .B1(n81), .B2(IN2[13]), .ZN(n136) );
  AOI22_X1 U35 ( .A1(n132), .A2(IN3[21]), .B1(n80), .B2(IN2[21]), .ZN(n142) );
  AOI22_X1 U36 ( .A1(n131), .A2(IN3[0]), .B1(n80), .B2(IN2[0]), .ZN(n134) );
  AOI22_X1 U37 ( .A1(n133), .A2(IN3[8]), .B1(n81), .B2(IN2[8]), .ZN(n154) );
  AOI22_X1 U38 ( .A1(n131), .A2(IN3[14]), .B1(n80), .B2(IN2[14]), .ZN(n87) );
  AOI22_X1 U39 ( .A1(n133), .A2(IN3[9]), .B1(n81), .B2(IN2[9]), .ZN(n89) );
  AOI22_X1 U40 ( .A1(n131), .A2(IN3[11]), .B1(n79), .B2(IN2[11]), .ZN(n91) );
  AOI22_X1 U41 ( .A1(n133), .A2(IN3[7]), .B1(n80), .B2(IN2[7]), .ZN(n95) );
  AOI22_X1 U42 ( .A1(n132), .A2(IN3[26]), .B1(n80), .B2(IN2[26]), .ZN(n99) );
  AOI22_X1 U43 ( .A1(n132), .A2(IN3[27]), .B1(n79), .B2(IN2[27]), .ZN(n101) );
  AOI22_X1 U44 ( .A1(n132), .A2(IN3[28]), .B1(n79), .B2(IN2[28]), .ZN(n148) );
  AOI22_X1 U45 ( .A1(n132), .A2(IN3[30]), .B1(n80), .B2(IN2[30]), .ZN(n150) );
  AOI22_X1 U46 ( .A1(n132), .A2(IN3[25]), .B1(n81), .B2(IN2[25]), .ZN(n146) );
  AOI22_X1 U47 ( .A1(n132), .A2(IN3[24]), .B1(n81), .B2(IN2[24]), .ZN(n144) );
  AOI22_X1 U48 ( .A1(n132), .A2(IN3[20]), .B1(n80), .B2(IN2[20]), .ZN(n140) );
  NAND2_X1 U49 ( .A1(n121), .A2(n122), .ZN(OUT1[17]) );
  NAND2_X1 U50 ( .A1(n92), .A2(n93), .ZN(OUT1[10]) );
  NAND2_X1 U51 ( .A1(n86), .A2(n87), .ZN(OUT1[14]) );
  NAND2_X1 U52 ( .A1(n111), .A2(n112), .ZN(OUT1[16]) );
  NAND2_X1 U53 ( .A1(n102), .A2(n103), .ZN(OUT1[18]) );
  NAND2_X1 U54 ( .A1(n82), .A2(n83), .ZN(OUT1[15]) );
  NAND2_X1 U55 ( .A1(n84), .A2(n85), .ZN(OUT1[31]) );
  AOI22_X1 U56 ( .A1(n130), .A2(IN1[15]), .B1(n125), .B2(IN0[15]), .ZN(n82) );
  AOI22_X1 U57 ( .A1(n130), .A2(IN1[31]), .B1(n126), .B2(IN0[31]), .ZN(n84) );
  NOR2_X1 U58 ( .A1(n110), .A2(CTRL[1]), .ZN(n157) );
  AOI22_X1 U59 ( .A1(n128), .A2(IN1[14]), .B1(n125), .B2(IN0[14]), .ZN(n86) );
  AOI22_X1 U60 ( .A1(n128), .A2(IN1[9]), .B1(n125), .B2(IN0[9]), .ZN(n88) );
  NAND2_X1 U61 ( .A1(n88), .A2(n89), .ZN(OUT1[9]) );
  AOI22_X1 U62 ( .A1(n128), .A2(IN1[11]), .B1(n126), .B2(IN0[11]), .ZN(n90) );
  AOI22_X1 U63 ( .A1(n128), .A2(IN1[10]), .B1(n125), .B2(IN0[10]), .ZN(n92) );
  AOI22_X1 U64 ( .A1(n129), .A2(IN1[7]), .B1(n126), .B2(IN0[7]), .ZN(n94) );
  NAND2_X1 U65 ( .A1(n94), .A2(n95), .ZN(OUT1[7]) );
  AOI22_X1 U66 ( .A1(n129), .A2(IN1[23]), .B1(n127), .B2(IN0[23]), .ZN(n96) );
  NAND2_X1 U67 ( .A1(n96), .A2(n97), .ZN(OUT1[23]) );
  AOI22_X1 U68 ( .A1(n128), .A2(IN1[26]), .B1(n127), .B2(IN0[26]), .ZN(n98) );
  NAND2_X1 U69 ( .A1(n98), .A2(n99), .ZN(OUT1[26]) );
  AOI22_X1 U70 ( .A1(n129), .A2(IN1[27]), .B1(n127), .B2(IN0[27]), .ZN(n100)
         );
  NAND2_X1 U71 ( .A1(n100), .A2(n101), .ZN(OUT1[27]) );
  AOI22_X1 U72 ( .A1(n129), .A2(IN1[18]), .B1(n126), .B2(IN0[18]), .ZN(n102)
         );
  AOI22_X1 U73 ( .A1(n128), .A2(IN1[29]), .B1(n127), .B2(IN0[29]), .ZN(n104)
         );
  NAND2_X1 U74 ( .A1(n104), .A2(n105), .ZN(OUT1[29]) );
  AOI22_X1 U75 ( .A1(n128), .A2(IN1[3]), .B1(n125), .B2(IN0[3]), .ZN(n106) );
  NAND2_X1 U76 ( .A1(n106), .A2(n107), .ZN(OUT1[3]) );
  AOI22_X1 U77 ( .A1(n130), .A2(IN1[2]), .B1(n127), .B2(IN0[2]), .ZN(n108) );
  NAND2_X1 U78 ( .A1(n108), .A2(n109), .ZN(OUT1[2]) );
  AOI22_X1 U79 ( .A1(n129), .A2(IN1[16]), .B1(n125), .B2(IN0[16]), .ZN(n111)
         );
  AOI22_X1 U80 ( .A1(n128), .A2(IN1[5]), .B1(n126), .B2(IN0[5]), .ZN(n113) );
  NAND2_X1 U81 ( .A1(n113), .A2(n114), .ZN(OUT1[5]) );
  AOI22_X1 U82 ( .A1(n129), .A2(IN1[22]), .B1(n126), .B2(IN0[22]), .ZN(n115)
         );
  NAND2_X1 U83 ( .A1(n115), .A2(n116), .ZN(OUT1[22]) );
  AOI22_X1 U84 ( .A1(n129), .A2(IN1[19]), .B1(n127), .B2(IN0[19]), .ZN(n117)
         );
  NAND2_X1 U85 ( .A1(n117), .A2(n118), .ZN(OUT1[19]) );
  AOI22_X1 U86 ( .A1(n128), .A2(IN1[12]), .B1(n125), .B2(IN0[12]), .ZN(n119)
         );
  NAND2_X1 U87 ( .A1(n119), .A2(n120), .ZN(OUT1[12]) );
  AOI22_X1 U88 ( .A1(n129), .A2(IN1[17]), .B1(n126), .B2(IN0[17]), .ZN(n121)
         );
  AOI22_X1 U89 ( .A1(n128), .A2(IN1[4]), .B1(n127), .B2(IN0[4]), .ZN(n123) );
  NAND2_X1 U90 ( .A1(n123), .A2(n124), .ZN(OUT1[4]) );
  NOR2_X1 U91 ( .A1(CTRL[0]), .A2(CTRL[1]), .ZN(n156) );
  NAND2_X1 U92 ( .A1(n151), .A2(n150), .ZN(OUT1[30]) );
  NAND2_X1 U93 ( .A1(n149), .A2(n148), .ZN(OUT1[28]) );
  NAND2_X1 U94 ( .A1(n153), .A2(n152), .ZN(OUT1[6]) );
  NAND2_X1 U95 ( .A1(n135), .A2(n134), .ZN(OUT1[0]) );
  NAND2_X1 U96 ( .A1(n139), .A2(n138), .ZN(OUT1[1]) );
  NAND2_X1 U97 ( .A1(n147), .A2(n146), .ZN(OUT1[25]) );
  NAND2_X1 U98 ( .A1(n141), .A2(n140), .ZN(OUT1[20]) );
  NAND2_X1 U99 ( .A1(n145), .A2(n144), .ZN(OUT1[24]) );
  NAND2_X1 U100 ( .A1(n143), .A2(n142), .ZN(OUT1[21]) );
  NAND2_X1 U101 ( .A1(n137), .A2(n136), .ZN(OUT1[13]) );
  NAND2_X1 U102 ( .A1(n155), .A2(n154), .ZN(OUT1[8]) );
  AOI22_X1 U103 ( .A1(n129), .A2(IN1[6]), .B1(n126), .B2(IN0[6]), .ZN(n153) );
  AOI22_X1 U104 ( .A1(n129), .A2(IN1[8]), .B1(n125), .B2(IN0[8]), .ZN(n155) );
  AOI22_X1 U105 ( .A1(n130), .A2(IN1[28]), .B1(n127), .B2(IN0[28]), .ZN(n149)
         );
  AOI22_X1 U106 ( .A1(n130), .A2(IN1[30]), .B1(n126), .B2(IN0[30]), .ZN(n151)
         );
  AOI22_X1 U107 ( .A1(n130), .A2(IN1[20]), .B1(n125), .B2(IN0[20]), .ZN(n141)
         );
  AOI22_X1 U108 ( .A1(n130), .A2(IN1[25]), .B1(n127), .B2(IN0[25]), .ZN(n147)
         );
  AOI22_X1 U109 ( .A1(n130), .A2(IN1[24]), .B1(n126), .B2(IN0[24]), .ZN(n145)
         );
  AOI22_X1 U110 ( .A1(n130), .A2(IN1[21]), .B1(n127), .B2(IN0[21]), .ZN(n143)
         );
  AOI22_X1 U111 ( .A1(n130), .A2(IN1[0]), .B1(n126), .B2(IN0[0]), .ZN(n135) );
  AOI22_X1 U112 ( .A1(n129), .A2(IN1[1]), .B1(n125), .B2(IN0[1]), .ZN(n139) );
  AOI22_X1 U113 ( .A1(n128), .A2(IN1[13]), .B1(n125), .B2(IN0[13]), .ZN(n137)
         );
endmodule


module booth_encoder_5 ( B_in, A_out );
  input [2:0] B_in;
  output [2:0] A_out;
  wire   N53, N55, N57, n18, n19, n20, n21;
  assign A_out[0] = N53;
  assign A_out[1] = N55;
  assign A_out[2] = N57;

  OAI33_X1 U9 ( .A1(B_in[0]), .A2(B_in[1]), .A3(n18), .B1(n21), .B2(n20), .B3(
        B_in[2]), .ZN(N53) );
  INV_X1 U6 ( .A(B_in[1]), .ZN(n20) );
  INV_X1 U3 ( .A(B_in[2]), .ZN(n18) );
  INV_X1 U4 ( .A(B_in[0]), .ZN(n21) );
  AOI21_X1 U5 ( .B1(B_in[0]), .B2(B_in[1]), .A(n18), .ZN(N55) );
  OAI221_X1 U7 ( .B1(B_in[1]), .B2(n21), .C1(n20), .C2(B_in[2]), .A(n19), .ZN(
        N57) );
  NAND2_X1 U8 ( .A1(B_in[2]), .A2(n21), .ZN(n19) );
endmodule


module booth_encoder_4 ( B_in, A_out );
  input [2:0] B_in;
  output [2:0] A_out;
  wire   N53, N55, N57, n18, n19, n20, n21;
  assign A_out[0] = N53;
  assign A_out[1] = N55;
  assign A_out[2] = N57;

  OAI33_X1 U9 ( .A1(B_in[0]), .A2(B_in[1]), .A3(n18), .B1(n21), .B2(n20), .B3(
        B_in[2]), .ZN(N53) );
  NAND2_X1 U4 ( .A1(B_in[2]), .A2(n21), .ZN(n19) );
  INV_X1 U8 ( .A(B_in[2]), .ZN(n18) );
  INV_X1 U3 ( .A(B_in[0]), .ZN(n21) );
  INV_X1 U5 ( .A(B_in[1]), .ZN(n20) );
  OAI221_X1 U6 ( .B1(B_in[1]), .B2(n21), .C1(n20), .C2(B_in[2]), .A(n19), .ZN(
        N57) );
  AOI21_X1 U7 ( .B1(B_in[0]), .B2(B_in[1]), .A(n18), .ZN(N55) );
endmodule


module booth_encoder_3 ( B_in, A_out );
  input [2:0] B_in;
  output [2:0] A_out;
  wire   N53, N55, N57, n18, n19, n20, n21;
  assign A_out[0] = N53;
  assign A_out[1] = N55;
  assign A_out[2] = N57;

  OAI33_X1 U9 ( .A1(B_in[0]), .A2(B_in[1]), .A3(n18), .B1(n21), .B2(n20), .B3(
        B_in[2]), .ZN(N53) );
  INV_X1 U7 ( .A(B_in[0]), .ZN(n21) );
  INV_X1 U3 ( .A(B_in[2]), .ZN(n18) );
  INV_X1 U4 ( .A(B_in[1]), .ZN(n20) );
  AOI21_X1 U5 ( .B1(B_in[0]), .B2(B_in[1]), .A(n18), .ZN(N55) );
  OAI221_X1 U6 ( .B1(B_in[1]), .B2(n21), .C1(n20), .C2(B_in[2]), .A(n19), .ZN(
        N57) );
  NAND2_X1 U8 ( .A1(B_in[2]), .A2(n21), .ZN(n19) );
endmodule


module booth_encoder_2 ( B_in, A_out );
  input [2:0] B_in;
  output [2:0] A_out;
  wire   N53, N55, N57, n18, n19, n20, n21;
  assign A_out[0] = N53;
  assign A_out[1] = N55;
  assign A_out[2] = N57;

  OAI33_X1 U9 ( .A1(B_in[0]), .A2(B_in[1]), .A3(n18), .B1(n21), .B2(n20), .B3(
        B_in[2]), .ZN(N53) );
  NAND2_X1 U4 ( .A1(B_in[2]), .A2(n21), .ZN(n19) );
  INV_X1 U3 ( .A(B_in[0]), .ZN(n21) );
  INV_X1 U5 ( .A(B_in[2]), .ZN(n18) );
  INV_X1 U6 ( .A(B_in[1]), .ZN(n20) );
  AOI21_X1 U7 ( .B1(B_in[0]), .B2(B_in[1]), .A(n18), .ZN(N55) );
  OAI221_X1 U8 ( .B1(B_in[1]), .B2(n21), .C1(n20), .C2(B_in[2]), .A(n19), .ZN(
        N57) );
endmodule


module FA_100 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n1) );
  XNOR2_X1 U1 ( .A(n1), .B(B), .ZN(S) );
endmodule


module FA_110 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n2, n3;

  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n1) );
  XNOR2_X1 U1 ( .A(Ci), .B(n1), .ZN(S) );
  OAI21_X1 U5 ( .B1(A), .B2(B), .A(Ci), .ZN(n2) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n3) );
  NAND2_X1 U3 ( .A1(n2), .A2(n3), .ZN(Co) );
endmodule


module FA_119 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(S) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Co) );
endmodule


module FA_124 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U2 ( .A(A), .B(Ci), .ZN(n1) );
  XNOR2_X1 U1 ( .A(n1), .B(B), .ZN(S) );
endmodule


module FA_126 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n2, n3;

  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n1) );
  XNOR2_X1 U1 ( .A(Ci), .B(n1), .ZN(S) );
  OAI21_X1 U5 ( .B1(A), .B2(B), .A(Ci), .ZN(n2) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n3) );
  NAND2_X1 U3 ( .A1(n2), .A2(n3), .ZN(Co) );
endmodule


module FA_0_0 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(S) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Co) );
endmodule


module RCA_N4_24 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_99 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(1'b1), .S(S[0]), .Co(CTMP[1]) );
  FA_98 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_97 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_96 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module RCA_N4_25 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_103 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(1'b0), .S(S[0]), .Co(CTMP[1]) );
  FA_102 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_101 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_100 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module RCA_N4_27 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;
  wire   n1;
  wire   [3:1] CTMP;

  FA_111 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(1'b0), .S(S[0]), .Co(n1) );
  FA_110 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(n1), .S(S[1]), .Co(CTMP[2]) );
  FA_109 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_108 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module mux21_SIZE4_14 ( IN0, IN1, CTRL, OUT1 );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] OUT1;
  input CTRL;


  MUX2_X1 U1 ( .A(IN0[3]), .B(IN1[3]), .S(CTRL), .Z(OUT1[3]) );
  MUX2_X1 U2 ( .A(IN0[2]), .B(IN1[2]), .S(CTRL), .Z(OUT1[2]) );
  MUX2_X1 U3 ( .A(IN0[1]), .B(IN1[1]), .S(CTRL), .Z(OUT1[1]) );
  MUX2_X1 U4 ( .A(IN0[0]), .B(IN1[0]), .S(CTRL), .Z(OUT1[0]) );
endmodule


module RCA_N4_29 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_119 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(1'b0), .S(S[0]), .Co(CTMP[1]) );
  FA_118 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_117 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_116 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module mux21_SIZE4_0_0 ( IN0, IN1, CTRL, OUT1 );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] OUT1;
  input CTRL;

  assign OUT1[3] = IN0[3];
  assign OUT1[2] = IN0[2];
  assign OUT1[1] = IN0[1];
  assign OUT1[0] = IN0[0];

endmodule


module RCA_N4_0_0 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_0_0 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(1'b0), .S(S[0]), .Co(CTMP[1]) );
  FA_126 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_125 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_124 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module shift_thirdLevel ( sel, A, Y );
  input [2:0] sel;
  input [38:0] A;
  output [31:0] Y;
  wire   n20, n21, n23, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n136, n137, n138, n139, n252,
         n253, n254, n255, n256, n257, n258, n259, n260;

  OAI22_X1 U138 ( .A1(A[3]), .A2(n257), .B1(A[1]), .B2(n30), .ZN(n137) );
  AOI21_X1 U137 ( .B1(n256), .B2(n38), .A(n137), .ZN(n136) );
  OAI21_X1 U136 ( .B1(A[5]), .B2(n40), .A(n136), .ZN(n98) );
  OAI22_X1 U43 ( .A1(A[30]), .A2(n30), .B1(A[34]), .B2(n40), .ZN(n66) );
  AOI21_X1 U42 ( .B1(n47), .B2(n65), .A(n66), .ZN(n64) );
  OAI21_X1 U41 ( .B1(A[36]), .B2(n255), .A(n64), .ZN(n56) );
  OAI22_X1 U34 ( .A1(A[33]), .A2(n257), .B1(A[35]), .B2(n40), .ZN(n59) );
  AOI21_X1 U33 ( .B1(n37), .B2(n58), .A(n59), .ZN(n57) );
  OAI21_X1 U32 ( .B1(A[37]), .B2(n255), .A(n57), .ZN(n54) );
  AOI22_X1 U31 ( .A1(n259), .A2(n56), .B1(n54), .B2(n260), .ZN(Y[30]) );
  OAI22_X1 U56 ( .A1(A[27]), .A2(n30), .B1(A[31]), .B2(n40), .ZN(n77) );
  AOI21_X1 U55 ( .B1(n47), .B2(n69), .A(n77), .ZN(n76) );
  OAI21_X1 U54 ( .B1(A[33]), .B2(n255), .A(n76), .ZN(n71) );
  NAND2_X1 U150 ( .A1(n139), .A2(sel[2]), .ZN(n29) );
  OAI22_X1 U52 ( .A1(A[30]), .A2(n29), .B1(A[32]), .B2(n40), .ZN(n74) );
  AOI21_X1 U51 ( .B1(n37), .B2(n73), .A(n74), .ZN(n72) );
  OAI21_X1 U50 ( .B1(A[34]), .B2(n255), .A(n72), .ZN(n67) );
  OAI22_X1 U74 ( .A1(A[25]), .A2(n257), .B1(A[27]), .B2(n40), .ZN(n90) );
  AOI21_X1 U73 ( .B1(n37), .B2(n89), .A(n90), .ZN(n88) );
  OAI21_X1 U72 ( .B1(A[29]), .B2(n255), .A(n88), .ZN(n84) );
  OAI22_X1 U69 ( .A1(A[24]), .A2(n30), .B1(A[26]), .B2(n257), .ZN(n86) );
  AOI21_X1 U68 ( .B1(n26), .B2(n73), .A(n86), .ZN(n85) );
  OAI21_X1 U67 ( .B1(A[30]), .B2(n255), .A(n85), .ZN(n81) );
  AOI22_X1 U66 ( .A1(n258), .A2(n84), .B1(n81), .B2(n260), .ZN(Y[23]) );
  OAI22_X1 U60 ( .A1(A[26]), .A2(n30), .B1(A[30]), .B2(n40), .ZN(n80) );
  AOI21_X1 U59 ( .B1(n47), .B2(n73), .A(n80), .ZN(n79) );
  OAI21_X1 U58 ( .B1(A[32]), .B2(n255), .A(n79), .ZN(n75) );
  AOI22_X1 U53 ( .A1(n258), .A2(n75), .B1(n71), .B2(n260), .ZN(Y[26]) );
  OAI22_X1 U78 ( .A1(A[24]), .A2(n29), .B1(A[26]), .B2(n40), .ZN(n94) );
  AOI21_X1 U77 ( .B1(n37), .B2(n93), .A(n94), .ZN(n92) );
  OAI21_X1 U76 ( .B1(A[28]), .B2(n255), .A(n92), .ZN(n87) );
  AOI22_X1 U71 ( .A1(n258), .A2(n87), .B1(n84), .B2(n260), .ZN(Y[22]) );
  OAI22_X1 U48 ( .A1(A[31]), .A2(n257), .B1(A[33]), .B2(n40), .ZN(n70) );
  AOI21_X1 U47 ( .B1(n37), .B2(n69), .A(n70), .ZN(n68) );
  OAI21_X1 U46 ( .B1(A[35]), .B2(n255), .A(n68), .ZN(n63) );
  AOI22_X1 U40 ( .A1(n259), .A2(n63), .B1(n56), .B2(n260), .ZN(Y[29]) );
  AOI22_X1 U45 ( .A1(n258), .A2(n67), .B1(n63), .B2(n260), .ZN(Y[28]) );
  OAI22_X1 U64 ( .A1(A[25]), .A2(n30), .B1(A[27]), .B2(n29), .ZN(n83) );
  AOI21_X1 U63 ( .B1(n26), .B2(n69), .A(n83), .ZN(n82) );
  OAI21_X1 U62 ( .B1(A[31]), .B2(n255), .A(n82), .ZN(n78) );
  AOI22_X1 U57 ( .A1(sel[0]), .A2(n78), .B1(n75), .B2(n260), .ZN(Y[25]) );
  OAI22_X1 U82 ( .A1(A[21]), .A2(n30), .B1(A[25]), .B2(n40), .ZN(n97) );
  AOI21_X1 U81 ( .B1(n47), .B2(n89), .A(n97), .ZN(n96) );
  OAI21_X1 U80 ( .B1(A[27]), .B2(n255), .A(n96), .ZN(n91) );
  AOI22_X1 U75 ( .A1(n258), .A2(n91), .B1(n87), .B2(n260), .ZN(Y[21]) );
  OAI22_X1 U91 ( .A1(A[20]), .A2(n30), .B1(A[24]), .B2(n40), .ZN(n103) );
  AOI21_X1 U90 ( .B1(n47), .B2(n93), .A(n103), .ZN(n102) );
  OAI21_X1 U89 ( .B1(A[26]), .B2(n255), .A(n102), .ZN(n95) );
  AOI22_X1 U79 ( .A1(n258), .A2(n95), .B1(n91), .B2(n260), .ZN(Y[20]) );
  AOI22_X1 U61 ( .A1(sel[0]), .A2(n81), .B1(n78), .B2(n260), .ZN(Y[24]) );
  AOI22_X1 U30 ( .A1(n47), .A2(A[34]), .B1(n37), .B2(A[32]), .ZN(n52) );
  AOI22_X1 U29 ( .A1(n256), .A2(A[38]), .B1(n26), .B2(A[36]), .ZN(n53) );
  OAI222_X1 U28 ( .A1(sel[0]), .A2(n52), .B1(sel[0]), .B2(n53), .C1(n54), .C2(
        n260), .ZN(Y[31]) );
  OAI22_X1 U95 ( .A1(A[19]), .A2(n30), .B1(A[21]), .B2(n257), .ZN(n106) );
  AOI21_X1 U94 ( .B1(n26), .B2(n89), .A(n106), .ZN(n105) );
  OAI21_X1 U93 ( .B1(A[25]), .B2(n255), .A(n105), .ZN(n101) );
  AOI22_X1 U88 ( .A1(n258), .A2(n101), .B1(n95), .B2(n260), .ZN(Y[19]) );
  OAI22_X1 U121 ( .A1(A[15]), .A2(n257), .B1(A[13]), .B2(n30), .ZN(n126) );
  AOI21_X1 U120 ( .B1(n26), .B2(n112), .A(n126), .ZN(n125) );
  OAI21_X1 U119 ( .B1(A[19]), .B2(n255), .A(n125), .ZN(n121) );
  OAI22_X1 U117 ( .A1(A[14]), .A2(n30), .B1(A[18]), .B2(n40), .ZN(n123) );
  AOI21_X1 U116 ( .B1(n47), .B2(n116), .A(n123), .ZN(n122) );
  OAI21_X1 U115 ( .B1(A[20]), .B2(n255), .A(n122), .ZN(n118) );
  AOI22_X1 U114 ( .A1(n259), .A2(n121), .B1(n118), .B2(n260), .ZN(Y[13]) );
  OAI22_X1 U113 ( .A1(A[15]), .A2(n30), .B1(A[19]), .B2(n40), .ZN(n120) );
  AOI21_X1 U112 ( .B1(n47), .B2(n112), .A(n120), .ZN(n119) );
  OAI21_X1 U111 ( .B1(A[21]), .B2(n255), .A(n119), .ZN(n114) );
  AOI22_X1 U110 ( .A1(n259), .A2(n118), .B1(n114), .B2(n260), .ZN(Y[14]) );
  OAI22_X1 U125 ( .A1(A[14]), .A2(n29), .B1(A[12]), .B2(n30), .ZN(n129) );
  AOI21_X1 U124 ( .B1(n26), .B2(n116), .A(n129), .ZN(n128) );
  OAI21_X1 U123 ( .B1(A[18]), .B2(n255), .A(n128), .ZN(n124) );
  AOI22_X1 U118 ( .A1(n259), .A2(n124), .B1(n121), .B2(n260), .ZN(Y[12]) );
  OAI22_X1 U129 ( .A1(A[13]), .A2(n257), .B1(A[11]), .B2(n30), .ZN(n131) );
  AOI21_X1 U128 ( .B1(n256), .B2(n112), .A(n131), .ZN(n130) );
  OAI21_X1 U127 ( .B1(A[15]), .B2(n40), .A(n130), .ZN(n127) );
  AOI22_X1 U122 ( .A1(n259), .A2(n127), .B1(n124), .B2(n260), .ZN(Y[11]) );
  OAI22_X1 U109 ( .A1(A[18]), .A2(n29), .B1(A[20]), .B2(n40), .ZN(n117) );
  AOI21_X1 U108 ( .B1(n37), .B2(n116), .A(n117), .ZN(n115) );
  OAI21_X1 U107 ( .B1(A[22]), .B2(n255), .A(n115), .ZN(n110) );
  AOI22_X1 U106 ( .A1(n259), .A2(n114), .B1(n110), .B2(n260), .ZN(Y[15]) );
  OAI22_X1 U15 ( .A1(A[11]), .A2(n40), .B1(A[9]), .B2(n29), .ZN(n39) );
  AOI21_X1 U14 ( .B1(n37), .B2(n38), .A(n39), .ZN(n36) );
  OAI21_X1 U13 ( .B1(A[13]), .B2(n255), .A(n36), .ZN(n31) );
  OAI22_X1 U10 ( .A1(A[10]), .A2(n29), .B1(A[8]), .B2(n30), .ZN(n34) );
  AOI21_X1 U9 ( .B1(n26), .B2(n33), .A(n34), .ZN(n32) );
  OAI21_X1 U8 ( .B1(A[14]), .B2(n255), .A(n32), .ZN(n23) );
  AOI22_X1 U7 ( .A1(n259), .A2(n31), .B1(n23), .B2(n260), .ZN(Y[7]) );
  OAI22_X1 U105 ( .A1(A[19]), .A2(n257), .B1(A[21]), .B2(n40), .ZN(n113) );
  AOI21_X1 U104 ( .B1(n37), .B2(n112), .A(n113), .ZN(n111) );
  OAI21_X1 U103 ( .B1(A[23]), .B2(n255), .A(n111), .ZN(n107) );
  OAI22_X1 U100 ( .A1(A[18]), .A2(n30), .B1(A[20]), .B2(n29), .ZN(n109) );
  AOI21_X1 U99 ( .B1(n26), .B2(n93), .A(n109), .ZN(n108) );
  OAI21_X1 U98 ( .B1(A[24]), .B2(n255), .A(n108), .ZN(n104) );
  AOI22_X1 U97 ( .A1(n259), .A2(n107), .B1(n104), .B2(n260), .ZN(Y[17]) );
  OAI22_X1 U133 ( .A1(A[12]), .A2(n29), .B1(A[10]), .B2(n30), .ZN(n133) );
  AOI21_X1 U132 ( .B1(n256), .B2(n116), .A(n133), .ZN(n132) );
  OAI21_X1 U131 ( .B1(A[14]), .B2(n40), .A(n132), .ZN(n21) );
  AOI22_X1 U126 ( .A1(n259), .A2(n21), .B1(n127), .B2(n260), .ZN(Y[10]) );
  OAI22_X1 U5 ( .A1(A[11]), .A2(n257), .B1(A[9]), .B2(n30), .ZN(n28) );
  AOI21_X1 U4 ( .B1(n26), .B2(n27), .A(n28), .ZN(n25) );
  OAI21_X1 U3 ( .B1(A[15]), .B2(n255), .A(n25), .ZN(n20) );
  AOI22_X1 U1 ( .A1(n258), .A2(n20), .B1(n21), .B2(n260), .ZN(Y[9]) );
  OAI22_X1 U39 ( .A1(A[5]), .A2(n29), .B1(A[3]), .B2(n30), .ZN(n62) );
  AOI21_X1 U38 ( .B1(n26), .B2(n38), .A(n62), .ZN(n61) );
  OAI21_X1 U37 ( .B1(A[9]), .B2(n255), .A(n61), .ZN(n49) );
  OAI22_X1 U27 ( .A1(A[4]), .A2(n30), .B1(A[8]), .B2(n40), .ZN(n51) );
  AOI21_X1 U26 ( .B1(n47), .B2(n43), .A(n51), .ZN(n50) );
  OAI21_X1 U25 ( .B1(A[10]), .B2(n255), .A(n50), .ZN(n45) );
  AOI22_X1 U24 ( .A1(sel[0]), .A2(n49), .B1(n45), .B2(n260), .ZN(Y[3]) );
  OAI22_X1 U86 ( .A1(A[2]), .A2(n30), .B1(A[4]), .B2(n29), .ZN(n100) );
  AOI21_X1 U85 ( .B1(n26), .B2(n43), .A(n100), .ZN(n99) );
  OAI21_X1 U84 ( .B1(A[8]), .B2(n255), .A(n99), .ZN(n60) );
  AOI22_X1 U83 ( .A1(n258), .A2(n98), .B1(n60), .B2(n260), .ZN(Y[1]) );
  AOI22_X1 U2 ( .A1(n259), .A2(n23), .B1(n20), .B2(n260), .ZN(Y[8]) );
  AOI22_X1 U92 ( .A1(n259), .A2(n104), .B1(n101), .B2(n260), .ZN(Y[18]) );
  AOI22_X1 U102 ( .A1(n259), .A2(n110), .B1(n107), .B2(n260), .ZN(Y[16]) );
  OAI22_X1 U23 ( .A1(A[5]), .A2(n30), .B1(A[9]), .B2(n40), .ZN(n48) );
  AOI21_X1 U22 ( .B1(n47), .B2(n38), .A(n48), .ZN(n46) );
  OAI21_X1 U21 ( .B1(A[11]), .B2(n255), .A(n46), .ZN(n41) );
  OAI22_X1 U19 ( .A1(A[10]), .A2(n40), .B1(A[8]), .B2(n257), .ZN(n44) );
  AOI21_X1 U18 ( .B1(n37), .B2(n43), .A(n44), .ZN(n42) );
  OAI21_X1 U17 ( .B1(A[12]), .B2(n255), .A(n42), .ZN(n35) );
  AOI22_X1 U16 ( .A1(sel[0]), .A2(n41), .B1(n35), .B2(n260), .ZN(Y[5]) );
  AOI22_X1 U20 ( .A1(n258), .A2(n45), .B1(n41), .B2(n260), .ZN(Y[4]) );
  AOI22_X1 U12 ( .A1(n259), .A2(n35), .B1(n31), .B2(n260), .ZN(Y[6]) );
  INV_X1 U148 ( .A(sel[2]), .ZN(n138) );
  INV_X1 U151 ( .A(sel[1]), .ZN(n139) );
  INV_X1 U142 ( .A(n40), .ZN(n26) );
  INV_X1 U149 ( .A(n257), .ZN(n47) );
  INV_X1 U139 ( .A(n37), .ZN(n30) );
  INV_X1 U35 ( .A(A[31]), .ZN(n58) );
  INV_X1 U44 ( .A(A[32]), .ZN(n65) );
  INV_X1 U101 ( .A(A[22]), .ZN(n93) );
  INV_X1 U65 ( .A(A[29]), .ZN(n69) );
  INV_X1 U96 ( .A(A[23]), .ZN(n89) );
  INV_X1 U70 ( .A(A[28]), .ZN(n73) );
  INV_X1 U6 ( .A(A[13]), .ZN(n27) );
  INV_X1 U87 ( .A(A[6]), .ZN(n43) );
  INV_X1 U130 ( .A(A[17]), .ZN(n112) );
  INV_X1 U134 ( .A(A[16]), .ZN(n116) );
  INV_X1 U11 ( .A(A[12]), .ZN(n33) );
  AOI22_X1 U36 ( .A1(A[4]), .A2(n26), .B1(A[6]), .B2(n256), .ZN(n252) );
  AOI22_X1 U49 ( .A1(A[0]), .A2(n37), .B1(A[2]), .B2(n47), .ZN(n253) );
  AND2_X1 U135 ( .A1(n252), .A2(n253), .ZN(n254) );
  OAI22_X1 U140 ( .A1(n260), .A2(n254), .B1(n259), .B2(n98), .ZN(Y[0]) );
  AOI22_X1 U141 ( .A1(n260), .A2(n49), .B1(n60), .B2(n259), .ZN(Y[2]) );
  INV_X1 U143 ( .A(A[7]), .ZN(n38) );
  AOI22_X1 U144 ( .A1(n260), .A2(n67), .B1(n71), .B2(n258), .ZN(Y[27]) );
  NAND2_X2 U145 ( .A1(n138), .A2(sel[1]), .ZN(n40) );
  CLKBUF_X1 U146 ( .A(sel[0]), .Z(n258) );
  INV_X2 U147 ( .A(sel[0]), .ZN(n260) );
  INV_X2 U152 ( .A(n256), .ZN(n255) );
  NOR2_X1 U153 ( .A1(n138), .A2(n139), .ZN(n37) );
  AND2_X1 U154 ( .A1(n138), .A2(n139), .ZN(n256) );
  BUF_X1 U155 ( .A(sel[0]), .Z(n259) );
  NAND2_X1 U156 ( .A1(n139), .A2(sel[2]), .ZN(n257) );
endmodule


module shift_secondLevel ( sel, mask00, mask08, mask16, Y );
  input [1:0] sel;
  input [38:0] mask00;
  input [38:0] mask08;
  input [38:0] mask16;
  output [38:0] Y;
  wire   n41, n42, n43, n44, n45, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n83, n136,
         n137, n138, n139, n140;

  AOI222_X1 U35 ( .A1(n139), .A2(mask00[2]), .B1(n43), .B2(mask08[2]), .C1(
        n138), .C2(mask16[2]), .ZN(n60) );
  AOI222_X1 U9 ( .A1(n139), .A2(mask00[6]), .B1(n43), .B2(mask08[6]), .C1(n138), .C2(mask16[6]), .ZN(n47) );
  AOI222_X1 U13 ( .A1(n139), .A2(mask00[4]), .B1(n43), .B2(mask08[4]), .C1(
        n138), .C2(mask16[4]), .ZN(n49) );
  AOI222_X1 U11 ( .A1(n139), .A2(mask00[5]), .B1(n43), .B2(mask08[5]), .C1(
        n138), .C2(mask16[5]), .ZN(n48) );
  AOI222_X1 U15 ( .A1(n139), .A2(mask00[3]), .B1(n43), .B2(mask08[3]), .C1(
        n138), .C2(mask16[3]), .ZN(n50) );
  AOI222_X1 U57 ( .A1(n139), .A2(mask00[1]), .B1(n140), .B2(mask08[1]), .C1(
        n138), .C2(mask16[1]), .ZN(n71) );
  AOI222_X1 U21 ( .A1(n139), .A2(mask00[36]), .B1(n43), .B2(mask08[36]), .C1(
        n138), .C2(mask16[36]), .ZN(n53) );
  AOI222_X1 U29 ( .A1(n139), .A2(mask00[32]), .B1(n43), .B2(mask08[32]), .C1(
        n138), .C2(mask16[32]), .ZN(n57) );
  AOI222_X1 U33 ( .A1(n139), .A2(mask00[30]), .B1(n43), .B2(mask08[30]), .C1(
        n138), .C2(mask16[30]), .ZN(n59) );
  AOI222_X1 U25 ( .A1(n139), .A2(mask00[34]), .B1(n43), .B2(mask08[34]), .C1(
        n138), .C2(mask16[34]), .ZN(n55) );
  AOI222_X1 U19 ( .A1(n139), .A2(mask00[37]), .B1(n43), .B2(mask08[37]), .C1(
        n138), .C2(mask16[37]), .ZN(n52) );
  AOI222_X1 U31 ( .A1(n139), .A2(mask00[31]), .B1(n43), .B2(mask08[31]), .C1(
        n138), .C2(mask16[31]), .ZN(n58) );
  AOI222_X1 U27 ( .A1(n139), .A2(mask00[33]), .B1(n43), .B2(mask08[33]), .C1(
        n138), .C2(mask16[33]), .ZN(n56) );
  AOI222_X1 U23 ( .A1(n139), .A2(mask00[35]), .B1(n43), .B2(mask08[35]), .C1(
        n138), .C2(mask16[35]), .ZN(n54) );
  AOI222_X1 U37 ( .A1(n139), .A2(mask00[29]), .B1(n43), .B2(mask08[29]), .C1(
        n138), .C2(mask16[29]), .ZN(n61) );
  AOI222_X1 U41 ( .A1(n139), .A2(mask00[27]), .B1(n43), .B2(mask08[27]), .C1(
        n138), .C2(mask16[27]), .ZN(n63) );
  AOI222_X1 U39 ( .A1(n139), .A2(mask00[28]), .B1(n43), .B2(mask08[28]), .C1(
        n138), .C2(mask16[28]), .ZN(n62) );
  AOI222_X1 U49 ( .A1(n139), .A2(mask00[23]), .B1(n43), .B2(mask08[23]), .C1(
        n138), .C2(mask16[23]), .ZN(n67) );
  AOI222_X1 U45 ( .A1(n139), .A2(mask00[25]), .B1(n140), .B2(mask08[25]), .C1(
        n138), .C2(mask16[25]), .ZN(n65) );
  AOI222_X1 U47 ( .A1(n139), .A2(mask00[24]), .B1(n43), .B2(mask08[24]), .C1(
        n138), .C2(mask16[24]), .ZN(n66) );
  AOI222_X1 U43 ( .A1(n139), .A2(mask00[26]), .B1(n43), .B2(mask08[26]), .C1(
        n138), .C2(mask16[26]), .ZN(n64) );
  AOI222_X1 U51 ( .A1(n139), .A2(mask00[22]), .B1(n43), .B2(mask08[22]), .C1(
        n138), .C2(mask16[22]), .ZN(n68) );
  AOI222_X1 U53 ( .A1(n139), .A2(mask00[21]), .B1(n43), .B2(mask08[21]), .C1(
        n138), .C2(mask16[21]), .ZN(n69) );
  AOI222_X1 U55 ( .A1(n139), .A2(mask00[20]), .B1(n43), .B2(mask08[20]), .C1(
        n138), .C2(mask16[20]), .ZN(n70) );
  AOI222_X1 U17 ( .A1(n139), .A2(mask00[38]), .B1(n140), .B2(mask08[38]), .C1(
        n138), .C2(mask16[38]), .ZN(n51) );
  AOI222_X1 U59 ( .A1(n139), .A2(mask00[19]), .B1(n140), .B2(mask08[19]), .C1(
        n138), .C2(mask16[19]), .ZN(n72) );
  AOI222_X1 U63 ( .A1(n139), .A2(mask00[17]), .B1(n140), .B2(mask08[17]), .C1(
        n138), .C2(mask16[17]), .ZN(n74) );
  AOI222_X1 U67 ( .A1(n139), .A2(mask00[15]), .B1(n140), .B2(mask08[15]), .C1(
        n138), .C2(mask16[15]), .ZN(n76) );
  AOI222_X1 U71 ( .A1(n139), .A2(mask00[13]), .B1(n140), .B2(mask08[13]), .C1(
        n138), .C2(mask16[13]), .ZN(n78) );
  AOI222_X1 U65 ( .A1(n139), .A2(mask00[16]), .B1(n140), .B2(mask08[16]), .C1(
        n138), .C2(mask16[16]), .ZN(n75) );
  AOI222_X1 U69 ( .A1(n139), .A2(mask00[14]), .B1(n140), .B2(mask08[14]), .C1(
        n138), .C2(mask16[14]), .ZN(n77) );
  AOI222_X1 U61 ( .A1(n139), .A2(mask00[18]), .B1(n140), .B2(mask08[18]), .C1(
        n138), .C2(mask16[18]), .ZN(n73) );
  AOI222_X1 U73 ( .A1(n139), .A2(mask00[12]), .B1(n140), .B2(mask08[12]), .C1(
        n138), .C2(mask16[12]), .ZN(n79) );
  AOI222_X1 U75 ( .A1(n139), .A2(mask00[11]), .B1(n140), .B2(mask08[11]), .C1(
        n138), .C2(mask16[11]), .ZN(n80) );
  AOI222_X1 U3 ( .A1(n139), .A2(mask00[9]), .B1(n43), .B2(mask08[9]), .C1(n138), .C2(mask16[9]), .ZN(n41) );
  AOI222_X1 U77 ( .A1(n139), .A2(mask00[10]), .B1(n140), .B2(mask08[10]), .C1(
        n138), .C2(mask16[10]), .ZN(n81) );
  AOI222_X1 U5 ( .A1(n139), .A2(mask00[8]), .B1(n43), .B2(mask08[8]), .C1(n138), .C2(mask16[8]), .ZN(n45) );
  INV_X1 U34 ( .A(n60), .ZN(Y[2]) );
  INV_X1 U58 ( .A(n72), .ZN(Y[19]) );
  INV_X1 U54 ( .A(n70), .ZN(Y[20]) );
  INV_X1 U52 ( .A(n69), .ZN(Y[21]) );
  INV_X1 U64 ( .A(n75), .ZN(Y[16]) );
  INV_X1 U10 ( .A(n48), .ZN(Y[5]) );
  INV_X1 U60 ( .A(n73), .ZN(Y[18]) );
  INV_X1 U68 ( .A(n77), .ZN(Y[14]) );
  INV_X1 U62 ( .A(n74), .ZN(Y[17]) );
  INV_X1 U56 ( .A(n71), .ZN(Y[1]) );
  INV_X1 U14 ( .A(n50), .ZN(Y[3]) );
  INV_X1 U70 ( .A(n78), .ZN(Y[13]) );
  INV_X1 U66 ( .A(n76), .ZN(Y[15]) );
  INV_X1 U12 ( .A(n49), .ZN(Y[4]) );
  INV_X1 U8 ( .A(n47), .ZN(Y[6]) );
  INV_X1 U22 ( .A(n54), .ZN(Y[35]) );
  INV_X1 U4 ( .A(n45), .ZN(Y[8]) );
  INV_X1 U76 ( .A(n81), .ZN(Y[10]) );
  INV_X1 U48 ( .A(n67), .ZN(Y[23]) );
  INV_X1 U26 ( .A(n56), .ZN(Y[33]) );
  INV_X1 U32 ( .A(n59), .ZN(Y[30]) );
  INV_X1 U46 ( .A(n66), .ZN(Y[24]) );
  INV_X1 U2 ( .A(n41), .ZN(Y[9]) );
  INV_X1 U42 ( .A(n64), .ZN(Y[26]) );
  INV_X1 U40 ( .A(n63), .ZN(Y[27]) );
  INV_X1 U20 ( .A(n53), .ZN(Y[36]) );
  INV_X1 U28 ( .A(n57), .ZN(Y[32]) );
  INV_X1 U74 ( .A(n80), .ZN(Y[11]) );
  INV_X1 U16 ( .A(n51), .ZN(Y[38]) );
  INV_X1 U24 ( .A(n55), .ZN(Y[34]) );
  INV_X1 U36 ( .A(n61), .ZN(Y[29]) );
  INV_X1 U44 ( .A(n65), .ZN(Y[25]) );
  INV_X1 U50 ( .A(n68), .ZN(Y[22]) );
  INV_X1 U18 ( .A(n52), .ZN(Y[37]) );
  INV_X1 U72 ( .A(n79), .ZN(Y[12]) );
  INV_X1 U38 ( .A(n62), .ZN(Y[28]) );
  INV_X1 U30 ( .A(n58), .ZN(Y[31]) );
  AOI222_X1 U6 ( .A1(mask00[0]), .A2(n139), .B1(mask16[0]), .B2(n138), .C1(
        mask08[0]), .C2(n140), .ZN(n136) );
  INV_X1 U7 ( .A(n136), .ZN(Y[0]) );
  AOI222_X1 U78 ( .A1(n43), .A2(mask08[7]), .B1(n138), .B2(mask16[7]), .C1(
        mask00[7]), .C2(n139), .ZN(n137) );
  INV_X1 U79 ( .A(n137), .ZN(Y[7]) );
  AND2_X2 U80 ( .A1(n83), .A2(sel[0]), .ZN(n43) );
  BUF_X2 U81 ( .A(n44), .Z(n138) );
  BUF_X2 U82 ( .A(n42), .Z(n139) );
  INV_X1 U83 ( .A(sel[1]), .ZN(n83) );
  BUF_X1 U84 ( .A(n43), .Z(n140) );
  NOR2_X1 U85 ( .A1(sel[0]), .A2(n83), .ZN(n44) );
  NOR2_X1 U86 ( .A1(sel[1]), .A2(sel[0]), .ZN(n42) );
endmodule


module shift_firstLevel ( A, sel, mask00, mask08, mask16 );
  input [31:0] A;
  input [1:0] sel;
  output [38:0] mask00;
  output [38:0] mask08;
  output [38:0] mask16;
  wire   n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n88, n89, n90, n91, n92, n93,
         n94, n95, n158, n159, \mask16[17] ;
  assign mask08[30] = mask16[38];
  assign mask08[29] = mask16[37];
  assign mask08[28] = mask16[36];
  assign mask08[27] = mask16[35];
  assign mask08[26] = mask16[34];
  assign mask08[25] = mask16[33];
  assign mask08[24] = mask16[32];
  assign mask08[14] = mask16[6];
  assign mask08[13] = mask16[5];
  assign mask08[12] = mask16[4];
  assign mask08[11] = mask16[3];
  assign mask08[10] = mask16[2];
  assign mask08[9] = mask16[1];
  assign mask08[8] = mask16[0];
  assign mask16[19] = \mask16[17] ;
  assign mask16[18] = \mask16[17] ;
  assign mask16[22] = \mask16[17] ;
  assign mask16[20] = \mask16[17] ;
  assign mask16[21] = \mask16[17] ;
  assign mask16[16] = \mask16[17] ;
  assign mask16[17] = \mask16[17] ;

  NAND2_X1 U155 ( .A1(sel[0]), .A2(A[10]), .ZN(n81) );
  NAND2_X1 U131 ( .A1(sel[0]), .A2(A[18]), .ZN(n53) );
  NAND2_X1 U62 ( .A1(sel[0]), .A2(A[8]), .ZN(n84) );
  NAND2_X1 U137 ( .A1(sel[0]), .A2(A[16]), .ZN(n67) );
  NAND2_X1 U143 ( .A1(sel[0]), .A2(A[14]), .ZN(n69) );
  NAND2_X1 U119 ( .A1(sel[0]), .A2(A[22]), .ZN(n39) );
  NAND2_X1 U149 ( .A1(sel[0]), .A2(A[12]), .ZN(n71) );
  NAND2_X1 U125 ( .A1(sel[0]), .A2(A[20]), .ZN(n41) );
  NAND2_X1 U146 ( .A1(sel[0]), .A2(A[13]), .ZN(n70) );
  NAND2_X1 U122 ( .A1(sel[0]), .A2(A[21]), .ZN(n40) );
  NOR2_X1 U157 ( .A1(sel[0]), .A2(sel[1]), .ZN(n85) );
  NAND2_X1 U67 ( .A1(n159), .A2(A[0]), .ZN(n60) );
  NAND2_X1 U140 ( .A1(sel[0]), .A2(A[15]), .ZN(n68) );
  NAND2_X1 U116 ( .A1(sel[0]), .A2(A[23]), .ZN(n38) );
  NAND2_X1 U152 ( .A1(sel[0]), .A2(A[11]), .ZN(n72) );
  NAND2_X1 U129 ( .A1(sel[0]), .A2(A[19]), .ZN(n42) );
  NAND2_X1 U59 ( .A1(sel[0]), .A2(A[9]), .ZN(n83) );
  NAND2_X1 U134 ( .A1(sel[0]), .A2(A[17]), .ZN(n61) );
  NAND2_X1 U91 ( .A1(sel[0]), .A2(A[31]), .ZN(n82) );
  AOI21_X1 U77 ( .B1(A[29]), .B2(n159), .A(\mask16[17] ), .ZN(n90) );
  NAND2_X1 U100 ( .A1(n159), .A2(A[21]), .ZN(n75) );
  NAND2_X1 U40 ( .A1(n75), .A2(n44), .ZN(mask08[36]) );
  NAND2_X1 U124 ( .A1(n159), .A2(A[13]), .ZN(n46) );
  NAND2_X1 U11 ( .A1(n46), .A2(n44), .ZN(mask16[36]) );
  AOI21_X1 U85 ( .B1(A[25]), .B2(n159), .A(\mask16[17] ), .ZN(n94) );
  NAND2_X1 U112 ( .A1(n159), .A2(A[17]), .ZN(n79) );
  NAND2_X1 U44 ( .A1(n79), .A2(n44), .ZN(mask08[32]) );
  NAND2_X1 U138 ( .A1(n85), .A2(A[9]), .ZN(n50) );
  NAND2_X1 U15 ( .A1(n50), .A2(n44), .ZN(mask16[32]) );
  NAND2_X1 U94 ( .A1(sel[0]), .A2(A[30]), .ZN(n62) );
  NAND2_X1 U93 ( .A1(n159), .A2(A[23]), .ZN(n73) );
  NAND2_X1 U92 ( .A1(n62), .A2(n73), .ZN(mask00[30]) );
  NAND2_X1 U118 ( .A1(n159), .A2(A[15]), .ZN(n43) );
  NAND2_X1 U9 ( .A1(n43), .A2(n44), .ZN(mask16[38]) );
  NAND2_X1 U144 ( .A1(n85), .A2(A[7]), .ZN(n52) );
  NAND2_X1 U17 ( .A1(n52), .A2(n44), .ZN(mask16[30]) );
  AOI21_X1 U81 ( .B1(A[27]), .B2(n159), .A(\mask16[17] ), .ZN(n92) );
  NAND2_X1 U106 ( .A1(n159), .A2(A[19]), .ZN(n77) );
  NAND2_X1 U42 ( .A1(n77), .A2(n44), .ZN(mask08[34]) );
  NAND2_X1 U132 ( .A1(n159), .A2(A[11]), .ZN(n48) );
  NAND2_X1 U13 ( .A1(n48), .A2(n44), .ZN(mask16[34]) );
  AOI21_X1 U75 ( .B1(A[30]), .B2(n159), .A(\mask16[17] ), .ZN(n89) );
  NAND2_X1 U97 ( .A1(n159), .A2(A[22]), .ZN(n74) );
  NAND2_X1 U39 ( .A1(n74), .A2(n44), .ZN(mask08[37]) );
  NAND2_X1 U121 ( .A1(n159), .A2(A[14]), .ZN(n45) );
  NAND2_X1 U10 ( .A1(n45), .A2(n44), .ZN(mask16[37]) );
  AOI21_X1 U89 ( .B1(A[24]), .B2(n159), .A(mask16[15]), .ZN(n95) );
  NAND2_X1 U115 ( .A1(n159), .A2(A[16]), .ZN(n80) );
  NAND2_X1 U45 ( .A1(n80), .A2(n44), .ZN(mask08[31]) );
  NAND2_X1 U141 ( .A1(n85), .A2(A[8]), .ZN(n51) );
  NAND2_X1 U16 ( .A1(n51), .A2(n44), .ZN(mask16[31]) );
  AOI21_X1 U83 ( .B1(A[26]), .B2(n159), .A(\mask16[17] ), .ZN(n93) );
  NAND2_X1 U109 ( .A1(n159), .A2(A[18]), .ZN(n78) );
  NAND2_X1 U43 ( .A1(n78), .A2(n44), .ZN(mask08[33]) );
  NAND2_X1 U135 ( .A1(n85), .A2(A[10]), .ZN(n49) );
  NAND2_X1 U14 ( .A1(n49), .A2(n44), .ZN(mask16[33]) );
  AOI21_X1 U79 ( .B1(A[28]), .B2(n159), .A(\mask16[17] ), .ZN(n91) );
  NAND2_X1 U103 ( .A1(n159), .A2(A[20]), .ZN(n76) );
  NAND2_X1 U41 ( .A1(n76), .A2(n44), .ZN(mask08[35]) );
  NAND2_X1 U128 ( .A1(n85), .A2(A[12]), .ZN(n47) );
  NAND2_X1 U12 ( .A1(n47), .A2(n44), .ZN(mask16[35]) );
  NAND2_X1 U98 ( .A1(sel[0]), .A2(A[29]), .ZN(n63) );
  NAND2_X1 U96 ( .A1(n63), .A2(n74), .ZN(mask00[29]) );
  NAND2_X1 U147 ( .A1(n159), .A2(A[6]), .ZN(n54) );
  NAND2_X1 U19 ( .A1(n54), .A2(n44), .ZN(mask16[29]) );
  NAND2_X1 U104 ( .A1(sel[0]), .A2(A[27]), .ZN(n65) );
  NAND2_X1 U102 ( .A1(n65), .A2(n76), .ZN(mask00[27]) );
  NAND2_X1 U153 ( .A1(n159), .A2(A[4]), .ZN(n56) );
  NAND2_X1 U21 ( .A1(n56), .A2(n44), .ZN(mask16[27]) );
  NAND2_X1 U101 ( .A1(sel[0]), .A2(A[28]), .ZN(n64) );
  NAND2_X1 U99 ( .A1(n64), .A2(n75), .ZN(mask00[28]) );
  NAND2_X1 U150 ( .A1(n159), .A2(A[5]), .ZN(n55) );
  NAND2_X1 U20 ( .A1(n55), .A2(n44), .ZN(mask16[28]) );
  NAND2_X1 U114 ( .A1(n38), .A2(n80), .ZN(mask00[23]) );
  NAND2_X1 U47 ( .A1(n51), .A2(n82), .ZN(mask08[23]) );
  NAND2_X1 U25 ( .A1(n44), .A2(n60), .ZN(mask16[23]) );
  NAND2_X1 U110 ( .A1(sel[0]), .A2(A[25]), .ZN(n36) );
  NAND2_X1 U108 ( .A1(n36), .A2(n78), .ZN(mask00[25]) );
  NAND2_X1 U60 ( .A1(n159), .A2(A[2]), .ZN(n58) );
  NAND2_X1 U23 ( .A1(n44), .A2(n58), .ZN(mask16[25]) );
  NAND2_X1 U113 ( .A1(sel[0]), .A2(A[24]), .ZN(n37) );
  NAND2_X1 U111 ( .A1(n37), .A2(n79), .ZN(mask00[24]) );
  NAND2_X1 U63 ( .A1(n159), .A2(A[1]), .ZN(n59) );
  NAND2_X1 U24 ( .A1(n44), .A2(n59), .ZN(mask16[24]) );
  NAND2_X1 U107 ( .A1(sel[0]), .A2(A[26]), .ZN(n66) );
  NAND2_X1 U105 ( .A1(n66), .A2(n77), .ZN(mask00[26]) );
  NAND2_X1 U156 ( .A1(n85), .A2(A[3]), .ZN(n57) );
  NAND2_X1 U22 ( .A1(n57), .A2(n44), .ZN(mask16[26]) );
  NAND2_X1 U117 ( .A1(n39), .A2(n43), .ZN(mask00[22]) );
  NAND2_X1 U48 ( .A1(n52), .A2(n62), .ZN(mask08[22]) );
  NAND2_X1 U120 ( .A1(n40), .A2(n45), .ZN(mask00[21]) );
  NAND2_X1 U49 ( .A1(n54), .A2(n63), .ZN(mask08[21]) );
  NAND2_X1 U123 ( .A1(n41), .A2(n46), .ZN(mask00[20]) );
  NAND2_X1 U50 ( .A1(n55), .A2(n64), .ZN(mask08[20]) );
  AOI21_X1 U73 ( .B1(A[31]), .B2(n159), .A(\mask16[17] ), .ZN(n88) );
  NAND2_X1 U38 ( .A1(n73), .A2(n44), .ZN(mask08[38]) );
  NAND2_X1 U127 ( .A1(n42), .A2(n47), .ZN(mask00[19]) );
  NAND2_X1 U52 ( .A1(n56), .A2(n65), .ZN(mask08[19]) );
  NAND2_X1 U133 ( .A1(n49), .A2(n61), .ZN(mask00[17]) );
  NAND2_X1 U54 ( .A1(n36), .A2(n58), .ZN(mask08[17]) );
  NAND2_X1 U139 ( .A1(n51), .A2(n68), .ZN(mask00[15]) );
  NAND2_X1 U56 ( .A1(n38), .A2(n60), .ZN(mask08[15]) );
  NAND2_X1 U145 ( .A1(n54), .A2(n70), .ZN(mask00[13]) );
  NAND2_X1 U136 ( .A1(n50), .A2(n67), .ZN(mask00[16]) );
  NAND2_X1 U55 ( .A1(n37), .A2(n59), .ZN(mask08[16]) );
  NAND2_X1 U142 ( .A1(n52), .A2(n69), .ZN(mask00[14]) );
  NAND2_X1 U130 ( .A1(n48), .A2(n53), .ZN(mask00[18]) );
  NAND2_X1 U53 ( .A1(n57), .A2(n66), .ZN(mask08[18]) );
  NAND2_X1 U148 ( .A1(n55), .A2(n71), .ZN(mask00[12]) );
  NAND2_X1 U151 ( .A1(n56), .A2(n72), .ZN(mask00[11]) );
  NAND2_X1 U58 ( .A1(n58), .A2(n83), .ZN(mask00[9]) );
  NAND2_X1 U154 ( .A1(n57), .A2(n81), .ZN(mask00[10]) );
  NAND2_X1 U61 ( .A1(n59), .A2(n84), .ZN(mask00[8]) );
  AND2_X1 U69 ( .A1(sel[0]), .A2(A[5]), .ZN(mask00[5]) );
  AND2_X1 U126 ( .A1(sel[0]), .A2(A[1]), .ZN(mask00[1]) );
  AND2_X1 U71 ( .A1(sel[0]), .A2(A[3]), .ZN(mask00[3]) );
  AND2_X1 U70 ( .A1(sel[0]), .A2(A[4]), .ZN(mask00[4]) );
  AND2_X1 U68 ( .A1(sel[0]), .A2(A[6]), .ZN(mask00[6]) );
  AND2_X1 U95 ( .A1(sel[0]), .A2(A[2]), .ZN(mask00[2]) );
  INV_X1 U51 ( .A(n83), .ZN(mask08[1]) );
  INV_X1 U31 ( .A(n66), .ZN(mask16[10]) );
  INV_X1 U3 ( .A(n37), .ZN(mask16[8]) );
  INV_X1 U26 ( .A(n61), .ZN(mask16[1]) );
  INV_X1 U30 ( .A(n65), .ZN(mask16[11]) );
  INV_X1 U18 ( .A(n53), .ZN(mask16[2]) );
  INV_X1 U6 ( .A(n40), .ZN(mask16[5]) );
  INV_X1 U46 ( .A(n81), .ZN(mask08[2]) );
  INV_X1 U35 ( .A(n70), .ZN(mask08[5]) );
  INV_X1 U90 ( .A(n82), .ZN(mask16[15]) );
  INV_X1 U2 ( .A(n36), .ZN(mask16[9]) );
  INV_X1 U28 ( .A(n63), .ZN(mask16[13]) );
  INV_X1 U29 ( .A(n64), .ZN(mask16[12]) );
  INV_X1 U37 ( .A(n72), .ZN(mask08[3]) );
  INV_X1 U34 ( .A(n69), .ZN(mask08[6]) );
  INV_X1 U5 ( .A(n39), .ZN(mask16[6]) );
  INV_X1 U8 ( .A(n42), .ZN(mask16[3]) );
  INV_X1 U27 ( .A(n62), .ZN(mask16[14]) );
  INV_X1 U36 ( .A(n71), .ZN(mask08[4]) );
  INV_X1 U32 ( .A(n67), .ZN(mask16[0]) );
  INV_X1 U7 ( .A(n41), .ZN(mask16[4]) );
  INV_X1 U88 ( .A(n95), .ZN(mask00[31]) );
  INV_X1 U74 ( .A(n89), .ZN(mask00[37]) );
  INV_X1 U78 ( .A(n91), .ZN(mask00[35]) );
  INV_X1 U76 ( .A(n90), .ZN(mask00[36]) );
  INV_X1 U72 ( .A(n88), .ZN(mask00[38]) );
  INV_X1 U82 ( .A(n93), .ZN(mask00[33]) );
  INV_X1 U80 ( .A(n92), .ZN(mask00[34]) );
  INV_X1 U84 ( .A(n94), .ZN(mask00[32]) );
  INV_X1 U4 ( .A(n84), .ZN(mask08[0]) );
  AND2_X1 U33 ( .A1(sel[0]), .A2(A[0]), .ZN(mask00[0]) );
  INV_X1 U57 ( .A(n38), .ZN(mask16[7]) );
  INV_X1 U64 ( .A(n68), .ZN(mask08[7]) );
  NAND2_X1 U65 ( .A1(sel[0]), .A2(A[7]), .ZN(n158) );
  NAND2_X1 U66 ( .A1(n60), .A2(n158), .ZN(mask00[7]) );
  NAND2_X1 U86 ( .A1(sel[1]), .A2(mask16[15]), .ZN(n44) );
  INV_X1 U87 ( .A(n44), .ZN(\mask16[17] ) );
  BUF_X1 U158 ( .A(n85), .Z(n159) );
endmodule


module mux21_1 ( IN0, IN1, CTRL, OUT1 );
  input [31:0] IN0;
  input [31:0] IN1;
  output [31:0] OUT1;
  input CTRL;
  wire   n2;

  MUX2_X1 U3 ( .A(IN0[9]), .B(IN1[9]), .S(CTRL), .Z(OUT1[9]) );
  MUX2_X1 U4 ( .A(IN0[8]), .B(IN1[8]), .S(CTRL), .Z(OUT1[8]) );
  MUX2_X1 U5 ( .A(IN0[7]), .B(IN1[7]), .S(CTRL), .Z(OUT1[7]) );
  MUX2_X1 U6 ( .A(IN0[6]), .B(IN1[6]), .S(CTRL), .Z(OUT1[6]) );
  MUX2_X1 U7 ( .A(IN0[5]), .B(IN1[5]), .S(CTRL), .Z(OUT1[5]) );
  MUX2_X1 U8 ( .A(IN0[4]), .B(IN1[4]), .S(CTRL), .Z(OUT1[4]) );
  MUX2_X1 U10 ( .A(IN0[31]), .B(IN1[31]), .S(CTRL), .Z(OUT1[31]) );
  MUX2_X1 U11 ( .A(IN0[30]), .B(IN1[30]), .S(CTRL), .Z(OUT1[30]) );
  MUX2_X1 U12 ( .A(IN0[2]), .B(IN1[2]), .S(CTRL), .Z(OUT1[2]) );
  MUX2_X1 U14 ( .A(IN0[28]), .B(IN1[28]), .S(CTRL), .Z(OUT1[28]) );
  MUX2_X1 U15 ( .A(IN0[27]), .B(IN1[27]), .S(CTRL), .Z(OUT1[27]) );
  MUX2_X1 U16 ( .A(IN0[26]), .B(IN1[26]), .S(CTRL), .Z(OUT1[26]) );
  MUX2_X1 U17 ( .A(IN0[25]), .B(IN1[25]), .S(CTRL), .Z(OUT1[25]) );
  MUX2_X1 U18 ( .A(IN0[24]), .B(IN1[24]), .S(CTRL), .Z(OUT1[24]) );
  MUX2_X1 U19 ( .A(IN0[23]), .B(IN1[23]), .S(CTRL), .Z(OUT1[23]) );
  MUX2_X1 U20 ( .A(IN0[22]), .B(IN1[22]), .S(CTRL), .Z(OUT1[22]) );
  MUX2_X1 U21 ( .A(IN0[21]), .B(IN1[21]), .S(CTRL), .Z(OUT1[21]) );
  MUX2_X1 U22 ( .A(IN0[20]), .B(IN1[20]), .S(CTRL), .Z(OUT1[20]) );
  MUX2_X1 U23 ( .A(IN0[1]), .B(IN1[1]), .S(CTRL), .Z(OUT1[1]) );
  MUX2_X1 U24 ( .A(IN0[19]), .B(IN1[19]), .S(CTRL), .Z(OUT1[19]) );
  MUX2_X1 U25 ( .A(IN0[18]), .B(IN1[18]), .S(CTRL), .Z(OUT1[18]) );
  MUX2_X1 U26 ( .A(IN0[17]), .B(IN1[17]), .S(CTRL), .Z(OUT1[17]) );
  MUX2_X1 U28 ( .A(IN0[15]), .B(IN1[15]), .S(CTRL), .Z(OUT1[15]) );
  MUX2_X1 U30 ( .A(IN0[13]), .B(IN1[13]), .S(CTRL), .Z(OUT1[13]) );
  MUX2_X1 U31 ( .A(IN0[12]), .B(IN1[12]), .S(CTRL), .Z(OUT1[12]) );
  MUX2_X1 U32 ( .A(IN0[11]), .B(IN1[11]), .S(CTRL), .Z(OUT1[11]) );
  MUX2_X1 U33 ( .A(IN0[10]), .B(IN1[10]), .S(CTRL), .Z(OUT1[10]) );
  INV_X1 U2 ( .A(IN0[0]), .ZN(n2) );
  NOR2_X1 U1 ( .A1(n2), .A2(CTRL), .ZN(OUT1[0]) );
  MUX2_X1 U9 ( .A(IN0[3]), .B(IN1[3]), .S(CTRL), .Z(OUT1[3]) );
  MUX2_X1 U13 ( .A(IN0[14]), .B(IN1[14]), .S(CTRL), .Z(OUT1[14]) );
  MUX2_X1 U27 ( .A(IN0[16]), .B(IN1[16]), .S(CTRL), .Z(OUT1[16]) );
  MUX2_X1 U29 ( .A(IN0[29]), .B(IN1[29]), .S(CTRL), .Z(OUT1[29]) );
endmodule


module piso_r_2_N32 ( Clock, ALOAD, D, SO );
  input [31:0] D;
  output [31:0] SO;
  input Clock, ALOAD;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17,
         N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31,
         N32, net645047, net645048, net645049, net645050, net645051, net645052,
         net645053, net645054, net645055, net645056, net645057, net645058,
         net645059, net645060, net645061, net645062, net645063, net645064,
         net645065, net645066, net645067, net645068, net645069, net645070,
         net645071, net645072, net645073, net645074, n1, n3, n4, n5, n6, n11,
         n12, n13, n16, n19, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30;

  DFF_X1 \tmp_reg[1]  ( .D(N4), .CK(Clock), .Q(SO[1]), .QN(net645074) );
  DFF_X1 \tmp_reg[3]  ( .D(N6), .CK(Clock), .Q(SO[3]), .QN(net645073) );
  DFF_X1 \tmp_reg[5]  ( .D(N8), .CK(Clock), .Q(SO[5]), .QN(net645072) );
  DFF_X1 \tmp_reg[7]  ( .D(N10), .CK(Clock), .Q(SO[7]), .QN(net645071) );
  DFF_X1 \tmp_reg[9]  ( .D(N12), .CK(Clock), .Q(SO[9]), .QN(net645070) );
  DFF_X1 \tmp_reg[11]  ( .D(N14), .CK(Clock), .Q(SO[11]), .QN(net645069) );
  DFF_X1 \tmp_reg[13]  ( .D(N16), .CK(Clock), .Q(SO[13]), .QN(net645068) );
  DFF_X1 \tmp_reg[15]  ( .D(N18), .CK(Clock), .Q(SO[15]), .QN(net645067) );
  DFF_X1 \tmp_reg[17]  ( .D(N20), .CK(Clock), .Q(SO[17]), .QN(net645066) );
  DFF_X1 \tmp_reg[19]  ( .D(N22), .CK(Clock), .Q(SO[19]), .QN(net645065) );
  DFF_X1 \tmp_reg[21]  ( .D(N24), .CK(Clock), .Q(SO[21]), .QN(net645064) );
  DFF_X1 \tmp_reg[23]  ( .D(N26), .CK(Clock), .Q(SO[23]), .QN(net645063) );
  DFF_X1 \tmp_reg[25]  ( .D(N28), .CK(Clock), .Q(SO[25]), .QN(net645062) );
  DFF_X1 \tmp_reg[27]  ( .D(N30), .CK(Clock), .Q(SO[27]), .QN(net645061) );
  DFF_X1 \tmp_reg[29]  ( .D(N32), .CK(Clock), .Q(SO[29]) );
  DFF_X1 \tmp_reg[0]  ( .D(N3), .CK(Clock), .Q(SO[0]), .QN(net645060) );
  DFF_X1 \tmp_reg[2]  ( .D(N5), .CK(Clock), .Q(SO[2]), .QN(net645059) );
  DFF_X1 \tmp_reg[4]  ( .D(N7), .CK(Clock), .Q(SO[4]), .QN(net645058) );
  DFF_X1 \tmp_reg[6]  ( .D(N9), .CK(Clock), .Q(SO[6]), .QN(net645057) );
  DFF_X1 \tmp_reg[8]  ( .D(N11), .CK(Clock), .Q(SO[8]), .QN(net645056) );
  DFF_X1 \tmp_reg[10]  ( .D(N13), .CK(Clock), .Q(SO[10]), .QN(net645055) );
  DFF_X1 \tmp_reg[12]  ( .D(N15), .CK(Clock), .Q(SO[12]), .QN(net645054) );
  DFF_X1 \tmp_reg[14]  ( .D(N17), .CK(Clock), .Q(SO[14]), .QN(net645053) );
  DFF_X1 \tmp_reg[16]  ( .D(N19), .CK(Clock), .Q(SO[16]), .QN(net645052) );
  DFF_X1 \tmp_reg[18]  ( .D(N21), .CK(Clock), .Q(SO[18]), .QN(net645051) );
  DFF_X1 \tmp_reg[20]  ( .D(N23), .CK(Clock), .Q(SO[20]), .QN(net645050) );
  DFF_X1 \tmp_reg[22]  ( .D(N25), .CK(Clock), .Q(SO[22]), .QN(net645049) );
  DFF_X1 \tmp_reg[24]  ( .D(N27), .CK(Clock), .Q(SO[24]), .QN(net645048) );
  DFF_X1 \tmp_reg[26]  ( .D(N29), .CK(Clock), .Q(SO[26]), .QN(net645047) );
  DFF_X1 \tmp_reg[28]  ( .D(N31), .CK(Clock), .Q(SO[28]) );
  SDFF_X1 \tmp_reg[31]  ( .D(SO[29]), .SI(D[31]), .SE(ALOAD), .CK(Clock), .Q(
        SO[31]) );
  SDFF_X1 \tmp_reg[30]  ( .D(SO[28]), .SI(D[30]), .SE(ALOAD), .CK(Clock), .Q(
        SO[30]) );
  OAI21_X1 U16 ( .B1(ALOAD), .B2(net645047), .A(n11), .ZN(N31) );
  NAND2_X1 U22 ( .A1(ALOAD), .A2(D[26]), .ZN(n11) );
  OAI21_X1 U21 ( .B1(ALOAD), .B2(net645048), .A(n11), .ZN(N29) );
  OAI21_X1 U18 ( .B1(ALOAD), .B2(net645062), .A(n12), .ZN(N30) );
  NAND2_X1 U38 ( .A1(ALOAD), .A2(D[18]), .ZN(n19) );
  OAI21_X1 U37 ( .B1(ALOAD), .B2(net645052), .A(n19), .ZN(N21) );
  OAI21_X1 U33 ( .B1(ALOAD), .B2(net645051), .A(n19), .ZN(N23) );
  NAND2_X1 U32 ( .A1(ALOAD), .A2(D[21]), .ZN(n16) );
  OAI21_X1 U31 ( .B1(ALOAD), .B2(net645065), .A(n16), .ZN(N24) );
  OAI21_X1 U39 ( .B1(ALOAD), .B2(net645067), .A(n16), .ZN(N20) );
  NAND2_X1 U42 ( .A1(ALOAD), .A2(D[16]), .ZN(n21) );
  OAI21_X1 U41 ( .B1(ALOAD), .B2(net645053), .A(n21), .ZN(N19) );
  OAI21_X1 U14 ( .B1(ALOAD), .B2(net645061), .A(n21), .ZN(N32) );
  NAND2_X1 U24 ( .A1(ALOAD), .A2(D[25]), .ZN(n12) );
  OAI21_X1 U23 ( .B1(ALOAD), .B2(net645063), .A(n12), .ZN(N28) );
  OAI21_X1 U29 ( .B1(ALOAD), .B2(net645050), .A(n13), .ZN(N25) );
  NAND2_X1 U26 ( .A1(ALOAD), .A2(D[24]), .ZN(n13) );
  OAI21_X1 U25 ( .B1(ALOAD), .B2(net645049), .A(n13), .ZN(N27) );
  OAI21_X1 U27 ( .B1(ALOAD), .B2(net645064), .A(n12), .ZN(N26) );
  OAI21_X1 U35 ( .B1(ALOAD), .B2(net645066), .A(n21), .ZN(N22) );
  NAND2_X1 U44 ( .A1(ALOAD), .A2(D[15]), .ZN(n22) );
  OAI21_X1 U43 ( .B1(ALOAD), .B2(net645068), .A(n22), .ZN(N18) );
  NAND2_X1 U52 ( .A1(ALOAD), .A2(D[11]), .ZN(n26) );
  OAI21_X1 U51 ( .B1(ALOAD), .B2(net645070), .A(n26), .ZN(N14) );
  NAND2_X1 U12 ( .A1(ALOAD), .A2(D[2]), .ZN(n6) );
  OAI21_X1 U11 ( .B1(ALOAD), .B2(net645060), .A(n6), .ZN(N5) );
  NAND2_X1 U54 ( .A1(ALOAD), .A2(D[10]), .ZN(n27) );
  OAI21_X1 U53 ( .B1(ALOAD), .B2(net645056), .A(n27), .ZN(N13) );
  NAND2_X1 U46 ( .A1(ALOAD), .A2(D[14]), .ZN(n23) );
  OAI21_X1 U45 ( .B1(ALOAD), .B2(net645054), .A(n23), .ZN(N17) );
  NAND2_X1 U50 ( .A1(ALOAD), .A2(D[12]), .ZN(n25) );
  OAI21_X1 U49 ( .B1(ALOAD), .B2(net645055), .A(n25), .ZN(N15) );
  NAND2_X1 U48 ( .A1(ALOAD), .A2(D[13]), .ZN(n24) );
  OAI21_X1 U47 ( .B1(ALOAD), .B2(net645069), .A(n24), .ZN(N16) );
  NAND2_X1 U58 ( .A1(ALOAD), .A2(D[8]), .ZN(n29) );
  OAI21_X1 U57 ( .B1(ALOAD), .B2(net645057), .A(n29), .ZN(N11) );
  NAND2_X1 U60 ( .A1(ALOAD), .A2(D[7]), .ZN(n30) );
  OAI21_X1 U59 ( .B1(ALOAD), .B2(net645072), .A(n30), .ZN(N10) );
  NAND2_X1 U56 ( .A1(ALOAD), .A2(D[9]), .ZN(n28) );
  OAI21_X1 U55 ( .B1(ALOAD), .B2(net645071), .A(n28), .ZN(N12) );
  NAND2_X1 U4 ( .A1(ALOAD), .A2(D[6]), .ZN(n1) );
  OAI21_X1 U3 ( .B1(ALOAD), .B2(net645058), .A(n1), .ZN(N9) );
  NAND2_X1 U8 ( .A1(ALOAD), .A2(D[4]), .ZN(n4) );
  OAI21_X1 U7 ( .B1(ALOAD), .B2(net645059), .A(n4), .ZN(N7) );
  NAND2_X1 U10 ( .A1(ALOAD), .A2(D[3]), .ZN(n5) );
  OAI21_X1 U9 ( .B1(ALOAD), .B2(net645074), .A(n5), .ZN(N6) );
  NAND2_X1 U6 ( .A1(ALOAD), .A2(D[5]), .ZN(n3) );
  OAI21_X1 U5 ( .B1(ALOAD), .B2(net645073), .A(n3), .ZN(N8) );
  AND2_X1 U13 ( .A1(ALOAD), .A2(D[1]), .ZN(N4) );
  AND2_X1 U15 ( .A1(ALOAD), .A2(D[0]), .ZN(N3) );
endmodule


module shift_N9_1 ( Clock, ALOAD, D, SO );
  input [8:0] D;
  input Clock, ALOAD;
  output SO;
  wire   n22;
  wire   [8:1] tmp;

  DFF_X1 \tmp_reg[8]  ( .D(n22), .CK(Clock), .Q(tmp[8]) );
  SDFF_X1 \tmp_reg[0]  ( .D(tmp[1]), .SI(D[0]), .SE(ALOAD), .CK(Clock), .Q(SO)
         );
  SDFF_X1 \tmp_reg[3]  ( .D(tmp[4]), .SI(D[3]), .SE(ALOAD), .CK(Clock), .Q(
        tmp[3]) );
  SDFF_X1 \tmp_reg[5]  ( .D(tmp[6]), .SI(D[5]), .SE(ALOAD), .CK(Clock), .Q(
        tmp[5]) );
  SDFF_X1 \tmp_reg[1]  ( .D(tmp[2]), .SI(D[1]), .SE(ALOAD), .CK(Clock), .Q(
        tmp[1]) );
  SDFF_X1 \tmp_reg[4]  ( .D(tmp[5]), .SI(D[4]), .SE(ALOAD), .CK(Clock), .Q(
        tmp[4]) );
  SDFF_X1 \tmp_reg[6]  ( .D(tmp[7]), .SI(D[6]), .SE(ALOAD), .CK(Clock), .Q(
        tmp[6]) );
  SDFF_X1 \tmp_reg[2]  ( .D(tmp[3]), .SI(D[2]), .SE(ALOAD), .CK(Clock), .Q(
        tmp[2]) );
  SDFF_X1 \tmp_reg[7]  ( .D(tmp[8]), .SI(D[7]), .SE(ALOAD), .CK(Clock), .Q(
        tmp[7]) );
  AND2_X1 U3 ( .A1(ALOAD), .A2(D[8]), .ZN(n22) );
endmodule


module shift_N9_2 ( Clock, ALOAD, D, SO );
  input [8:0] D;
  input Clock, ALOAD;
  output SO;
  wire   n22;
  wire   [8:1] tmp;

  DFF_X1 \tmp_reg[8]  ( .D(n22), .CK(Clock), .Q(tmp[8]) );
  SDFF_X1 \tmp_reg[0]  ( .D(tmp[1]), .SI(D[0]), .SE(ALOAD), .CK(Clock), .Q(SO)
         );
  SDFF_X1 \tmp_reg[2]  ( .D(tmp[3]), .SI(D[2]), .SE(ALOAD), .CK(Clock), .Q(
        tmp[2]) );
  SDFF_X1 \tmp_reg[4]  ( .D(tmp[5]), .SI(D[4]), .SE(ALOAD), .CK(Clock), .Q(
        tmp[4]) );
  SDFF_X1 \tmp_reg[3]  ( .D(tmp[4]), .SI(D[3]), .SE(ALOAD), .CK(Clock), .Q(
        tmp[3]) );
  SDFF_X1 \tmp_reg[5]  ( .D(tmp[6]), .SI(D[5]), .SE(ALOAD), .CK(Clock), .Q(
        tmp[5]) );
  SDFF_X1 \tmp_reg[7]  ( .D(tmp[8]), .SI(D[7]), .SE(ALOAD), .CK(Clock), .Q(
        tmp[7]) );
  SDFF_X1 \tmp_reg[1]  ( .D(tmp[2]), .SI(D[1]), .SE(ALOAD), .CK(Clock), .Q(
        tmp[1]) );
  SDFF_X1 \tmp_reg[6]  ( .D(tmp[7]), .SI(D[6]), .SE(ALOAD), .CK(Clock), .Q(
        tmp[6]) );
  AND2_X1 U3 ( .A1(ALOAD), .A2(D[8]), .ZN(n22) );
endmodule


module shift_N9_0 ( Clock, ALOAD, D, SO );
  input [8:0] D;
  input Clock, ALOAD;
  output SO;
  wire   n22;
  wire   [8:1] tmp;

  DFF_X1 \tmp_reg[8]  ( .D(n22), .CK(Clock), .Q(tmp[8]) );
  SDFF_X1 \tmp_reg[3]  ( .D(tmp[4]), .SI(D[3]), .SE(ALOAD), .CK(Clock), .Q(
        tmp[3]) );
  SDFF_X1 \tmp_reg[5]  ( .D(tmp[6]), .SI(D[5]), .SE(ALOAD), .CK(Clock), .Q(
        tmp[5]) );
  SDFF_X1 \tmp_reg[4]  ( .D(tmp[5]), .SI(D[4]), .SE(ALOAD), .CK(Clock), .Q(
        tmp[4]) );
  SDFF_X1 \tmp_reg[1]  ( .D(tmp[2]), .SI(D[1]), .SE(ALOAD), .CK(Clock), .Q(
        tmp[1]) );
  SDFF_X1 \tmp_reg[2]  ( .D(tmp[3]), .SI(D[2]), .SE(ALOAD), .CK(Clock), .Q(
        tmp[2]) );
  SDFF_X1 \tmp_reg[7]  ( .D(tmp[8]), .SI(D[7]), .SE(ALOAD), .CK(Clock), .Q(
        tmp[7]) );
  SDFF_X1 \tmp_reg[6]  ( .D(tmp[7]), .SI(D[6]), .SE(ALOAD), .CK(Clock), .Q(
        tmp[6]) );
  SDFF_X2 \tmp_reg[0]  ( .D(tmp[1]), .SI(D[0]), .SE(ALOAD), .CK(Clock), .Q(SO)
         );
  AND2_X1 U3 ( .A1(ALOAD), .A2(D[8]), .ZN(n22) );
endmodule


module booth_encoder_1 ( B_in, A_out );
  input [2:0] B_in;
  output [2:0] A_out;
  wire   N53, N55, N57, n3, n4, n5;
  assign A_out[0] = N53;
  assign A_out[1] = N55;
  assign A_out[2] = N57;

  NAND2_X1 U7 ( .A1(B_in[1]), .A2(n3), .ZN(n5) );
  OAI221_X1 U3 ( .B1(B_in[0]), .B2(n3), .C1(n4), .C2(B_in[1]), .A(n5), .ZN(N57) );
  NOR2_X1 U5 ( .A1(n5), .A2(n4), .ZN(N53) );
  INV_X1 U8 ( .A(B_in[2]), .ZN(n3) );
  AND2_X1 U4 ( .A1(n4), .A2(B_in[1]), .ZN(N55) );
  INV_X1 U6 ( .A(B_in[0]), .ZN(n4) );
endmodule


module booth_encoder_6 ( B_in, A_out );
  input [2:0] B_in;
  output [2:0] A_out;
  wire   N53, N55, N57, n4, n5, n6, n7;
  assign A_out[0] = N53;
  assign A_out[1] = N55;
  assign A_out[2] = N57;

  OAI33_X1 U9 ( .A1(B_in[0]), .A2(B_in[1]), .A3(n7), .B1(n4), .B2(n5), .B3(
        B_in[2]), .ZN(N53) );
  INV_X1 U3 ( .A(B_in[1]), .ZN(n5) );
  INV_X1 U4 ( .A(B_in[0]), .ZN(n4) );
  INV_X1 U5 ( .A(B_in[2]), .ZN(n7) );
  NAND2_X1 U6 ( .A1(B_in[2]), .A2(n4), .ZN(n6) );
  OAI221_X1 U7 ( .B1(B_in[1]), .B2(n4), .C1(n5), .C2(B_in[2]), .A(n6), .ZN(N57) );
  AOI21_X1 U8 ( .B1(B_in[0]), .B2(B_in[1]), .A(n7), .ZN(N55) );
endmodule


module booth_encoder_7 ( B_in, A_out );
  input [2:0] B_in;
  output [2:0] A_out;
  wire   N53, N55, N57, n4, n5, n6, n7;
  assign A_out[0] = N53;
  assign A_out[1] = N55;
  assign A_out[2] = N57;

  OAI33_X1 U9 ( .A1(B_in[0]), .A2(B_in[1]), .A3(n7), .B1(n4), .B2(n5), .B3(
        B_in[2]), .ZN(N53) );
  INV_X1 U3 ( .A(B_in[1]), .ZN(n5) );
  INV_X1 U4 ( .A(B_in[0]), .ZN(n4) );
  INV_X1 U5 ( .A(B_in[2]), .ZN(n7) );
  AOI21_X1 U6 ( .B1(B_in[0]), .B2(B_in[1]), .A(n7), .ZN(N55) );
  OAI221_X1 U7 ( .B1(B_in[1]), .B2(n4), .C1(n5), .C2(B_in[2]), .A(n6), .ZN(N57) );
  NAND2_X1 U8 ( .A1(B_in[2]), .A2(n4), .ZN(n6) );
endmodule


module booth_encoder_8 ( B_in, A_out );
  input [2:0] B_in;
  output [2:0] A_out;
  wire   N53, N55, N57, n4, n5, n6, n7;
  assign A_out[0] = N53;
  assign A_out[1] = N55;
  assign A_out[2] = N57;

  OAI33_X1 U9 ( .A1(B_in[0]), .A2(B_in[1]), .A3(n7), .B1(n4), .B2(n5), .B3(
        B_in[2]), .ZN(N53) );
  INV_X1 U3 ( .A(B_in[2]), .ZN(n7) );
  INV_X1 U4 ( .A(B_in[1]), .ZN(n5) );
  INV_X1 U5 ( .A(B_in[0]), .ZN(n4) );
  AOI21_X1 U6 ( .B1(B_in[0]), .B2(B_in[1]), .A(n7), .ZN(N55) );
  NAND2_X1 U7 ( .A1(B_in[2]), .A2(n4), .ZN(n6) );
  OAI221_X1 U8 ( .B1(B_in[1]), .B2(n4), .C1(n5), .C2(B_in[2]), .A(n6), .ZN(N57) );
endmodule


module booth_encoder_0 ( B_in, A_out );
  input [2:0] B_in;
  output [2:0] A_out;
  wire   N53, N57, n2;
  assign A_out[1] = B_in[2];
  assign A_out[0] = N53;
  assign A_out[2] = N57;

  INV_X1 U3 ( .A(B_in[2]), .ZN(n2) );
  OR2_X1 U4 ( .A1(B_in[1]), .A2(B_in[2]), .ZN(N57) );
  NOR2_X1 U5 ( .A1(B_in[1]), .A2(n2), .ZN(N53) );
endmodule


module carry_sel_gen_N4_11 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:0] nocarry_sum_to_mux;
  wire   [3:0] carry_sum_to_mux;

  RCA_N4_23 rca_nocarry ( .A(A), .B(B), .Ci(1'b0), .S(nocarry_sum_to_mux) );
  RCA_N4_22 rca_carry ( .A(A), .B(B), .Ci(1'b1), .S(carry_sum_to_mux) );
  mux21_SIZE4_11 outmux ( .IN0(nocarry_sum_to_mux), .IN1(carry_sum_to_mux), 
        .CTRL(Ci), .OUT1(S) );
endmodule


module carry_sel_gen_N4_12 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:0] nocarry_sum_to_mux;
  wire   [3:0] carry_sum_to_mux;

  RCA_N4_25 rca_nocarry ( .A(A), .B(B), .Ci(1'b0), .S(nocarry_sum_to_mux) );
  RCA_N4_24 rca_carry ( .A(A), .B(B), .Ci(1'b1), .S(carry_sum_to_mux) );
  mux21_SIZE4_12 outmux ( .IN0(nocarry_sum_to_mux), .IN1(carry_sum_to_mux), 
        .CTRL(Ci), .OUT1(S) );
endmodule


module carry_sel_gen_N4_13 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:0] nocarry_sum_to_mux;
  wire   [3:0] carry_sum_to_mux;

  RCA_N4_27 rca_nocarry ( .A(A), .B(B), .Ci(1'b0), .S(nocarry_sum_to_mux) );
  RCA_N4_26 rca_carry ( .A(A), .B(B), .Ci(1'b1), .S(carry_sum_to_mux) );
  mux21_SIZE4_13 outmux ( .IN0(nocarry_sum_to_mux), .IN1(carry_sum_to_mux), 
        .CTRL(Ci), .OUT1(S) );
endmodule


module carry_sel_gen_N4_14 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:0] nocarry_sum_to_mux;
  wire   [3:0] carry_sum_to_mux;

  RCA_N4_29 rca_nocarry ( .A(A), .B(B), .Ci(1'b0), .S(nocarry_sum_to_mux) );
  RCA_N4_28 rca_carry ( .A(A), .B(B), .Ci(1'b1), .S(carry_sum_to_mux) );
  mux21_SIZE4_14 outmux ( .IN0(nocarry_sum_to_mux), .IN1(carry_sum_to_mux), 
        .CTRL(Ci), .OUT1(S) );
endmodule


module carry_sel_gen_N4_0_0 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:0] nocarry_sum_to_mux;

  RCA_N4_0_0 rca_nocarry ( .A(A), .B(B), .Ci(1'b0), .S(nocarry_sum_to_mux) );
  mux21_SIZE4_0_0 outmux ( .IN0(nocarry_sum_to_mux), .IN1({1'b0, 1'b0, 1'b0, 
        1'b0}), .CTRL(1'b0), .OUT1(S) );
endmodule


module pg_37 ( p, g_prec, p_prec, g_out, p_out, g_BAR );
  input p, g_prec, p_prec, g_BAR;
  output g_out, p_out;
  wire   g, n1;
  assign g = g_BAR;

  NAND2_X1 U3 ( .A1(p), .A2(g_prec), .ZN(n1) );
  NAND2_X1 U2 ( .A1(g), .A2(n1), .ZN(g_out) );
  AND2_X1 U1 ( .A1(p), .A2(p_prec), .ZN(p_out) );
endmodule


module pg_38 ( p, g_prec, p_prec, g_out, p_out, g_BAR );
  input p, g_prec, p_prec, g_BAR;
  output g_out, p_out;
  wire   g, n1;
  assign g = g_BAR;

  NAND2_X1 U3 ( .A1(p), .A2(g_prec), .ZN(n1) );
  NAND2_X1 U2 ( .A1(g), .A2(n1), .ZN(g_out) );
  AND2_X1 U1 ( .A1(p), .A2(p_prec), .ZN(p_out) );
endmodule


module g_17 ( g, p, g_prec, g_out );
  input g, p, g_prec;
  output g_out;
  wire   n2;

  AOI21_X1 U2 ( .B1(p), .B2(g_prec), .A(g), .ZN(n2) );
  INV_X1 U1 ( .A(n2), .ZN(g_out) );
endmodule


module pg_46 ( g, p, g_prec, p_prec, g_out, p_out );
  input g, p, g_prec, p_prec;
  output g_out, p_out;
  wire   n6, n7;

  INV_X1 U1 ( .A(g), .ZN(n7) );
  AND2_X1 U2 ( .A1(p), .A2(p_prec), .ZN(p_out) );
  NAND2_X1 U3 ( .A1(p), .A2(g_prec), .ZN(n6) );
  NAND2_X1 U4 ( .A1(n6), .A2(n7), .ZN(g_out) );
endmodule


module pg_51 ( g, p, g_prec, p_prec, p_out, g_out_BAR );
  input g, p, g_prec, p_prec;
  output p_out, g_out_BAR;


  AOI21_X1 U2 ( .B1(g_prec), .B2(p), .A(g), .ZN(g_out_BAR) );
  AND2_X1 U1 ( .A1(p), .A2(p_prec), .ZN(p_out) );
endmodule


module pg_52 ( g, p, g_prec, p_prec, g_out, p_out );
  input g, p, g_prec, p_prec;
  output g_out, p_out;
  wire   n2;

  AOI21_X1 U3 ( .B1(g_prec), .B2(p), .A(g), .ZN(n2) );
  AND2_X1 U1 ( .A1(p), .A2(p_prec), .ZN(p_out) );
  INV_X1 U2 ( .A(n2), .ZN(g_out) );
endmodule


module pg_0_0 ( g, p, g_prec, p_prec, g_out, p_out );
  input g, p, g_prec, p_prec;
  output g_out, p_out;
  wire   n2;

  AOI21_X1 U3 ( .B1(g_prec), .B2(p), .A(g), .ZN(n2) );
  AND2_X1 U1 ( .A1(p), .A2(p_prec), .ZN(p_out) );
  INV_X1 U2 ( .A(n2), .ZN(g_out) );
endmodule


module g_18 ( g, p, g_prec, g_out );
  input g, p, g_prec;
  output g_out;
  wire   n2;

  AOI21_X1 U2 ( .B1(p), .B2(g_prec), .A(g), .ZN(n2) );
  INV_X1 U1 ( .A(n2), .ZN(g_out) );
endmodule


module g_0_0 ( g, p, g_prec, g_out );
  input g, p, g_prec;
  output g_out;
  wire   g;
  assign g_out = g;

endmodule


module pg_net_49 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p_out) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g_out) );
endmodule


module pg_net_62 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p_out) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g_out) );
endmodule


module pg_net_0_0 ( a, b, g_out, p_out );
  input a, b;
  output g_out, p_out;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p_out) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g_out) );
endmodule


module logic_unit_SIZE32 ( IN1, IN2, CTRL, OUT1 );
  input [31:0] IN1;
  input [31:0] IN2;
  input [1:0] CTRL;
  output [31:0] OUT1;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n22, n23, n24, n25, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n268, n269, n270, n271, n272, n273;

  XOR2_X1 U98 ( .A(n273), .B(CTRL[0]), .Z(n3) );
  OAI21_X1 U95 ( .B1(n273), .B2(n64), .A(n65), .ZN(OUT1[0]) );
  NAND2_X1 U28 ( .A1(IN2[30]), .A2(IN1[30]), .ZN(n18) );
  OAI211_X1 U27 ( .C1(IN2[30]), .C2(IN1[30]), .A(n272), .B(n18), .ZN(n19) );
  OAI21_X1 U26 ( .B1(CTRL[1]), .B2(n18), .A(n19), .ZN(OUT1[30]) );
  NAND2_X1 U52 ( .A1(IN2[23]), .A2(IN1[23]), .ZN(n34) );
  OAI211_X1 U51 ( .C1(IN2[23]), .C2(IN1[23]), .A(n272), .B(n34), .ZN(n35) );
  OAI21_X1 U50 ( .B1(CTRL[1]), .B2(n34), .A(n35), .ZN(OUT1[23]) );
  NAND2_X1 U43 ( .A1(IN2[26]), .A2(IN1[26]), .ZN(n28) );
  OAI211_X1 U42 ( .C1(IN2[26]), .C2(IN1[26]), .A(n272), .B(n28), .ZN(n29) );
  OAI21_X1 U41 ( .B1(CTRL[1]), .B2(n28), .A(n29), .ZN(OUT1[26]) );
  NAND2_X1 U55 ( .A1(IN2[22]), .A2(IN1[22]), .ZN(n36) );
  OAI211_X1 U54 ( .C1(IN2[22]), .C2(IN1[22]), .A(n272), .B(n36), .ZN(n37) );
  OAI21_X1 U53 ( .B1(CTRL[1]), .B2(n36), .A(n37), .ZN(OUT1[22]) );
  NAND2_X1 U34 ( .A1(IN2[29]), .A2(IN1[29]), .ZN(n22) );
  OAI211_X1 U33 ( .C1(IN2[29]), .C2(IN1[29]), .A(n272), .B(n22), .ZN(n23) );
  OAI21_X1 U32 ( .B1(n273), .B2(n22), .A(n23), .ZN(OUT1[29]) );
  NAND2_X1 U37 ( .A1(IN2[28]), .A2(IN1[28]), .ZN(n24) );
  OAI211_X1 U36 ( .C1(IN2[28]), .C2(IN1[28]), .A(n272), .B(n24), .ZN(n25) );
  OAI21_X1 U35 ( .B1(n273), .B2(n24), .A(n25), .ZN(OUT1[28]) );
  NAND2_X1 U46 ( .A1(IN2[25]), .A2(IN1[25]), .ZN(n30) );
  OAI211_X1 U45 ( .C1(IN2[25]), .C2(IN1[25]), .A(n272), .B(n30), .ZN(n31) );
  OAI21_X1 U44 ( .B1(CTRL[1]), .B2(n30), .A(n31), .ZN(OUT1[25]) );
  NAND2_X1 U58 ( .A1(IN2[21]), .A2(IN1[21]), .ZN(n38) );
  OAI211_X1 U57 ( .C1(IN2[21]), .C2(IN1[21]), .A(n272), .B(n38), .ZN(n39) );
  OAI21_X1 U56 ( .B1(n273), .B2(n38), .A(n39), .ZN(OUT1[21]) );
  NAND2_X1 U61 ( .A1(IN2[20]), .A2(IN1[20]), .ZN(n40) );
  OAI211_X1 U60 ( .C1(IN2[20]), .C2(IN1[20]), .A(n272), .B(n40), .ZN(n41) );
  OAI21_X1 U59 ( .B1(n273), .B2(n40), .A(n41), .ZN(OUT1[20]) );
  NAND2_X1 U49 ( .A1(IN2[24]), .A2(IN1[24]), .ZN(n32) );
  OAI211_X1 U48 ( .C1(IN2[24]), .C2(IN1[24]), .A(n272), .B(n32), .ZN(n33) );
  OAI21_X1 U47 ( .B1(n273), .B2(n32), .A(n33), .ZN(OUT1[24]) );
  NAND2_X1 U25 ( .A1(IN2[31]), .A2(IN1[31]), .ZN(n16) );
  OAI211_X1 U24 ( .C1(IN2[31]), .C2(IN1[31]), .A(n272), .B(n16), .ZN(n17) );
  OAI21_X1 U23 ( .B1(n273), .B2(n16), .A(n17), .ZN(OUT1[31]) );
  NAND2_X1 U67 ( .A1(IN2[19]), .A2(IN1[19]), .ZN(n44) );
  OAI211_X1 U66 ( .C1(IN2[19]), .C2(IN1[19]), .A(n272), .B(n44), .ZN(n45) );
  OAI21_X1 U65 ( .B1(n273), .B2(n44), .A(n45), .ZN(OUT1[19]) );
  OAI21_X1 U83 ( .B1(CTRL[1]), .B2(n56), .A(n57), .ZN(OUT1[13]) );
  OAI21_X1 U80 ( .B1(CTRL[1]), .B2(n54), .A(n55), .ZN(OUT1[14]) );
  OAI21_X1 U86 ( .B1(CTRL[1]), .B2(n58), .A(n59), .ZN(OUT1[12]) );
  NAND2_X1 U91 ( .A1(IN2[11]), .A2(IN1[11]), .ZN(n60) );
  OAI211_X1 U90 ( .C1(IN2[11]), .C2(IN1[11]), .A(n272), .B(n60), .ZN(n61) );
  OAI21_X1 U89 ( .B1(n273), .B2(n60), .A(n61), .ZN(OUT1[11]) );
  NAND2_X1 U79 ( .A1(IN2[15]), .A2(IN1[15]), .ZN(n52) );
  OAI211_X1 U78 ( .C1(IN2[15]), .C2(IN1[15]), .A(n272), .B(n52), .ZN(n53) );
  OAI21_X1 U77 ( .B1(CTRL[1]), .B2(n52), .A(n53), .ZN(OUT1[15]) );
  OAI21_X1 U8 ( .B1(n273), .B2(n6), .A(n7), .ZN(OUT1[7]) );
  OAI21_X1 U71 ( .B1(CTRL[1]), .B2(n48), .A(n49), .ZN(OUT1[17]) );
  OAI21_X1 U92 ( .B1(CTRL[1]), .B2(n62), .A(n63), .ZN(OUT1[10]) );
  OAI21_X1 U2 ( .B1(n273), .B2(n1), .A(n2), .ZN(OUT1[9]) );
  OAI21_X1 U20 ( .B1(n273), .B2(n14), .A(n15), .ZN(OUT1[3]) );
  OAI21_X1 U62 ( .B1(CTRL[1]), .B2(n42), .A(n43), .ZN(OUT1[1]) );
  NAND2_X1 U7 ( .A1(IN2[8]), .A2(IN1[8]), .ZN(n4) );
  OAI211_X1 U6 ( .C1(IN2[8]), .C2(IN1[8]), .A(n3), .B(n4), .ZN(n5) );
  OAI21_X1 U5 ( .B1(n273), .B2(n4), .A(n5), .ZN(OUT1[8]) );
  NAND2_X1 U70 ( .A1(IN2[18]), .A2(IN1[18]), .ZN(n46) );
  OAI211_X1 U69 ( .C1(IN2[18]), .C2(IN1[18]), .A(n272), .B(n46), .ZN(n47) );
  OAI21_X1 U68 ( .B1(n273), .B2(n46), .A(n47), .ZN(OUT1[18]) );
  NAND2_X1 U76 ( .A1(IN2[16]), .A2(IN1[16]), .ZN(n50) );
  OAI211_X1 U75 ( .C1(IN2[16]), .C2(IN1[16]), .A(n272), .B(n50), .ZN(n51) );
  OAI21_X1 U74 ( .B1(CTRL[1]), .B2(n50), .A(n51), .ZN(OUT1[16]) );
  OAI21_X1 U14 ( .B1(n273), .B2(n10), .A(n11), .ZN(OUT1[5]) );
  OAI21_X1 U17 ( .B1(n273), .B2(n12), .A(n13), .ZN(OUT1[4]) );
  OAI21_X1 U11 ( .B1(n273), .B2(n8), .A(n9), .ZN(OUT1[6]) );
  NAND2_X1 U3 ( .A1(IN2[2]), .A2(IN1[2]), .ZN(n268) );
  OAI211_X1 U4 ( .C1(IN2[2]), .C2(IN1[2]), .A(n272), .B(n268), .ZN(n269) );
  OAI21_X1 U9 ( .B1(CTRL[1]), .B2(n268), .A(n269), .ZN(OUT1[2]) );
  NAND2_X1 U10 ( .A1(IN2[27]), .A2(IN1[27]), .ZN(n270) );
  OAI211_X1 U12 ( .C1(IN2[27]), .C2(IN1[27]), .A(n272), .B(n270), .ZN(n271) );
  OAI21_X1 U13 ( .B1(CTRL[1]), .B2(n270), .A(n271), .ZN(OUT1[27]) );
  BUF_X2 U15 ( .A(n3), .Z(n272) );
  BUF_X1 U16 ( .A(CTRL[1]), .Z(n273) );
  OAI211_X1 U18 ( .C1(IN2[10]), .C2(IN1[10]), .A(n272), .B(n62), .ZN(n63) );
  NAND2_X1 U19 ( .A1(IN2[10]), .A2(IN1[10]), .ZN(n62) );
  OAI211_X1 U21 ( .C1(IN2[12]), .C2(IN1[12]), .A(n272), .B(n58), .ZN(n59) );
  NAND2_X1 U22 ( .A1(IN2[12]), .A2(IN1[12]), .ZN(n58) );
  OAI211_X1 U29 ( .C1(IN2[4]), .C2(IN1[4]), .A(n272), .B(n12), .ZN(n13) );
  NAND2_X1 U30 ( .A1(IN2[4]), .A2(IN1[4]), .ZN(n12) );
  OAI211_X1 U31 ( .C1(IN2[17]), .C2(IN1[17]), .A(n272), .B(n48), .ZN(n49) );
  NAND2_X1 U38 ( .A1(IN2[17]), .A2(IN1[17]), .ZN(n48) );
  OAI211_X1 U39 ( .C1(IN2[1]), .C2(IN1[1]), .A(n272), .B(n42), .ZN(n43) );
  NAND2_X1 U40 ( .A1(IN2[1]), .A2(IN1[1]), .ZN(n42) );
  OAI211_X1 U63 ( .C1(IN2[13]), .C2(IN1[13]), .A(n272), .B(n56), .ZN(n57) );
  NAND2_X1 U64 ( .A1(IN2[13]), .A2(IN1[13]), .ZN(n56) );
  OAI211_X1 U72 ( .C1(IN2[7]), .C2(IN1[7]), .A(n272), .B(n6), .ZN(n7) );
  NAND2_X1 U73 ( .A1(IN2[7]), .A2(IN1[7]), .ZN(n6) );
  OAI211_X1 U81 ( .C1(IN2[3]), .C2(IN1[3]), .A(n272), .B(n14), .ZN(n15) );
  NAND2_X1 U82 ( .A1(IN2[3]), .A2(IN1[3]), .ZN(n14) );
  OAI211_X1 U84 ( .C1(IN2[14]), .C2(IN1[14]), .A(n272), .B(n54), .ZN(n55) );
  NAND2_X1 U85 ( .A1(IN2[14]), .A2(IN1[14]), .ZN(n54) );
  OAI211_X1 U87 ( .C1(IN2[6]), .C2(IN1[6]), .A(n3), .B(n8), .ZN(n9) );
  NAND2_X1 U88 ( .A1(IN2[6]), .A2(IN1[6]), .ZN(n8) );
  OAI211_X1 U93 ( .C1(IN2[0]), .C2(IN1[0]), .A(n272), .B(n64), .ZN(n65) );
  NAND2_X1 U94 ( .A1(IN2[0]), .A2(IN1[0]), .ZN(n64) );
  OAI211_X1 U96 ( .C1(IN2[9]), .C2(IN1[9]), .A(n272), .B(n1), .ZN(n2) );
  NAND2_X1 U97 ( .A1(IN2[9]), .A2(IN1[9]), .ZN(n1) );
  OAI211_X1 U99 ( .C1(IN2[5]), .C2(IN1[5]), .A(n3), .B(n10), .ZN(n11) );
  NAND2_X1 U100 ( .A1(IN2[5]), .A2(IN1[5]), .ZN(n10) );
endmodule


module shifter ( A, B, LOGIC_ARITH, LEFT_RIGHT, OUTPUT );
  input [31:0] A;
  input [4:0] B;
  output [31:0] OUTPUT;
  input LOGIC_ARITH, LEFT_RIGHT;
  wire   n2, n3, n4, n6, n10, n11, n12, n9, n14, n15, n16, n17;
  wire   [2:0] s3;
  wire   [38:0] m0;
  wire   [38:0] m8;
  wire   [38:0] m16;
  wire   [38:0] y;

  shift_firstLevel IL ( .A(A), .sel({LOGIC_ARITH, LEFT_RIGHT}), .mask00(m0), 
        .mask08(m8), .mask16({m16[38:23], n3, n11, n6, n2, n12, n4, n10, 
        m16[15:0]}) );
  shift_secondLevel IIL ( .sel(B[4:3]), .mask00(m0), .mask08(m8), .mask16({
        m16[38:23], n3, n11, n6, n2, n12, n4, n10, m16[15:0]}), .Y(y) );
  shift_thirdLevel IIIL ( .sel(s3), .A(y), .Y(OUTPUT) );
  OR2_X1 U8 ( .A1(LOGIC_ARITH), .A2(LEFT_RIGHT), .ZN(n9) );
  INV_X1 U1 ( .A(LEFT_RIGHT), .ZN(n17) );
  INV_X1 U2 ( .A(B[0]), .ZN(n16) );
  INV_X1 U3 ( .A(B[2]), .ZN(n14) );
  INV_X1 U4 ( .A(B[1]), .ZN(n15) );
  AOI22_X1 U5 ( .A1(B[0]), .A2(n9), .B1(n17), .B2(n16), .ZN(s3[0]) );
  AOI22_X1 U6 ( .A1(B[2]), .A2(n9), .B1(n17), .B2(n14), .ZN(s3[2]) );
  AOI22_X1 U7 ( .A1(B[1]), .A2(n9), .B1(n17), .B2(n15), .ZN(s3[1]) );
endmodule


module comparator_M32 ( C, V, SUM, sel, sign, S );
  input [31:0] SUM;
  input [2:0] sel;
  input C, V, sign;
  output S;
  wire   n6, n24, n23, n22, n21, n20, n19, n18, n17, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83;

  NOR4_X1 U14 ( .A1(SUM[9]), .A2(SUM[8]), .A3(SUM[7]), .A4(SUM[6]), .ZN(n18)
         );
  NOR4_X1 U17 ( .A1(SUM[16]), .A2(SUM[15]), .A3(SUM[14]), .A4(SUM[13]), .ZN(
        n24) );
  NOR4_X1 U18 ( .A1(SUM[12]), .A2(SUM[11]), .A3(SUM[10]), .A4(SUM[0]), .ZN(n23) );
  NOR4_X1 U20 ( .A1(SUM[1]), .A2(SUM[19]), .A3(SUM[18]), .A4(SUM[17]), .ZN(n21) );
  XNOR2_X1 U1 ( .A(n83), .B(V), .ZN(n66) );
  MUX2_X1 U2 ( .A(C), .B(n66), .S(sign), .Z(n6) );
  INV_X1 U3 ( .A(sel[0]), .ZN(n77) );
  INV_X1 U4 ( .A(sel[1]), .ZN(n80) );
  INV_X1 U5 ( .A(sel[2]), .ZN(n79) );
  AND3_X1 U6 ( .A1(n21), .A2(n68), .A3(n22), .ZN(n69) );
  AND2_X1 U7 ( .A1(n24), .A2(n23), .ZN(n68) );
  CLKBUF_X1 U8 ( .A(SUM[31]), .Z(n83) );
  AND2_X1 U9 ( .A1(n67), .A2(n69), .ZN(n71) );
  AND2_X1 U10 ( .A1(n67), .A2(n69), .ZN(n70) );
  AND4_X1 U11 ( .A1(n17), .A2(n18), .A3(n19), .A4(n20), .ZN(n67) );
  NOR2_X1 U12 ( .A1(sel[0]), .A2(sel[1]), .ZN(n76) );
  NAND2_X1 U13 ( .A1(n79), .A2(n80), .ZN(n78) );
  AOI21_X1 U15 ( .B1(n71), .B2(n77), .A(n78), .ZN(n74) );
  XNOR2_X1 U16 ( .A(n70), .B(n76), .ZN(n75) );
  NAND2_X1 U19 ( .A1(n71), .A2(sel[0]), .ZN(n82) );
  NAND2_X1 U21 ( .A1(n73), .A2(n72), .ZN(S) );
  NOR4_X1 U22 ( .A1(SUM[23]), .A2(SUM[22]), .A3(SUM[21]), .A4(SUM[20]), .ZN(
        n22) );
  NOR4_X1 U23 ( .A1(SUM[30]), .A2(SUM[28]), .A3(SUM[29]), .A4(SUM[2]), .ZN(n20) );
  NOR4_X1 U24 ( .A1(SUM[27]), .A2(SUM[26]), .A3(SUM[25]), .A4(SUM[24]), .ZN(
        n19) );
  NOR4_X1 U25 ( .A1(SUM[31]), .A2(SUM[5]), .A3(SUM[3]), .A4(SUM[4]), .ZN(n17)
         );
  NAND3_X1 U26 ( .A1(n81), .A2(n79), .A3(sel[1]), .ZN(n72) );
  NAND2_X1 U27 ( .A1(n6), .A2(n82), .ZN(n81) );
  AOI22_X1 U28 ( .A1(n6), .A2(n74), .B1(n75), .B2(sel[2]), .ZN(n73) );
endmodule


module simple_booth_add_ext_N16 ( Clock, Reset, sign, enable, valid, A, B, 
        A_to_add, B_to_add, sign_to_add, final_out, ACC_from_add );
  input [15:0] A;
  input [15:0] B;
  output [31:0] A_to_add;
  output [31:0] B_to_add;
  output [31:0] final_out;
  input [31:0] ACC_from_add;
  input Clock, Reset, sign, enable;
  output valid, sign_to_add;
  wire   \enc_N2_in[2] , \extend_vector[15] , \input_mux_sel[2] ,
         input_mux_sel_0, reg_enable, n50, n51, n52, n54, n22, n37, n40,
         net645046, n49, n53, n55, n56, n57, n58, n59, n60, n61, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n90, n91, n92, n93, n41, n42,
         n46, n47, n48, n62, n78;
  wire   [8:0] piso_0_in;
  wire   [8:0] piso_1_in;
  wire   [8:0] piso_2_in;
  wire   [31:0] A_to_mux;
  wire   [31:0] next_accumulate;

  DFFR_X1 \count_reg[1]  ( .D(n51), .CK(Clock), .RN(n78), .Q(n48), .QN(
        net645046) );
  DFFR_X1 \count_reg[2]  ( .D(n50), .CK(Clock), .RN(n78), .QN(n37) );
  DFFS_X1 \count_reg[0]  ( .D(n54), .CK(Clock), .SN(n78), .QN(n40) );
  DFFS_X1 \count_reg[3]  ( .D(n52), .CK(Clock), .SN(n78), .QN(n47) );
  MUX2_X1 U85 ( .A(n49), .B(n48), .S(n86), .Z(n51) );
  MUX2_X1 U87 ( .A(A_to_add[9]), .B(ACC_from_add[9]), .S(n62), .Z(final_out[9]) );
  MUX2_X1 U88 ( .A(A_to_add[8]), .B(ACC_from_add[8]), .S(\input_mux_sel[2] ), 
        .Z(final_out[8]) );
  MUX2_X1 U89 ( .A(A_to_add[7]), .B(ACC_from_add[7]), .S(\input_mux_sel[2] ), 
        .Z(final_out[7]) );
  MUX2_X1 U90 ( .A(A_to_add[6]), .B(ACC_from_add[6]), .S(n62), .Z(final_out[6]) );
  MUX2_X1 U91 ( .A(A_to_add[5]), .B(ACC_from_add[5]), .S(\input_mux_sel[2] ), 
        .Z(final_out[5]) );
  MUX2_X1 U92 ( .A(A_to_add[4]), .B(ACC_from_add[4]), .S(\input_mux_sel[2] ), 
        .Z(final_out[4]) );
  MUX2_X1 U93 ( .A(A_to_add[3]), .B(ACC_from_add[3]), .S(\input_mux_sel[2] ), 
        .Z(final_out[3]) );
  MUX2_X1 U94 ( .A(A_to_add[31]), .B(ACC_from_add[31]), .S(\input_mux_sel[2] ), 
        .Z(final_out[31]) );
  MUX2_X1 U95 ( .A(A_to_add[30]), .B(ACC_from_add[30]), .S(\input_mux_sel[2] ), 
        .Z(final_out[30]) );
  MUX2_X1 U97 ( .A(A_to_add[29]), .B(ACC_from_add[29]), .S(\input_mux_sel[2] ), 
        .Z(final_out[29]) );
  MUX2_X1 U98 ( .A(A_to_add[28]), .B(ACC_from_add[28]), .S(\input_mux_sel[2] ), 
        .Z(final_out[28]) );
  MUX2_X1 U100 ( .A(A_to_add[26]), .B(ACC_from_add[26]), .S(\input_mux_sel[2] ), .Z(final_out[26]) );
  MUX2_X1 U101 ( .A(A_to_add[25]), .B(ACC_from_add[25]), .S(\input_mux_sel[2] ), .Z(final_out[25]) );
  MUX2_X1 U102 ( .A(A_to_add[24]), .B(ACC_from_add[24]), .S(\input_mux_sel[2] ), .Z(final_out[24]) );
  MUX2_X1 U103 ( .A(A_to_add[23]), .B(ACC_from_add[23]), .S(\input_mux_sel[2] ), .Z(final_out[23]) );
  MUX2_X1 U104 ( .A(A_to_add[22]), .B(ACC_from_add[22]), .S(\input_mux_sel[2] ), .Z(final_out[22]) );
  MUX2_X1 U105 ( .A(A_to_add[21]), .B(ACC_from_add[21]), .S(\input_mux_sel[2] ), .Z(final_out[21]) );
  MUX2_X1 U106 ( .A(A_to_add[20]), .B(ACC_from_add[20]), .S(\input_mux_sel[2] ), .Z(final_out[20]) );
  MUX2_X1 U107 ( .A(A_to_add[1]), .B(ACC_from_add[1]), .S(n62), .Z(
        final_out[1]) );
  MUX2_X1 U108 ( .A(A_to_add[19]), .B(ACC_from_add[19]), .S(n62), .Z(
        final_out[19]) );
  MUX2_X1 U109 ( .A(A_to_add[18]), .B(ACC_from_add[18]), .S(n62), .Z(
        final_out[18]) );
  MUX2_X1 U110 ( .A(A_to_add[17]), .B(ACC_from_add[17]), .S(n62), .Z(
        final_out[17]) );
  MUX2_X1 U111 ( .A(A_to_add[16]), .B(ACC_from_add[16]), .S(n62), .Z(
        final_out[16]) );
  MUX2_X1 U112 ( .A(A_to_add[15]), .B(ACC_from_add[15]), .S(n62), .Z(
        final_out[15]) );
  MUX2_X1 U113 ( .A(A_to_add[14]), .B(ACC_from_add[14]), .S(n62), .Z(
        final_out[14]) );
  MUX2_X1 U114 ( .A(A_to_add[13]), .B(ACC_from_add[13]), .S(n62), .Z(
        final_out[13]) );
  MUX2_X1 U115 ( .A(A_to_add[12]), .B(ACC_from_add[12]), .S(n62), .Z(
        final_out[12]) );
  MUX2_X1 U116 ( .A(A_to_add[11]), .B(ACC_from_add[11]), .S(n62), .Z(
        final_out[11]) );
  MUX2_X1 U117 ( .A(A_to_add[10]), .B(ACC_from_add[10]), .S(n62), .Z(
        final_out[10]) );
  booth_encoder_0 encod_0_0 ( .B_in({B[1:0], 1'b0}), .A_out({piso_2_in[0], 
        piso_1_in[0], piso_0_in[0]}) );
  booth_encoder_8 encod_i_1 ( .B_in(B[3:1]), .A_out({piso_2_in[1], 
        piso_1_in[1], piso_0_in[1]}) );
  booth_encoder_7 encod_i_2 ( .B_in(B[5:3]), .A_out({piso_2_in[2], 
        piso_1_in[2], piso_0_in[2]}) );
  booth_encoder_6 encod_i_3 ( .B_in(B[7:5]), .A_out({piso_2_in[3], 
        piso_1_in[3], piso_0_in[3]}) );
  booth_encoder_5 encod_i_4 ( .B_in(B[9:7]), .A_out({piso_2_in[4], 
        piso_1_in[4], piso_0_in[4]}) );
  booth_encoder_4 encod_i_5 ( .B_in(B[11:9]), .A_out({piso_2_in[5], 
        piso_1_in[5], piso_0_in[5]}) );
  booth_encoder_3 encod_i_6 ( .B_in(B[13:11]), .A_out({piso_2_in[6], 
        piso_1_in[6], piso_0_in[6]}) );
  booth_encoder_2 encod_i_7 ( .B_in(B[15:13]), .A_out({piso_2_in[7], 
        piso_1_in[7], piso_0_in[7]}) );
  booth_encoder_1 encod_i_8 ( .B_in({\enc_N2_in[2] , \enc_N2_in[2] , B[15]}), 
        .A_out({piso_2_in[8], piso_1_in[8], piso_0_in[8]}) );
  shift_N9_0 piso_0 ( .Clock(Clock), .ALOAD(n46), .D(piso_0_in), .SO(
        input_mux_sel_0) );
  shift_N9_2 piso_1 ( .Clock(Clock), .ALOAD(n46), .D(piso_1_in), .SO(
        sign_to_add) );
  shift_N9_1 piso_2 ( .Clock(Clock), .ALOAD(n46), .D(piso_2_in), .SO(
        \input_mux_sel[2] ) );
  piso_r_2_N32 A_reg ( .Clock(Clock), .ALOAD(n46), .D({\extend_vector[15] , 
        \extend_vector[15] , \extend_vector[15] , \extend_vector[15] , 
        \extend_vector[15] , \extend_vector[15] , \extend_vector[15] , 
        \extend_vector[15] , \extend_vector[15] , \extend_vector[15] , 
        \extend_vector[15] , \extend_vector[15] , \extend_vector[15] , 
        \extend_vector[15] , \extend_vector[15] , \extend_vector[15] , A}), 
        .SO(A_to_mux) );
  mux21_1 INPUTMUX ( .IN0(A_to_mux), .IN1({A_to_mux[30:0], 1'b0}), .CTRL(
        input_mux_sel_0), .OUT1(B_to_add) );
  ff32_en_SIZE32_1 ACCUMULATOR ( .D(next_accumulate), .en(reg_enable), .clk(
        Clock), .rst(Reset), .Q(A_to_add) );
  NOR2_X1 U20 ( .A1(n46), .A2(n61), .ZN(next_accumulate[31]) );
  NOR2_X1 U38 ( .A1(n46), .A2(n70), .ZN(next_accumulate[23]) );
  NOR2_X1 U30 ( .A1(n46), .A2(n66), .ZN(next_accumulate[27]) );
  NOR2_X1 U40 ( .A1(n46), .A2(n71), .ZN(next_accumulate[22]) );
  NOR2_X1 U32 ( .A1(n46), .A2(n67), .ZN(next_accumulate[26]) );
  NOR2_X1 U26 ( .A1(n46), .A2(n64), .ZN(next_accumulate[29]) );
  NOR2_X1 U28 ( .A1(n46), .A2(n65), .ZN(next_accumulate[28]) );
  NOR2_X1 U34 ( .A1(n46), .A2(n68), .ZN(next_accumulate[25]) );
  NOR2_X1 U42 ( .A1(n46), .A2(n72), .ZN(next_accumulate[21]) );
  NOR2_X1 U44 ( .A1(n46), .A2(n73), .ZN(next_accumulate[20]) );
  NOR2_X1 U36 ( .A1(n46), .A2(n69), .ZN(next_accumulate[24]) );
  NOR2_X1 U48 ( .A1(n46), .A2(n75), .ZN(next_accumulate[19]) );
  NOR2_X1 U60 ( .A1(n46), .A2(n81), .ZN(next_accumulate[13]) );
  NOR2_X1 U58 ( .A1(n46), .A2(n80), .ZN(next_accumulate[14]) );
  NOR2_X1 U62 ( .A1(n46), .A2(n82), .ZN(next_accumulate[12]) );
  NOR2_X1 U56 ( .A1(n46), .A2(n79), .ZN(next_accumulate[15]) );
  NOR2_X1 U10 ( .A1(n46), .A2(n56), .ZN(next_accumulate[7]) );
  NOR2_X1 U64 ( .A1(n46), .A2(n83), .ZN(next_accumulate[11]) );
  NOR2_X1 U8 ( .A1(n46), .A2(n55), .ZN(next_accumulate[8]) );
  NOR2_X1 U6 ( .A1(n46), .A2(n53), .ZN(next_accumulate[9]) );
  NOR2_X1 U52 ( .A1(n46), .A2(n77), .ZN(next_accumulate[17]) );
  NOR2_X1 U50 ( .A1(n46), .A2(n76), .ZN(next_accumulate[18]) );
  NOR2_X1 U66 ( .A1(n46), .A2(n84), .ZN(next_accumulate[10]) );
  NOR2_X1 U18 ( .A1(n46), .A2(n60), .ZN(next_accumulate[3]) );
  NOR2_X1 U12 ( .A1(n46), .A2(n57), .ZN(next_accumulate[6]) );
  NOR2_X1 U14 ( .A1(n46), .A2(n58), .ZN(next_accumulate[5]) );
  NOR2_X1 U16 ( .A1(n46), .A2(n59), .ZN(next_accumulate[4]) );
  NOR2_X1 U24 ( .A1(n46), .A2(n63), .ZN(next_accumulate[2]) );
  NOR2_X1 U46 ( .A1(n46), .A2(n74), .ZN(next_accumulate[1]) );
  NOR2_X1 U68 ( .A1(n46), .A2(n85), .ZN(next_accumulate[0]) );
  NOR2_X1 U4 ( .A1(valid), .A2(n48), .ZN(n49) );
  NAND2_X1 U78 ( .A1(n40), .A2(enable), .ZN(n86) );
  NOR2_X1 U76 ( .A1(n93), .A2(n86), .ZN(n88) );
  NAND2_X1 U74 ( .A1(n88), .A2(n87), .ZN(n91) );
  OAI221_X1 U73 ( .B1(n37), .B2(net645046), .C1(n37), .C2(n90), .A(n91), .ZN(
        n50) );
  OAI211_X1 U70 ( .C1(n40), .C2(enable), .A(n86), .B(n87), .ZN(n54) );
  OAI21_X1 U71 ( .B1(n88), .B2(n47), .A(n87), .ZN(n52) );
  NOR3_X1 U80 ( .A1(n40), .A2(n47), .A3(n93), .ZN(n22) );
  NAND2_X1 U81 ( .A1(n37), .A2(net645046), .ZN(n93) );
  NAND3_X1 U86 ( .A1(n47), .A2(n92), .A3(n40), .ZN(n87) );
  INV_X1 U77 ( .A(n86), .ZN(n90) );
  INV_X1 U75 ( .A(n93), .ZN(n92) );
  INV_X1 U72 ( .A(n87), .ZN(valid) );
  INV_X1 U69 ( .A(ACC_from_add[0]), .ZN(n85) );
  INV_X1 U47 ( .A(ACC_from_add[1]), .ZN(n74) );
  INV_X1 U25 ( .A(ACC_from_add[2]), .ZN(n63) );
  INV_X1 U15 ( .A(ACC_from_add[5]), .ZN(n58) );
  INV_X1 U19 ( .A(ACC_from_add[3]), .ZN(n60) );
  INV_X1 U13 ( .A(ACC_from_add[6]), .ZN(n57) );
  INV_X1 U17 ( .A(ACC_from_add[4]), .ZN(n59) );
  INV_X1 U11 ( .A(ACC_from_add[7]), .ZN(n56) );
  INV_X1 U65 ( .A(ACC_from_add[11]), .ZN(n83) );
  INV_X1 U67 ( .A(ACC_from_add[10]), .ZN(n84) );
  INV_X1 U7 ( .A(ACC_from_add[9]), .ZN(n53) );
  INV_X1 U9 ( .A(ACC_from_add[8]), .ZN(n55) );
  INV_X1 U53 ( .A(ACC_from_add[17]), .ZN(n77) );
  INV_X1 U49 ( .A(ACC_from_add[19]), .ZN(n75) );
  INV_X1 U63 ( .A(ACC_from_add[12]), .ZN(n82) );
  INV_X1 U51 ( .A(ACC_from_add[18]), .ZN(n76) );
  INV_X1 U31 ( .A(ACC_from_add[27]), .ZN(n66) );
  INV_X1 U39 ( .A(ACC_from_add[23]), .ZN(n70) );
  INV_X1 U41 ( .A(ACC_from_add[22]), .ZN(n71) );
  MUX2_X1 U3 ( .A(A_to_add[0]), .B(ACC_from_add[0]), .S(n62), .Z(final_out[0])
         );
  MUX2_X1 U5 ( .A(A_to_add[2]), .B(ACC_from_add[2]), .S(\input_mux_sel[2] ), 
        .Z(final_out[2]) );
  MUX2_X1 U21 ( .A(A_to_add[27]), .B(ACC_from_add[27]), .S(\input_mux_sel[2] ), 
        .Z(final_out[27]) );
  INV_X1 U22 ( .A(ACC_from_add[16]), .ZN(n41) );
  NOR2_X1 U23 ( .A1(n46), .A2(n41), .ZN(next_accumulate[16]) );
  INV_X1 U27 ( .A(ACC_from_add[30]), .ZN(n42) );
  NOR2_X1 U29 ( .A1(n46), .A2(n42), .ZN(next_accumulate[30]) );
  OR2_X2 U33 ( .A1(n46), .A2(\input_mux_sel[2] ), .ZN(reg_enable) );
  AND2_X1 U35 ( .A1(sign), .A2(A[15]), .ZN(\extend_vector[15] ) );
  BUF_X8 U37 ( .A(n22), .Z(n46) );
  INV_X1 U43 ( .A(Reset), .ZN(n78) );
  INV_X1 U45 ( .A(ACC_from_add[14]), .ZN(n80) );
  INV_X1 U54 ( .A(ACC_from_add[21]), .ZN(n72) );
  INV_X1 U55 ( .A(ACC_from_add[26]), .ZN(n67) );
  INV_X1 U57 ( .A(ACC_from_add[20]), .ZN(n73) );
  INV_X1 U59 ( .A(ACC_from_add[15]), .ZN(n79) );
  INV_X1 U61 ( .A(ACC_from_add[13]), .ZN(n81) );
  INV_X1 U79 ( .A(ACC_from_add[29]), .ZN(n64) );
  INV_X1 U82 ( .A(ACC_from_add[25]), .ZN(n68) );
  AND2_X1 U83 ( .A1(sign), .A2(B[15]), .ZN(\enc_N2_in[2] ) );
  INV_X1 U84 ( .A(ACC_from_add[31]), .ZN(n61) );
  INV_X1 U96 ( .A(ACC_from_add[24]), .ZN(n69) );
  INV_X1 U99 ( .A(ACC_from_add[28]), .ZN(n65) );
  BUF_X1 U118 ( .A(\input_mux_sel[2] ), .Z(n62) );
endmodule


module sum_gen_N32_0 ( A, B, Cin, S );
  input [31:0] A;
  input [31:0] B;
  input [8:0] Cin;
  output [31:0] S;


  carry_sel_gen_N4_0_0 csel_N_0 ( .A(A[3:0]), .B(B[3:0]), .Ci(1'b0), .S(S[3:0]) );
  carry_sel_gen_N4_14 csel_N_1 ( .A(A[7:4]), .B(B[7:4]), .Ci(Cin[1]), .S(
        S[7:4]) );
  carry_sel_gen_N4_13 csel_N_2 ( .A(A[11:8]), .B(B[11:8]), .Ci(Cin[2]), .S(
        S[11:8]) );
  carry_sel_gen_N4_12 csel_N_3 ( .A(A[15:12]), .B(B[15:12]), .Ci(Cin[3]), .S(
        S[15:12]) );
  carry_sel_gen_N4_11 csel_N_4 ( .A(A[19:16]), .B(B[19:16]), .Ci(Cin[4]), .S(
        S[19:16]) );
  carry_sel_gen_N4_10 csel_N_5 ( .A(A[23:20]), .B(B[23:20]), .Ci(Cin[5]), .S(
        S[23:20]) );
  carry_sel_gen_N4_9 csel_N_6 ( .A(A[27:24]), .B(B[27:24]), .Ci(Cin[6]), .S(
        S[27:24]) );
  carry_sel_gen_N4_8 csel_N_7 ( .A(A[31:28]), .B(B[31:28]), .Ci(Cin[7]), .S(
        S[31:28]) );
endmodule


module carry_tree_N32_logN5_0 ( A, B, Cin, Cout );
  input [31:0] A;
  input [31:0] B;
  output [7:0] Cout;
  input Cin;
  wire   \magic_pro[0] , \pg_1[13][1] , \pg_1[13][0] , \pg_1[12][1] ,
         \pg_1[12][0] , \pg_1[11][1] , \pg_1[11][0] , \pg_1[10][1] ,
         \pg_1[10][0] , \pg_1[9][1] , \pg_1[9][0] , \pg_1[8][1] , \pg_1[8][0] ,
         \pg_1[7][1] , \pg_1[7][0] , \pg_1[6][1] , \pg_1[6][0] , \pg_1[5][1] ,
         \pg_1[5][0] , \pg_1[4][1] , \pg_1[4][0] , \pg_1[3][1] , \pg_1[3][0] ,
         \pg_1[2][1] , \pg_1[2][0] , \pg_1[1][1] , \pg_1[1][0] , \pg_1[0][0] ,
         \pg_n[4][6][1] , \pg_n[4][6][0] , \pg_n[3][5][1] , \pg_n[3][3][1] ,
         \pg_n[3][3][0] , \pg_n[2][6][1] , \pg_n[2][6][0] , \pg_n[2][5][1] ,
         \pg_n[2][5][0] , \pg_n[2][4][1] , \pg_n[2][3][1] , \pg_n[2][3][0] ,
         \pg_n[2][2][1] , \pg_n[2][2][0] , \pg_n[2][1][1] , \pg_n[2][1][0] ,
         n1, n5, n7, n8;
  wire   [31:1] p_net;
  wire   [31:0] g_net;
  assign Cout[3] = n1;
  assign Cout[1] = n8;

  pg_net_0_0 pg_net_x_1 ( .a(A[1]), .b(B[1]), .g_out(g_net[1]), .p_out(
        p_net[1]) );
  pg_net_62 pg_net_x_2 ( .a(A[2]), .b(B[2]), .g_out(g_net[2]), .p_out(p_net[2]) );
  pg_net_61 pg_net_x_3 ( .a(A[3]), .b(B[3]), .g_out(g_net[3]), .p_out(p_net[3]) );
  pg_net_60 pg_net_x_4 ( .a(A[4]), .b(B[4]), .g_out(g_net[4]), .p_out(p_net[4]) );
  pg_net_59 pg_net_x_5 ( .a(A[5]), .b(B[5]), .g_out(g_net[5]), .p_out(p_net[5]) );
  pg_net_58 pg_net_x_6 ( .a(A[6]), .b(B[6]), .g_out(g_net[6]), .p_out(p_net[6]) );
  pg_net_57 pg_net_x_7 ( .a(A[7]), .b(B[7]), .g_out(g_net[7]), .p_out(p_net[7]) );
  pg_net_56 pg_net_x_8 ( .a(A[8]), .b(B[8]), .g_out(g_net[8]), .p_out(p_net[8]) );
  pg_net_55 pg_net_x_9 ( .a(A[9]), .b(B[9]), .g_out(g_net[9]), .p_out(p_net[9]) );
  pg_net_54 pg_net_x_10 ( .a(A[10]), .b(B[10]), .g_out(g_net[10]), .p_out(
        p_net[10]) );
  pg_net_53 pg_net_x_11 ( .a(A[11]), .b(B[11]), .g_out(g_net[11]), .p_out(
        p_net[11]) );
  pg_net_52 pg_net_x_12 ( .a(A[12]), .b(B[12]), .g_out(g_net[12]), .p_out(
        p_net[12]) );
  pg_net_51 pg_net_x_13 ( .a(A[13]), .b(B[13]), .g_out(g_net[13]), .p_out(
        p_net[13]) );
  pg_net_50 pg_net_x_14 ( .a(A[14]), .b(B[14]), .g_out(g_net[14]), .p_out(
        p_net[14]) );
  pg_net_49 pg_net_x_15 ( .a(A[15]), .b(B[15]), .g_out(g_net[15]), .p_out(
        p_net[15]) );
  pg_net_48 pg_net_x_16 ( .a(A[16]), .b(B[16]), .g_out(g_net[16]), .p_out(
        p_net[16]) );
  pg_net_47 pg_net_x_17 ( .a(A[17]), .b(B[17]), .g_out(g_net[17]), .p_out(
        p_net[17]) );
  pg_net_46 pg_net_x_18 ( .a(A[18]), .b(B[18]), .g_out(g_net[18]), .p_out(
        p_net[18]) );
  pg_net_45 pg_net_x_19 ( .a(A[19]), .b(B[19]), .g_out(g_net[19]), .p_out(
        p_net[19]) );
  pg_net_44 pg_net_x_20 ( .a(A[20]), .b(B[20]), .g_out(g_net[20]), .p_out(
        p_net[20]) );
  pg_net_43 pg_net_x_21 ( .a(A[21]), .b(B[21]), .g_out(g_net[21]), .p_out(
        p_net[21]) );
  pg_net_42 pg_net_x_22 ( .a(A[22]), .b(B[22]), .g_out(g_net[22]), .p_out(
        p_net[22]) );
  pg_net_41 pg_net_x_23 ( .a(A[23]), .b(B[23]), .g_out(g_net[23]), .p_out(
        p_net[23]) );
  pg_net_40 pg_net_x_24 ( .a(A[24]), .b(B[24]), .g_out(g_net[24]), .p_out(
        p_net[24]) );
  pg_net_39 pg_net_x_25 ( .a(A[25]), .b(B[25]), .g_out(g_net[25]), .p_out(
        p_net[25]) );
  pg_net_38 pg_net_x_26 ( .a(A[26]), .b(B[26]), .g_out(g_net[26]), .p_out(
        p_net[26]) );
  pg_net_37 pg_net_x_27 ( .a(A[27]), .b(B[27]), .g_out(g_net[27]), .p_out(
        p_net[27]) );
  pg_net_32 pg_net_0_MAGIC ( .a(A[0]), .b(B[0]), .g_out(\magic_pro[0] ) );
  g_0_0 xG_0_0_MAGIC ( .g(\magic_pro[0] ), .p(1'b0), .g_prec(1'b0), .g_out(
        g_net[0]) );
  g_18 xG_1_0 ( .g(g_net[1]), .p(p_net[1]), .g_prec(g_net[0]), .g_out(
        \pg_1[0][0] ) );
  pg_0_0 xPG_1_1 ( .g(g_net[3]), .p(p_net[3]), .g_prec(g_net[2]), .p_prec(
        p_net[2]), .g_out(\pg_1[1][0] ), .p_out(\pg_1[1][1] ) );
  pg_52 xPG_1_2 ( .g(g_net[5]), .p(p_net[5]), .g_prec(g_net[4]), .p_prec(
        p_net[4]), .g_out(\pg_1[2][0] ), .p_out(\pg_1[2][1] ) );
  pg_51 xPG_1_3 ( .g(g_net[7]), .p(p_net[7]), .g_prec(g_net[6]), .p_prec(
        p_net[6]), .p_out(\pg_1[3][1] ), .g_out_BAR(\pg_1[3][0] ) );
  pg_50 xPG_1_4 ( .g(g_net[9]), .p(p_net[9]), .g_prec(g_net[8]), .p_prec(
        p_net[8]), .g_out(\pg_1[4][0] ), .p_out(\pg_1[4][1] ) );
  pg_49 xPG_1_5 ( .g(g_net[11]), .p(p_net[11]), .g_prec(g_net[10]), .p_prec(
        p_net[10]), .p_out(\pg_1[5][1] ), .g_out_BAR(\pg_1[5][0] ) );
  pg_48 xPG_1_6 ( .g(g_net[13]), .p(p_net[13]), .g_prec(g_net[12]), .p_prec(
        p_net[12]), .g_out(\pg_1[6][0] ), .p_out(\pg_1[6][1] ) );
  pg_47 xPG_1_7 ( .g(g_net[15]), .p(p_net[15]), .g_prec(g_net[14]), .p_prec(
        p_net[14]), .p_out(\pg_1[7][1] ), .g_out_BAR(\pg_1[7][0] ) );
  pg_46 xPG_1_8 ( .g(g_net[17]), .p(p_net[17]), .g_prec(g_net[16]), .p_prec(
        p_net[16]), .g_out(\pg_1[8][0] ), .p_out(\pg_1[8][1] ) );
  pg_45 xPG_1_9 ( .g(g_net[19]), .p(p_net[19]), .g_prec(g_net[18]), .p_prec(
        p_net[18]), .p_out(\pg_1[9][1] ), .g_out_BAR(\pg_1[9][0] ) );
  pg_44 xPG_1_10 ( .g(g_net[21]), .p(p_net[21]), .g_prec(g_net[20]), .p_prec(
        p_net[20]), .g_out(\pg_1[10][0] ), .p_out(\pg_1[10][1] ) );
  pg_43 xPG_1_11 ( .g(g_net[23]), .p(p_net[23]), .g_prec(g_net[22]), .p_prec(
        p_net[22]), .g_out(\pg_1[11][0] ), .p_out(\pg_1[11][1] ) );
  pg_42 xPG_1_12 ( .g(g_net[25]), .p(p_net[25]), .g_prec(g_net[24]), .p_prec(
        p_net[24]), .g_out(\pg_1[12][0] ), .p_out(\pg_1[12][1] ) );
  pg_41 xPG_1_13 ( .g(g_net[27]), .p(p_net[27]), .g_prec(g_net[26]), .p_prec(
        p_net[26]), .p_out(\pg_1[13][1] ), .g_out_BAR(\pg_1[13][0] ) );
  g_17 xG_2_0 ( .g(\pg_1[1][0] ), .p(\pg_1[1][1] ), .g_prec(\pg_1[0][0] ), 
        .g_out(Cout[0]) );
  pg_38 xPG_2_1 ( .p(\pg_1[3][1] ), .g_prec(\pg_1[2][0] ), .p_prec(
        \pg_1[2][1] ), .g_out(\pg_n[2][1][0] ), .p_out(\pg_n[2][1][1] ), 
        .g_BAR(\pg_1[3][0] ) );
  pg_37 xPG_2_2 ( .p(\pg_1[5][1] ), .g_prec(\pg_1[4][0] ), .p_prec(
        \pg_1[4][1] ), .g_out(\pg_n[2][2][0] ), .p_out(\pg_n[2][2][1] ), 
        .g_BAR(\pg_1[5][0] ) );
  pg_36 xPG_2_3 ( .p(\pg_1[7][1] ), .g_prec(\pg_1[6][0] ), .p_prec(
        \pg_1[6][1] ), .g_out(\pg_n[2][3][0] ), .p_out(\pg_n[2][3][1] ), 
        .g_BAR(\pg_1[7][0] ) );
  pg_35 xPG_2_4 ( .p(\pg_1[9][1] ), .g_prec(\pg_1[8][0] ), .p_prec(
        \pg_1[8][1] ), .g_out(n5), .p_out(\pg_n[2][4][1] ), .g_BAR(
        \pg_1[9][0] ) );
  pg_34 xPG_2_5 ( .g(\pg_1[11][0] ), .p(\pg_1[11][1] ), .g_prec(\pg_1[10][0] ), 
        .p_prec(\pg_1[10][1] ), .p_out(\pg_n[2][5][1] ), .g_out_BAR(
        \pg_n[2][5][0] ) );
  pg_33 xPG_2_6 ( .p(\pg_1[13][1] ), .g_prec(\pg_1[12][0] ), .p_prec(
        \pg_1[12][1] ), .g_out(\pg_n[2][6][0] ), .p_out(\pg_n[2][6][1] ), 
        .g_BAR(\pg_1[13][0] ) );
  g_16 xG_3_1 ( .g(\pg_n[2][1][0] ), .p(\pg_n[2][1][1] ), .g_prec(Cout[0]), 
        .g_out(n8) );
  g_15 xG_4_2 ( .g(\pg_n[2][2][0] ), .p(\pg_n[2][2][1] ), .g_prec(n8), .g_out(
        Cout[2]) );
  g_14 xG_4_3 ( .g(\pg_n[3][3][0] ), .p(\pg_n[3][3][1] ), .g_prec(n8), .g_out(
        n1) );
  g_13 xG_5_4 ( .g(n5), .p(\pg_n[2][4][1] ), .g_prec(n1), .g_out(Cout[4]) );
  g_12 xG_5_5 ( .g(n7), .p(\pg_n[3][5][1] ), .g_prec(n1), .g_out(Cout[5]) );
  g_11 xG_5_6 ( .g(\pg_n[4][6][0] ), .p(\pg_n[4][6][1] ), .g_prec(n1), .g_out(
        Cout[6]) );
  pg_31 xPG_3_3 ( .g(\pg_n[2][3][0] ), .p(\pg_n[2][3][1] ), .g_prec(
        \pg_n[2][2][0] ), .p_prec(\pg_n[2][2][1] ), .g_out(\pg_n[3][3][0] ), 
        .p_out(\pg_n[3][3][1] ) );
  pg_30 xPG_3_5 ( .p(\pg_n[2][5][1] ), .g_prec(n5), .p_prec(\pg_n[2][4][1] ), 
        .g_out(n7), .p_out(\pg_n[3][5][1] ), .g_BAR(\pg_n[2][5][0] ) );
  pg_28 xPG_4_6 ( .g(\pg_n[2][6][0] ), .p(\pg_n[2][6][1] ), .g_prec(n7), 
        .p_prec(\pg_n[3][5][1] ), .g_out(\pg_n[4][6][0] ), .p_out(
        \pg_n[4][6][1] ) );
endmodule


module xor_gen_N32_0 ( A, B, S );
  input [31:0] A;
  output [31:0] S;
  input B;
  wire   \A[21] , \A[19] ;
  assign S[31] = A[31];
  assign S[30] = A[30];
  assign S[29] = A[29];
  assign S[28] = A[28];
  assign S[27] = A[27];
  assign S[26] = A[26];
  assign S[25] = A[25];
  assign S[24] = A[24];
  assign S[23] = A[23];
  assign S[22] = A[22];
  assign S[20] = A[20];
  assign S[18] = A[18];
  assign S[17] = A[17];
  assign S[16] = A[16];
  assign S[15] = A[15];
  assign S[14] = A[14];
  assign S[13] = A[13];
  assign S[12] = A[12];
  assign S[11] = A[11];
  assign S[10] = A[10];
  assign S[9] = A[9];
  assign S[8] = A[8];
  assign S[7] = A[7];
  assign S[6] = A[6];
  assign S[5] = A[5];
  assign S[4] = A[4];
  assign S[3] = A[3];
  assign S[2] = A[2];
  assign S[1] = A[1];
  assign S[0] = A[0];
  assign S[21] = \A[21] ;
  assign \A[21]  = A[21];
  assign S[19] = \A[19] ;
  assign \A[19]  = A[19];

endmodule


module ff32_SIZE5 ( D, clk, rst, Q );
  input [4:0] D;
  output [4:0] Q;
  input clk, rst;
  wire   n1, n4, n6, n8, n10;

  DFFR_X1 \Q_reg[4]  ( .D(D[4]), .CK(clk), .RN(n10), .Q(Q[4]) );
  DFFR_X1 \Q_reg[3]  ( .D(D[3]), .CK(clk), .RN(n10), .QN(n4) );
  DFFR_X1 \Q_reg[2]  ( .D(D[2]), .CK(clk), .RN(n10), .QN(n6) );
  DFFR_X1 \Q_reg[1]  ( .D(D[1]), .CK(clk), .RN(n10), .QN(n1) );
  DFFR_X1 \Q_reg[0]  ( .D(D[0]), .CK(clk), .RN(n10), .QN(n8) );
  INV_X1 U3 ( .A(n1), .ZN(Q[1]) );
  INV_X1 U4 ( .A(n4), .ZN(Q[3]) );
  INV_X1 U5 ( .A(n6), .ZN(Q[2]) );
  INV_X1 U6 ( .A(rst), .ZN(n10) );
  INV_X1 U7 ( .A(n8), .ZN(Q[0]) );
endmodule


module ff32_SIZE32 ( D, clk, rst, Q );
  input [31:0] D;
  output [31:0] Q;
  input clk, rst;
  wire   n32;

  DFFR_X1 \Q_reg[31]  ( .D(D[31]), .CK(clk), .RN(n32), .Q(Q[31]) );
  DFFR_X1 \Q_reg[30]  ( .D(D[30]), .CK(clk), .RN(n32), .Q(Q[30]) );
  DFFR_X1 \Q_reg[29]  ( .D(D[29]), .CK(clk), .RN(n32), .Q(Q[29]) );
  DFFR_X1 \Q_reg[28]  ( .D(D[28]), .CK(clk), .RN(n32), .Q(Q[28]) );
  DFFR_X1 \Q_reg[27]  ( .D(D[27]), .CK(clk), .RN(n32), .Q(Q[27]) );
  DFFR_X1 \Q_reg[26]  ( .D(D[26]), .CK(clk), .RN(n32), .Q(Q[26]) );
  DFFR_X1 \Q_reg[25]  ( .D(D[25]), .CK(clk), .RN(n32), .Q(Q[25]) );
  DFFR_X1 \Q_reg[24]  ( .D(D[24]), .CK(clk), .RN(n32), .Q(Q[24]) );
  DFFR_X1 \Q_reg[23]  ( .D(D[23]), .CK(clk), .RN(n32), .Q(Q[23]) );
  DFFR_X1 \Q_reg[22]  ( .D(D[22]), .CK(clk), .RN(n32), .Q(Q[22]) );
  DFFR_X1 \Q_reg[21]  ( .D(D[21]), .CK(clk), .RN(n32), .Q(Q[21]) );
  DFFR_X1 \Q_reg[20]  ( .D(D[20]), .CK(clk), .RN(n32), .Q(Q[20]) );
  DFFR_X1 \Q_reg[19]  ( .D(D[19]), .CK(clk), .RN(n32), .Q(Q[19]) );
  DFFR_X1 \Q_reg[18]  ( .D(D[18]), .CK(clk), .RN(n32), .Q(Q[18]) );
  DFFR_X1 \Q_reg[17]  ( .D(D[17]), .CK(clk), .RN(n32), .Q(Q[17]) );
  DFFR_X1 \Q_reg[16]  ( .D(D[16]), .CK(clk), .RN(n32), .Q(Q[16]) );
  DFFR_X1 \Q_reg[15]  ( .D(D[15]), .CK(clk), .RN(n32), .Q(Q[15]) );
  DFFR_X1 \Q_reg[14]  ( .D(D[14]), .CK(clk), .RN(n32), .Q(Q[14]) );
  DFFR_X1 \Q_reg[13]  ( .D(D[13]), .CK(clk), .RN(n32), .Q(Q[13]) );
  DFFR_X1 \Q_reg[12]  ( .D(D[12]), .CK(clk), .RN(n32), .Q(Q[12]) );
  DFFR_X1 \Q_reg[11]  ( .D(D[11]), .CK(clk), .RN(n32), .Q(Q[11]) );
  DFFR_X1 \Q_reg[10]  ( .D(D[10]), .CK(clk), .RN(n32), .Q(Q[10]) );
  DFFR_X1 \Q_reg[9]  ( .D(D[9]), .CK(clk), .RN(n32), .Q(Q[9]) );
  DFFR_X1 \Q_reg[8]  ( .D(D[8]), .CK(clk), .RN(n32), .Q(Q[8]) );
  DFFR_X1 \Q_reg[7]  ( .D(D[7]), .CK(clk), .RN(n32), .Q(Q[7]) );
  DFFR_X1 \Q_reg[6]  ( .D(D[6]), .CK(clk), .RN(n32), .Q(Q[6]) );
  DFFR_X1 \Q_reg[5]  ( .D(D[5]), .CK(clk), .RN(n32), .Q(Q[5]) );
  DFFR_X1 \Q_reg[4]  ( .D(D[4]), .CK(clk), .RN(n32), .Q(Q[4]) );
  DFFR_X1 \Q_reg[3]  ( .D(D[3]), .CK(clk), .RN(n32), .Q(Q[3]) );
  DFFR_X1 \Q_reg[2]  ( .D(D[2]), .CK(clk), .RN(n32), .Q(Q[2]) );
  DFFR_X1 \Q_reg[1]  ( .D(D[1]), .CK(clk), .RN(n32), .Q(Q[1]) );
  DFFR_X1 \Q_reg[0]  ( .D(D[0]), .CK(clk), .RN(n32), .Q(Q[0]) );
  INV_X2 U3 ( .A(rst), .ZN(n32) );
endmodule


module mux41_MUX_SIZE32_1 ( IN0, IN1, IN2, IN3, CTRL, OUT1 );
  input [31:0] IN0;
  input [31:0] IN1;
  input [31:0] IN2;
  input [31:0] IN3;
  input [1:0] CTRL;
  output [31:0] OUT1;
  wire   n35, n36, n38, n39, n40, n42, n44, n45, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n58, n61, n65, n66, n67, n37, n69, n186, n187,
         n188, n189, n190, n191, n192, n194, n195, n196, n197, n199, n202,
         n203, n204, n205, n206, n207, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n220, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236;

  INV_X1 U23 ( .A(n48), .ZN(OUT1[28]) );
  INV_X1 U31 ( .A(n52), .ZN(OUT1[24]) );
  INV_X1 U25 ( .A(n49), .ZN(OUT1[27]) );
  INV_X1 U21 ( .A(n47), .ZN(OUT1[29]) );
  INV_X1 U15 ( .A(n44), .ZN(OUT1[31]) );
  INV_X1 U17 ( .A(n45), .ZN(OUT1[30]) );
  INV_X1 U39 ( .A(n56), .ZN(OUT1[20]) );
  BUF_X2 U1 ( .A(n35), .Z(n234) );
  BUF_X2 U2 ( .A(n36), .Z(n233) );
  BUF_X2 U3 ( .A(n36), .Z(n231) );
  OR3_X1 U4 ( .A1(n205), .A2(n206), .A3(n207), .ZN(OUT1[2]) );
  OR3_X1 U5 ( .A1(n225), .A2(n224), .A3(n223), .ZN(OUT1[13]) );
  NAND2_X1 U6 ( .A1(IN1[3]), .A2(n233), .ZN(n186) );
  AOI21_X1 U7 ( .B1(n236), .B2(IN0[3]), .A(n220), .ZN(n187) );
  NAND2_X1 U8 ( .A1(n186), .A2(n187), .ZN(OUT1[3]) );
  NAND2_X1 U9 ( .A1(IN2[15]), .A2(n229), .ZN(n188) );
  AOI21_X1 U10 ( .B1(n234), .B2(IN0[15]), .A(n194), .ZN(n189) );
  NAND2_X1 U11 ( .A1(n188), .A2(n189), .ZN(OUT1[15]) );
  NAND2_X1 U12 ( .A1(IN1[17]), .A2(n231), .ZN(n190) );
  AOI21_X1 U13 ( .B1(n234), .B2(IN0[17]), .A(n199), .ZN(n191) );
  NAND2_X1 U14 ( .A1(n190), .A2(n191), .ZN(OUT1[17]) );
  NAND2_X1 U16 ( .A1(IN0[18]), .A2(n234), .ZN(n192) );
  NAND3_X1 U18 ( .A1(n192), .A2(n196), .A3(n197), .ZN(OUT1[18]) );
  BUF_X2 U19 ( .A(n36), .Z(n232) );
  BUF_X2 U20 ( .A(n37), .Z(n230) );
  AND2_X1 U22 ( .A1(n231), .A2(IN1[15]), .ZN(n194) );
  BUF_X2 U24 ( .A(n37), .Z(n195) );
  NAND2_X1 U26 ( .A1(n231), .A2(IN1[18]), .ZN(n196) );
  NAND2_X1 U27 ( .A1(n195), .A2(IN2[18]), .ZN(n197) );
  BUF_X1 U28 ( .A(n37), .Z(n229) );
  BUF_X1 U29 ( .A(n37), .Z(n210) );
  AND2_X1 U30 ( .A1(n210), .A2(IN2[17]), .ZN(n199) );
  NAND3_X1 U32 ( .A1(n202), .A2(n203), .A3(n204), .ZN(OUT1[14]) );
  BUF_X1 U33 ( .A(n35), .Z(n235) );
  INV_X1 U34 ( .A(n50), .ZN(OUT1[26]) );
  AND2_X1 U35 ( .A1(n234), .A2(IN0[13]), .ZN(n223) );
  BUF_X1 U36 ( .A(n35), .Z(n236) );
  INV_X1 U37 ( .A(n61), .ZN(OUT1[16]) );
  INV_X1 U38 ( .A(n55), .ZN(OUT1[21]) );
  INV_X1 U40 ( .A(n53), .ZN(OUT1[23]) );
  INV_X1 U41 ( .A(n58), .ZN(OUT1[19]) );
  INV_X1 U42 ( .A(n54), .ZN(OUT1[22]) );
  INV_X1 U43 ( .A(n66), .ZN(OUT1[11]) );
  AND2_X1 U44 ( .A1(n233), .A2(IN1[13]), .ZN(n224) );
  NAND2_X1 U45 ( .A1(n234), .A2(IN0[14]), .ZN(n202) );
  NAND2_X1 U46 ( .A1(n233), .A2(IN1[14]), .ZN(n203) );
  NAND2_X1 U47 ( .A1(n230), .A2(IN2[14]), .ZN(n204) );
  AND2_X1 U48 ( .A1(n235), .A2(IN0[2]), .ZN(n205) );
  AND2_X1 U49 ( .A1(n232), .A2(IN1[2]), .ZN(n206) );
  AND2_X1 U50 ( .A1(n229), .A2(IN2[2]), .ZN(n207) );
  INV_X1 U51 ( .A(n39), .ZN(OUT1[7]) );
  INV_X1 U52 ( .A(n51), .ZN(OUT1[25]) );
  AND2_X1 U53 ( .A1(n69), .A2(CTRL[0]), .ZN(n36) );
  INV_X1 U54 ( .A(n38), .ZN(OUT1[8]) );
  INV_X1 U55 ( .A(n65), .ZN(OUT1[12]) );
  INV_X1 U56 ( .A(n67), .ZN(OUT1[10]) );
  NOR2_X1 U57 ( .A1(n69), .A2(CTRL[0]), .ZN(n37) );
  INV_X1 U58 ( .A(n40), .ZN(OUT1[6]) );
  INV_X1 U59 ( .A(n42), .ZN(OUT1[4]) );
  AND2_X1 U60 ( .A1(n210), .A2(IN2[13]), .ZN(n225) );
  AND2_X1 U61 ( .A1(n210), .A2(IN2[3]), .ZN(n220) );
  NAND3_X1 U62 ( .A1(n227), .A2(n226), .A3(n228), .ZN(OUT1[9]) );
  INV_X1 U63 ( .A(CTRL[1]), .ZN(n69) );
  NAND2_X1 U64 ( .A1(n230), .A2(IN2[5]), .ZN(n211) );
  NAND2_X1 U65 ( .A1(n195), .A2(IN2[0]), .ZN(n216) );
  AOI222_X1 U66 ( .A1(n235), .A2(IN0[30]), .B1(n233), .B2(IN1[30]), .C1(n210), 
        .C2(IN2[30]), .ZN(n45) );
  AOI222_X1 U67 ( .A1(n235), .A2(IN0[22]), .B1(n233), .B2(IN1[22]), .C1(n210), 
        .C2(IN2[22]), .ZN(n54) );
  AOI222_X1 U68 ( .A1(n234), .A2(IN0[16]), .B1(n233), .B2(IN1[16]), .C1(n210), 
        .C2(IN2[16]), .ZN(n61) );
  AOI222_X1 U69 ( .A1(n235), .A2(IN0[26]), .B1(n231), .B2(IN1[26]), .C1(n195), 
        .C2(IN2[26]), .ZN(n50) );
  NAND2_X1 U70 ( .A1(n230), .A2(IN2[9]), .ZN(n228) );
  AOI222_X1 U71 ( .A1(n235), .A2(IN0[25]), .B1(n231), .B2(IN1[25]), .C1(n230), 
        .C2(IN2[25]), .ZN(n51) );
  AOI222_X1 U72 ( .A1(n236), .A2(IN0[6]), .B1(n232), .B2(IN1[6]), .C1(n210), 
        .C2(IN2[6]), .ZN(n40) );
  AOI222_X1 U73 ( .A1(n236), .A2(IN0[7]), .B1(n232), .B2(IN1[7]), .C1(n195), 
        .C2(IN2[7]), .ZN(n39) );
  NAND3_X1 U74 ( .A1(n216), .A2(n215), .A3(n214), .ZN(OUT1[0]) );
  NAND3_X1 U75 ( .A1(n212), .A2(n211), .A3(n213), .ZN(OUT1[5]) );
  NAND2_X1 U76 ( .A1(n232), .A2(IN1[5]), .ZN(n212) );
  NAND2_X1 U77 ( .A1(n236), .A2(IN0[5]), .ZN(n213) );
  NAND2_X1 U78 ( .A1(n234), .A2(IN0[0]), .ZN(n214) );
  NAND2_X1 U79 ( .A1(n232), .A2(IN1[0]), .ZN(n215) );
  NAND2_X1 U80 ( .A1(n195), .A2(IN2[1]), .ZN(n217) );
  NAND2_X1 U81 ( .A1(n217), .A2(n218), .ZN(OUT1[1]) );
  AOI22_X1 U82 ( .A1(n231), .A2(IN1[1]), .B1(n234), .B2(IN0[1]), .ZN(n218) );
  AOI222_X1 U83 ( .A1(n236), .A2(IN0[31]), .B1(n231), .B2(IN1[31]), .C1(n230), 
        .C2(IN2[31]), .ZN(n44) );
  AOI222_X1 U84 ( .A1(n236), .A2(IN0[4]), .B1(n232), .B2(IN1[4]), .C1(n230), 
        .C2(IN2[4]), .ZN(n42) );
  AOI222_X1 U85 ( .A1(n236), .A2(IN0[8]), .B1(n233), .B2(IN1[8]), .C1(n229), 
        .C2(IN2[8]), .ZN(n38) );
  AOI222_X1 U86 ( .A1(n235), .A2(IN0[24]), .B1(n232), .B2(IN1[24]), .C1(n230), 
        .C2(IN2[24]), .ZN(n52) );
  NAND2_X1 U87 ( .A1(n236), .A2(IN0[9]), .ZN(n226) );
  NAND2_X1 U88 ( .A1(n233), .A2(IN1[9]), .ZN(n227) );
  AOI222_X1 U89 ( .A1(n235), .A2(IN0[20]), .B1(n232), .B2(IN1[20]), .C1(n229), 
        .C2(IN2[20]), .ZN(n56) );
  AOI222_X1 U90 ( .A1(n235), .A2(IN0[28]), .B1(n233), .B2(IN1[28]), .C1(n210), 
        .C2(IN2[28]), .ZN(n48) );
  AOI222_X1 U91 ( .A1(n235), .A2(IN0[29]), .B1(n232), .B2(IN1[29]), .C1(n195), 
        .C2(IN2[29]), .ZN(n47) );
  AOI222_X1 U92 ( .A1(n235), .A2(IN0[23]), .B1(n231), .B2(IN1[23]), .C1(n230), 
        .C2(IN2[23]), .ZN(n53) );
  AOI222_X1 U93 ( .A1(n235), .A2(IN0[27]), .B1(n232), .B2(IN1[27]), .C1(n229), 
        .C2(IN2[27]), .ZN(n49) );
  AOI222_X1 U94 ( .A1(n235), .A2(IN0[21]), .B1(n231), .B2(IN1[21]), .C1(n210), 
        .C2(IN2[21]), .ZN(n55) );
  AOI222_X1 U95 ( .A1(n234), .A2(IN0[19]), .B1(n233), .B2(IN1[19]), .C1(n230), 
        .C2(IN2[19]), .ZN(n58) );
  AOI222_X1 U96 ( .A1(n234), .A2(IN0[12]), .B1(n231), .B2(IN1[12]), .C1(n229), 
        .C2(IN2[12]), .ZN(n65) );
  AOI222_X1 U97 ( .A1(n234), .A2(IN0[11]), .B1(n233), .B2(IN1[11]), .C1(n230), 
        .C2(IN2[11]), .ZN(n66) );
  AOI222_X1 U98 ( .A1(n234), .A2(IN0[10]), .B1(n231), .B2(IN1[10]), .C1(n230), 
        .C2(IN2[10]), .ZN(n67) );
  NOR2_X1 U99 ( .A1(CTRL[0]), .A2(CTRL[1]), .ZN(n35) );
endmodule


module mux41_MUX_SIZE32_0 ( IN0, IN1, IN2, IN3, CTRL, OUT1 );
  input [31:0] IN0;
  input [31:0] IN1;
  input [31:0] IN2;
  input [31:0] IN3;
  input [1:0] CTRL;
  output [31:0] OUT1;
  wire   n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n69, n114, n116, n117, n118, n119, n120,
         n121, n122, n123;

  AOI222_X1 U18 ( .A1(n122), .A2(IN2[30]), .B1(n114), .B2(IN0[30]), .C1(n120), 
        .C2(IN1[30]), .ZN(n45) );
  AOI222_X1 U22 ( .A1(n122), .A2(IN2[29]), .B1(n114), .B2(IN0[29]), .C1(n120), 
        .C2(IN1[29]), .ZN(n47) );
  AOI222_X1 U24 ( .A1(n123), .A2(IN2[28]), .B1(n114), .B2(IN0[28]), .C1(n120), 
        .C2(IN1[28]), .ZN(n48) );
  AOI222_X1 U16 ( .A1(n123), .A2(IN2[31]), .B1(n114), .B2(IN0[31]), .C1(n119), 
        .C2(IN1[31]), .ZN(n44) );
  AOI222_X1 U42 ( .A1(n35), .A2(IN2[1]), .B1(n121), .B2(IN0[1]), .C1(n119), 
        .C2(IN1[1]), .ZN(n57) );
  AOI222_X1 U20 ( .A1(n35), .A2(IN2[2]), .B1(n114), .B2(IN0[2]), .C1(n119), 
        .C2(IN1[2]), .ZN(n46) );
  AOI222_X1 U14 ( .A1(n122), .A2(IN2[3]), .B1(n114), .B2(IN0[3]), .C1(n120), 
        .C2(IN1[3]), .ZN(n43) );
  AOI222_X1 U8 ( .A1(n123), .A2(IN2[6]), .B1(n114), .B2(IN0[6]), .C1(n119), 
        .C2(IN1[6]), .ZN(n40) );
  AOI222_X1 U6 ( .A1(n122), .A2(IN2[7]), .B1(n114), .B2(IN0[7]), .C1(n120), 
        .C2(IN1[7]), .ZN(n39) );
  AOI222_X1 U10 ( .A1(n123), .A2(IN2[5]), .B1(n114), .B2(IN0[5]), .C1(n119), 
        .C2(IN1[5]), .ZN(n41) );
  AOI222_X1 U12 ( .A1(n122), .A2(IN2[4]), .B1(n114), .B2(IN0[4]), .C1(n120), 
        .C2(IN1[4]), .ZN(n42) );
  AOI222_X1 U56 ( .A1(n122), .A2(IN2[13]), .B1(n121), .B2(IN0[13]), .C1(n119), 
        .C2(IN1[13]), .ZN(n64) );
  AOI222_X1 U62 ( .A1(n122), .A2(IN2[10]), .B1(n121), .B2(IN0[10]), .C1(n119), 
        .C2(IN1[10]), .ZN(n67) );
  AOI222_X1 U2 ( .A1(n123), .A2(IN2[9]), .B1(n114), .B2(IN0[9]), .C1(n119), 
        .C2(IN1[9]), .ZN(n34) );
  AOI222_X1 U4 ( .A1(n123), .A2(IN2[8]), .B1(n114), .B2(IN0[8]), .C1(n120), 
        .C2(IN1[8]), .ZN(n38) );
  AOI222_X1 U26 ( .A1(n123), .A2(IN2[27]), .B1(n114), .B2(IN0[27]), .C1(n120), 
        .C2(IN1[27]), .ZN(n49) );
  AOI222_X1 U28 ( .A1(n122), .A2(IN2[26]), .B1(n114), .B2(IN0[26]), .C1(n120), 
        .C2(IN1[26]), .ZN(n50) );
  AOI222_X1 U30 ( .A1(n122), .A2(IN2[25]), .B1(n114), .B2(IN0[25]), .C1(n120), 
        .C2(IN1[25]), .ZN(n51) );
  AOI222_X1 U32 ( .A1(n123), .A2(IN2[24]), .B1(n114), .B2(IN0[24]), .C1(n119), 
        .C2(IN1[24]), .ZN(n52) );
  AOI222_X1 U38 ( .A1(n122), .A2(IN2[21]), .B1(n114), .B2(IN0[21]), .C1(n120), 
        .C2(IN1[21]), .ZN(n55) );
  AOI222_X1 U40 ( .A1(n123), .A2(IN2[20]), .B1(n114), .B2(IN0[20]), .C1(n119), 
        .C2(IN1[20]), .ZN(n56) );
  AOI222_X1 U34 ( .A1(n123), .A2(IN2[23]), .B1(n114), .B2(IN0[23]), .C1(n120), 
        .C2(IN1[23]), .ZN(n53) );
  AOI222_X1 U36 ( .A1(n122), .A2(IN2[22]), .B1(n114), .B2(IN0[22]), .C1(n120), 
        .C2(IN1[22]), .ZN(n54) );
  AOI222_X1 U46 ( .A1(n123), .A2(IN2[18]), .B1(n121), .B2(IN0[18]), .C1(n120), 
        .C2(IN1[18]), .ZN(n59) );
  AOI222_X1 U48 ( .A1(n123), .A2(IN2[17]), .B1(n121), .B2(IN0[17]), .C1(n120), 
        .C2(IN1[17]), .ZN(n60) );
  AND2_X1 U67 ( .A1(CTRL[1]), .A2(n69), .ZN(n35) );
  INV_X1 U57 ( .A(n65), .ZN(OUT1[12]) );
  INV_X1 U49 ( .A(n61), .ZN(OUT1[16]) );
  INV_X1 U53 ( .A(n63), .ZN(OUT1[14]) );
  INV_X1 U47 ( .A(n60), .ZN(OUT1[17]) );
  INV_X1 U51 ( .A(n62), .ZN(OUT1[15]) );
  INV_X1 U45 ( .A(n59), .ZN(OUT1[18]) );
  INV_X1 U55 ( .A(n64), .ZN(OUT1[13]) );
  INV_X1 U11 ( .A(n42), .ZN(OUT1[4]) );
  INV_X1 U15 ( .A(n44), .ZN(OUT1[31]) );
  INV_X1 U17 ( .A(n45), .ZN(OUT1[30]) );
  INV_X1 U21 ( .A(n47), .ZN(OUT1[29]) );
  INV_X1 U23 ( .A(n48), .ZN(OUT1[28]) );
  INV_X1 U5 ( .A(n39), .ZN(OUT1[7]) );
  INV_X1 U25 ( .A(n49), .ZN(OUT1[27]) );
  INV_X1 U3 ( .A(n38), .ZN(OUT1[8]) );
  INV_X1 U27 ( .A(n50), .ZN(OUT1[26]) );
  INV_X1 U1 ( .A(n34), .ZN(OUT1[9]) );
  INV_X1 U29 ( .A(n51), .ZN(OUT1[25]) );
  INV_X1 U31 ( .A(n52), .ZN(OUT1[24]) );
  INV_X1 U33 ( .A(n53), .ZN(OUT1[23]) );
  INV_X1 U35 ( .A(n54), .ZN(OUT1[22]) );
  INV_X1 U37 ( .A(n55), .ZN(OUT1[21]) );
  INV_X1 U7 ( .A(n40), .ZN(OUT1[6]) );
  INV_X1 U39 ( .A(n56), .ZN(OUT1[20]) );
  INV_X1 U43 ( .A(n58), .ZN(OUT1[19]) );
  INV_X1 U61 ( .A(n67), .ZN(OUT1[10]) );
  INV_X1 U59 ( .A(n66), .ZN(OUT1[11]) );
  BUF_X2 U9 ( .A(n37), .Z(n120) );
  BUF_X2 U13 ( .A(n37), .Z(n119) );
  BUF_X2 U19 ( .A(n35), .Z(n123) );
  BUF_X1 U41 ( .A(n35), .Z(n122) );
  BUF_X1 U44 ( .A(n36), .Z(n121) );
  BUF_X2 U50 ( .A(n36), .Z(n114) );
  AND2_X1 U52 ( .A1(n119), .A2(IN1[0]), .ZN(n117) );
  INV_X1 U54 ( .A(n43), .ZN(OUT1[3]) );
  INV_X1 U58 ( .A(n57), .ZN(OUT1[1]) );
  INV_X1 U60 ( .A(n46), .ZN(OUT1[2]) );
  INV_X1 U63 ( .A(n41), .ZN(OUT1[5]) );
  AOI222_X1 U64 ( .A1(n123), .A2(IN2[11]), .B1(n121), .B2(IN0[11]), .C1(n120), 
        .C2(IN1[11]), .ZN(n66) );
  AOI222_X1 U65 ( .A1(n123), .A2(IN2[12]), .B1(n121), .B2(IN0[12]), .C1(n120), 
        .C2(IN1[12]), .ZN(n65) );
  AOI222_X1 U66 ( .A1(n123), .A2(IN2[19]), .B1(n121), .B2(IN0[19]), .C1(n120), 
        .C2(IN1[19]), .ZN(n58) );
  AOI222_X1 U68 ( .A1(n122), .A2(IN2[14]), .B1(n121), .B2(IN0[14]), .C1(n120), 
        .C2(IN1[14]), .ZN(n63) );
  AOI222_X1 U69 ( .A1(n122), .A2(IN2[15]), .B1(n121), .B2(IN0[15]), .C1(n120), 
        .C2(IN1[15]), .ZN(n62) );
  AOI222_X1 U70 ( .A1(n122), .A2(IN2[16]), .B1(n121), .B2(IN0[16]), .C1(n120), 
        .C2(IN1[16]), .ZN(n61) );
  AND2_X1 U71 ( .A1(n121), .A2(IN0[0]), .ZN(n118) );
  AND2_X1 U72 ( .A1(n35), .A2(IN2[0]), .ZN(n116) );
  OR3_X2 U73 ( .A1(n118), .A2(n117), .A3(n116), .ZN(OUT1[0]) );
  NOR2_X1 U74 ( .A1(CTRL[1]), .A2(CTRL[0]), .ZN(n36) );
  NOR2_X1 U75 ( .A1(CTRL[1]), .A2(n69), .ZN(n37) );
  INV_X1 U76 ( .A(CTRL[0]), .ZN(n69) );
endmodule


module mux41_MUX_SIZE5 ( IN0, IN1, IN2, IN3, CTRL, OUT1 );
  input [4:0] IN0;
  input [4:0] IN1;
  input [4:0] IN2;
  input [4:0] IN3;
  input [1:0] CTRL;
  output [4:0] OUT1;
  wire   n1, n2, n3, n4, n5, n6;

  AOI22_X1 U6 ( .A1(CTRL[0]), .A2(IN1[2]), .B1(CTRL[1]), .B2(IN2[2]), .ZN(n4)
         );
  AOI22_X1 U8 ( .A1(CTRL[0]), .A2(IN1[1]), .B1(CTRL[1]), .B2(IN2[1]), .ZN(n5)
         );
  AOI22_X1 U4 ( .A1(CTRL[0]), .A2(IN1[3]), .B1(CTRL[1]), .B2(IN2[3]), .ZN(n3)
         );
  AOI22_X1 U2 ( .A1(CTRL[0]), .A2(IN1[4]), .B1(CTRL[1]), .B2(IN2[4]), .ZN(n1)
         );
  AOI22_X1 U11 ( .A1(CTRL[0]), .A2(IN1[0]), .B1(CTRL[1]), .B2(IN2[0]), .ZN(n6)
         );
  NAND2_X1 U9 ( .A1(n6), .A2(n2), .ZN(OUT1[0]) );
  NAND2_X1 U3 ( .A1(n3), .A2(n2), .ZN(OUT1[3]) );
  NAND2_X1 U1 ( .A1(n1), .A2(n2), .ZN(OUT1[4]) );
  NAND2_X1 U5 ( .A1(n4), .A2(n2), .ZN(OUT1[2]) );
  NAND2_X1 U7 ( .A1(n5), .A2(n2), .ZN(OUT1[1]) );
  NAND2_X1 U10 ( .A1(CTRL[0]), .A2(CTRL[1]), .ZN(n2) );
endmodule


module real_alu_DATA_SIZE32 ( IN1, IN2, ALUW_i, DOUT, stall_o, Clock, Reset );
  input [31:0] IN1;
  input [31:0] IN2;
  input [12:0] ALUW_i;
  output [31:0] DOUT;
  input Clock, Reset;
  output stall_o;
  wire   mux_sign, sign_booth_to_add, valid_from_booth, carry_from_adder,
         overflow, comp_out, n120, n146, n147, n148, n149, n150, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n183, n184, n185, n186, n8, n10, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n38, n39, n40, n41, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n84, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364;
  wire   [31:0] mux_A;
  wire   [31:0] A_booth_to_add;
  wire   [31:0] mux_B;
  wire   [31:0] B_booth_to_add;
  wire   [31:0] mult_out;
  wire   [31:0] sum_out;
  wire   [31:0] shift_out;
  wire   [31:0] lu_out;
  assign n146 = IN2[17];
  assign n147 = IN2[10];
  assign n148 = IN2[19];
  assign n170 = IN2[12];
  assign n171 = IN2[7];
  assign n173 = IN2[6];
  assign n175 = IN2[11];
  assign n176 = IN2[9];
  assign n177 = IN2[15];
  assign n178 = IN2[4];
  assign n180 = IN2[3];
  assign n181 = IN2[1];
  assign n183 = IN2[5];
  assign n184 = IN2[0];
  assign n186 = IN2[2];

  MUX2_X1 U120 ( .A(B_booth_to_add[31]), .B(IN2[31]), .S(n8), .Z(mux_B[31]) );
  MUX2_X1 U121 ( .A(B_booth_to_add[30]), .B(IN2[30]), .S(n8), .Z(mux_B[30]) );
  MUX2_X1 U124 ( .A(B_booth_to_add[28]), .B(IN2[28]), .S(n8), .Z(mux_B[28]) );
  MUX2_X1 U126 ( .A(B_booth_to_add[26]), .B(IN2[26]), .S(n8), .Z(mux_B[26]) );
  MUX2_X1 U127 ( .A(B_booth_to_add[25]), .B(IN2[25]), .S(n8), .Z(mux_B[25]) );
  MUX2_X1 U128 ( .A(B_booth_to_add[24]), .B(IN2[24]), .S(n8), .Z(mux_B[24]) );
  MUX2_X1 U129 ( .A(B_booth_to_add[23]), .B(IN2[23]), .S(n8), .Z(mux_B[23]) );
  MUX2_X1 U130 ( .A(B_booth_to_add[22]), .B(IN2[22]), .S(n8), .Z(mux_B[22]) );
  MUX2_X1 U132 ( .A(B_booth_to_add[20]), .B(IN2[20]), .S(n8), .Z(mux_B[20]) );
  MUX2_X1 U145 ( .A(A_booth_to_add[9]), .B(IN1[9]), .S(n282), .Z(mux_A[9]) );
  MUX2_X1 U146 ( .A(A_booth_to_add[8]), .B(IN1[8]), .S(n282), .Z(mux_A[8]) );
  MUX2_X1 U147 ( .A(A_booth_to_add[7]), .B(IN1[7]), .S(n282), .Z(mux_A[7]) );
  MUX2_X1 U150 ( .A(A_booth_to_add[4]), .B(IN1[4]), .S(n282), .Z(mux_A[4]) );
  MUX2_X1 U151 ( .A(A_booth_to_add[3]), .B(IN1[3]), .S(n282), .Z(mux_A[3]) );
  MUX2_X1 U152 ( .A(A_booth_to_add[31]), .B(IN1[31]), .S(n282), .Z(mux_A[31])
         );
  MUX2_X1 U153 ( .A(A_booth_to_add[30]), .B(IN1[30]), .S(n282), .Z(mux_A[30])
         );
  MUX2_X1 U155 ( .A(A_booth_to_add[29]), .B(IN1[29]), .S(n282), .Z(mux_A[29])
         );
  MUX2_X1 U156 ( .A(A_booth_to_add[28]), .B(IN1[28]), .S(n282), .Z(mux_A[28])
         );
  MUX2_X1 U157 ( .A(A_booth_to_add[27]), .B(IN1[27]), .S(n282), .Z(mux_A[27])
         );
  MUX2_X1 U158 ( .A(A_booth_to_add[26]), .B(IN1[26]), .S(n282), .Z(mux_A[26])
         );
  MUX2_X1 U159 ( .A(A_booth_to_add[25]), .B(IN1[25]), .S(n282), .Z(mux_A[25])
         );
  MUX2_X1 U160 ( .A(A_booth_to_add[24]), .B(IN1[24]), .S(n282), .Z(mux_A[24])
         );
  MUX2_X1 U161 ( .A(A_booth_to_add[23]), .B(IN1[23]), .S(n282), .Z(mux_A[23])
         );
  MUX2_X1 U162 ( .A(A_booth_to_add[22]), .B(IN1[22]), .S(n282), .Z(mux_A[22])
         );
  MUX2_X1 U163 ( .A(A_booth_to_add[21]), .B(IN1[21]), .S(n282), .Z(mux_A[21])
         );
  MUX2_X1 U164 ( .A(A_booth_to_add[20]), .B(IN1[20]), .S(n282), .Z(mux_A[20])
         );
  MUX2_X1 U165 ( .A(A_booth_to_add[1]), .B(IN1[1]), .S(n282), .Z(mux_A[1]) );
  MUX2_X1 U166 ( .A(A_booth_to_add[19]), .B(IN1[19]), .S(n282), .Z(mux_A[19])
         );
  MUX2_X1 U167 ( .A(A_booth_to_add[18]), .B(IN1[18]), .S(n282), .Z(mux_A[18])
         );
  MUX2_X1 U168 ( .A(A_booth_to_add[17]), .B(IN1[17]), .S(n282), .Z(mux_A[17])
         );
  MUX2_X1 U169 ( .A(A_booth_to_add[16]), .B(IN1[16]), .S(n282), .Z(mux_A[16])
         );
  MUX2_X1 U170 ( .A(A_booth_to_add[15]), .B(IN1[15]), .S(n282), .Z(mux_A[15])
         );
  MUX2_X1 U171 ( .A(A_booth_to_add[14]), .B(IN1[14]), .S(n282), .Z(mux_A[14])
         );
  MUX2_X1 U172 ( .A(A_booth_to_add[13]), .B(IN1[13]), .S(n282), .Z(mux_A[13])
         );
  MUX2_X1 U173 ( .A(A_booth_to_add[12]), .B(IN1[12]), .S(n282), .Z(mux_A[12])
         );
  MUX2_X1 U174 ( .A(A_booth_to_add[11]), .B(IN1[11]), .S(n282), .Z(mux_A[11])
         );
  MUX2_X1 U175 ( .A(A_booth_to_add[10]), .B(IN1[10]), .S(n282), .Z(mux_A[10])
         );
  NAND3_X1 U178 ( .A1(n84), .A2(n80), .A3(ALUW_i[12]), .ZN(n31) );
  simple_booth_add_ext_N16 MULT ( .Clock(Clock), .Reset(Reset), .sign(
        ALUW_i[0]), .enable(ALUW_i[1]), .valid(valid_from_booth), .A(IN1[15:0]), .B({n286, IN2[14], n288, n287, n363, n300, n362, n291, n289, n285, n299, 
        n293, n297, n186, n298, n292}), .A_to_add(A_booth_to_add), .B_to_add(
        B_booth_to_add), .sign_to_add(sign_booth_to_add), .final_out(mult_out), 
        .ACC_from_add({n185, sum_out[30], n296, n290, sum_out[27:26], n294, 
        n295, sum_out[23], n169, n174, n179, n120, sum_out[18:14], n283, 
        sum_out[12:0]}) );
  p4add_N32_logN5_1 ADDER ( .A(mux_A), .B(mux_B), .Cin(1'b0), .sign(mux_sign), 
        .S({n185, sum_out[30], n168, n172, sum_out[27:26], n149, n150, 
        sum_out[23], n169, n174, n179, n120, sum_out[18:0]}), .Cout(
        carry_from_adder) );
  comparator_M32 COMP ( .C(carry_from_adder), .V(overflow), .SUM({n185, 
        sum_out[30], n168, n172, sum_out[27:26], n149, n150, sum_out[23], n169, 
        n174, n179, n120, sum_out[18:0]}), .sel(ALUW_i[4:2]), .sign(ALUW_i[0]), 
        .S(comp_out) );
  shifter SHIFT ( .A(IN1), .B({n293, n297, n186, n298, n292}), .LOGIC_ARITH(
        ALUW_i[8]), .LEFT_RIGHT(ALUW_i[9]), .OUTPUT(shift_out) );
  logic_unit_SIZE32 LU ( .IN1(IN1), .IN2({IN2[31:20], n148, IN2[18], n284, 
        IN2[16], n286, IN2[14], n288, n287, n363, n300, n362, n291, n289, n173, 
        n299, n293, n297, n186, n298, n292}), .CTRL(ALUW_i[6:5]), .OUT1(lu_out) );
  MUX2_X1 U134 ( .A(B_booth_to_add[19]), .B(n148), .S(n8), .Z(mux_B[19]) );
  AOI222_X1 U33 ( .A1(IN2[30]), .A2(n16), .B1(n17), .B2(mult_out[30]), .C1(
        n280), .C2(shift_out[30]), .ZN(n34) );
  AOI22_X1 U32 ( .A1(n281), .A2(lu_out[30]), .B1(n15), .B2(sum_out[30]), .ZN(
        n35) );
  NAND2_X1 U31 ( .A1(n34), .A2(n35), .ZN(DOUT[30]) );
  AOI222_X1 U57 ( .A1(IN2[23]), .A2(n16), .B1(n17), .B2(mult_out[23]), .C1(
        n280), .C2(shift_out[23]), .ZN(n50) );
  AOI22_X1 U56 ( .A1(n281), .A2(lu_out[23]), .B1(n364), .B2(sum_out[23]), .ZN(
        n51) );
  NAND2_X1 U55 ( .A1(n50), .A2(n51), .ZN(DOUT[23]) );
  AOI222_X1 U48 ( .A1(IN2[26]), .A2(n16), .B1(n17), .B2(mult_out[26]), .C1(
        n280), .C2(shift_out[26]), .ZN(n44) );
  AOI22_X1 U47 ( .A1(n281), .A2(lu_out[26]), .B1(sum_out[26]), .B2(n15), .ZN(
        n45) );
  NAND2_X1 U46 ( .A1(n44), .A2(n45), .ZN(DOUT[26]) );
  AOI222_X1 U60 ( .A1(IN2[22]), .A2(n16), .B1(n17), .B2(mult_out[22]), .C1(
        n280), .C2(shift_out[22]), .ZN(n52) );
  AOI22_X1 U59 ( .A1(n281), .A2(lu_out[22]), .B1(n364), .B2(n169), .ZN(n53) );
  NAND2_X1 U58 ( .A1(n52), .A2(n53), .ZN(DOUT[22]) );
  AOI222_X1 U39 ( .A1(IN2[29]), .A2(n16), .B1(n17), .B2(mult_out[29]), .C1(
        n280), .C2(shift_out[29]), .ZN(n38) );
  NAND2_X1 U37 ( .A1(n38), .A2(n39), .ZN(DOUT[29]) );
  AOI222_X1 U42 ( .A1(IN2[28]), .A2(n16), .B1(n17), .B2(mult_out[28]), .C1(
        n280), .C2(shift_out[28]), .ZN(n40) );
  NAND2_X1 U40 ( .A1(n40), .A2(n41), .ZN(DOUT[28]) );
  NAND2_X1 U49 ( .A1(n46), .A2(n47), .ZN(DOUT[25]) );
  AOI222_X1 U63 ( .A1(IN2[21]), .A2(n16), .B1(n17), .B2(mult_out[21]), .C1(
        n280), .C2(shift_out[21]), .ZN(n54) );
  NAND2_X1 U61 ( .A1(n54), .A2(n55), .ZN(DOUT[21]) );
  AOI222_X1 U66 ( .A1(IN2[20]), .A2(n16), .B1(n17), .B2(mult_out[20]), .C1(
        n280), .C2(shift_out[20]), .ZN(n56) );
  NAND2_X1 U64 ( .A1(n56), .A2(n57), .ZN(DOUT[20]) );
  AOI222_X1 U54 ( .A1(IN2[24]), .A2(n16), .B1(n17), .B2(mult_out[24]), .C1(
        n280), .C2(shift_out[24]), .ZN(n48) );
  NAND2_X1 U52 ( .A1(n48), .A2(n49), .ZN(DOUT[24]) );
  AOI22_X1 U28 ( .A1(n17), .A2(mult_out[31]), .B1(n280), .B2(shift_out[31]), 
        .ZN(n33) );
  OAI211_X1 U27 ( .C1(n31), .C2(n10), .A(n32), .B(n33), .ZN(DOUT[31]) );
  AOI222_X1 U72 ( .A1(n148), .A2(n16), .B1(n17), .B2(mult_out[19]), .C1(n280), 
        .C2(shift_out[19]), .ZN(n60) );
  AOI22_X1 U71 ( .A1(n281), .A2(lu_out[19]), .B1(n364), .B2(n120), .ZN(n61) );
  NAND2_X1 U70 ( .A1(n60), .A2(n61), .ZN(DOUT[19]) );
  AOI22_X1 U89 ( .A1(n281), .A2(lu_out[13]), .B1(n364), .B2(n283), .ZN(n73) );
  NAND2_X1 U88 ( .A1(n72), .A2(n73), .ZN(DOUT[13]) );
  AOI22_X1 U86 ( .A1(n281), .A2(lu_out[14]), .B1(n364), .B2(sum_out[14]), .ZN(
        n71) );
  NAND2_X1 U85 ( .A1(n70), .A2(n71), .ZN(DOUT[14]) );
  AOI22_X1 U92 ( .A1(n281), .A2(lu_out[12]), .B1(n364), .B2(sum_out[12]), .ZN(
        n75) );
  NAND2_X1 U91 ( .A1(n74), .A2(n75), .ZN(DOUT[12]) );
  AOI222_X1 U96 ( .A1(n363), .A2(n16), .B1(n17), .B2(mult_out[11]), .C1(n280), 
        .C2(shift_out[11]), .ZN(n76) );
  AOI22_X1 U95 ( .A1(n281), .A2(lu_out[11]), .B1(n364), .B2(sum_out[11]), .ZN(
        n77) );
  NAND2_X1 U94 ( .A1(n76), .A2(n77), .ZN(DOUT[11]) );
  AOI222_X1 U84 ( .A1(n286), .A2(n16), .B1(n17), .B2(mult_out[15]), .C1(n18), 
        .C2(shift_out[15]), .ZN(n68) );
  AOI22_X1 U83 ( .A1(n281), .A2(lu_out[15]), .B1(n364), .B2(sum_out[15]), .ZN(
        n69) );
  NAND2_X1 U82 ( .A1(n68), .A2(n69), .ZN(DOUT[15]) );
  AOI22_X1 U13 ( .A1(n281), .A2(lu_out[7]), .B1(n15), .B2(sum_out[7]), .ZN(n22) );
  NAND2_X1 U12 ( .A1(n21), .A2(n22), .ZN(DOUT[7]) );
  AOI22_X1 U77 ( .A1(n281), .A2(lu_out[17]), .B1(n364), .B2(sum_out[17]), .ZN(
        n65) );
  NAND2_X1 U76 ( .A1(n64), .A2(n65), .ZN(DOUT[17]) );
  AOI22_X1 U98 ( .A1(n281), .A2(lu_out[10]), .B1(n364), .B2(sum_out[10]), .ZN(
        n79) );
  NAND2_X1 U97 ( .A1(n78), .A2(n79), .ZN(DOUT[10]) );
  AOI22_X1 U7 ( .A1(n281), .A2(lu_out[9]), .B1(n364), .B2(sum_out[9]), .ZN(n13) );
  NAND2_X1 U6 ( .A1(n12), .A2(n13), .ZN(DOUT[9]) );
  AOI22_X1 U25 ( .A1(n14), .A2(lu_out[3]), .B1(n364), .B2(sum_out[3]), .ZN(n30) );
  NAND2_X1 U24 ( .A1(n29), .A2(n30), .ZN(DOUT[3]) );
  AOI22_X1 U68 ( .A1(n281), .A2(lu_out[1]), .B1(n364), .B2(sum_out[1]), .ZN(
        n59) );
  NAND2_X1 U67 ( .A1(n58), .A2(n59), .ZN(DOUT[1]) );
  AOI222_X1 U11 ( .A1(n291), .A2(n16), .B1(n17), .B2(mult_out[8]), .C1(n280), 
        .C2(shift_out[8]), .ZN(n19) );
  AOI22_X1 U10 ( .A1(n281), .A2(lu_out[8]), .B1(n364), .B2(sum_out[8]), .ZN(
        n20) );
  NAND2_X1 U9 ( .A1(n19), .A2(n20), .ZN(DOUT[8]) );
  AOI222_X1 U75 ( .A1(IN2[18]), .A2(n16), .B1(n17), .B2(mult_out[18]), .C1(
        n280), .C2(shift_out[18]), .ZN(n62) );
  AOI22_X1 U74 ( .A1(n281), .A2(lu_out[18]), .B1(n364), .B2(sum_out[18]), .ZN(
        n63) );
  NAND2_X1 U73 ( .A1(n62), .A2(n63), .ZN(DOUT[18]) );
  AOI222_X1 U81 ( .A1(IN2[16]), .A2(n16), .B1(n17), .B2(mult_out[16]), .C1(n18), .C2(shift_out[16]), .ZN(n66) );
  AOI22_X1 U80 ( .A1(n281), .A2(lu_out[16]), .B1(n364), .B2(sum_out[16]), .ZN(
        n67) );
  NAND2_X1 U79 ( .A1(n66), .A2(n67), .ZN(DOUT[16]) );
  AOI22_X1 U19 ( .A1(n281), .A2(lu_out[5]), .B1(n364), .B2(sum_out[5]), .ZN(
        n26) );
  NAND2_X1 U18 ( .A1(n25), .A2(n26), .ZN(DOUT[5]) );
  AOI22_X1 U22 ( .A1(n281), .A2(lu_out[4]), .B1(n364), .B2(sum_out[4]), .ZN(
        n28) );
  NAND2_X1 U21 ( .A1(n27), .A2(n28), .ZN(DOUT[4]) );
  AOI22_X1 U16 ( .A1(n281), .A2(lu_out[6]), .B1(n364), .B2(sum_out[6]), .ZN(
        n24) );
  NAND2_X1 U15 ( .A1(n23), .A2(n24), .ZN(DOUT[6]) );
  MUX2_X1 U154 ( .A(A_booth_to_add[2]), .B(IN1[2]), .S(n282), .Z(mux_A[2]) );
  MUX2_X1 U149 ( .A(A_booth_to_add[5]), .B(IN1[5]), .S(n282), .Z(mux_A[5]) );
  MUX2_X1 U148 ( .A(A_booth_to_add[6]), .B(IN1[6]), .S(n282), .Z(mux_A[6]) );
  INV_X1 U109 ( .A(ALUW_i[10]), .ZN(n80) );
  NOR2_X1 U2 ( .A1(valid_from_booth), .A2(n282), .ZN(stall_o) );
  NAND2_X1 U3 ( .A1(n329), .A2(n317), .ZN(mux_A[0]) );
  MUX2_X1 U4 ( .A(B_booth_to_add[0]), .B(n184), .S(n282), .Z(mux_B[0]) );
  NAND2_X1 U5 ( .A1(n315), .A2(n349), .ZN(mux_B[3]) );
  AOI22_X1 U8 ( .A1(sum_out[0]), .A2(n364), .B1(n280), .B2(shift_out[0]), .ZN(
        n267) );
  AOI22_X1 U14 ( .A1(n16), .A2(n292), .B1(n17), .B2(mult_out[0]), .ZN(n268) );
  AND2_X1 U17 ( .A1(n267), .A2(n268), .ZN(n359) );
  MUX2_X1 U20 ( .A(B_booth_to_add[5]), .B(n183), .S(n282), .Z(mux_B[5]) );
  OAI21_X1 U23 ( .B1(n282), .B2(n319), .A(n318), .ZN(mux_B[9]) );
  INV_X1 U26 ( .A(n186), .ZN(n269) );
  INV_X1 U29 ( .A(n16), .ZN(n270) );
  AOI22_X1 U30 ( .A1(shift_out[2]), .A2(n280), .B1(mult_out[2]), .B2(n17), 
        .ZN(n271) );
  AOI22_X1 U34 ( .A1(sum_out[2]), .A2(n364), .B1(lu_out[2]), .B2(n281), .ZN(
        n272) );
  OAI211_X1 U35 ( .C1(n269), .C2(n270), .A(n271), .B(n272), .ZN(DOUT[2]) );
  INV_X1 U36 ( .A(n282), .ZN(n273) );
  NAND2_X1 U38 ( .A1(B_booth_to_add[3]), .A2(n273), .ZN(n315) );
  MUX2_X1 U41 ( .A(B_booth_to_add[14]), .B(IN2[14]), .S(n8), .Z(mux_B[14]) );
  MUX2_X1 U43 ( .A(B_booth_to_add[21]), .B(IN2[21]), .S(n8), .Z(mux_B[21]) );
  INV_X1 U44 ( .A(n8), .ZN(n274) );
  NAND2_X1 U45 ( .A1(B_booth_to_add[16]), .A2(n274), .ZN(n304) );
  MUX2_X1 U50 ( .A(B_booth_to_add[29]), .B(IN2[29]), .S(n8), .Z(mux_B[29]) );
  INV_X1 U51 ( .A(IN2[27]), .ZN(n275) );
  INV_X1 U53 ( .A(n16), .ZN(n276) );
  AOI22_X1 U62 ( .A1(shift_out[27]), .A2(n280), .B1(mult_out[27]), .B2(n17), 
        .ZN(n277) );
  AOI22_X1 U65 ( .A1(sum_out[27]), .A2(n364), .B1(lu_out[27]), .B2(n281), .ZN(
        n278) );
  OAI211_X1 U69 ( .C1(n275), .C2(n276), .A(n277), .B(n278), .ZN(DOUT[27]) );
  CLKBUF_X1 U78 ( .A(n177), .Z(n279) );
  CLKBUF_X1 U87 ( .A(n170), .Z(n287) );
  AOI222_X1 U90 ( .A1(IN2[25]), .A2(n16), .B1(n17), .B2(mult_out[25]), .C1(
        n280), .C2(shift_out[25]), .ZN(n46) );
  BUF_X1 U93 ( .A(n149), .Z(n294) );
  AOI222_X1 U99 ( .A1(n284), .A2(n16), .B1(n17), .B2(mult_out[17]), .C1(n280), 
        .C2(shift_out[17]), .ZN(n64) );
  AOI222_X1 U100 ( .A1(n300), .A2(n16), .B1(n17), .B2(mult_out[10]), .C1(n280), 
        .C2(shift_out[10]), .ZN(n78) );
  AOI222_X1 U101 ( .A1(n299), .A2(n16), .B1(n17), .B2(mult_out[5]), .C1(n280), 
        .C2(shift_out[5]), .ZN(n25) );
  AOI222_X1 U102 ( .A1(n289), .A2(n16), .B1(n17), .B2(mult_out[7]), .C1(n280), 
        .C2(shift_out[7]), .ZN(n21) );
  AOI222_X1 U103 ( .A1(n298), .A2(n16), .B1(n17), .B2(mult_out[1]), .C1(n280), 
        .C2(shift_out[1]), .ZN(n58) );
  BUF_X1 U104 ( .A(n184), .Z(n292) );
  BUF_X1 U105 ( .A(n147), .Z(n300) );
  BUF_X1 U106 ( .A(n181), .Z(n298) );
  BUF_X1 U107 ( .A(n146), .Z(n284) );
  OR2_X1 U108 ( .A1(n282), .A2(n330), .ZN(n317) );
  OR2_X1 U110 ( .A1(n282), .A2(n332), .ZN(n311) );
  OR2_X1 U111 ( .A1(n282), .A2(n342), .ZN(n312) );
  OR2_X1 U112 ( .A1(n282), .A2(n340), .ZN(n316) );
  OR2_X1 U113 ( .A1(n282), .A2(n346), .ZN(n313) );
  OR2_X1 U114 ( .A1(n282), .A2(n328), .ZN(n310) );
  OR2_X1 U115 ( .A1(n282), .A2(n348), .ZN(n314) );
  AND2_X2 U116 ( .A1(n31), .A2(ALUW_i[12]), .ZN(n17) );
  CLKBUF_X3 U117 ( .A(n8), .Z(n282) );
  INV_X2 U118 ( .A(ALUW_i[1]), .ZN(n8) );
  AOI222_X1 U119 ( .A1(IN2[14]), .A2(n16), .B1(n17), .B2(mult_out[14]), .C1(
        n18), .C2(shift_out[14]), .ZN(n70) );
  BUF_X1 U122 ( .A(n172), .Z(n290) );
  INV_X1 U123 ( .A(n359), .ZN(n358) );
  INV_X1 U125 ( .A(n360), .ZN(n357) );
  BUF_X1 U131 ( .A(n173), .Z(n285) );
  BUF_X1 U133 ( .A(n171), .Z(n289) );
  INV_X1 U135 ( .A(IN2[31]), .ZN(n10) );
  BUF_X1 U136 ( .A(n178), .Z(n293) );
  BUF_X1 U137 ( .A(IN2[8]), .Z(n291) );
  OR2_X1 U138 ( .A1(n8), .A2(n336), .ZN(n306) );
  OR2_X1 U139 ( .A1(n8), .A2(n338), .ZN(n307) );
  OR2_X1 U140 ( .A1(n8), .A2(n323), .ZN(n302) );
  OR2_X1 U141 ( .A1(n8), .A2(n344), .ZN(n308) );
  OR2_X1 U142 ( .A1(n8), .A2(n325), .ZN(n303) );
  OR2_X1 U143 ( .A1(n8), .A2(n321), .ZN(n301) );
  OR2_X1 U144 ( .A1(n8), .A2(n334), .ZN(n305) );
  OR2_X1 U176 ( .A1(n8), .A2(n351), .ZN(n309) );
  INV_X1 U177 ( .A(B_booth_to_add[9]), .ZN(n319) );
  INV_X1 U179 ( .A(B_booth_to_add[4]), .ZN(n346) );
  INV_X1 U180 ( .A(B_booth_to_add[8]), .ZN(n342) );
  INV_X1 U181 ( .A(B_booth_to_add[6]), .ZN(n328) );
  INV_X1 U182 ( .A(B_booth_to_add[7]), .ZN(n348) );
  BUF_X2 U183 ( .A(n15), .Z(n364) );
  INV_X1 U184 ( .A(B_booth_to_add[13]), .ZN(n338) );
  INV_X1 U185 ( .A(B_booth_to_add[12]), .ZN(n323) );
  BUF_X2 U186 ( .A(n18), .Z(n280) );
  INV_X1 U187 ( .A(B_booth_to_add[11]), .ZN(n334) );
  INV_X1 U188 ( .A(B_booth_to_add[1]), .ZN(n351) );
  INV_X1 U189 ( .A(B_booth_to_add[10]), .ZN(n340) );
  INV_X1 U190 ( .A(B_booth_to_add[15]), .ZN(n336) );
  INV_X1 U191 ( .A(B_booth_to_add[2]), .ZN(n332) );
  INV_X1 U192 ( .A(B_booth_to_add[17]), .ZN(n344) );
  BUF_X2 U193 ( .A(n14), .Z(n281) );
  INV_X1 U194 ( .A(B_booth_to_add[27]), .ZN(n321) );
  INV_X1 U195 ( .A(B_booth_to_add[18]), .ZN(n325) );
  INV_X1 U196 ( .A(ALUW_i[11]), .ZN(n84) );
  INV_X1 U197 ( .A(A_booth_to_add[0]), .ZN(n330) );
  BUF_X1 U198 ( .A(sum_out[13]), .Z(n283) );
  CLKBUF_X1 U199 ( .A(n176), .Z(n362) );
  BUF_X1 U200 ( .A(n279), .Z(n286) );
  CLKBUF_X1 U201 ( .A(IN2[13]), .Z(n288) );
  CLKBUF_X1 U202 ( .A(n150), .Z(n295) );
  CLKBUF_X1 U203 ( .A(n168), .Z(n296) );
  BUF_X1 U204 ( .A(n180), .Z(n297) );
  BUF_X1 U205 ( .A(n183), .Z(n299) );
  AOI222_X1 U206 ( .A1(n285), .A2(n16), .B1(n17), .B2(mult_out[6]), .C1(n280), 
        .C2(shift_out[6]), .ZN(n23) );
  INV_X1 U207 ( .A(n355), .ZN(DOUT[0]) );
  NOR3_X1 U208 ( .A1(ALUW_i[12]), .A2(ALUW_i[11]), .A3(ALUW_i[10]), .ZN(n15)
         );
  NOR3_X1 U209 ( .A1(ALUW_i[12]), .A2(ALUW_i[10]), .A3(n84), .ZN(n18) );
  BUF_X1 U210 ( .A(n175), .Z(n363) );
  INV_X2 U211 ( .A(n31), .ZN(n16) );
  MUX2_X2 U212 ( .A(sign_booth_to_add), .B(ALUW_i[7]), .S(n8), .Z(mux_sign) );
  AOI222_X1 U213 ( .A1(n293), .A2(n16), .B1(n17), .B2(mult_out[4]), .C1(n280), 
        .C2(shift_out[4]), .ZN(n27) );
  AOI222_X1 U214 ( .A1(n297), .A2(n16), .B1(n17), .B2(mult_out[3]), .C1(n280), 
        .C2(shift_out[3]), .ZN(n29) );
  AOI222_X1 U215 ( .A1(n362), .A2(n16), .B1(n17), .B2(mult_out[9]), .C1(n280), 
        .C2(shift_out[9]), .ZN(n12) );
  AOI222_X1 U216 ( .A1(n287), .A2(n16), .B1(n17), .B2(mult_out[12]), .C1(n18), 
        .C2(shift_out[12]), .ZN(n74) );
  AOI222_X1 U217 ( .A1(n288), .A2(n16), .B1(n17), .B2(mult_out[13]), .C1(n280), 
        .C2(shift_out[13]), .ZN(n72) );
  OAI21_X1 U218 ( .B1(lu_out[0]), .B2(ALUW_i[11]), .A(n361), .ZN(n360) );
  NOR2_X1 U219 ( .A1(n80), .A2(ALUW_i[12]), .ZN(n361) );
  NAND2_X1 U220 ( .A1(n359), .A2(ALUW_i[11]), .ZN(n356) );
  NOR2_X1 U221 ( .A1(n10), .A2(IN1[31]), .ZN(n354) );
  NAND2_X1 U222 ( .A1(n10), .A2(IN1[31]), .ZN(n352) );
  NOR3_X1 U223 ( .A1(ALUW_i[12]), .A2(ALUW_i[11]), .A3(n80), .ZN(n14) );
  NAND2_X1 U224 ( .A1(n176), .A2(n282), .ZN(n318) );
  NAND2_X1 U225 ( .A1(IN2[27]), .A2(n8), .ZN(n320) );
  NAND2_X1 U226 ( .A1(n320), .A2(n301), .ZN(mux_B[27]) );
  NAND2_X1 U227 ( .A1(n170), .A2(n8), .ZN(n322) );
  NAND2_X1 U228 ( .A1(n322), .A2(n302), .ZN(mux_B[12]) );
  NAND2_X1 U229 ( .A1(IN2[18]), .A2(n8), .ZN(n324) );
  NAND2_X1 U230 ( .A1(n324), .A2(n303), .ZN(mux_B[18]) );
  NAND2_X1 U231 ( .A1(IN2[16]), .A2(n8), .ZN(n326) );
  NAND2_X1 U232 ( .A1(n326), .A2(n304), .ZN(mux_B[16]) );
  NAND2_X1 U233 ( .A1(n173), .A2(n282), .ZN(n327) );
  NAND2_X1 U234 ( .A1(n327), .A2(n310), .ZN(mux_B[6]) );
  NAND2_X1 U235 ( .A1(IN1[0]), .A2(n282), .ZN(n329) );
  NAND2_X1 U236 ( .A1(n186), .A2(n282), .ZN(n331) );
  NAND2_X1 U237 ( .A1(n331), .A2(n311), .ZN(mux_B[2]) );
  NAND2_X1 U238 ( .A1(n175), .A2(n8), .ZN(n333) );
  NAND2_X1 U239 ( .A1(n333), .A2(n305), .ZN(mux_B[11]) );
  NAND2_X1 U240 ( .A1(n177), .A2(n8), .ZN(n335) );
  NAND2_X1 U241 ( .A1(n335), .A2(n306), .ZN(mux_B[15]) );
  NAND2_X1 U242 ( .A1(IN2[13]), .A2(n8), .ZN(n337) );
  NAND2_X1 U243 ( .A1(n337), .A2(n307), .ZN(mux_B[13]) );
  NAND2_X1 U244 ( .A1(n147), .A2(n282), .ZN(n339) );
  NAND2_X1 U245 ( .A1(n339), .A2(n316), .ZN(mux_B[10]) );
  NAND2_X1 U246 ( .A1(IN2[8]), .A2(n282), .ZN(n341) );
  NAND2_X1 U247 ( .A1(n341), .A2(n312), .ZN(mux_B[8]) );
  NAND2_X1 U248 ( .A1(n146), .A2(n8), .ZN(n343) );
  NAND2_X1 U249 ( .A1(n343), .A2(n308), .ZN(mux_B[17]) );
  NAND2_X1 U250 ( .A1(n178), .A2(n282), .ZN(n345) );
  NAND2_X1 U251 ( .A1(n345), .A2(n313), .ZN(mux_B[4]) );
  NAND2_X1 U252 ( .A1(n171), .A2(n282), .ZN(n347) );
  NAND2_X1 U253 ( .A1(n347), .A2(n314), .ZN(mux_B[7]) );
  NAND2_X1 U254 ( .A1(n180), .A2(n282), .ZN(n349) );
  NAND2_X1 U255 ( .A1(n181), .A2(n8), .ZN(n350) );
  NAND2_X1 U256 ( .A1(n350), .A2(n309), .ZN(mux_B[1]) );
  NAND2_X1 U257 ( .A1(n185), .A2(n354), .ZN(n353) );
  OAI21_X1 U258 ( .B1(n185), .B2(n352), .A(n353), .ZN(overflow) );
  OAI22_X1 U259 ( .A1(comp_out), .A2(n356), .B1(n357), .B2(n358), .ZN(n355) );
  AOI22_X1 U260 ( .A1(n281), .A2(lu_out[25]), .B1(n15), .B2(n294), .ZN(n47) );
  AOI22_X1 U261 ( .A1(n281), .A2(lu_out[21]), .B1(n364), .B2(n174), .ZN(n55)
         );
  AOI22_X1 U262 ( .A1(n281), .A2(lu_out[29]), .B1(n364), .B2(n296), .ZN(n39)
         );
  AOI22_X1 U263 ( .A1(n281), .A2(lu_out[28]), .B1(n364), .B2(n290), .ZN(n41)
         );
  AOI22_X1 U264 ( .A1(n281), .A2(lu_out[24]), .B1(n364), .B2(n295), .ZN(n49)
         );
  AOI22_X1 U265 ( .A1(n281), .A2(lu_out[20]), .B1(n364), .B2(n179), .ZN(n57)
         );
  AOI22_X1 U266 ( .A1(n281), .A2(lu_out[31]), .B1(n185), .B2(n364), .ZN(n32)
         );
endmodule


module mux21_0 ( IN0, IN1, CTRL, OUT1 );
  input [31:0] IN0;
  input [31:0] IN1;
  output [31:0] OUT1;
  input CTRL;
  wire   n15, n16, n17, n18, n19, n20, n21;

  MUX2_X1 U8 ( .A(IN0[31]), .B(IN1[31]), .S(CTRL), .Z(OUT1[31]) );
  MUX2_X1 U9 ( .A(IN0[30]), .B(IN1[30]), .S(CTRL), .Z(OUT1[30]) );
  MUX2_X1 U11 ( .A(IN0[29]), .B(IN1[29]), .S(CTRL), .Z(OUT1[29]) );
  MUX2_X1 U12 ( .A(IN0[28]), .B(IN1[28]), .S(CTRL), .Z(OUT1[28]) );
  MUX2_X1 U14 ( .A(IN0[26]), .B(IN1[26]), .S(CTRL), .Z(OUT1[26]) );
  MUX2_X1 U16 ( .A(IN0[24]), .B(IN1[24]), .S(CTRL), .Z(OUT1[24]) );
  MUX2_X1 U18 ( .A(IN0[22]), .B(IN1[22]), .S(CTRL), .Z(OUT1[22]) );
  MUX2_X1 U19 ( .A(IN0[21]), .B(IN1[21]), .S(CTRL), .Z(OUT1[21]) );
  MUX2_X1 U20 ( .A(IN0[20]), .B(IN1[20]), .S(CTRL), .Z(OUT1[20]) );
  MUX2_X1 U22 ( .A(IN0[19]), .B(IN1[19]), .S(CTRL), .Z(OUT1[19]) );
  MUX2_X1 U1 ( .A(IN0[13]), .B(IN1[13]), .S(CTRL), .Z(OUT1[13]) );
  MUX2_X1 U2 ( .A(IN0[17]), .B(IN1[17]), .S(CTRL), .Z(OUT1[17]) );
  MUX2_X1 U3 ( .A(IN0[12]), .B(IN1[12]), .S(CTRL), .Z(OUT1[12]) );
  MUX2_X1 U4 ( .A(IN0[18]), .B(IN1[18]), .S(CTRL), .Z(OUT1[18]) );
  MUX2_X1 U5 ( .A(IN0[14]), .B(IN1[14]), .S(CTRL), .Z(OUT1[14]) );
  MUX2_X1 U6 ( .A(IN0[15]), .B(IN1[15]), .S(CTRL), .Z(OUT1[15]) );
  MUX2_X2 U7 ( .A(IN0[27]), .B(IN1[27]), .S(CTRL), .Z(OUT1[27]) );
  MUX2_X2 U10 ( .A(IN0[16]), .B(IN1[16]), .S(CTRL), .Z(OUT1[16]) );
  MUX2_X1 U13 ( .A(IN0[8]), .B(IN1[8]), .S(CTRL), .Z(OUT1[8]) );
  MUX2_X1 U15 ( .A(IN0[10]), .B(IN1[10]), .S(CTRL), .Z(OUT1[10]) );
  MUX2_X1 U17 ( .A(IN0[4]), .B(IN1[4]), .S(CTRL), .Z(OUT1[4]) );
  MUX2_X2 U21 ( .A(IN0[23]), .B(IN1[23]), .S(CTRL), .Z(OUT1[23]) );
  NAND2_X1 U23 ( .A1(n16), .A2(n17), .ZN(OUT1[6]) );
  NAND2_X1 U24 ( .A1(n20), .A2(n21), .ZN(OUT1[7]) );
  NAND2_X1 U25 ( .A1(n18), .A2(n19), .ZN(OUT1[0]) );
  MUX2_X1 U26 ( .A(IN0[3]), .B(IN1[3]), .S(CTRL), .Z(OUT1[3]) );
  NAND2_X1 U27 ( .A1(IN0[6]), .A2(n15), .ZN(n16) );
  NAND2_X1 U28 ( .A1(IN1[6]), .A2(CTRL), .ZN(n17) );
  INV_X1 U29 ( .A(CTRL), .ZN(n15) );
  MUX2_X2 U30 ( .A(IN0[2]), .B(IN1[2]), .S(CTRL), .Z(OUT1[2]) );
  MUX2_X1 U31 ( .A(IN0[1]), .B(IN1[1]), .S(CTRL), .Z(OUT1[1]) );
  MUX2_X1 U32 ( .A(IN0[5]), .B(IN1[5]), .S(CTRL), .Z(OUT1[5]) );
  MUX2_X1 U33 ( .A(IN0[25]), .B(IN1[25]), .S(CTRL), .Z(OUT1[25]) );
  MUX2_X1 U34 ( .A(IN0[11]), .B(IN1[11]), .S(CTRL), .Z(OUT1[11]) );
  NAND2_X1 U35 ( .A1(CTRL), .A2(IN1[7]), .ZN(n21) );
  NAND2_X1 U36 ( .A1(IN1[0]), .A2(CTRL), .ZN(n19) );
  NAND2_X1 U37 ( .A1(IN0[0]), .A2(n15), .ZN(n18) );
  NAND2_X1 U38 ( .A1(IN0[7]), .A2(n15), .ZN(n20) );
  MUX2_X1 U39 ( .A(IN0[9]), .B(IN1[9]), .S(CTRL), .Z(OUT1[9]) );
endmodule


module ff32_en_SIZE13 ( D, en, clk, rst, Q );
  input [12:0] D;
  output [12:0] Q;
  input en, clk, rst;
  wire   n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n40, n1,
         n2, net645036, net645037, net645038, net645039, net645040, net645041,
         net645042, net645043, net645044, net645045, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n18;

  DFFR_X1 \Q_reg[12]  ( .D(n40), .CK(clk), .RN(n18), .Q(Q[12]), .QN(net645045)
         );
  DFFR_X1 \Q_reg[11]  ( .D(n38), .CK(clk), .RN(n18), .Q(Q[11]), .QN(net645044)
         );
  DFFR_X1 \Q_reg[10]  ( .D(n37), .CK(clk), .RN(n18), .Q(Q[10]), .QN(net645043)
         );
  DFFR_X1 \Q_reg[8]  ( .D(n35), .CK(clk), .RN(n18), .Q(Q[8]), .QN(net645042)
         );
  DFFR_X1 \Q_reg[7]  ( .D(n34), .CK(clk), .RN(n18), .Q(Q[7]), .QN(net645041)
         );
  DFFR_X1 \Q_reg[5]  ( .D(n32), .CK(clk), .RN(n18), .Q(Q[5]), .QN(net645040)
         );
  DFFR_X1 \Q_reg[4]  ( .D(n31), .CK(clk), .RN(n18), .Q(Q[4]), .QN(net645039)
         );
  DFFR_X1 \Q_reg[3]  ( .D(n30), .CK(clk), .RN(n18), .Q(Q[3]), .QN(net645038)
         );
  DFFR_X1 \Q_reg[2]  ( .D(n29), .CK(clk), .RN(n18), .Q(Q[2]), .QN(net645037)
         );
  DFFR_X1 \Q_reg[1]  ( .D(n28), .CK(clk), .RN(n18), .Q(Q[1]) );
  DFFR_X1 \Q_reg[0]  ( .D(n27), .CK(clk), .RN(n18), .Q(Q[0]), .QN(net645036)
         );
  MUX2_X1 U27 ( .A(Q[1]), .B(D[1]), .S(en), .Z(n28) );
  DFFR_X1 \Q_reg[6]  ( .D(n33), .CK(clk), .RN(n18), .Q(Q[6]), .QN(n1) );
  NAND2_X1 U8 ( .A1(en), .A2(D[10]), .ZN(n7) );
  OAI21_X1 U7 ( .B1(en), .B2(net645043), .A(n7), .ZN(n37) );
  NAND2_X1 U6 ( .A1(en), .A2(D[11]), .ZN(n6) );
  OAI21_X1 U5 ( .B1(en), .B2(net645044), .A(n6), .ZN(n38) );
  NAND2_X1 U3 ( .A1(en), .A2(D[12]), .ZN(n5) );
  OAI21_X1 U2 ( .B1(en), .B2(net645045), .A(n5), .ZN(n40) );
  NAND2_X1 U12 ( .A1(en), .A2(D[8]), .ZN(n9) );
  OAI21_X1 U11 ( .B1(en), .B2(net645042), .A(n9), .ZN(n35) );
  NAND2_X1 U10 ( .A1(en), .A2(D[9]), .ZN(n8) );
  OAI21_X1 U9 ( .B1(en), .B2(n2), .A(n8), .ZN(n36) );
  NAND2_X1 U24 ( .A1(en), .A2(D[2]), .ZN(n15) );
  OAI21_X1 U23 ( .B1(en), .B2(net645037), .A(n15), .ZN(n29) );
  NAND2_X1 U22 ( .A1(en), .A2(D[3]), .ZN(n14) );
  OAI21_X1 U21 ( .B1(en), .B2(net645038), .A(n14), .ZN(n30) );
  NAND2_X1 U16 ( .A1(en), .A2(D[6]), .ZN(n11) );
  OAI21_X1 U15 ( .B1(en), .B2(n1), .A(n11), .ZN(n33) );
  NAND2_X1 U14 ( .A1(en), .A2(D[7]), .ZN(n10) );
  OAI21_X1 U13 ( .B1(en), .B2(net645041), .A(n10), .ZN(n34) );
  NAND2_X1 U18 ( .A1(en), .A2(D[5]), .ZN(n12) );
  OAI21_X1 U17 ( .B1(en), .B2(net645040), .A(n12), .ZN(n32) );
  NAND2_X1 U26 ( .A1(en), .A2(D[0]), .ZN(n16) );
  OAI21_X1 U25 ( .B1(en), .B2(net645036), .A(n16), .ZN(n27) );
  NAND2_X1 U20 ( .A1(en), .A2(D[4]), .ZN(n13) );
  OAI21_X1 U19 ( .B1(en), .B2(net645039), .A(n13), .ZN(n31) );
  DFFR_X2 \Q_reg[9]  ( .D(n36), .CK(clk), .RN(n18), .Q(Q[9]), .QN(n2) );
  INV_X1 U4 ( .A(rst), .ZN(n18) );
endmodule


module ff32_en_SIZE5_3 ( D, en, clk, rst, Q );
  input [4:0] D;
  output [4:0] Q;
  input en, clk, rst;
  wire   n1, n3, n4, n5, n6, net645267, net645268, net645269, net645270,
         net645271, n8, n9, n10, n11, n12, n13;

  DFFR_X1 \Q_reg[4]  ( .D(n1), .CK(clk), .RN(n13), .Q(Q[4]), .QN(net645271) );
  DFFR_X1 \Q_reg[3]  ( .D(n3), .CK(clk), .RN(n13), .Q(Q[3]), .QN(net645270) );
  DFFR_X1 \Q_reg[2]  ( .D(n4), .CK(clk), .RN(n13), .Q(Q[2]), .QN(net645269) );
  DFFR_X1 \Q_reg[0]  ( .D(n6), .CK(clk), .RN(n13), .Q(Q[0]), .QN(net645267) );
  DFFR_X1 \Q_reg[1]  ( .D(n5), .CK(clk), .RN(n13), .Q(Q[1]), .QN(net645268) );
  NAND2_X1 U7 ( .A1(en), .A2(D[2]), .ZN(n10) );
  OAI21_X1 U6 ( .B1(en), .B2(net645269), .A(n10), .ZN(n4) );
  NAND2_X1 U9 ( .A1(en), .A2(D[3]), .ZN(n11) );
  OAI21_X1 U8 ( .B1(en), .B2(net645270), .A(n11), .ZN(n3) );
  NAND2_X1 U12 ( .A1(en), .A2(D[4]), .ZN(n12) );
  OAI21_X1 U11 ( .B1(en), .B2(net645271), .A(n12), .ZN(n1) );
  NAND2_X1 U5 ( .A1(en), .A2(D[1]), .ZN(n9) );
  OAI21_X1 U4 ( .B1(en), .B2(net645268), .A(n9), .ZN(n5) );
  NAND2_X1 U3 ( .A1(en), .A2(D[0]), .ZN(n8) );
  OAI21_X1 U2 ( .B1(en), .B2(net645267), .A(n8), .ZN(n6) );
  INV_X1 U10 ( .A(rst), .ZN(n13) );
endmodule


module ff32_en_SIZE5_0 ( D, en, clk, rst, Q );
  input [4:0] D;
  output [4:0] Q;
  input en, clk, rst;
  wire   n11, n12, n13, n14, n16, net645031, net645032, net645033, net645034,
         net645035, n2, n3, n4, n5, n6, n7;

  DFFR_X1 \Q_reg[4]  ( .D(n16), .CK(clk), .RN(n7), .Q(Q[4]), .QN(net645035) );
  DFFR_X1 \Q_reg[3]  ( .D(n14), .CK(clk), .RN(n7), .Q(Q[3]), .QN(net645034) );
  DFFR_X1 \Q_reg[2]  ( .D(n13), .CK(clk), .RN(n7), .Q(Q[2]), .QN(net645033) );
  DFFR_X1 \Q_reg[1]  ( .D(n12), .CK(clk), .RN(n7), .Q(Q[1]), .QN(net645032) );
  DFFR_X1 \Q_reg[0]  ( .D(n11), .CK(clk), .RN(n7), .Q(Q[0]), .QN(net645031) );
  NAND2_X1 U10 ( .A1(en), .A2(D[1]), .ZN(n5) );
  OAI21_X1 U9 ( .B1(en), .B2(net645032), .A(n5), .ZN(n12) );
  NAND2_X1 U8 ( .A1(en), .A2(D[2]), .ZN(n4) );
  OAI21_X1 U7 ( .B1(en), .B2(net645033), .A(n4), .ZN(n13) );
  NAND2_X1 U6 ( .A1(en), .A2(D[3]), .ZN(n3) );
  OAI21_X1 U5 ( .B1(en), .B2(net645034), .A(n3), .ZN(n14) );
  NAND2_X1 U12 ( .A1(en), .A2(D[0]), .ZN(n6) );
  OAI21_X1 U11 ( .B1(en), .B2(net645031), .A(n6), .ZN(n11) );
  NAND2_X1 U3 ( .A1(en), .A2(D[4]), .ZN(n2) );
  OAI21_X1 U2 ( .B1(en), .B2(net645035), .A(n2), .ZN(n16) );
  INV_X1 U4 ( .A(rst), .ZN(n7) );
endmodule


module ff32_en_SIZE32_0 ( D, en, clk, rst, Q );
  input [31:0] D;
  output [31:0] Q;
  input en, clk, rst;
  wire   n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n97, net645107, net645108, net645109, net645110,
         net645111, net645112, net645113, net645114, net645115, net645116,
         net645117, net645118, net645119, net645120, net645121, net645122,
         net645123, net645124, net645125, net645126, net645127, net645128,
         net645129, net645130, net645131, net645132, net645133, net645134,
         net645135, net645136, net645137, net645138, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n36, n37,
         n38;

  DFFR_X1 \Q_reg[31]  ( .D(n97), .CK(clk), .RN(n38), .Q(Q[31]), .QN(net645138)
         );
  DFFR_X1 \Q_reg[30]  ( .D(n95), .CK(clk), .RN(n38), .Q(Q[30]), .QN(net645137)
         );
  DFFR_X1 \Q_reg[29]  ( .D(n94), .CK(clk), .RN(n38), .Q(Q[29]), .QN(net645136)
         );
  DFFR_X1 \Q_reg[28]  ( .D(n93), .CK(clk), .RN(n38), .Q(Q[28]), .QN(net645135)
         );
  DFFR_X1 \Q_reg[27]  ( .D(n92), .CK(clk), .RN(n38), .Q(Q[27]), .QN(net645134)
         );
  DFFR_X1 \Q_reg[26]  ( .D(n91), .CK(clk), .RN(n38), .Q(Q[26]), .QN(net645133)
         );
  DFFR_X1 \Q_reg[25]  ( .D(n90), .CK(clk), .RN(n38), .Q(Q[25]), .QN(net645132)
         );
  DFFR_X1 \Q_reg[24]  ( .D(n89), .CK(clk), .RN(n38), .Q(Q[24]), .QN(net645131)
         );
  DFFR_X1 \Q_reg[23]  ( .D(n88), .CK(clk), .RN(n38), .Q(Q[23]), .QN(net645130)
         );
  DFFR_X1 \Q_reg[22]  ( .D(n87), .CK(clk), .RN(n38), .Q(Q[22]), .QN(net645129)
         );
  DFFR_X1 \Q_reg[21]  ( .D(n86), .CK(clk), .RN(n38), .Q(Q[21]), .QN(net645128)
         );
  DFFR_X1 \Q_reg[19]  ( .D(n84), .CK(clk), .RN(n38), .Q(Q[19]), .QN(net645127)
         );
  DFFR_X1 \Q_reg[18]  ( .D(n83), .CK(clk), .RN(n38), .Q(Q[18]), .QN(net645126)
         );
  DFFR_X1 \Q_reg[17]  ( .D(n82), .CK(clk), .RN(n38), .Q(Q[17]), .QN(net645125)
         );
  DFFR_X1 \Q_reg[16]  ( .D(n81), .CK(clk), .RN(n38), .Q(Q[16]), .QN(net645124)
         );
  DFFR_X1 \Q_reg[15]  ( .D(n80), .CK(clk), .RN(n38), .Q(Q[15]), .QN(net645123)
         );
  DFFR_X1 \Q_reg[14]  ( .D(n79), .CK(clk), .RN(n38), .Q(Q[14]), .QN(net645122)
         );
  DFFR_X1 \Q_reg[13]  ( .D(n78), .CK(clk), .RN(n38), .Q(Q[13]), .QN(net645121)
         );
  DFFR_X1 \Q_reg[12]  ( .D(n77), .CK(clk), .RN(n38), .Q(Q[12]), .QN(net645120)
         );
  DFFR_X1 \Q_reg[11]  ( .D(n76), .CK(clk), .RN(n38), .Q(Q[11]), .QN(net645119)
         );
  DFFR_X1 \Q_reg[10]  ( .D(n75), .CK(clk), .RN(n38), .Q(Q[10]), .QN(net645118)
         );
  DFFR_X1 \Q_reg[9]  ( .D(n74), .CK(clk), .RN(n38), .Q(Q[9]), .QN(net645117)
         );
  DFFR_X1 \Q_reg[8]  ( .D(n73), .CK(clk), .RN(n38), .Q(Q[8]), .QN(net645116)
         );
  DFFR_X1 \Q_reg[7]  ( .D(n72), .CK(clk), .RN(n38), .Q(Q[7]), .QN(net645115)
         );
  DFFR_X1 \Q_reg[6]  ( .D(n71), .CK(clk), .RN(n38), .Q(Q[6]), .QN(net645114)
         );
  DFFR_X1 \Q_reg[5]  ( .D(n70), .CK(clk), .RN(n38), .Q(Q[5]), .QN(net645113)
         );
  DFFR_X1 \Q_reg[4]  ( .D(n69), .CK(clk), .RN(n38), .Q(Q[4]), .QN(net645112)
         );
  DFFR_X1 \Q_reg[3]  ( .D(n68), .CK(clk), .RN(n38), .Q(Q[3]), .QN(net645111)
         );
  DFFR_X1 \Q_reg[2]  ( .D(n67), .CK(clk), .RN(n38), .Q(Q[2]), .QN(net645110)
         );
  DFFR_X1 \Q_reg[1]  ( .D(n66), .CK(clk), .RN(n38), .Q(Q[1]), .QN(net645109)
         );
  DFFR_X1 \Q_reg[0]  ( .D(n65), .CK(clk), .RN(n38), .Q(Q[0]), .QN(net645108)
         );
  DFFR_X1 \Q_reg[20]  ( .D(n85), .CK(clk), .RN(n38), .Q(Q[20]), .QN(net645107)
         );
  NAND2_X1 U39 ( .A1(n36), .A2(D[13]), .ZN(n20) );
  OAI21_X1 U38 ( .B1(en), .B2(net645121), .A(n20), .ZN(n78) );
  NAND2_X1 U37 ( .A1(n36), .A2(D[14]), .ZN(n19) );
  OAI21_X1 U36 ( .B1(en), .B2(net645122), .A(n19), .ZN(n79) );
  NAND2_X1 U45 ( .A1(n36), .A2(D[10]), .ZN(n23) );
  OAI21_X1 U44 ( .B1(en), .B2(net645118), .A(n23), .ZN(n75) );
  NAND2_X1 U43 ( .A1(n36), .A2(D[11]), .ZN(n22) );
  OAI21_X1 U42 ( .B1(en), .B2(net645119), .A(n22), .ZN(n76) );
  NAND2_X1 U59 ( .A1(n37), .A2(D[3]), .ZN(n30) );
  OAI21_X1 U58 ( .B1(n36), .B2(net645111), .A(n30), .ZN(n68) );
  NAND2_X1 U23 ( .A1(n37), .A2(D[21]), .ZN(n12) );
  OAI21_X1 U22 ( .B1(n36), .B2(net645128), .A(n12), .ZN(n86) );
  NAND2_X1 U57 ( .A1(n37), .A2(D[4]), .ZN(n29) );
  OAI21_X1 U56 ( .B1(n36), .B2(net645112), .A(n29), .ZN(n69) );
  NAND2_X1 U55 ( .A1(en), .A2(D[5]), .ZN(n28) );
  OAI21_X1 U54 ( .B1(n36), .B2(net645113), .A(n28), .ZN(n70) );
  NAND2_X1 U61 ( .A1(n37), .A2(D[2]), .ZN(n31) );
  OAI21_X1 U60 ( .B1(n36), .B2(net645110), .A(n31), .ZN(n67) );
  NAND2_X1 U49 ( .A1(en), .A2(D[8]), .ZN(n25) );
  OAI21_X1 U48 ( .B1(n36), .B2(net645116), .A(n25), .ZN(n73) );
  NAND2_X1 U53 ( .A1(n37), .A2(D[6]), .ZN(n27) );
  OAI21_X1 U52 ( .B1(n36), .B2(net645114), .A(n27), .ZN(n71) );
  NAND2_X1 U25 ( .A1(en), .A2(D[20]), .ZN(n13) );
  OAI21_X1 U24 ( .B1(n37), .B2(net645107), .A(n13), .ZN(n85) );
  NAND2_X1 U27 ( .A1(en), .A2(D[19]), .ZN(n14) );
  OAI21_X1 U26 ( .B1(en), .B2(net645127), .A(n14), .ZN(n84) );
  NAND2_X1 U47 ( .A1(en), .A2(D[9]), .ZN(n24) );
  OAI21_X1 U46 ( .B1(en), .B2(net645117), .A(n24), .ZN(n74) );
  NAND2_X1 U51 ( .A1(en), .A2(D[7]), .ZN(n26) );
  OAI21_X1 U50 ( .B1(en), .B2(net645115), .A(n26), .ZN(n72) );
  NAND2_X1 U19 ( .A1(n37), .A2(D[23]), .ZN(n10) );
  OAI21_X1 U18 ( .B1(en), .B2(net645130), .A(n10), .ZN(n88) );
  NAND2_X1 U9 ( .A1(n37), .A2(D[28]), .ZN(n5) );
  OAI21_X1 U8 ( .B1(en), .B2(net645135), .A(n5), .ZN(n93) );
  NAND2_X1 U7 ( .A1(n37), .A2(D[29]), .ZN(n4) );
  OAI21_X1 U6 ( .B1(en), .B2(net645136), .A(n4), .ZN(n94) );
  NAND2_X1 U41 ( .A1(en), .A2(D[12]), .ZN(n21) );
  OAI21_X1 U40 ( .B1(en), .B2(net645120), .A(n21), .ZN(n77) );
  NAND2_X1 U21 ( .A1(en), .A2(D[22]), .ZN(n11) );
  OAI21_X1 U20 ( .B1(en), .B2(net645129), .A(n11), .ZN(n87) );
  NAND2_X1 U29 ( .A1(en), .A2(D[18]), .ZN(n15) );
  OAI21_X1 U28 ( .B1(en), .B2(net645126), .A(n15), .ZN(n83) );
  NAND2_X1 U11 ( .A1(n37), .A2(D[27]), .ZN(n6) );
  OAI21_X1 U10 ( .B1(en), .B2(net645134), .A(n6), .ZN(n92) );
  NAND2_X1 U31 ( .A1(en), .A2(D[17]), .ZN(n16) );
  OAI21_X1 U30 ( .B1(en), .B2(net645125), .A(n16), .ZN(n82) );
  NAND2_X1 U35 ( .A1(en), .A2(D[15]), .ZN(n18) );
  OAI21_X1 U34 ( .B1(en), .B2(net645123), .A(n18), .ZN(n80) );
  NAND2_X1 U33 ( .A1(en), .A2(D[16]), .ZN(n17) );
  OAI21_X1 U32 ( .B1(en), .B2(net645124), .A(n17), .ZN(n81) );
  NAND2_X1 U15 ( .A1(n37), .A2(D[25]), .ZN(n8) );
  OAI21_X1 U14 ( .B1(en), .B2(net645132), .A(n8), .ZN(n90) );
  NAND2_X1 U13 ( .A1(n37), .A2(D[26]), .ZN(n7) );
  OAI21_X1 U12 ( .B1(en), .B2(net645133), .A(n7), .ZN(n91) );
  NAND2_X1 U17 ( .A1(n37), .A2(D[24]), .ZN(n9) );
  OAI21_X1 U16 ( .B1(en), .B2(net645131), .A(n9), .ZN(n89) );
  NAND2_X1 U63 ( .A1(en), .A2(D[1]), .ZN(n32) );
  OAI21_X1 U62 ( .B1(n36), .B2(net645109), .A(n32), .ZN(n66) );
  NAND2_X1 U65 ( .A1(en), .A2(D[0]), .ZN(n33) );
  OAI21_X1 U64 ( .B1(n36), .B2(net645108), .A(n33), .ZN(n65) );
  NAND2_X1 U5 ( .A1(en), .A2(D[30]), .ZN(n3) );
  OAI21_X1 U4 ( .B1(en), .B2(net645137), .A(n3), .ZN(n95) );
  NAND2_X1 U3 ( .A1(en), .A2(D[31]), .ZN(n2) );
  OAI21_X1 U2 ( .B1(en), .B2(net645138), .A(n2), .ZN(n97) );
  INV_X2 U66 ( .A(rst), .ZN(n38) );
  BUF_X1 U67 ( .A(en), .Z(n37) );
  BUF_X1 U68 ( .A(en), .Z(n36) );
endmodule


module alu_ctrl ( .OP({\OP[4] , \OP[3] , \OP[2] , \OP[1] , \OP[0] }), ALU_WORD
 );
  output [12:0] ALU_WORD;
  input \OP[4] , \OP[3] , \OP[2] , \OP[1] , \OP[0] ;
  wire   N20, N21, N22, N23, N24, N25, N26, N27, N29, N30, N31, N32, N33, n37,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n38, n39, n40;

  DLH_X1 \comp_sel_reg[2]  ( .G(N32), .D(N33), .Q(ALU_WORD[4]) );
  DLH_X1 \comp_sel_reg[1]  ( .G(N32), .D(N31), .Q(ALU_WORD[3]) );
  DLH_X1 \comp_sel_reg[0]  ( .G(N32), .D(N30), .Q(ALU_WORD[2]) );
  DLH_X1 sign_to_booth_reg ( .G(N20), .D(N21), .Q(ALU_WORD[0]) );
  DLH_X1 left_right_reg ( .G(N23), .D(N22), .Q(ALU_WORD[9]) );
  DLH_X1 logic_arith_reg ( .G(N23), .D(N24), .Q(ALU_WORD[8]) );
  DLH_X1 sign_to_adder_reg ( .G(N25), .D(N26), .Q(ALU_WORD[7]) );
  DLL_X1 \lu_ctrl_reg[1]  ( .D(N29), .GN(n37), .Q(ALU_WORD[6]) );
  DLL_X1 \lu_ctrl_reg[0]  ( .D(N27), .GN(n37), .Q(ALU_WORD[5]) );
  NAND3_X1 U43 ( .A1(n21), .A2(n37), .A3(n27), .ZN(ALU_WORD[10]) );
  NAND3_X1 U44 ( .A1(n17), .A2(n29), .A3(OP[2]), .ZN(n13) );
  OAI33_X1 U45 ( .A1(n14), .A2(n17), .A3(n19), .B1(n26), .B2(n30), .B3(OP[3]), 
        .ZN(n25) );
  NAND3_X1 U46 ( .A1(n15), .A2(OP[0]), .A3(OP[1]), .ZN(n12) );
  NAND3_X1 U47 ( .A1(OP[1]), .A2(n17), .A3(n15), .ZN(n35) );
  NAND2_X1 U42 ( .A1(OP[4]), .A2(OP[3]), .ZN(n16) );
  NOR2_X1 U36 ( .A1(OP[2]), .A2(OP[1]), .ZN(n33) );
  NAND2_X1 U35 ( .A1(OP[0]), .A2(n33), .ZN(n18) );
  NOR2_X1 U34 ( .A1(n18), .A2(n16), .ZN(n39) );
  NAND2_X1 U32 ( .A1(OP[2]), .A2(OP[1]), .ZN(n19) );
  NAND2_X1 U31 ( .A1(n33), .A2(n17), .ZN(n26) );
  AOI221_X1 U28 ( .B1(n13), .B2(n30), .C1(n13), .C2(n12), .A(n31), .ZN(n40) );
  AOI211_X1 U26 ( .C1(n38), .C2(n34), .A(n39), .B(N30), .ZN(n36) );
  OAI221_X1 U25 ( .B1(n17), .B2(n29), .C1(OP[0]), .C2(OP[1]), .A(OP[2]), .ZN(
        n32) );
  OAI211_X1 U23 ( .C1(n16), .C2(n35), .A(n36), .B(n23), .ZN(N32) );
  NOR2_X1 U21 ( .A1(n14), .A2(n35), .ZN(N29) );
  AOI21_X1 U20 ( .B1(n33), .B2(n34), .A(N29), .ZN(n37) );
  NOR2_X1 U19 ( .A1(n16), .A2(n32), .ZN(ALU_WORD[1]) );
  NOR3_X1 U16 ( .A1(OP[2]), .A2(n29), .A3(n20), .ZN(N22) );
  OAI21_X1 U14 ( .B1(n18), .B2(n20), .A(n28), .ZN(N23) );
  OAI21_X1 U12 ( .B1(n26), .B2(n20), .A(n27), .ZN(ALU_WORD[12]) );
  NOR2_X1 U4 ( .A1(n14), .A2(n18), .ZN(N27) );
  NOR2_X1 U7 ( .A1(n12), .A2(n20), .ZN(N24) );
  OAI21_X1 U5 ( .B1(n19), .B2(n20), .A(n21), .ZN(N26) );
  AOI21_X1 U2 ( .B1(n12), .B2(n13), .A(n14), .ZN(N33) );
  OAI211_X1 U8 ( .C1(n19), .C2(n22), .A(n23), .B(n24), .ZN(N21) );
  AOI221_X1 U3 ( .B1(OP[2]), .B2(n14), .C1(n15), .C2(n16), .A(n17), .ZN(N31)
         );
  OAI21_X1 U6 ( .B1(n15), .B2(n20), .A(n21), .ZN(N25) );
  NOR2_X1 U37 ( .A1(n31), .A2(OP[4]), .ZN(n34) );
  NAND2_X1 U17 ( .A1(n30), .A2(n31), .ZN(n20) );
  INV_X1 U29 ( .A(OP[1]), .ZN(n29) );
  INV_X1 U41 ( .A(OP[0]), .ZN(n17) );
  INV_X1 U40 ( .A(OP[2]), .ZN(n15) );
  INV_X1 U30 ( .A(OP[4]), .ZN(n30) );
  INV_X1 U38 ( .A(OP[3]), .ZN(n31) );
  OR2_X1 U10 ( .A1(OP[0]), .A2(n16), .ZN(n22) );
  INV_X1 U39 ( .A(n12), .ZN(n38) );
  INV_X1 U33 ( .A(n34), .ZN(n14) );
  INV_X1 U18 ( .A(ALU_WORD[1]), .ZN(n27) );
  OR2_X1 U24 ( .A1(n14), .A2(n32), .ZN(n23) );
  INV_X1 U15 ( .A(N22), .ZN(n28) );
  INV_X1 U9 ( .A(n25), .ZN(n24) );
  OR2_X1 U27 ( .A1(n25), .A2(n40), .ZN(N30) );
  OR2_X1 U13 ( .A1(N32), .A2(N23), .ZN(ALU_WORD[11]) );
  OR2_X1 U11 ( .A1(N32), .A2(ALU_WORD[12]), .ZN(N20) );
  INV_X1 U22 ( .A(N32), .ZN(n21) );
endmodule


module cw_mem_MICROCODE_MEM_SIZE64_OP_CODE_SIZE6_CW_SIZE13 ( OPCODE_IN, CW_OUT
 );
  input [5:0] OPCODE_IN;
  output [12:0] CW_OUT;
  wire   CW_OUT_4, CW_OUT_3, CW_OUT_2, CW_OUT_1, CW_OUT_0, n9, n10, n11, n12,
         n13, n14, n15, n16, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n17, n30, n31, n32, n33, n34, n35, n36, n37;
  assign CW_OUT[4] = CW_OUT_4;
  assign CW_OUT[3] = CW_OUT_3;
  assign CW_OUT[2] = CW_OUT_2;
  assign CW_OUT[1] = CW_OUT_1;
  assign CW_OUT[0] = CW_OUT_0;

  NAND2_X1 U29 ( .A1(n29), .A2(n28), .ZN(n14) );
  AOI21_X1 U11 ( .B1(n20), .B2(n26), .A(CW_OUT[7]), .ZN(n25) );
  INV_X1 U19 ( .A(OPCODE_IN[0]), .ZN(n12) );
  OR3_X1 U2 ( .A1(CW_OUT_1), .A2(CW_OUT_4), .A3(n13), .ZN(CW_OUT_0) );
  OR2_X1 U9 ( .A1(CW_OUT_3), .A2(n13), .ZN(CW_OUT[6]) );
  OAI21_X1 U1 ( .B1(n14), .B2(n30), .A(n35), .ZN(CW_OUT[11]) );
  OR2_X1 U3 ( .A1(n22), .A2(n27), .ZN(n30) );
  OAI221_X1 U4 ( .B1(n22), .B2(n23), .C1(n22), .C2(n24), .A(n25), .ZN(n13) );
  NAND2_X1 U5 ( .A1(n16), .A2(n21), .ZN(CW_OUT[12]) );
  CLKBUF_X1 U6 ( .A(n21), .Z(n35) );
  OR2_X1 U7 ( .A1(n33), .A2(CW_OUT[12]), .ZN(CW_OUT[9]) );
  NOR2_X1 U8 ( .A1(n11), .A2(n31), .ZN(CW_OUT[10]) );
  NOR2_X1 U10 ( .A1(n10), .A2(OPCODE_IN[5]), .ZN(n20) );
  INV_X1 U12 ( .A(OPCODE_IN[1]), .ZN(n27) );
  NAND2_X1 U13 ( .A1(OPCODE_IN[1]), .A2(n19), .ZN(n11) );
  INV_X1 U14 ( .A(OPCODE_IN[4]), .ZN(n22) );
  NOR2_X1 U15 ( .A1(OPCODE_IN[4]), .A2(OPCODE_IN[2]), .ZN(n19) );
  INV_X1 U16 ( .A(OPCODE_IN[3]), .ZN(n10) );
  INV_X1 U17 ( .A(OPCODE_IN[2]), .ZN(n28) );
  OR2_X1 U18 ( .A1(OPCODE_IN[3]), .A2(OPCODE_IN[5]), .ZN(n37) );
  INV_X1 U20 ( .A(CW_OUT[10]), .ZN(n16) );
  BUF_X1 U21 ( .A(n11), .Z(n36) );
  OR3_X2 U22 ( .A1(n15), .A2(n28), .A3(n37), .ZN(n21) );
  OR2_X1 U23 ( .A1(OPCODE_IN[5]), .A2(OPCODE_IN[3]), .ZN(n31) );
  NOR2_X1 U24 ( .A1(OPCODE_IN[2]), .A2(OPCODE_IN[4]), .ZN(n32) );
  NAND2_X1 U25 ( .A1(n32), .A2(n20), .ZN(n17) );
  NOR2_X1 U26 ( .A1(OPCODE_IN[0]), .A2(n17), .ZN(n33) );
  NAND2_X1 U27 ( .A1(n22), .A2(n27), .ZN(n34) );
  OAI22_X1 U28 ( .A1(n14), .A2(n34), .B1(n16), .B2(n12), .ZN(CW_OUT_4) );
  INV_X1 U30 ( .A(OPCODE_IN[5]), .ZN(n9) );
  NOR2_X1 U31 ( .A1(OPCODE_IN[5]), .A2(OPCODE_IN[3]), .ZN(n29) );
  NOR4_X1 U32 ( .A1(n9), .A2(n10), .A3(n36), .A4(n12), .ZN(CW_OUT_2) );
  NOR3_X1 U33 ( .A1(n9), .A2(n36), .A3(n12), .ZN(CW_OUT_3) );
  NOR4_X1 U34 ( .A1(OPCODE_IN[3]), .A2(n9), .A3(n36), .A4(n12), .ZN(CW_OUT_1)
         );
  NOR2_X1 U35 ( .A1(n12), .A2(n35), .ZN(CW_OUT[8]) );
  OAI221_X1 U36 ( .B1(OPCODE_IN[2]), .B2(OPCODE_IN[1]), .C1(n28), .C2(n27), 
        .A(OPCODE_IN[3]), .ZN(n24) );
  OAI211_X1 U37 ( .C1(OPCODE_IN[1]), .C2(n12), .A(n29), .B(OPCODE_IN[2]), .ZN(
        n23) );
  OAI211_X1 U38 ( .C1(OPCODE_IN[4]), .C2(OPCODE_IN[0]), .A(OPCODE_IN[2]), .B(
        OPCODE_IN[1]), .ZN(n26) );
  NOR3_X1 U39 ( .A1(n14), .A2(n27), .A3(n12), .ZN(CW_OUT[7]) );
  NAND2_X1 U40 ( .A1(n22), .A2(n27), .ZN(n15) );
endmodule


module stall_logic_FUNC_SIZE11_OP_CODE_SIZE6 ( OPCODE_i, FUNC_i, rA_i, rB_i, 
        D1_i, D2_i, S_mem_LOAD_i, S_exe_LOAD_i, S_MUX_PC_BUS_i, mispredict_i, 
        bubble_dec_o, bubble_exe_o, stall_exe_o, stall_dec_o, stall_btb_o, 
        stall_fetch_o, S_exe_WRITE_i_BAR );
  input [5:0] OPCODE_i;
  input [10:0] FUNC_i;
  input [4:0] rA_i;
  input [4:0] rB_i;
  input [4:0] D1_i;
  input [4:0] D2_i;
  input [1:0] S_MUX_PC_BUS_i;
  input S_mem_LOAD_i, S_exe_LOAD_i, mispredict_i, S_exe_WRITE_i_BAR;
  output bubble_dec_o, bubble_exe_o, stall_exe_o, stall_dec_o, stall_btb_o,
         stall_fetch_o;
  wire   S_exe_WRITE_i, n16, n27, n28, n29, n30, n31, n32, n33, n34, n41, n43,
         n44, n45, n46, n47, n48, n50, n51, n52, n53, n54, n55, n56, n42, n49,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73;
  assign S_exe_WRITE_i = S_exe_WRITE_i_BAR;

  OAI22_X1 U38 ( .A1(n54), .A2(D1_i[2]), .B1(n55), .B2(D1_i[1]), .ZN(n56) );
  AOI221_X1 U37 ( .B1(n54), .B2(D1_i[2]), .C1(D1_i[1]), .C2(n55), .A(n56), 
        .ZN(n50) );
  OAI22_X1 U34 ( .A1(n44), .A2(D1_i[3]), .B1(n46), .B2(D1_i[4]), .ZN(n53) );
  AOI221_X1 U33 ( .B1(n44), .B2(D1_i[3]), .C1(D1_i[4]), .C2(n46), .A(n53), 
        .ZN(n51) );
  XNOR2_X1 U32 ( .A(rA_i[0]), .B(D1_i[0]), .ZN(n52) );
  OAI22_X1 U12 ( .A1(n33), .A2(rB_i[2]), .B1(n32), .B2(rB_i[1]), .ZN(n34) );
  AOI221_X1 U11 ( .B1(rB_i[1]), .B2(n32), .C1(n33), .C2(rB_i[2]), .A(n34), 
        .ZN(n27) );
  OAI22_X1 U8 ( .A1(n30), .A2(rB_i[3]), .B1(n29), .B2(rB_i[4]), .ZN(n31) );
  AOI221_X1 U7 ( .B1(rB_i[4]), .B2(n29), .C1(n30), .C2(rB_i[3]), .A(n31), .ZN(
        n28) );
  NOR2_X1 U2 ( .A1(stall_fetch_o), .A2(n16), .ZN(bubble_dec_o) );
  INV_X1 U40 ( .A(rA_i[2]), .ZN(n54) );
  INV_X1 U39 ( .A(rA_i[1]), .ZN(n55) );
  INV_X1 U36 ( .A(rA_i[3]), .ZN(n44) );
  INV_X1 U22 ( .A(D2_i[2]), .ZN(n43) );
  INV_X1 U9 ( .A(D1_i[3]), .ZN(n30) );
  INV_X1 U10 ( .A(D1_i[4]), .ZN(n29) );
  INV_X1 U13 ( .A(D1_i[2]), .ZN(n33) );
  INV_X1 U14 ( .A(D1_i[1]), .ZN(n32) );
  INV_X1 U35 ( .A(rA_i[4]), .ZN(n46) );
  INV_X1 U3 ( .A(S_exe_LOAD_i), .ZN(n42) );
  NOR2_X1 U4 ( .A1(OPCODE_i[4]), .A2(OPCODE_i[1]), .ZN(n49) );
  INV_X1 U5 ( .A(OPCODE_i[2]), .ZN(n57) );
  NAND2_X1 U6 ( .A1(OPCODE_i[4]), .A2(OPCODE_i[1]), .ZN(n58) );
  OAI221_X1 U15 ( .B1(n57), .B2(OPCODE_i[0]), .C1(n57), .C2(OPCODE_i[4]), .A(
        n58), .ZN(n59) );
  NOR4_X1 U16 ( .A1(n49), .A2(OPCODE_i[5]), .A3(OPCODE_i[3]), .A4(n59), .ZN(
        n60) );
  NAND3_X1 U17 ( .A1(n50), .A2(n52), .A3(n51), .ZN(n61) );
  INV_X1 U18 ( .A(n49), .ZN(n62) );
  AOI22_X1 U19 ( .A1(OPCODE_i[2]), .A2(n62), .B1(n58), .B2(n57), .ZN(n63) );
  INV_X1 U20 ( .A(rA_i[1]), .ZN(n64) );
  AOI22_X1 U21 ( .A1(n47), .A2(D2_i[0]), .B1(n46), .B2(D2_i[4]), .ZN(n65) );
  OAI21_X1 U23 ( .B1(n64), .B2(D2_i[1]), .A(n65), .ZN(n66) );
  AOI211_X1 U24 ( .C1(n64), .C2(D2_i[1]), .A(n48), .B(n66), .ZN(n67) );
  NAND3_X1 U25 ( .A1(n41), .A2(S_mem_LOAD_i), .A3(n67), .ZN(n68) );
  OAI21_X1 U26 ( .B1(S_exe_WRITE_i), .B2(n61), .A(n68), .ZN(n69) );
  XOR2_X1 U27 ( .A(D1_i[0]), .B(rB_i[0]), .Z(n70) );
  NAND4_X1 U28 ( .A1(S_exe_LOAD_i), .A2(n49), .A3(n28), .A4(n27), .ZN(n71) );
  NOR4_X1 U29 ( .A1(OPCODE_i[0]), .A2(OPCODE_i[2]), .A3(n70), .A4(n71), .ZN(
        n72) );
  AOI21_X1 U30 ( .B1(n63), .B2(n69), .A(n72), .ZN(n73) );
  OAI33_X1 U31 ( .A1(n42), .A2(n60), .A3(n61), .B1(OPCODE_i[5]), .B2(n73), 
        .B3(OPCODE_i[3]), .ZN(stall_fetch_o) );
  INV_X1 U41 ( .A(mispredict_i), .ZN(n16) );
  INV_X1 U42 ( .A(rA_i[0]), .ZN(n47) );
  AOI221_X1 U43 ( .B1(rA_i[2]), .B2(n43), .C1(n44), .C2(D2_i[3]), .A(n45), 
        .ZN(n41) );
  OAI22_X1 U44 ( .A1(n47), .A2(D2_i[0]), .B1(n46), .B2(D2_i[4]), .ZN(n48) );
  OAI22_X1 U45 ( .A1(n44), .A2(D2_i[3]), .B1(n43), .B2(rA_i[2]), .ZN(n45) );
endmodule


module mux41_MUX_SIZE32 ( IN0, IN1, IN2, IN3, CTRL, OUT1 );
  input [31:0] IN0;
  input [31:0] IN1;
  input [31:0] IN2;
  input [31:0] IN3;
  input [1:0] CTRL;
  output [31:0] OUT1;
  wire   n2, n3, n5, n6, n7, n8, n9, n10, n11, n12, n13, n16, n17, n18, n19,
         n20, n21, n24, n25, n28, n29, n30, n31, n34, n35, n36, n37, n44, n45,
         n46, n47, n60, n61, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126;

  NAND2_X1 U61 ( .A1(n46), .A2(n47), .ZN(OUT1[1]) );
  BUF_X1 U1 ( .A(n6), .Z(n71) );
  BUF_X1 U2 ( .A(n6), .Z(n73) );
  BUF_X2 U3 ( .A(n6), .Z(n72) );
  AND2_X2 U4 ( .A1(n70), .A2(CTRL[0]), .ZN(n6) );
  BUF_X1 U5 ( .A(n7), .Z(n119) );
  BUF_X2 U6 ( .A(n5), .Z(n125) );
  BUF_X2 U7 ( .A(n7), .Z(n121) );
  BUF_X2 U8 ( .A(n7), .Z(n120) );
  BUF_X2 U9 ( .A(n6), .Z(n123) );
  NOR2_X1 U10 ( .A1(CTRL[0]), .A2(n70), .ZN(n5) );
  NOR2_X1 U11 ( .A1(CTRL[0]), .A2(n118), .ZN(n7) );
  BUF_X2 U12 ( .A(n6), .Z(n122) );
  BUF_X2 U13 ( .A(n5), .Z(n126) );
  BUF_X2 U14 ( .A(n5), .Z(n124) );
  BUF_X1 U15 ( .A(CTRL[1]), .Z(n118) );
  NAND2_X1 U16 ( .A1(n126), .A2(IN2[28]), .ZN(n29) );
  NAND2_X1 U17 ( .A1(n125), .A2(IN2[24]), .ZN(n37) );
  NAND2_X1 U18 ( .A1(n126), .A2(IN2[20]), .ZN(n45) );
  NAND3_X1 U19 ( .A1(n75), .A2(n74), .A3(n76), .ZN(OUT1[12]) );
  NAND2_X1 U20 ( .A1(n6), .A2(IN1[12]), .ZN(n75) );
  NAND2_X1 U21 ( .A1(n119), .A2(IN0[12]), .ZN(n76) );
  NAND2_X1 U22 ( .A1(n125), .A2(IN2[12]), .ZN(n74) );
  NAND3_X1 U23 ( .A1(n79), .A2(n78), .A3(n77), .ZN(OUT1[29]) );
  NAND2_X1 U24 ( .A1(n123), .A2(IN1[29]), .ZN(n79) );
  NAND2_X1 U25 ( .A1(n120), .A2(IN0[29]), .ZN(n78) );
  NAND2_X1 U26 ( .A1(n125), .A2(IN2[29]), .ZN(n77) );
  NAND3_X1 U27 ( .A1(n82), .A2(n81), .A3(n80), .ZN(OUT1[26]) );
  NAND2_X1 U28 ( .A1(n72), .A2(IN1[26]), .ZN(n82) );
  NAND2_X1 U29 ( .A1(n120), .A2(IN0[26]), .ZN(n81) );
  NAND2_X1 U30 ( .A1(n126), .A2(IN2[26]), .ZN(n80) );
  NAND3_X1 U31 ( .A1(n84), .A2(n83), .A3(n85), .ZN(OUT1[14]) );
  NAND2_X1 U32 ( .A1(n72), .A2(IN1[14]), .ZN(n84) );
  NAND2_X1 U33 ( .A1(n119), .A2(IN0[14]), .ZN(n85) );
  NAND2_X1 U34 ( .A1(n124), .A2(IN2[14]), .ZN(n83) );
  NAND3_X1 U35 ( .A1(n88), .A2(n87), .A3(n86), .ZN(OUT1[18]) );
  NAND2_X1 U36 ( .A1(n123), .A2(IN1[18]), .ZN(n88) );
  NAND2_X1 U37 ( .A1(n120), .A2(IN0[18]), .ZN(n87) );
  NAND2_X1 U38 ( .A1(n124), .A2(IN2[18]), .ZN(n86) );
  AOI22_X1 U39 ( .A1(n120), .A2(IN0[5]), .B1(n73), .B2(IN1[5]), .ZN(n90) );
  NAND2_X1 U40 ( .A1(n90), .A2(n89), .ZN(OUT1[5]) );
  NAND2_X1 U41 ( .A1(n125), .A2(IN2[5]), .ZN(n89) );
  NAND3_X1 U42 ( .A1(n93), .A2(n92), .A3(n91), .ZN(OUT1[22]) );
  NAND2_X1 U43 ( .A1(n72), .A2(IN1[22]), .ZN(n93) );
  NAND2_X1 U44 ( .A1(n120), .A2(IN0[22]), .ZN(n92) );
  NAND2_X1 U45 ( .A1(n124), .A2(IN2[22]), .ZN(n91) );
  NAND3_X1 U46 ( .A1(n95), .A2(n94), .A3(n96), .ZN(OUT1[30]) );
  NAND2_X1 U47 ( .A1(n122), .A2(IN1[30]), .ZN(n95) );
  NAND2_X1 U48 ( .A1(n120), .A2(IN0[30]), .ZN(n96) );
  NAND2_X1 U49 ( .A1(n124), .A2(IN2[30]), .ZN(n94) );
  NAND3_X1 U50 ( .A1(n98), .A2(n97), .A3(n99), .ZN(OUT1[19]) );
  NAND2_X1 U51 ( .A1(n71), .A2(IN1[19]), .ZN(n98) );
  NAND2_X1 U52 ( .A1(n120), .A2(IN0[19]), .ZN(n99) );
  NAND2_X1 U53 ( .A1(n124), .A2(IN2[19]), .ZN(n97) );
  NAND3_X1 U54 ( .A1(n101), .A2(n100), .A3(n102), .ZN(OUT1[11]) );
  NAND2_X1 U55 ( .A1(n71), .A2(IN1[11]), .ZN(n101) );
  NAND2_X1 U56 ( .A1(n120), .A2(IN0[11]), .ZN(n102) );
  NAND2_X1 U57 ( .A1(n125), .A2(IN2[11]), .ZN(n100) );
  NAND3_X1 U58 ( .A1(n105), .A2(n104), .A3(n103), .ZN(OUT1[17]) );
  NAND2_X1 U59 ( .A1(n122), .A2(IN1[17]), .ZN(n105) );
  NAND2_X1 U60 ( .A1(n120), .A2(IN0[17]), .ZN(n104) );
  NAND2_X1 U62 ( .A1(n124), .A2(IN2[17]), .ZN(n103) );
  NAND3_X1 U63 ( .A1(n107), .A2(n106), .A3(n108), .ZN(OUT1[15]) );
  NAND2_X1 U64 ( .A1(n122), .A2(IN1[15]), .ZN(n107) );
  NAND2_X1 U65 ( .A1(n119), .A2(IN0[15]), .ZN(n108) );
  NAND2_X1 U66 ( .A1(n125), .A2(IN2[15]), .ZN(n106) );
  NAND3_X1 U67 ( .A1(n110), .A2(n109), .A3(n111), .ZN(OUT1[21]) );
  NAND2_X1 U68 ( .A1(n72), .A2(IN1[21]), .ZN(n110) );
  NAND2_X1 U69 ( .A1(n119), .A2(IN0[21]), .ZN(n111) );
  NAND2_X1 U70 ( .A1(n124), .A2(IN2[21]), .ZN(n109) );
  NAND3_X1 U71 ( .A1(n114), .A2(n113), .A3(n112), .ZN(OUT1[23]) );
  NAND2_X1 U72 ( .A1(n123), .A2(IN1[23]), .ZN(n114) );
  NAND2_X1 U73 ( .A1(n119), .A2(IN0[23]), .ZN(n113) );
  NAND2_X1 U74 ( .A1(n125), .A2(IN2[23]), .ZN(n112) );
  NAND3_X1 U75 ( .A1(n117), .A2(n116), .A3(n115), .ZN(OUT1[16]) );
  NAND2_X1 U76 ( .A1(n122), .A2(IN1[16]), .ZN(n117) );
  NAND2_X1 U77 ( .A1(n120), .A2(IN0[16]), .ZN(n116) );
  NAND2_X1 U78 ( .A1(n126), .A2(IN2[16]), .ZN(n115) );
  NAND2_X1 U79 ( .A1(n66), .A2(n67), .ZN(OUT1[10]) );
  NAND2_X1 U80 ( .A1(n60), .A2(n61), .ZN(OUT1[13]) );
  AOI22_X1 U81 ( .A1(n71), .A2(IN1[9]), .B1(n121), .B2(IN0[9]), .ZN(n2) );
  AOI22_X1 U82 ( .A1(n123), .A2(IN1[4]), .B1(n121), .B2(IN0[4]), .ZN(n16) );
  AOI22_X1 U83 ( .A1(n73), .A2(IN1[8]), .B1(n121), .B2(IN0[8]), .ZN(n8) );
  AOI22_X1 U84 ( .A1(n123), .A2(IN1[3]), .B1(n120), .B2(IN0[3]), .ZN(n18) );
  AOI22_X1 U85 ( .A1(n72), .A2(IN1[7]), .B1(n119), .B2(IN0[7]), .ZN(n10) );
  NAND2_X1 U86 ( .A1(n68), .A2(n69), .ZN(OUT1[0]) );
  NAND2_X1 U87 ( .A1(n126), .A2(IN2[27]), .ZN(n31) );
  NAND2_X1 U88 ( .A1(n126), .A2(IN2[2]), .ZN(n25) );
  NAND2_X1 U89 ( .A1(n126), .A2(IN2[25]), .ZN(n35) );
  NAND2_X1 U90 ( .A1(n12), .A2(n13), .ZN(OUT1[6]) );
  NAND2_X1 U91 ( .A1(n2), .A2(n3), .ZN(OUT1[9]) );
  AOI22_X1 U92 ( .A1(n123), .A2(IN1[27]), .B1(n121), .B2(IN0[27]), .ZN(n30) );
  AOI22_X1 U93 ( .A1(n122), .A2(IN1[2]), .B1(n120), .B2(IN0[2]), .ZN(n24) );
  AOI22_X1 U94 ( .A1(n123), .A2(IN1[25]), .B1(n121), .B2(IN0[25]), .ZN(n34) );
  AOI22_X1 U95 ( .A1(n73), .A2(IN1[28]), .B1(n121), .B2(IN0[28]), .ZN(n28) );
  AOI22_X1 U96 ( .A1(n72), .A2(IN1[20]), .B1(n121), .B2(IN0[20]), .ZN(n44) );
  AOI22_X1 U97 ( .A1(n72), .A2(IN1[24]), .B1(n121), .B2(IN0[24]), .ZN(n36) );
  NAND2_X1 U98 ( .A1(n30), .A2(n31), .ZN(OUT1[27]) );
  NAND2_X1 U99 ( .A1(n125), .A2(IN2[1]), .ZN(n47) );
  NAND2_X1 U100 ( .A1(n125), .A2(IN2[10]), .ZN(n67) );
  AOI22_X1 U101 ( .A1(n122), .A2(IN1[6]), .B1(n121), .B2(IN0[6]), .ZN(n12) );
  NAND2_X1 U102 ( .A1(n10), .A2(n11), .ZN(OUT1[7]) );
  NAND2_X1 U103 ( .A1(n8), .A2(n9), .ZN(OUT1[8]) );
  AOI22_X1 U104 ( .A1(n71), .A2(IN1[1]), .B1(n119), .B2(IN0[1]), .ZN(n46) );
  AOI22_X1 U105 ( .A1(n71), .A2(IN1[10]), .B1(n121), .B2(IN0[10]), .ZN(n66) );
  AOI22_X1 U106 ( .A1(n71), .A2(IN1[0]), .B1(n119), .B2(IN0[0]), .ZN(n68) );
  AOI22_X1 U107 ( .A1(n122), .A2(IN1[13]), .B1(n120), .B2(IN0[13]), .ZN(n60)
         );
  AOI22_X1 U108 ( .A1(n73), .A2(IN1[31]), .B1(n121), .B2(IN0[31]), .ZN(n20) );
  NAND2_X1 U109 ( .A1(n125), .A2(IN2[31]), .ZN(n21) );
  NAND2_X1 U110 ( .A1(n18), .A2(n19), .ZN(OUT1[3]) );
  NAND2_X1 U111 ( .A1(n34), .A2(n35), .ZN(OUT1[25]) );
  NAND2_X1 U112 ( .A1(n20), .A2(n21), .ZN(OUT1[31]) );
  NAND2_X1 U113 ( .A1(n16), .A2(n17), .ZN(OUT1[4]) );
  NAND2_X1 U114 ( .A1(n28), .A2(n29), .ZN(OUT1[28]) );
  NAND2_X1 U115 ( .A1(n24), .A2(n25), .ZN(OUT1[2]) );
  NAND2_X1 U116 ( .A1(n36), .A2(n37), .ZN(OUT1[24]) );
  NAND2_X1 U117 ( .A1(n44), .A2(n45), .ZN(OUT1[20]) );
  NAND2_X1 U118 ( .A1(n125), .A2(IN2[9]), .ZN(n3) );
  NAND2_X1 U119 ( .A1(n125), .A2(IN2[4]), .ZN(n17) );
  NAND2_X1 U120 ( .A1(n126), .A2(IN2[8]), .ZN(n9) );
  NAND2_X1 U121 ( .A1(n126), .A2(IN2[3]), .ZN(n19) );
  NAND2_X1 U122 ( .A1(n126), .A2(IN2[7]), .ZN(n11) );
  NAND2_X1 U123 ( .A1(n126), .A2(IN2[6]), .ZN(n13) );
  NAND2_X1 U124 ( .A1(n126), .A2(IN2[0]), .ZN(n69) );
  NAND2_X1 U125 ( .A1(n126), .A2(IN2[13]), .ZN(n61) );
  INV_X1 U126 ( .A(CTRL[1]), .ZN(n70) );
endmodule


module zerocheck ( IN0, CTRL, OUT1 );
  input [31:0] IN0;
  input CTRL;
  output OUT1;
  wire   n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42;

  INV_X1 U1 ( .A(IN0[7]), .ZN(n32) );
  INV_X1 U2 ( .A(IN0[13]), .ZN(n28) );
  INV_X1 U3 ( .A(IN0[12]), .ZN(n21) );
  INV_X1 U4 ( .A(IN0[1]), .ZN(n20) );
  NOR2_X1 U5 ( .A1(n25), .A2(n26), .ZN(n15) );
  AND3_X1 U6 ( .A1(n14), .A2(n16), .A3(n15), .ZN(n42) );
  XNOR2_X1 U7 ( .A(n42), .B(CTRL), .ZN(OUT1) );
  INV_X1 U8 ( .A(IN0[3]), .ZN(n31) );
  INV_X1 U9 ( .A(IN0[0]), .ZN(n29) );
  NAND3_X1 U10 ( .A1(n19), .A2(n20), .A3(n21), .ZN(n18) );
  NAND3_X1 U11 ( .A1(n23), .A2(n24), .A3(n22), .ZN(n17) );
  NAND3_X1 U12 ( .A1(n27), .A2(n28), .A3(n29), .ZN(n26) );
  NAND3_X1 U13 ( .A1(n30), .A2(n31), .A3(n32), .ZN(n25) );
  NAND3_X1 U14 ( .A1(n35), .A2(n36), .A3(n37), .ZN(n34) );
  NOR2_X1 U15 ( .A1(IN0[31]), .A2(IN0[14]), .ZN(n38) );
  NAND4_X1 U16 ( .A1(n38), .A2(n39), .A3(n40), .A4(n41), .ZN(n33) );
  NOR2_X1 U17 ( .A1(IN0[18]), .A2(IN0[19]), .ZN(n39) );
  NOR2_X1 U18 ( .A1(IN0[22]), .A2(IN0[17]), .ZN(n40) );
  NOR2_X1 U19 ( .A1(IN0[30]), .A2(IN0[21]), .ZN(n41) );
  NOR2_X1 U20 ( .A1(IN0[20]), .A2(IN0[15]), .ZN(n35) );
  NOR2_X1 U21 ( .A1(IN0[27]), .A2(IN0[29]), .ZN(n36) );
  NOR2_X1 U22 ( .A1(IN0[25]), .A2(IN0[26]), .ZN(n37) );
  NOR2_X1 U23 ( .A1(IN0[11]), .A2(IN0[23]), .ZN(n19) );
  NOR2_X1 U24 ( .A1(IN0[5]), .A2(IN0[16]), .ZN(n27) );
  NOR2_X1 U25 ( .A1(IN0[10]), .A2(IN0[6]), .ZN(n30) );
  NOR2_X1 U26 ( .A1(IN0[24]), .A2(IN0[28]), .ZN(n22) );
  NOR2_X1 U27 ( .A1(IN0[4]), .A2(IN0[9]), .ZN(n23) );
  NOR2_X1 U28 ( .A1(IN0[2]), .A2(IN0[8]), .ZN(n24) );
  NOR2_X1 U29 ( .A1(n17), .A2(n18), .ZN(n16) );
  NOR2_X1 U30 ( .A1(n33), .A2(n34), .ZN(n14) );
endmodule


module mux21_2 ( IN0, IN1, CTRL, OUT1 );
  input [31:0] IN0;
  input [31:0] IN1;
  output [31:0] OUT1;
  input CTRL;
  wire   n1, n2, n3, n4, n5, n6, n7, n8;

  MUX2_X1 U1 ( .A(IN0[9]), .B(IN1[9]), .S(n8), .Z(OUT1[9]) );
  MUX2_X1 U3 ( .A(IN0[7]), .B(IN1[7]), .S(n8), .Z(OUT1[7]) );
  MUX2_X1 U5 ( .A(IN0[5]), .B(IN1[5]), .S(n8), .Z(OUT1[5]) );
  MUX2_X1 U10 ( .A(IN0[2]), .B(IN1[2]), .S(n3), .Z(OUT1[2]) );
  MUX2_X1 U17 ( .A(IN0[23]), .B(IN1[23]), .S(n3), .Z(OUT1[23]) );
  MUX2_X1 U20 ( .A(IN0[20]), .B(IN1[20]), .S(n7), .Z(OUT1[20]) );
  MUX2_X1 U22 ( .A(IN0[19]), .B(IN1[19]), .S(n7), .Z(OUT1[19]) );
  MUX2_X1 U23 ( .A(IN0[18]), .B(IN1[18]), .S(n8), .Z(OUT1[18]) );
  MUX2_X1 U24 ( .A(IN0[17]), .B(IN1[17]), .S(n7), .Z(OUT1[17]) );
  MUX2_X1 U25 ( .A(IN0[16]), .B(IN1[16]), .S(n7), .Z(OUT1[16]) );
  MUX2_X1 U26 ( .A(IN0[15]), .B(IN1[15]), .S(n8), .Z(OUT1[15]) );
  MUX2_X1 U28 ( .A(IN0[13]), .B(IN1[13]), .S(n3), .Z(OUT1[13]) );
  MUX2_X1 U29 ( .A(IN0[12]), .B(IN1[12]), .S(n3), .Z(OUT1[12]) );
  MUX2_X1 U14 ( .A(IN0[26]), .B(IN1[26]), .S(n7), .Z(OUT1[26]) );
  MUX2_X1 U4 ( .A(IN0[6]), .B(IN1[6]), .S(n3), .Z(OUT1[6]) );
  MUX2_X1 U6 ( .A(IN0[4]), .B(IN1[4]), .S(n3), .Z(OUT1[4]) );
  MUX2_X1 U7 ( .A(IN0[3]), .B(IN1[3]), .S(n7), .Z(OUT1[3]) );
  MUX2_X1 U9 ( .A(IN0[30]), .B(IN1[30]), .S(n7), .Z(OUT1[30]) );
  MUX2_X1 U32 ( .A(IN0[0]), .B(IN1[0]), .S(n3), .Z(OUT1[0]) );
  MUX2_X1 U13 ( .A(IN0[27]), .B(IN1[27]), .S(n3), .Z(OUT1[27]) );
  MUX2_X1 U19 ( .A(IN0[21]), .B(IN1[21]), .S(n3), .Z(OUT1[21]) );
  MUX2_X1 U21 ( .A(IN0[1]), .B(IN1[1]), .S(n7), .Z(OUT1[1]) );
  MUX2_X1 U16 ( .A(IN0[24]), .B(IN1[24]), .S(n7), .Z(OUT1[24]) );
  MUX2_X1 U30 ( .A(IN0[11]), .B(IN1[11]), .S(n8), .Z(OUT1[11]) );
  MUX2_X1 U2 ( .A(IN0[10]), .B(IN1[10]), .S(n7), .Z(OUT1[10]) );
  MUX2_X1 U8 ( .A(IN0[8]), .B(IN1[8]), .S(n7), .Z(OUT1[8]) );
  MUX2_X1 U11 ( .A(IN0[14]), .B(IN1[14]), .S(n7), .Z(OUT1[14]) );
  MUX2_X1 U12 ( .A(IN0[25]), .B(IN1[25]), .S(n3), .Z(OUT1[25]) );
  MUX2_X1 U15 ( .A(IN0[22]), .B(IN1[22]), .S(n7), .Z(OUT1[22]) );
  CLKBUF_X2 U18 ( .A(CTRL), .Z(n8) );
  CLKBUF_X3 U27 ( .A(CTRL), .Z(n3) );
  CLKBUF_X3 U31 ( .A(CTRL), .Z(n7) );
  INV_X1 U33 ( .A(n7), .ZN(n4) );
  NAND2_X1 U34 ( .A1(n3), .A2(IN1[31]), .ZN(n2) );
  NAND2_X1 U35 ( .A1(IN0[31]), .A2(n4), .ZN(n1) );
  NAND2_X1 U36 ( .A1(n1), .A2(n2), .ZN(OUT1[31]) );
  NAND2_X1 U37 ( .A1(IN1[28]), .A2(n3), .ZN(n6) );
  NAND2_X1 U38 ( .A1(IN0[28]), .A2(n4), .ZN(n5) );
  NAND2_X1 U39 ( .A1(n5), .A2(n6), .ZN(OUT1[28]) );
  MUX2_X1 U40 ( .A(IN0[29]), .B(IN1[29]), .S(n3), .Z(OUT1[29]) );
endmodule


module p4add_N32_logN5_0 ( A, B, Cin, sign, S, Cout );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input Cin, sign;
  output Cout;
  wire   n1, n2, n3, n5, n6, n8, n10, n11, n12, n14, n15, n16, n17, n19, n22,
         n23, n24, n25, n27;
  wire   [31:0] new_B;
  wire   [7:0] carry_pro;
  wire   SYNOPSYS_UNCONNECTED__0;

  xor_gen_N32_0 xor32 ( .A(B), .B(1'b0), .S({new_B[31:27], n1, n14, 
        new_B[24:20], n27, n8, n22, new_B[16], n3, n16, n6, new_B[12], n2, n17, 
        n15, n5, n25, new_B[6], n19, n23, n12, n11, n24, n10}) );
  carry_tree_N32_logN5_0 ct ( .A({1'b0, 1'b0, 1'b0, 1'b0, A[27:0]}), .B({1'b0, 
        1'b0, 1'b0, 1'b0, new_B[27], n1, n14, new_B[24:20], n27, n8, n22, 
        new_B[16], n3, n16, n6, new_B[12], n2, n17, n15, n5, n25, new_B[6], 
        n19, n23, n12, n11, n24, n10}), .Cin(1'b0), .Cout({
        SYNOPSYS_UNCONNECTED__0, carry_pro[7:1]}) );
  sum_gen_N32_0 add ( .A(A), .B({new_B[31:27], n1, n14, new_B[24:20], n27, n8, 
        n22, new_B[16], n3, n16, n6, new_B[12], n2, n17, n15, n5, n25, 
        new_B[6], n19, n23, n12, n11, n24, n10}), .Cin({1'b0, carry_pro[7:1], 
        1'b0}), .S(S) );
endmodule


module extender_32 ( IN1, CTRL, SIGN, OUT1 );
  input [31:0] IN1;
  output [31:0] OUT1;
  input CTRL, SIGN;
  wire   OUT1_25, n2, n3, n4, n5, n7, n8, n9, n10, n12, n11, n13, n14, n15,
         n16, \OUT1[28] , \OUT1[27] , \OUT1[26] ;
  assign OUT1[15] = IN1[15];
  assign OUT1[14] = IN1[14];
  assign OUT1[13] = IN1[13];
  assign OUT1[12] = IN1[12];
  assign OUT1[11] = IN1[11];
  assign OUT1[10] = IN1[10];
  assign OUT1[9] = IN1[9];
  assign OUT1[8] = IN1[8];
  assign OUT1[7] = IN1[7];
  assign OUT1[6] = IN1[6];
  assign OUT1[5] = IN1[5];
  assign OUT1[4] = IN1[4];
  assign OUT1[3] = IN1[3];
  assign OUT1[2] = IN1[2];
  assign OUT1[1] = IN1[1];
  assign OUT1[0] = IN1[0];
  assign OUT1[30] = \OUT1[28] ;
  assign OUT1[29] = \OUT1[28] ;
  assign OUT1[28] = \OUT1[28] ;
  assign OUT1[25] = \OUT1[27] ;
  assign OUT1[27] = \OUT1[27] ;
  assign OUT1[31] = \OUT1[26] ;
  assign OUT1[26] = \OUT1[26] ;

  BUF_X2 U2 ( .A(OUT1_25), .Z(\OUT1[28] ) );
  NAND2_X1 U3 ( .A1(IN1[22]), .A2(CTRL), .ZN(n14) );
  NAND2_X1 U4 ( .A1(n15), .A2(n14), .ZN(OUT1[22]) );
  INV_X1 U5 ( .A(CTRL), .ZN(n13) );
  NAND3_X1 U6 ( .A1(SIGN), .A2(IN1[15]), .A3(n13), .ZN(n16) );
  NAND3_X1 U7 ( .A1(SIGN), .A2(IN1[15]), .A3(n13), .ZN(n15) );
  NAND3_X1 U8 ( .A1(SIGN), .A2(IN1[15]), .A3(n13), .ZN(n2) );
  NAND2_X1 U9 ( .A1(n2), .A2(n10), .ZN(OUT1[18]) );
  NAND2_X1 U10 ( .A1(n2), .A2(n11), .ZN(OUT1[17]) );
  NAND2_X1 U11 ( .A1(n2), .A2(n3), .ZN(OUT1_25) );
  BUF_X2 U12 ( .A(OUT1_25), .Z(\OUT1[27] ) );
  CLKBUF_X2 U13 ( .A(OUT1_25), .Z(\OUT1[26] ) );
  NAND2_X1 U14 ( .A1(n16), .A2(n7), .ZN(OUT1[21]) );
  NAND2_X1 U15 ( .A1(CTRL), .A2(IN1[17]), .ZN(n11) );
  NAND2_X1 U16 ( .A1(CTRL), .A2(IN1[24]), .ZN(n4) );
  NAND2_X1 U17 ( .A1(CTRL), .A2(IN1[20]), .ZN(n8) );
  NAND2_X1 U18 ( .A1(CTRL), .A2(IN1[16]), .ZN(n12) );
  NAND2_X1 U19 ( .A1(CTRL), .A2(IN1[23]), .ZN(n5) );
  NAND2_X1 U20 ( .A1(CTRL), .A2(IN1[19]), .ZN(n9) );
  NAND2_X1 U21 ( .A1(CTRL), .A2(IN1[21]), .ZN(n7) );
  NAND2_X1 U22 ( .A1(CTRL), .A2(IN1[18]), .ZN(n10) );
  NAND2_X1 U23 ( .A1(CTRL), .A2(IN1[25]), .ZN(n3) );
  NAND2_X1 U24 ( .A1(n15), .A2(n4), .ZN(OUT1[24]) );
  NAND2_X1 U25 ( .A1(n15), .A2(n8), .ZN(OUT1[20]) );
  NAND2_X1 U26 ( .A1(n15), .A2(n5), .ZN(OUT1[23]) );
  NAND2_X1 U27 ( .A1(n16), .A2(n9), .ZN(OUT1[19]) );
  NAND2_X1 U28 ( .A1(n16), .A2(n12), .ZN(OUT1[16]) );
endmodule


module ff32_en_IR ( D, en, clk, rst, Q );
  input [31:0] D;
  output [31:0] Q;
  input en, clk, rst;
  wire   n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n97, net644967, net644968, net644969, net644970,
         net644971, net644972, net644973, net644974, net644975, net644976,
         net644977, net644978, net644979, net644980, net644981, net644982,
         net644983, net644984, net644985, net644986, net644987, net644988,
         net644989, net644990, net644991, net644992, net644993, net644994,
         net644995, net644996, net644997, net644998, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35;

  DFFR_X1 \Q_reg[24]  ( .D(n89), .CK(clk), .RN(n35), .Q(Q[24]), .QN(net644991)
         );
  DFFR_X1 \Q_reg[23]  ( .D(n88), .CK(clk), .RN(n35), .Q(Q[23]), .QN(net644990)
         );
  DFFR_X1 \Q_reg[22]  ( .D(n87), .CK(clk), .RN(n35), .Q(Q[22]), .QN(net644989)
         );
  DFFR_X1 \Q_reg[20]  ( .D(n85), .CK(clk), .RN(n35), .Q(Q[20]), .QN(net644987)
         );
  DFFR_X1 \Q_reg[19]  ( .D(n84), .CK(clk), .RN(n35), .Q(Q[19]), .QN(net644986)
         );
  DFFR_X1 \Q_reg[18]  ( .D(n83), .CK(clk), .RN(n35), .Q(Q[18]), .QN(net644985)
         );
  DFFR_X1 \Q_reg[17]  ( .D(n82), .CK(clk), .RN(n35), .Q(Q[17]), .QN(net644984)
         );
  DFFR_X1 \Q_reg[16]  ( .D(n81), .CK(clk), .RN(n35), .Q(Q[16]), .QN(net644983)
         );
  DFFR_X1 \Q_reg[15]  ( .D(n80), .CK(clk), .RN(n35), .Q(Q[15]), .QN(net644982)
         );
  DFFR_X1 \Q_reg[14]  ( .D(n79), .CK(clk), .RN(n35), .Q(Q[14]), .QN(net644981)
         );
  DFFR_X1 \Q_reg[13]  ( .D(n78), .CK(clk), .RN(n35), .Q(Q[13]), .QN(net644980)
         );
  DFFR_X1 \Q_reg[12]  ( .D(n77), .CK(clk), .RN(n35), .Q(Q[12]), .QN(net644979)
         );
  DFFR_X1 \Q_reg[11]  ( .D(n76), .CK(clk), .RN(n35), .Q(Q[11]), .QN(net644978)
         );
  DFFR_X1 \Q_reg[10]  ( .D(n75), .CK(clk), .RN(n35), .Q(Q[10]), .QN(net644977)
         );
  DFFR_X1 \Q_reg[9]  ( .D(n74), .CK(clk), .RN(n35), .Q(Q[9]), .QN(net644976)
         );
  DFFR_X1 \Q_reg[8]  ( .D(n73), .CK(clk), .RN(n35), .Q(Q[8]), .QN(net644975)
         );
  DFFR_X1 \Q_reg[7]  ( .D(n72), .CK(clk), .RN(n35), .Q(Q[7]), .QN(net644974)
         );
  DFFR_X1 \Q_reg[6]  ( .D(n71), .CK(clk), .RN(n35), .Q(Q[6]), .QN(net644973)
         );
  DFFR_X1 \Q_reg[5]  ( .D(n70), .CK(clk), .RN(n35), .Q(Q[5]), .QN(net644972)
         );
  DFFR_X1 \Q_reg[4]  ( .D(n69), .CK(clk), .RN(n35), .Q(Q[4]), .QN(net644971)
         );
  DFFR_X1 \Q_reg[3]  ( .D(n68), .CK(clk), .RN(n35), .Q(Q[3]), .QN(net644970)
         );
  DFFR_X1 \Q_reg[2]  ( .D(n67), .CK(clk), .RN(n35), .Q(Q[2]), .QN(net644969)
         );
  DFFR_X1 \Q_reg[1]  ( .D(n66), .CK(clk), .RN(n35), .Q(Q[1]), .QN(net644968)
         );
  DFFR_X1 \Q_reg[0]  ( .D(n65), .CK(clk), .RN(n35), .Q(Q[0]), .QN(net644967)
         );
  DFFR_X2 \Q_reg[31]  ( .D(n97), .CK(clk), .RN(n35), .Q(Q[31]), .QN(net644998)
         );
  NAND2_X1 U6 ( .A1(en), .A2(D[30]), .ZN(n3) );
  OAI21_X1 U5 ( .B1(en), .B2(net644997), .A(n3), .ZN(n95) );
  NAND2_X1 U3 ( .A1(en), .A2(D[31]), .ZN(n2) );
  OAI21_X1 U2 ( .B1(en), .B2(net644998), .A(n2), .ZN(n97) );
  NAND2_X1 U48 ( .A1(en), .A2(D[9]), .ZN(n24) );
  OAI21_X1 U47 ( .B1(en), .B2(net644976), .A(n24), .ZN(n74) );
  NAND2_X1 U52 ( .A1(en), .A2(D[7]), .ZN(n26) );
  OAI21_X1 U51 ( .B1(en), .B2(net644974), .A(n26), .ZN(n72) );
  NAND2_X1 U34 ( .A1(en), .A2(D[16]), .ZN(n17) );
  OAI21_X1 U33 ( .B1(en), .B2(net644983), .A(n17), .ZN(n81) );
  NAND2_X1 U64 ( .A1(en), .A2(D[1]), .ZN(n32) );
  OAI21_X1 U63 ( .B1(n34), .B2(net644968), .A(n32), .ZN(n66) );
  NAND2_X1 U66 ( .A1(en), .A2(D[0]), .ZN(n33) );
  OAI21_X1 U65 ( .B1(en), .B2(net644967), .A(n33), .ZN(n65) );
  NAND2_X1 U50 ( .A1(en), .A2(D[8]), .ZN(n25) );
  OAI21_X1 U49 ( .B1(en), .B2(net644975), .A(n25), .ZN(n73) );
  NAND2_X1 U54 ( .A1(n34), .A2(D[6]), .ZN(n27) );
  OAI21_X1 U53 ( .B1(en), .B2(net644973), .A(n27), .ZN(n71) );
  NAND2_X1 U62 ( .A1(n34), .A2(D[2]), .ZN(n31) );
  OAI21_X1 U61 ( .B1(en), .B2(net644969), .A(n31), .ZN(n67) );
  NAND2_X1 U60 ( .A1(n34), .A2(D[3]), .ZN(n30) );
  OAI21_X1 U59 ( .B1(en), .B2(net644970), .A(n30), .ZN(n68) );
  NAND2_X1 U56 ( .A1(en), .A2(D[5]), .ZN(n28) );
  OAI21_X1 U55 ( .B1(en), .B2(net644972), .A(n28), .ZN(n70) );
  NAND2_X1 U16 ( .A1(n34), .A2(D[25]), .ZN(n8) );
  OAI21_X1 U15 ( .B1(en), .B2(net644992), .A(n8), .ZN(n90) );
  NAND2_X1 U24 ( .A1(n34), .A2(D[21]), .ZN(n12) );
  OAI21_X1 U23 ( .B1(en), .B2(net644988), .A(n12), .ZN(n86) );
  NAND2_X1 U18 ( .A1(n34), .A2(D[24]), .ZN(n9) );
  OAI21_X1 U17 ( .B1(en), .B2(net644991), .A(n9), .ZN(n89) );
  NAND2_X1 U20 ( .A1(n34), .A2(D[23]), .ZN(n10) );
  OAI21_X1 U19 ( .B1(en), .B2(net644990), .A(n10), .ZN(n88) );
  NAND2_X1 U8 ( .A1(n34), .A2(D[29]), .ZN(n4) );
  OAI21_X1 U7 ( .B1(en), .B2(net644996), .A(n4), .ZN(n94) );
  NAND2_X1 U14 ( .A1(n34), .A2(D[26]), .ZN(n7) );
  OAI21_X1 U13 ( .B1(en), .B2(net644993), .A(n7), .ZN(n91) );
  NAND2_X1 U58 ( .A1(n34), .A2(D[4]), .ZN(n29) );
  OAI21_X1 U57 ( .B1(n34), .B2(net644971), .A(n29), .ZN(n69) );
  NAND2_X1 U12 ( .A1(n34), .A2(D[27]), .ZN(n6) );
  NAND2_X1 U10 ( .A1(n34), .A2(D[28]), .ZN(n5) );
  NAND2_X1 U36 ( .A1(en), .A2(D[15]), .ZN(n18) );
  OAI21_X1 U35 ( .B1(n34), .B2(net644982), .A(n18), .ZN(n80) );
  NAND2_X1 U32 ( .A1(en), .A2(D[17]), .ZN(n16) );
  OAI21_X1 U31 ( .B1(n34), .B2(net644984), .A(n16), .ZN(n82) );
  NAND2_X1 U30 ( .A1(en), .A2(D[18]), .ZN(n15) );
  OAI21_X1 U29 ( .B1(en), .B2(net644985), .A(n15), .ZN(n83) );
  NAND2_X1 U26 ( .A1(en), .A2(D[20]), .ZN(n13) );
  OAI21_X1 U25 ( .B1(en), .B2(net644987), .A(n13), .ZN(n85) );
  NAND2_X1 U40 ( .A1(en), .A2(D[13]), .ZN(n20) );
  OAI21_X1 U39 ( .B1(en), .B2(net644980), .A(n20), .ZN(n78) );
  NAND2_X1 U38 ( .A1(en), .A2(D[14]), .ZN(n19) );
  OAI21_X1 U37 ( .B1(en), .B2(net644981), .A(n19), .ZN(n79) );
  NAND2_X1 U42 ( .A1(en), .A2(D[12]), .ZN(n21) );
  OAI21_X1 U41 ( .B1(en), .B2(net644979), .A(n21), .ZN(n77) );
  NAND2_X1 U22 ( .A1(en), .A2(D[22]), .ZN(n11) );
  OAI21_X1 U21 ( .B1(en), .B2(net644989), .A(n11), .ZN(n87) );
  NAND2_X1 U46 ( .A1(en), .A2(D[10]), .ZN(n23) );
  OAI21_X1 U45 ( .B1(en), .B2(net644977), .A(n23), .ZN(n75) );
  NAND2_X1 U28 ( .A1(en), .A2(D[19]), .ZN(n14) );
  OAI21_X1 U27 ( .B1(en), .B2(net644986), .A(n14), .ZN(n84) );
  NAND2_X1 U44 ( .A1(en), .A2(D[11]), .ZN(n22) );
  OAI21_X1 U43 ( .B1(en), .B2(net644978), .A(n22), .ZN(n76) );
  DFFR_X2 \Q_reg[21]  ( .D(n86), .CK(clk), .RN(n35), .Q(Q[21]), .QN(net644988)
         );
  DFFS_X1 \Q_reg[28]  ( .D(n93), .CK(clk), .SN(n35), .Q(Q[28]), .QN(net644995)
         );
  DFFS_X1 \Q_reg[26]  ( .D(n91), .CK(clk), .SN(n35), .Q(Q[26]), .QN(net644993)
         );
  DFFR_X1 \Q_reg[29]  ( .D(n94), .CK(clk), .RN(n35), .Q(Q[29]), .QN(net644996)
         );
  DFFR_X1 \Q_reg[27]  ( .D(n92), .CK(clk), .RN(n35), .Q(Q[27]), .QN(net644994)
         );
  DFFS_X2 \Q_reg[30]  ( .D(n95), .CK(clk), .SN(n35), .Q(Q[30]), .QN(net644997)
         );
  DFFR_X1 \Q_reg[25]  ( .D(n90), .CK(clk), .RN(n35), .Q(Q[25]), .QN(net644992)
         );
  INV_X2 U4 ( .A(rst), .ZN(n35) );
  BUF_X1 U9 ( .A(en), .Z(n34) );
  OAI21_X1 U11 ( .B1(en), .B2(net644994), .A(n6), .ZN(n92) );
  OAI21_X1 U67 ( .B1(en), .B2(net644995), .A(n5), .ZN(n93) );
endmodule


module ff32_en_1 ( D, en, clk, rst, Q );
  input [31:0] D;
  output [31:0] Q;
  input en, clk, rst;
  wire   n1, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, net645075, net645076, net645077, net645078, net645079,
         net645080, net645081, net645082, net645083, net645084, net645085,
         net645086, net645087, net645088, net645089, net645090, net645091,
         net645092, net645093, net645094, net645095, net645096, net645097,
         net645098, net645099, net645100, net645101, net645102, net645103,
         net645104, net645105, net645106, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68;

  DFFR_X1 \Q_reg[31]  ( .D(n1), .CK(clk), .RN(n68), .Q(Q[31]), .QN(net645106)
         );
  DFFR_X1 \Q_reg[30]  ( .D(n3), .CK(clk), .RN(n68), .Q(Q[30]), .QN(net645105)
         );
  DFFR_X1 \Q_reg[29]  ( .D(n4), .CK(clk), .RN(n68), .Q(Q[29]), .QN(net645104)
         );
  DFFR_X1 \Q_reg[28]  ( .D(n5), .CK(clk), .RN(n68), .Q(Q[28]), .QN(net645103)
         );
  DFFR_X1 \Q_reg[27]  ( .D(n6), .CK(clk), .RN(n68), .Q(Q[27]), .QN(net645102)
         );
  DFFR_X1 \Q_reg[26]  ( .D(n7), .CK(clk), .RN(n68), .Q(Q[26]), .QN(net645101)
         );
  DFFR_X1 \Q_reg[25]  ( .D(n8), .CK(clk), .RN(n68), .Q(Q[25]), .QN(net645100)
         );
  DFFR_X1 \Q_reg[24]  ( .D(n9), .CK(clk), .RN(n68), .Q(Q[24]), .QN(net645099)
         );
  DFFR_X1 \Q_reg[23]  ( .D(n10), .CK(clk), .RN(n68), .Q(Q[23]), .QN(net645098)
         );
  DFFR_X1 \Q_reg[22]  ( .D(n11), .CK(clk), .RN(n68), .Q(Q[22]), .QN(net645097)
         );
  DFFR_X1 \Q_reg[21]  ( .D(n12), .CK(clk), .RN(n68), .Q(Q[21]), .QN(net645096)
         );
  DFFR_X1 \Q_reg[20]  ( .D(n13), .CK(clk), .RN(n68), .Q(Q[20]), .QN(net645095)
         );
  DFFR_X1 \Q_reg[19]  ( .D(n14), .CK(clk), .RN(n68), .Q(Q[19]), .QN(net645094)
         );
  DFFR_X1 \Q_reg[18]  ( .D(n15), .CK(clk), .RN(n68), .Q(Q[18]), .QN(net645093)
         );
  DFFR_X1 \Q_reg[17]  ( .D(n16), .CK(clk), .RN(n68), .Q(Q[17]), .QN(net645092)
         );
  DFFR_X1 \Q_reg[16]  ( .D(n17), .CK(clk), .RN(n68), .Q(Q[16]), .QN(net645091)
         );
  DFFR_X1 \Q_reg[15]  ( .D(n18), .CK(clk), .RN(n68), .Q(Q[15]), .QN(net645090)
         );
  DFFR_X1 \Q_reg[14]  ( .D(n19), .CK(clk), .RN(n68), .Q(Q[14]), .QN(net645089)
         );
  DFFR_X1 \Q_reg[13]  ( .D(n20), .CK(clk), .RN(n68), .Q(Q[13]), .QN(net645088)
         );
  DFFR_X1 \Q_reg[12]  ( .D(n21), .CK(clk), .RN(n68), .Q(Q[12]), .QN(net645087)
         );
  DFFR_X1 \Q_reg[11]  ( .D(n22), .CK(clk), .RN(n68), .Q(Q[11]), .QN(net645086)
         );
  DFFR_X1 \Q_reg[10]  ( .D(n23), .CK(clk), .RN(n68), .Q(Q[10]), .QN(net645085)
         );
  DFFR_X1 \Q_reg[9]  ( .D(n24), .CK(clk), .RN(n68), .Q(Q[9]), .QN(net645084)
         );
  DFFR_X1 \Q_reg[8]  ( .D(n25), .CK(clk), .RN(n68), .Q(Q[8]), .QN(net645083)
         );
  DFFR_X1 \Q_reg[7]  ( .D(n26), .CK(clk), .RN(n68), .Q(Q[7]), .QN(net645082)
         );
  DFFR_X1 \Q_reg[6]  ( .D(n27), .CK(clk), .RN(n68), .Q(Q[6]), .QN(net645081)
         );
  DFFR_X1 \Q_reg[5]  ( .D(n28), .CK(clk), .RN(n68), .Q(Q[5]), .QN(net645080)
         );
  DFFR_X1 \Q_reg[4]  ( .D(n29), .CK(clk), .RN(n68), .Q(Q[4]), .QN(net645079)
         );
  DFFR_X1 \Q_reg[3]  ( .D(n30), .CK(clk), .RN(n68), .Q(Q[3]), .QN(net645078)
         );
  DFFR_X1 \Q_reg[2]  ( .D(n31), .CK(clk), .RN(n68), .Q(Q[2]), .QN(net645077)
         );
  DFFR_X1 \Q_reg[1]  ( .D(n32), .CK(clk), .RN(n68), .Q(Q[1]), .QN(net645076)
         );
  DFFR_X1 \Q_reg[0]  ( .D(n33), .CK(clk), .RN(n68), .Q(Q[0]), .QN(net645075)
         );
  NAND2_X1 U66 ( .A1(en), .A2(D[31]), .ZN(n66) );
  OAI21_X1 U65 ( .B1(en), .B2(net645106), .A(n66), .ZN(n1) );
  NAND2_X1 U23 ( .A1(n67), .A2(D[30]), .ZN(n45) );
  OAI21_X1 U22 ( .B1(en), .B2(net645105), .A(n45), .ZN(n3) );
  NAND2_X1 U13 ( .A1(en), .A2(D[29]), .ZN(n40) );
  OAI21_X1 U12 ( .B1(en), .B2(net645104), .A(n40), .ZN(n4) );
  NAND2_X1 U11 ( .A1(en), .A2(D[28]), .ZN(n39) );
  OAI21_X1 U10 ( .B1(en), .B2(net645103), .A(n39), .ZN(n5) );
  NAND2_X1 U9 ( .A1(n67), .A2(D[27]), .ZN(n38) );
  OAI21_X1 U8 ( .B1(en), .B2(net645102), .A(n38), .ZN(n6) );
  NAND2_X1 U7 ( .A1(en), .A2(D[26]), .ZN(n37) );
  OAI21_X1 U6 ( .B1(en), .B2(net645101), .A(n37), .ZN(n7) );
  NAND2_X1 U5 ( .A1(en), .A2(D[25]), .ZN(n36) );
  OAI21_X1 U4 ( .B1(en), .B2(net645100), .A(n36), .ZN(n8) );
  NAND2_X1 U19 ( .A1(en), .A2(D[2]), .ZN(n43) );
  OAI21_X1 U18 ( .B1(en), .B2(net645077), .A(n43), .ZN(n31) );
  NAND2_X1 U3 ( .A1(en), .A2(D[24]), .ZN(n35) );
  OAI21_X1 U2 ( .B1(en), .B2(net645099), .A(n35), .ZN(n9) );
  NAND2_X1 U62 ( .A1(en), .A2(D[22]), .ZN(n64) );
  OAI21_X1 U61 ( .B1(n67), .B2(net645097), .A(n64), .ZN(n11) );
  NAND2_X1 U64 ( .A1(en), .A2(D[23]), .ZN(n65) );
  OAI21_X1 U63 ( .B1(en), .B2(net645098), .A(n65), .ZN(n10) );
  NAND2_X1 U17 ( .A1(n67), .A2(D[1]), .ZN(n42) );
  OAI21_X1 U16 ( .B1(en), .B2(net645076), .A(n42), .ZN(n32) );
  NAND2_X1 U52 ( .A1(n67), .A2(D[17]), .ZN(n59) );
  OAI21_X1 U51 ( .B1(en), .B2(net645092), .A(n59), .ZN(n16) );
  NAND2_X1 U39 ( .A1(n67), .A2(D[11]), .ZN(n53) );
  OAI21_X1 U38 ( .B1(en), .B2(net645086), .A(n53), .ZN(n22) );
  NAND2_X1 U41 ( .A1(n67), .A2(D[12]), .ZN(n54) );
  OAI21_X1 U40 ( .B1(en), .B2(net645087), .A(n54), .ZN(n21) );
  NAND2_X1 U35 ( .A1(n67), .A2(D[9]), .ZN(n51) );
  OAI21_X1 U34 ( .B1(en), .B2(net645084), .A(n51), .ZN(n24) );
  NAND2_X1 U31 ( .A1(n67), .A2(D[7]), .ZN(n49) );
  OAI21_X1 U30 ( .B1(en), .B2(net645082), .A(n49), .ZN(n26) );
  NAND2_X1 U33 ( .A1(n67), .A2(D[8]), .ZN(n50) );
  OAI21_X1 U32 ( .B1(en), .B2(net645083), .A(n50), .ZN(n25) );
  NAND2_X1 U48 ( .A1(n67), .A2(D[15]), .ZN(n57) );
  OAI21_X1 U47 ( .B1(en), .B2(net645090), .A(n57), .ZN(n18) );
  NAND2_X1 U25 ( .A1(n67), .A2(D[4]), .ZN(n46) );
  OAI21_X1 U24 ( .B1(en), .B2(net645079), .A(n46), .ZN(n29) );
  NAND2_X1 U43 ( .A1(n67), .A2(D[13]), .ZN(n55) );
  OAI21_X1 U42 ( .B1(en), .B2(net645088), .A(n55), .ZN(n20) );
  NAND2_X1 U29 ( .A1(n67), .A2(D[6]), .ZN(n48) );
  OAI21_X1 U28 ( .B1(en), .B2(net645081), .A(n48), .ZN(n27) );
  NAND2_X1 U37 ( .A1(n67), .A2(D[10]), .ZN(n52) );
  OAI21_X1 U36 ( .B1(en), .B2(net645085), .A(n52), .ZN(n23) );
  NAND2_X1 U21 ( .A1(n67), .A2(D[3]), .ZN(n44) );
  OAI21_X1 U20 ( .B1(en), .B2(net645078), .A(n44), .ZN(n30) );
  NAND2_X1 U46 ( .A1(n67), .A2(D[14]), .ZN(n56) );
  OAI21_X1 U45 ( .B1(en), .B2(net645089), .A(n56), .ZN(n19) );
  NAND2_X1 U27 ( .A1(n67), .A2(D[5]), .ZN(n47) );
  OAI21_X1 U26 ( .B1(en), .B2(net645080), .A(n47), .ZN(n28) );
  NAND2_X1 U50 ( .A1(n67), .A2(D[16]), .ZN(n58) );
  OAI21_X1 U49 ( .B1(n67), .B2(net645091), .A(n58), .ZN(n17) );
  NAND2_X1 U58 ( .A1(n67), .A2(D[20]), .ZN(n62) );
  OAI21_X1 U57 ( .B1(n67), .B2(net645095), .A(n62), .ZN(n13) );
  NAND2_X1 U54 ( .A1(n67), .A2(D[18]), .ZN(n60) );
  OAI21_X1 U53 ( .B1(n67), .B2(net645093), .A(n60), .ZN(n15) );
  NAND2_X1 U60 ( .A1(n67), .A2(D[21]), .ZN(n63) );
  OAI21_X1 U59 ( .B1(n67), .B2(net645096), .A(n63), .ZN(n12) );
  NAND2_X1 U56 ( .A1(n67), .A2(D[19]), .ZN(n61) );
  OAI21_X1 U55 ( .B1(en), .B2(net645094), .A(n61), .ZN(n14) );
  NAND2_X1 U15 ( .A1(en), .A2(D[0]), .ZN(n41) );
  OAI21_X1 U14 ( .B1(en), .B2(net645075), .A(n41), .ZN(n33) );
  INV_X2 U44 ( .A(rst), .ZN(n68) );
  BUF_X2 U67 ( .A(en), .Z(n67) );
endmodule


module predictor_2_15 ( clock, reset, enable, taken_i, prediction_o );
  input clock, reset, enable, taken_i;
  output prediction_o;
  wire   N11, N12, n5, n6, n8, n9, n11, n10, n12;
  wire   [1:0] next_STATE;

  DLH_X1 \next_STATE_reg[0]  ( .G(enable), .D(N11), .Q(next_STATE[0]) );
  DFFR_X1 \STATE_reg[0]  ( .D(n6), .CK(clock), .RN(n12), .Q(n5), .QN(n10) );
  DLH_X1 \next_STATE_reg[1]  ( .G(enable), .D(N12), .Q(next_STATE[1]) );
  DFFR_X1 \STATE_reg[1]  ( .D(n8), .CK(clock), .RN(n12), .Q(prediction_o) );
  MUX2_X1 U8 ( .A(prediction_o), .B(next_STATE[1]), .S(enable), .Z(n8) );
  MUX2_X1 U9 ( .A(n5), .B(next_STATE[0]), .S(enable), .Z(n6) );
  NOR2_X1 U7 ( .A1(prediction_o), .A2(taken_i), .ZN(n9) );
  NAND2_X1 U6 ( .A1(prediction_o), .A2(taken_i), .ZN(n11) );
  OAI21_X1 U3 ( .B1(n9), .B2(n10), .A(n11), .ZN(N12) );
  OAI21_X1 U5 ( .B1(n5), .B2(n9), .A(n11), .ZN(N11) );
  INV_X1 U2 ( .A(reset), .ZN(n12) );
endmodule


module predictor_2_0 ( clock, reset, enable, taken_i, prediction_o );
  input clock, reset, enable, taken_i;
  output prediction_o;
  wire   N11, N12, n9, n11, n5, n6, n8, n7, n10;
  wire   [1:0] next_STATE;

  DLH_X1 \next_STATE_reg[0]  ( .G(enable), .D(N11), .Q(next_STATE[0]) );
  DFFR_X1 \STATE_reg[0]  ( .D(n11), .CK(clock), .RN(n10), .Q(n5), .QN(n7) );
  DLH_X1 \next_STATE_reg[1]  ( .G(enable), .D(N12), .Q(next_STATE[1]) );
  DFFR_X1 \STATE_reg[1]  ( .D(n9), .CK(clock), .RN(n10), .Q(prediction_o) );
  MUX2_X1 U8 ( .A(prediction_o), .B(next_STATE[1]), .S(enable), .Z(n9) );
  MUX2_X1 U9 ( .A(n5), .B(next_STATE[0]), .S(enable), .Z(n11) );
  NOR2_X1 U7 ( .A1(prediction_o), .A2(taken_i), .ZN(n6) );
  NAND2_X1 U6 ( .A1(prediction_o), .A2(taken_i), .ZN(n8) );
  OAI21_X1 U3 ( .B1(n6), .B2(n7), .A(n8), .ZN(N12) );
  OAI21_X1 U5 ( .B1(n5), .B2(n6), .A(n8), .ZN(N11) );
  INV_X1 U2 ( .A(reset), .ZN(n10) );
endmodule


module mux41_0 ( IN0, IN1, IN2, IN3, CTRL, OUT1 );
  input [31:0] IN0;
  input [31:0] IN1;
  input [31:0] IN2;
  input [31:0] IN3;
  input [1:0] CTRL;
  output [31:0] OUT1;
  wire   n194, n4, n5, n6, n7, n10, n11, n18, n19, n60, n61, n62, n63, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n166, n167, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193;

  AOI22_X1 U87 ( .A1(n6), .A2(IN1[12]), .B1(n193), .B2(IN0[12]), .ZN(n62) );
  AOI22_X1 U86 ( .A1(n89), .A2(IN3[12]), .B1(n90), .B2(IN2[12]), .ZN(n63) );
  AOI22_X1 U84 ( .A1(n6), .A2(IN1[13]), .B1(n193), .B2(IN0[13]), .ZN(n60) );
  AOI22_X1 U83 ( .A1(n89), .A2(IN3[13]), .B1(n90), .B2(IN2[13]), .ZN(n61) );
  AOI22_X1 U9 ( .A1(n6), .A2(IN1[7]), .B1(n193), .B2(IN0[7]), .ZN(n10) );
  AOI22_X1 U8 ( .A1(IN3[7]), .A2(n89), .B1(n90), .B2(IN2[7]), .ZN(n11) );
  AOI22_X1 U98 ( .A1(n6), .A2(IN1[0]), .B1(n193), .B2(IN0[0]), .ZN(n68) );
  AOI22_X1 U95 ( .A1(n89), .A2(IN3[0]), .B1(n90), .B2(IN2[0]), .ZN(n69) );
  AOI22_X1 U21 ( .A1(n6), .A2(IN1[3]), .B1(n193), .B2(IN0[3]), .ZN(n18) );
  AOI22_X1 U20 ( .A1(n89), .A2(IN3[3]), .B1(n90), .B2(IN2[3]), .ZN(n19) );
  NOR2_X1 U96 ( .A1(CTRL[0]), .A2(n70), .ZN(n5) );
  NOR2_X1 U99 ( .A1(CTRL[0]), .A2(CTRL[1]), .ZN(n7) );
  INV_X1 U101 ( .A(CTRL[1]), .ZN(n70) );
  AND2_X2 U100 ( .A1(n70), .A2(CTRL[0]), .ZN(n6) );
  NAND3_X1 U1 ( .A1(n169), .A2(n170), .A3(n171), .ZN(OUT1[1]) );
  BUF_X2 U2 ( .A(n194), .Z(OUT1[7]) );
  OR2_X2 U3 ( .A1(n134), .A2(n135), .ZN(OUT1[5]) );
  NAND2_X1 U4 ( .A1(n89), .A2(IN3[10]), .ZN(n71) );
  NAND2_X1 U5 ( .A1(n90), .A2(IN2[10]), .ZN(n72) );
  NAND2_X1 U6 ( .A1(n6), .A2(IN1[10]), .ZN(n73) );
  NAND4_X1 U7 ( .A1(n181), .A2(n71), .A3(n72), .A4(n73), .ZN(OUT1[10]) );
  AOI222_X1 U10 ( .A1(n90), .A2(IN2[8]), .B1(IN0[8]), .B2(n193), .C1(n6), .C2(
        IN1[8]), .ZN(n74) );
  NAND2_X1 U11 ( .A1(n89), .A2(IN3[8]), .ZN(n75) );
  NAND2_X1 U12 ( .A1(n74), .A2(n75), .ZN(OUT1[8]) );
  NAND2_X1 U13 ( .A1(n89), .A2(IN3[14]), .ZN(n76) );
  NAND2_X1 U14 ( .A1(n90), .A2(IN2[14]), .ZN(n77) );
  NAND2_X1 U15 ( .A1(n6), .A2(IN1[14]), .ZN(n78) );
  NAND4_X1 U16 ( .A1(n121), .A2(n76), .A3(n77), .A4(n78), .ZN(OUT1[14]) );
  AOI222_X1 U17 ( .A1(n7), .A2(IN0[4]), .B1(n6), .B2(IN1[4]), .C1(n5), .C2(
        IN2[4]), .ZN(n187) );
  AOI222_X1 U18 ( .A1(n90), .A2(IN2[25]), .B1(IN0[25]), .B2(n193), .C1(n6), 
        .C2(IN1[25]), .ZN(n79) );
  NAND2_X1 U19 ( .A1(n89), .A2(IN3[25]), .ZN(n80) );
  NAND2_X1 U22 ( .A1(n79), .A2(n80), .ZN(OUT1[25]) );
  AOI22_X1 U23 ( .A1(IN0[29]), .A2(n193), .B1(n6), .B2(IN1[29]), .ZN(n81) );
  INV_X1 U24 ( .A(n81), .ZN(n162) );
  AOI22_X1 U25 ( .A1(IN0[18]), .A2(n193), .B1(n6), .B2(IN1[18]), .ZN(n82) );
  INV_X1 U26 ( .A(n82), .ZN(n153) );
  AOI22_X1 U27 ( .A1(IN0[5]), .A2(n7), .B1(IN2[5]), .B2(n5), .ZN(n83) );
  INV_X1 U28 ( .A(n83), .ZN(n133) );
  NAND2_X1 U29 ( .A1(n89), .A2(IN3[22]), .ZN(n84) );
  NAND2_X1 U30 ( .A1(n90), .A2(IN2[22]), .ZN(n85) );
  NAND2_X1 U31 ( .A1(n6), .A2(IN1[22]), .ZN(n86) );
  NAND4_X1 U32 ( .A1(n154), .A2(n84), .A3(n85), .A4(n86), .ZN(OUT1[22]) );
  NAND2_X1 U33 ( .A1(n89), .A2(IN3[4]), .ZN(n87) );
  NAND2_X1 U34 ( .A1(n187), .A2(n87), .ZN(OUT1[4]) );
  NAND2_X4 U35 ( .A1(n151), .A2(n152), .ZN(OUT1[18]) );
  NAND2_X1 U36 ( .A1(n11), .A2(n10), .ZN(n194) );
  NAND2_X2 U37 ( .A1(n122), .A2(n123), .ZN(OUT1[15]) );
  OR3_X2 U38 ( .A1(n174), .A2(n175), .A3(n173), .ZN(OUT1[2]) );
  BUF_X2 U39 ( .A(n4), .Z(n89) );
  NAND2_X1 U40 ( .A1(n91), .A2(n92), .ZN(OUT1[24]) );
  AND2_X1 U41 ( .A1(IN3[5]), .A2(n89), .ZN(n134) );
  AND2_X1 U42 ( .A1(IN3[2]), .A2(n89), .ZN(n174) );
  INV_X1 U43 ( .A(n132), .ZN(n135) );
  INV_X1 U44 ( .A(n172), .ZN(n175) );
  BUF_X2 U45 ( .A(n7), .Z(n193) );
  BUF_X2 U46 ( .A(n5), .Z(n90) );
  AND2_X1 U47 ( .A1(CTRL[0]), .A2(CTRL[1]), .ZN(n4) );
  NAND2_X1 U48 ( .A1(n127), .A2(n128), .ZN(OUT1[17]) );
  NAND2_X1 U49 ( .A1(n160), .A2(n161), .ZN(OUT1[29]) );
  NAND2_X1 U50 ( .A1(n182), .A2(n183), .ZN(OUT1[16]) );
  NAND2_X1 U51 ( .A1(n136), .A2(n137), .ZN(OUT1[20]) );
  AND2_X1 U52 ( .A1(IN1[2]), .A2(n6), .ZN(n173) );
  NAND2_X1 U53 ( .A1(n111), .A2(n112), .ZN(OUT1[21]) );
  NAND2_X1 U54 ( .A1(n106), .A2(n107), .ZN(OUT1[23]) );
  NAND2_X1 U55 ( .A1(n146), .A2(n147), .ZN(OUT1[11]) );
  NAND2_X1 U56 ( .A1(n141), .A2(n142), .ZN(OUT1[19]) );
  NAND2_X1 U57 ( .A1(n62), .A2(n63), .ZN(OUT1[12]) );
  NAND2_X1 U58 ( .A1(n101), .A2(n102), .ZN(OUT1[31]) );
  NAND2_X1 U59 ( .A1(n68), .A2(n69), .ZN(OUT1[0]) );
  NAND2_X1 U60 ( .A1(n116), .A2(n117), .ZN(OUT1[26]) );
  NAND2_X1 U61 ( .A1(n60), .A2(n61), .ZN(OUT1[13]) );
  NAND2_X1 U62 ( .A1(n18), .A2(n19), .ZN(OUT1[3]) );
  NAND2_X1 U63 ( .A1(n155), .A2(n156), .ZN(OUT1[27]) );
  NAND2_X1 U64 ( .A1(n163), .A2(n164), .ZN(OUT1[30]) );
  NAND2_X1 U65 ( .A1(n177), .A2(n176), .ZN(OUT1[28]) );
  NAND2_X1 U66 ( .A1(IN3[28]), .A2(n89), .ZN(n176) );
  NAND2_X2 U67 ( .A1(n188), .A2(n189), .ZN(OUT1[6]) );
  NAND2_X2 U68 ( .A1(n96), .A2(n97), .ZN(OUT1[9]) );
  AOI21_X1 U69 ( .B1(IN2[17]), .B2(n90), .A(n129), .ZN(n128) );
  NAND2_X1 U70 ( .A1(n130), .A2(n131), .ZN(n129) );
  NAND2_X1 U71 ( .A1(n193), .A2(IN0[17]), .ZN(n131) );
  NAND2_X1 U72 ( .A1(IN1[17]), .A2(n6), .ZN(n130) );
  AOI21_X1 U73 ( .B1(IN2[16]), .B2(n90), .A(n184), .ZN(n183) );
  NAND2_X1 U74 ( .A1(n185), .A2(n186), .ZN(n184) );
  NAND2_X1 U75 ( .A1(n193), .A2(IN0[16]), .ZN(n186) );
  NAND2_X1 U76 ( .A1(IN1[16]), .A2(n6), .ZN(n185) );
  AOI21_X1 U77 ( .B1(IN2[19]), .B2(n90), .A(n143), .ZN(n142) );
  NAND2_X1 U78 ( .A1(n144), .A2(n145), .ZN(n143) );
  NAND2_X1 U79 ( .A1(n193), .A2(IN0[19]), .ZN(n145) );
  NAND2_X1 U80 ( .A1(IN1[19]), .A2(n6), .ZN(n144) );
  AOI21_X1 U81 ( .B1(IN2[18]), .B2(n90), .A(n153), .ZN(n152) );
  NAND2_X1 U82 ( .A1(n179), .A2(n180), .ZN(n178) );
  NAND2_X1 U85 ( .A1(n193), .A2(IN0[28]), .ZN(n180) );
  NAND2_X1 U88 ( .A1(IN1[28]), .A2(n6), .ZN(n179) );
  AOI21_X1 U89 ( .B1(IN2[27]), .B2(n90), .A(n157), .ZN(n156) );
  NAND2_X1 U90 ( .A1(n158), .A2(n159), .ZN(n157) );
  NAND2_X1 U91 ( .A1(n193), .A2(IN0[27]), .ZN(n159) );
  NAND2_X1 U92 ( .A1(IN1[27]), .A2(n6), .ZN(n158) );
  AOI21_X1 U93 ( .B1(IN2[30]), .B2(n90), .A(n165), .ZN(n164) );
  NAND2_X1 U94 ( .A1(n166), .A2(n167), .ZN(n165) );
  NAND2_X1 U97 ( .A1(n193), .A2(IN0[30]), .ZN(n167) );
  NAND2_X1 U102 ( .A1(IN1[30]), .A2(n6), .ZN(n166) );
  AOI21_X1 U103 ( .B1(IN2[23]), .B2(n90), .A(n108), .ZN(n107) );
  NAND2_X1 U104 ( .A1(n109), .A2(n110), .ZN(n108) );
  NAND2_X1 U105 ( .A1(n193), .A2(IN0[23]), .ZN(n110) );
  NAND2_X1 U106 ( .A1(IN1[23]), .A2(n6), .ZN(n109) );
  NAND2_X1 U107 ( .A1(n193), .A2(IN0[22]), .ZN(n154) );
  AOI21_X1 U108 ( .B1(IN2[21]), .B2(n90), .A(n113), .ZN(n112) );
  NAND2_X1 U109 ( .A1(n114), .A2(n115), .ZN(n113) );
  NAND2_X1 U110 ( .A1(n193), .A2(IN0[21]), .ZN(n115) );
  NAND2_X1 U111 ( .A1(IN1[21]), .A2(n6), .ZN(n114) );
  AOI21_X1 U112 ( .B1(IN2[20]), .B2(n90), .A(n138), .ZN(n137) );
  NAND2_X1 U113 ( .A1(n139), .A2(n140), .ZN(n138) );
  NAND2_X1 U114 ( .A1(n193), .A2(IN0[20]), .ZN(n140) );
  NAND2_X1 U115 ( .A1(IN1[20]), .A2(n6), .ZN(n139) );
  AOI21_X1 U116 ( .B1(IN2[26]), .B2(n90), .A(n118), .ZN(n117) );
  NAND2_X1 U117 ( .A1(n119), .A2(n120), .ZN(n118) );
  NAND2_X1 U118 ( .A1(n193), .A2(IN0[26]), .ZN(n120) );
  NAND2_X1 U119 ( .A1(IN1[26]), .A2(n6), .ZN(n119) );
  AOI21_X1 U120 ( .B1(IN2[24]), .B2(n90), .A(n93), .ZN(n92) );
  NAND2_X1 U121 ( .A1(n94), .A2(n95), .ZN(n93) );
  NAND2_X1 U122 ( .A1(n193), .A2(IN0[24]), .ZN(n95) );
  NAND2_X1 U123 ( .A1(IN1[24]), .A2(n6), .ZN(n94) );
  AOI21_X1 U124 ( .B1(IN2[31]), .B2(n90), .A(n103), .ZN(n102) );
  NAND2_X1 U125 ( .A1(n104), .A2(n105), .ZN(n103) );
  NAND2_X1 U126 ( .A1(n193), .A2(IN0[31]), .ZN(n105) );
  NAND2_X1 U127 ( .A1(IN1[31]), .A2(n6), .ZN(n104) );
  AOI22_X1 U128 ( .A1(n90), .A2(IN2[2]), .B1(n7), .B2(IN0[2]), .ZN(n172) );
  NAND2_X1 U129 ( .A1(IN1[1]), .A2(n6), .ZN(n171) );
  AOI22_X1 U130 ( .A1(n90), .A2(IN2[1]), .B1(n193), .B2(IN0[1]), .ZN(n170) );
  AOI21_X1 U131 ( .B1(IN1[6]), .B2(n6), .A(n190), .ZN(n189) );
  NAND2_X1 U132 ( .A1(n191), .A2(n192), .ZN(n190) );
  NAND2_X1 U133 ( .A1(n193), .A2(IN0[6]), .ZN(n192) );
  NAND2_X1 U134 ( .A1(n90), .A2(IN2[6]), .ZN(n191) );
  AOI21_X1 U135 ( .B1(IN1[5]), .B2(n6), .A(n133), .ZN(n132) );
  AOI21_X1 U136 ( .B1(IN2[11]), .B2(n90), .A(n148), .ZN(n147) );
  NAND2_X1 U137 ( .A1(n149), .A2(n150), .ZN(n148) );
  NAND2_X1 U138 ( .A1(n193), .A2(IN0[11]), .ZN(n150) );
  NAND2_X1 U139 ( .A1(IN1[11]), .A2(n6), .ZN(n149) );
  NAND2_X1 U140 ( .A1(n193), .A2(IN0[10]), .ZN(n181) );
  AOI21_X1 U141 ( .B1(IN2[9]), .B2(n90), .A(n98), .ZN(n97) );
  NAND2_X1 U142 ( .A1(n99), .A2(n100), .ZN(n98) );
  NAND2_X1 U143 ( .A1(n193), .A2(IN0[9]), .ZN(n100) );
  NAND2_X1 U144 ( .A1(IN1[9]), .A2(n6), .ZN(n99) );
  AOI21_X1 U145 ( .B1(IN2[15]), .B2(n90), .A(n124), .ZN(n123) );
  NAND2_X1 U146 ( .A1(n125), .A2(n126), .ZN(n124) );
  NAND2_X1 U147 ( .A1(n193), .A2(IN0[15]), .ZN(n126) );
  NAND2_X1 U148 ( .A1(IN1[15]), .A2(n6), .ZN(n125) );
  NAND2_X1 U149 ( .A1(n193), .A2(IN0[14]), .ZN(n121) );
  NAND2_X1 U150 ( .A1(IN3[24]), .A2(n4), .ZN(n91) );
  NAND2_X1 U151 ( .A1(IN3[9]), .A2(n89), .ZN(n96) );
  NAND2_X1 U152 ( .A1(IN3[31]), .A2(n89), .ZN(n101) );
  NAND2_X1 U153 ( .A1(IN3[23]), .A2(n89), .ZN(n106) );
  NAND2_X1 U154 ( .A1(IN3[21]), .A2(n89), .ZN(n111) );
  NAND2_X1 U155 ( .A1(IN3[26]), .A2(n89), .ZN(n116) );
  NAND2_X1 U156 ( .A1(IN3[15]), .A2(n89), .ZN(n122) );
  NAND2_X1 U157 ( .A1(IN3[17]), .A2(n89), .ZN(n127) );
  NAND2_X1 U158 ( .A1(IN3[20]), .A2(n89), .ZN(n136) );
  NAND2_X1 U159 ( .A1(IN3[19]), .A2(n89), .ZN(n141) );
  NAND2_X1 U160 ( .A1(IN3[11]), .A2(n89), .ZN(n146) );
  NAND2_X1 U161 ( .A1(IN3[18]), .A2(n89), .ZN(n151) );
  NAND2_X1 U162 ( .A1(IN3[27]), .A2(n89), .ZN(n155) );
  NAND2_X1 U163 ( .A1(IN3[29]), .A2(n4), .ZN(n160) );
  AOI21_X1 U164 ( .B1(IN2[29]), .B2(n90), .A(n162), .ZN(n161) );
  NAND2_X1 U165 ( .A1(IN3[30]), .A2(n4), .ZN(n163) );
  NAND2_X1 U166 ( .A1(IN3[1]), .A2(n89), .ZN(n169) );
  AOI21_X1 U167 ( .B1(IN2[28]), .B2(n90), .A(n178), .ZN(n177) );
  NAND2_X1 U168 ( .A1(IN3[16]), .A2(n89), .ZN(n182) );
  NAND2_X1 U169 ( .A1(IN3[6]), .A2(n89), .ZN(n188) );
endmodule


module add4 ( IN1, OUT1 );
  input [31:0] IN1;
  output [31:0] OUT1;
  wire   \IN1[1] , \IN1[0] , \add_27/carry[4] , \add_27/carry[5] ,
         \add_27/carry[6] , \add_27/carry[7] , \add_27/carry[8] ,
         \add_27/carry[9] , \add_27/carry[10] , \add_27/carry[11] ,
         \add_27/carry[12] , \add_27/carry[13] , \add_27/carry[14] ,
         \add_27/carry[15] , \add_27/carry[16] , \add_27/carry[17] ,
         \add_27/carry[18] , \add_27/carry[19] , \add_27/carry[20] ,
         \add_27/carry[21] , \add_27/carry[22] , \add_27/carry[23] ,
         \add_27/carry[24] , \add_27/carry[25] , \add_27/carry[26] ,
         \add_27/carry[27] , \add_27/carry[28] , \add_27/carry[29] ,
         \add_27/carry[30] , n1;
  assign OUT1[1] = \IN1[1] ;
  assign \IN1[1]  = IN1[1];
  assign OUT1[0] = \IN1[0] ;
  assign \IN1[0]  = IN1[0];

  XOR2_X1 \add_27/U57  ( .A(IN1[3]), .B(IN1[2]), .Z(OUT1[3]) );
  XOR2_X1 \add_27/U55  ( .A(IN1[4]), .B(\add_27/carry[4] ), .Z(OUT1[4]) );
  XOR2_X1 \add_27/U53  ( .A(IN1[5]), .B(\add_27/carry[5] ), .Z(OUT1[5]) );
  XOR2_X1 \add_27/U51  ( .A(IN1[6]), .B(\add_27/carry[6] ), .Z(OUT1[6]) );
  XOR2_X1 \add_27/U49  ( .A(IN1[7]), .B(\add_27/carry[7] ), .Z(OUT1[7]) );
  XOR2_X1 \add_27/U47  ( .A(IN1[8]), .B(\add_27/carry[8] ), .Z(OUT1[8]) );
  XOR2_X1 \add_27/U45  ( .A(IN1[9]), .B(\add_27/carry[9] ), .Z(OUT1[9]) );
  XOR2_X1 \add_27/U43  ( .A(IN1[10]), .B(\add_27/carry[10] ), .Z(OUT1[10]) );
  XOR2_X1 \add_27/U41  ( .A(IN1[11]), .B(\add_27/carry[11] ), .Z(OUT1[11]) );
  XOR2_X1 \add_27/U39  ( .A(IN1[12]), .B(\add_27/carry[12] ), .Z(OUT1[12]) );
  XOR2_X1 \add_27/U37  ( .A(IN1[13]), .B(\add_27/carry[13] ), .Z(OUT1[13]) );
  XOR2_X1 \add_27/U35  ( .A(IN1[14]), .B(\add_27/carry[14] ), .Z(OUT1[14]) );
  XOR2_X1 \add_27/U33  ( .A(IN1[15]), .B(\add_27/carry[15] ), .Z(OUT1[15]) );
  XOR2_X1 \add_27/U31  ( .A(IN1[16]), .B(\add_27/carry[16] ), .Z(OUT1[16]) );
  XOR2_X1 \add_27/U29  ( .A(IN1[17]), .B(\add_27/carry[17] ), .Z(OUT1[17]) );
  XOR2_X1 \add_27/U27  ( .A(IN1[18]), .B(\add_27/carry[18] ), .Z(OUT1[18]) );
  XOR2_X1 \add_27/U25  ( .A(IN1[19]), .B(\add_27/carry[19] ), .Z(OUT1[19]) );
  XOR2_X1 \add_27/U23  ( .A(IN1[20]), .B(\add_27/carry[20] ), .Z(OUT1[20]) );
  XOR2_X1 \add_27/U21  ( .A(IN1[21]), .B(\add_27/carry[21] ), .Z(OUT1[21]) );
  XOR2_X1 \add_27/U19  ( .A(IN1[22]), .B(\add_27/carry[22] ), .Z(OUT1[22]) );
  XOR2_X1 \add_27/U17  ( .A(IN1[23]), .B(\add_27/carry[23] ), .Z(OUT1[23]) );
  XOR2_X1 \add_27/U15  ( .A(IN1[24]), .B(\add_27/carry[24] ), .Z(OUT1[24]) );
  XOR2_X1 \add_27/U13  ( .A(IN1[25]), .B(\add_27/carry[25] ), .Z(OUT1[25]) );
  XOR2_X1 \add_27/U11  ( .A(IN1[26]), .B(\add_27/carry[26] ), .Z(OUT1[26]) );
  XOR2_X1 \add_27/U9  ( .A(IN1[27]), .B(\add_27/carry[27] ), .Z(OUT1[27]) );
  XOR2_X1 \add_27/U7  ( .A(IN1[28]), .B(\add_27/carry[28] ), .Z(OUT1[28]) );
  XOR2_X1 \add_27/U5  ( .A(IN1[29]), .B(\add_27/carry[29] ), .Z(OUT1[29]) );
  XOR2_X1 \add_27/U3  ( .A(IN1[30]), .B(\add_27/carry[30] ), .Z(OUT1[30]) );
  INV_X1 \add_27/U58  ( .A(IN1[2]), .ZN(OUT1[2]) );
  AND2_X1 \add_27/U36  ( .A1(\add_27/carry[13] ), .A2(IN1[13]), .ZN(
        \add_27/carry[14] ) );
  AND2_X1 \add_27/U34  ( .A1(\add_27/carry[14] ), .A2(IN1[14]), .ZN(
        \add_27/carry[15] ) );
  AND2_X1 \add_27/U32  ( .A1(\add_27/carry[15] ), .A2(IN1[15]), .ZN(
        \add_27/carry[16] ) );
  AND2_X1 \add_27/U30  ( .A1(\add_27/carry[16] ), .A2(IN1[16]), .ZN(
        \add_27/carry[17] ) );
  AND2_X1 \add_27/U28  ( .A1(\add_27/carry[17] ), .A2(IN1[17]), .ZN(
        \add_27/carry[18] ) );
  AND2_X1 \add_27/U26  ( .A1(\add_27/carry[18] ), .A2(IN1[18]), .ZN(
        \add_27/carry[19] ) );
  AND2_X1 \add_27/U12  ( .A1(\add_27/carry[25] ), .A2(IN1[25]), .ZN(
        \add_27/carry[26] ) );
  AND2_X1 \add_27/U10  ( .A1(\add_27/carry[26] ), .A2(IN1[26]), .ZN(
        \add_27/carry[27] ) );
  AND2_X1 \add_27/U8  ( .A1(\add_27/carry[27] ), .A2(IN1[27]), .ZN(
        \add_27/carry[28] ) );
  AND2_X1 \add_27/U6  ( .A1(\add_27/carry[28] ), .A2(IN1[28]), .ZN(
        \add_27/carry[29] ) );
  AND2_X1 \add_27/U4  ( .A1(\add_27/carry[29] ), .A2(IN1[29]), .ZN(
        \add_27/carry[30] ) );
  AND2_X1 U3 ( .A1(IN1[2]), .A2(IN1[3]), .ZN(\add_27/carry[4] ) );
  AND2_X1 U4 ( .A1(\add_27/carry[4] ), .A2(IN1[4]), .ZN(\add_27/carry[5] ) );
  AND2_X1 U5 ( .A1(\add_27/carry[19] ), .A2(IN1[19]), .ZN(\add_27/carry[20] )
         );
  AND2_X1 U6 ( .A1(\add_27/carry[24] ), .A2(IN1[24]), .ZN(\add_27/carry[25] )
         );
  NAND2_X1 U7 ( .A1(\add_27/carry[30] ), .A2(IN1[30]), .ZN(n1) );
  XNOR2_X1 U8 ( .A(n1), .B(IN1[31]), .ZN(OUT1[31]) );
  AND2_X2 U9 ( .A1(\add_27/carry[23] ), .A2(IN1[23]), .ZN(\add_27/carry[24] )
         );
  AND2_X2 U10 ( .A1(\add_27/carry[22] ), .A2(IN1[22]), .ZN(\add_27/carry[23] )
         );
  AND2_X2 U11 ( .A1(\add_27/carry[20] ), .A2(IN1[20]), .ZN(\add_27/carry[21] )
         );
  AND2_X2 U12 ( .A1(\add_27/carry[21] ), .A2(IN1[21]), .ZN(\add_27/carry[22] )
         );
  AND2_X2 U13 ( .A1(\add_27/carry[6] ), .A2(IN1[6]), .ZN(\add_27/carry[7] ) );
  AND2_X2 U14 ( .A1(\add_27/carry[5] ), .A2(IN1[5]), .ZN(\add_27/carry[6] ) );
  AND2_X2 U15 ( .A1(\add_27/carry[8] ), .A2(IN1[8]), .ZN(\add_27/carry[9] ) );
  AND2_X2 U16 ( .A1(\add_27/carry[7] ), .A2(IN1[7]), .ZN(\add_27/carry[8] ) );
  AND2_X2 U17 ( .A1(\add_27/carry[10] ), .A2(IN1[10]), .ZN(\add_27/carry[11] )
         );
  AND2_X2 U18 ( .A1(\add_27/carry[9] ), .A2(IN1[9]), .ZN(\add_27/carry[10] )
         );
  AND2_X2 U19 ( .A1(\add_27/carry[12] ), .A2(IN1[12]), .ZN(\add_27/carry[13] )
         );
  AND2_X2 U20 ( .A1(\add_27/carry[11] ), .A2(IN1[11]), .ZN(\add_27/carry[12] )
         );
endmodule


module ff32_en_0 ( D, en, clk, rst, Q );
  input [31:0] D;
  output [31:0] Q;
  input en, clk, rst;
  wire   n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n97, net644934, net644935, net644936, net644937,
         net644938, net644939, net644940, net644941, net644942, net644943,
         net644944, net644945, net644947, net644948, net644949, net644950,
         net644951, net644952, net644953, net644954, net644955, net644956,
         net644957, net644958, net644959, net644960, net644961, net644962,
         net644963, net644964, net644965, n3, n5, n8, n9, n12, n13, n20, n25,
         n27, n32, n33, n29, n11, n14, n16, n28, n17, n31, n30, n10, n15, n23,
         n4, n6, n19, n26, n7, n24, n2, n18, n1, n21, n22, n34, n36, n37, n38,
         n39;

  DFFR_X1 \Q_reg[30]  ( .D(n95), .CK(clk), .RN(n39), .Q(Q[30]), .QN(net644964)
         );
  DFFR_X1 \Q_reg[29]  ( .D(n94), .CK(clk), .RN(n39), .Q(Q[29]), .QN(net644963)
         );
  DFFR_X1 \Q_reg[28]  ( .D(n93), .CK(clk), .RN(n39), .Q(Q[28]), .QN(net644962)
         );
  DFFR_X1 \Q_reg[27]  ( .D(n92), .CK(clk), .RN(n39), .Q(Q[27]), .QN(net644961)
         );
  DFFR_X1 \Q_reg[26]  ( .D(n91), .CK(clk), .RN(n39), .Q(Q[26]), .QN(net644960)
         );
  DFFR_X1 \Q_reg[25]  ( .D(n90), .CK(clk), .RN(n39), .Q(Q[25]), .QN(net644959)
         );
  DFFR_X1 \Q_reg[24]  ( .D(n89), .CK(clk), .RN(n39), .Q(Q[24]), .QN(net644958)
         );
  DFFR_X1 \Q_reg[23]  ( .D(n88), .CK(clk), .RN(n39), .Q(Q[23]), .QN(net644957)
         );
  DFFR_X1 \Q_reg[22]  ( .D(n87), .CK(clk), .RN(n39), .Q(Q[22]), .QN(net644956)
         );
  DFFR_X1 \Q_reg[21]  ( .D(n86), .CK(clk), .RN(n39), .Q(Q[21]), .QN(net644955)
         );
  DFFR_X1 \Q_reg[20]  ( .D(n85), .CK(clk), .RN(n39), .Q(Q[20]), .QN(net644954)
         );
  DFFR_X1 \Q_reg[19]  ( .D(n84), .CK(clk), .RN(n39), .Q(Q[19]), .QN(net644953)
         );
  DFFR_X1 \Q_reg[18]  ( .D(n83), .CK(clk), .RN(n39), .Q(Q[18]), .QN(net644952)
         );
  DFFR_X1 \Q_reg[17]  ( .D(n82), .CK(clk), .RN(n39), .Q(Q[17]), .QN(net644951)
         );
  DFFR_X1 \Q_reg[16]  ( .D(n81), .CK(clk), .RN(n39), .Q(Q[16]), .QN(net644950)
         );
  DFFR_X1 \Q_reg[15]  ( .D(n80), .CK(clk), .RN(n39), .Q(Q[15]), .QN(net644949)
         );
  DFFR_X1 \Q_reg[14]  ( .D(n79), .CK(clk), .RN(n39), .Q(Q[14]), .QN(net644948)
         );
  DFFR_X1 \Q_reg[12]  ( .D(n77), .CK(clk), .RN(n39), .Q(Q[12]) );
  DFFR_X1 \Q_reg[10]  ( .D(n75), .CK(clk), .RN(n39), .Q(Q[10]), .QN(net644944)
         );
  DFFR_X1 \Q_reg[9]  ( .D(n74), .CK(clk), .RN(n39), .Q(Q[9]), .QN(net644943)
         );
  DFFR_X1 \Q_reg[8]  ( .D(n73), .CK(clk), .RN(n39), .Q(Q[8]), .QN(net644942)
         );
  DFFR_X1 \Q_reg[7]  ( .D(n72), .CK(clk), .RN(n39), .Q(Q[7]), .QN(net644941)
         );
  DFFR_X1 \Q_reg[6]  ( .D(n71), .CK(clk), .RN(n39), .Q(Q[6]), .QN(net644940)
         );
  DFFR_X1 \Q_reg[5]  ( .D(n70), .CK(clk), .RN(n39), .Q(Q[5]), .QN(net644939)
         );
  DFFR_X1 \Q_reg[4]  ( .D(n69), .CK(clk), .RN(n39), .Q(Q[4]), .QN(net644938)
         );
  DFFR_X1 \Q_reg[3]  ( .D(n68), .CK(clk), .RN(n39), .Q(Q[3]), .QN(net644937)
         );
  DFFR_X1 \Q_reg[2]  ( .D(n67), .CK(clk), .RN(n39), .Q(Q[2]), .QN(net644936)
         );
  DFFR_X1 \Q_reg[1]  ( .D(n66), .CK(clk), .RN(n39), .Q(Q[1]), .QN(net644935)
         );
  DFFR_X1 \Q_reg[0]  ( .D(n65), .CK(clk), .RN(n39), .Q(Q[0]), .QN(net644934)
         );
  DFFR_X1 \Q_reg[13]  ( .D(n78), .CK(clk), .RN(n39), .Q(Q[13]), .QN(net644947)
         );
  DFFR_X1 \Q_reg[31]  ( .D(n97), .CK(clk), .RN(n39), .Q(Q[31]), .QN(net644965)
         );
  DFFR_X1 \Q_reg[11]  ( .D(n76), .CK(clk), .RN(n39), .Q(Q[11]), .QN(net644945)
         );
  NAND2_X1 U2 ( .A1(n37), .A2(D[11]), .ZN(n1) );
  OAI21_X1 U3 ( .B1(en), .B2(net644945), .A(n1), .ZN(n76) );
  INV_X1 U4 ( .A(Q[12]), .ZN(n21) );
  NAND2_X1 U5 ( .A1(D[12]), .A2(n36), .ZN(n22) );
  OAI21_X1 U6 ( .B1(n21), .B2(en), .A(n22), .ZN(n77) );
  OR2_X1 U7 ( .A1(en), .A2(net644965), .ZN(n34) );
  NAND2_X1 U8 ( .A1(n34), .A2(n2), .ZN(n97) );
  INV_X2 U9 ( .A(rst), .ZN(n39) );
  BUF_X1 U10 ( .A(en), .Z(n36) );
  BUF_X1 U11 ( .A(en), .Z(n37) );
  BUF_X1 U12 ( .A(en), .Z(n38) );
  OAI21_X1 U13 ( .B1(en), .B2(net644949), .A(n18), .ZN(n80) );
  OAI21_X1 U14 ( .B1(en), .B2(net644944), .A(n23), .ZN(n75) );
  OAI21_X1 U15 ( .B1(en), .B2(net644952), .A(n15), .ZN(n83) );
  OAI21_X1 U16 ( .B1(en), .B2(net644948), .A(n19), .ZN(n79) );
  OAI21_X1 U17 ( .B1(en), .B2(net644950), .A(n17), .ZN(n81) );
  OAI21_X1 U18 ( .B1(en), .B2(net644951), .A(n16), .ZN(n82) );
  NAND2_X1 U19 ( .A1(D[15]), .A2(en), .ZN(n18) );
  NAND2_X1 U20 ( .A1(en), .A2(D[31]), .ZN(n2) );
  NAND2_X1 U21 ( .A1(D[9]), .A2(en), .ZN(n24) );
  OAI21_X1 U22 ( .B1(en), .B2(net644943), .A(n24), .ZN(n74) );
  NAND2_X1 U23 ( .A1(n38), .A2(D[26]), .ZN(n7) );
  OAI21_X1 U24 ( .B1(n36), .B2(net644960), .A(n7), .ZN(n91) );
  NAND2_X1 U25 ( .A1(D[7]), .A2(en), .ZN(n26) );
  OAI21_X1 U26 ( .B1(en), .B2(net644941), .A(n26), .ZN(n72) );
  NAND2_X1 U27 ( .A1(D[14]), .A2(n37), .ZN(n19) );
  NAND2_X1 U28 ( .A1(n38), .A2(D[27]), .ZN(n6) );
  OAI21_X1 U29 ( .B1(n36), .B2(net644961), .A(n6), .ZN(n92) );
  NAND2_X1 U30 ( .A1(D[29]), .A2(n38), .ZN(n4) );
  OAI21_X1 U31 ( .B1(n36), .B2(net644963), .A(n4), .ZN(n94) );
  NAND2_X1 U32 ( .A1(D[10]), .A2(n37), .ZN(n23) );
  NAND2_X1 U33 ( .A1(D[18]), .A2(en), .ZN(n15) );
  NAND2_X1 U34 ( .A1(n38), .A2(D[23]), .ZN(n10) );
  OAI21_X1 U35 ( .B1(n36), .B2(net644957), .A(n10), .ZN(n88) );
  NAND2_X1 U36 ( .A1(D[3]), .A2(n38), .ZN(n30) );
  OAI21_X1 U37 ( .B1(n37), .B2(net644937), .A(n30), .ZN(n68) );
  NAND2_X1 U38 ( .A1(n38), .A2(D[2]), .ZN(n31) );
  OAI21_X1 U39 ( .B1(n37), .B2(net644936), .A(n31), .ZN(n67) );
  NAND2_X1 U40 ( .A1(D[16]), .A2(en), .ZN(n17) );
  NAND2_X1 U41 ( .A1(D[5]), .A2(n38), .ZN(n28) );
  OAI21_X1 U42 ( .B1(n37), .B2(net644939), .A(n28), .ZN(n70) );
  NAND2_X1 U43 ( .A1(D[17]), .A2(en), .ZN(n16) );
  NAND2_X1 U44 ( .A1(D[19]), .A2(n38), .ZN(n14) );
  OAI21_X1 U45 ( .B1(n36), .B2(net644953), .A(n14), .ZN(n84) );
  NAND2_X1 U46 ( .A1(D[22]), .A2(en), .ZN(n11) );
  OAI21_X1 U47 ( .B1(n36), .B2(net644956), .A(n11), .ZN(n87) );
  NAND2_X1 U48 ( .A1(n38), .A2(D[4]), .ZN(n29) );
  OAI21_X1 U49 ( .B1(n37), .B2(net644938), .A(n29), .ZN(n69) );
  OAI21_X1 U50 ( .B1(n37), .B2(net644934), .A(n33), .ZN(n65) );
  OAI21_X1 U51 ( .B1(n36), .B2(net644955), .A(n12), .ZN(n86) );
  OAI21_X1 U52 ( .B1(n36), .B2(net644962), .A(n5), .ZN(n93) );
  NAND2_X1 U53 ( .A1(n38), .A2(D[28]), .ZN(n5) );
  OAI21_X1 U54 ( .B1(n36), .B2(net644964), .A(n3), .ZN(n95) );
  NAND2_X1 U55 ( .A1(en), .A2(D[30]), .ZN(n3) );
  OAI21_X1 U56 ( .B1(n36), .B2(net644958), .A(n9), .ZN(n89) );
  NAND2_X1 U57 ( .A1(D[24]), .A2(n38), .ZN(n9) );
  OAI21_X1 U58 ( .B1(n36), .B2(net644959), .A(n8), .ZN(n90) );
  NAND2_X1 U59 ( .A1(n38), .A2(D[25]), .ZN(n8) );
  OAI21_X1 U60 ( .B1(n36), .B2(net644954), .A(n13), .ZN(n85) );
  NAND2_X1 U61 ( .A1(D[20]), .A2(n36), .ZN(n13) );
  OAI21_X1 U62 ( .B1(n37), .B2(net644942), .A(n25), .ZN(n73) );
  NAND2_X1 U63 ( .A1(D[8]), .A2(n37), .ZN(n25) );
  NAND2_X1 U64 ( .A1(en), .A2(D[0]), .ZN(n33) );
  OAI21_X1 U65 ( .B1(n37), .B2(net644940), .A(n27), .ZN(n71) );
  NAND2_X1 U66 ( .A1(D[6]), .A2(n38), .ZN(n27) );
  OAI21_X1 U67 ( .B1(n37), .B2(net644935), .A(n32), .ZN(n66) );
  NAND2_X1 U68 ( .A1(en), .A2(D[1]), .ZN(n32) );
  NAND2_X1 U69 ( .A1(n38), .A2(D[21]), .ZN(n12) );
  OAI21_X1 U70 ( .B1(en), .B2(net644947), .A(n20), .ZN(n78) );
  NAND2_X1 U71 ( .A1(D[13]), .A2(n37), .ZN(n20) );
endmodule


module fw_logic ( D1_i, rAdec_i, D2_i, D3_i, rA_i, rB_i, S_mem_W, S_wb_W, 
        S_exe_W, S_FWAdec, S_FWA, S_FWB, S_mem_LOAD_BAR );
  input [4:0] D1_i;
  input [4:0] rAdec_i;
  input [4:0] D2_i;
  input [4:0] D3_i;
  input [4:0] rA_i;
  input [4:0] rB_i;
  output [1:0] S_FWAdec;
  output [1:0] S_FWA;
  output [1:0] S_FWB;
  input S_mem_W, S_wb_W, S_exe_W, S_mem_LOAD_BAR;
  wire   S_mem_LOAD, n102, n103, n22, n24, n25, n28, n29, n30, n31, n32, n34,
         n35, n36, n37, n38, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n44, n43, n42, n41,
         n40, n39, n101, n65, n66, n67, n69, n70, n71, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n99, n100;
  assign S_mem_LOAD = S_mem_LOAD_BAR;

  XOR2_X1 U53 ( .A(D2_i[2]), .B(rB_i[2]), .Z(n29) );
  XOR2_X1 U54 ( .A(D2_i[2]), .B(rAdec_i[2]), .Z(n45) );
  XOR2_X1 U55 ( .A(D2_i[2]), .B(rA_i[2]), .Z(n60) );
  OAI221_X1 U39 ( .B1(rA_i[3]), .B2(n28), .C1(n59), .C2(n67), .A(S_wb_W), .ZN(
        n50) );
  INV_X1 U24 ( .A(rAdec_i[3]), .ZN(n44) );
  INV_X1 U40 ( .A(rA_i[3]), .ZN(n59) );
  INV_X1 U37 ( .A(rA_i[2]), .ZN(n57) );
  INV_X1 U38 ( .A(rA_i[1]), .ZN(n56) );
  INV_X1 U33 ( .A(rA_i[0]), .ZN(n54) );
  INV_X1 U34 ( .A(rA_i[4]), .ZN(n53) );
  OR2_X1 U2 ( .A1(n94), .A2(rB_i[1]), .ZN(n99) );
  CLKBUF_X1 U3 ( .A(n66), .Z(n73) );
  INV_X1 U4 ( .A(D2_i[1]), .ZN(n97) );
  OR2_X1 U5 ( .A1(n34), .A2(rB_i[3]), .ZN(n100) );
  INV_X1 U6 ( .A(n90), .ZN(n76) );
  CLKBUF_X1 U7 ( .A(D3_i[1]), .Z(n65) );
  INV_X1 U8 ( .A(D3_i[2]), .ZN(n25) );
  CLKBUF_X1 U9 ( .A(D3_i[0]), .Z(n91) );
  OR2_X1 U10 ( .A1(n96), .A2(rAdec_i[4]), .ZN(n92) );
  INV_X1 U11 ( .A(D3_i[4]), .ZN(n66) );
  INV_X1 U12 ( .A(n28), .ZN(n67) );
  INV_X1 U13 ( .A(D3_i[3]), .ZN(n28) );
  NOR4_X1 U14 ( .A1(n60), .A2(n62), .A3(n61), .A4(n30), .ZN(S_FWA[0]) );
  NOR4_X1 U15 ( .A1(n60), .A2(n62), .A3(n61), .A4(n30), .ZN(n102) );
  INV_X1 U16 ( .A(n91), .ZN(n69) );
  OR2_X1 U17 ( .A1(n37), .A2(rAdec_i[0]), .ZN(n93) );
  AOI22_X1 U18 ( .A1(n36), .A2(rAdec_i[4]), .B1(rAdec_i[0]), .B2(n37), .ZN(n49) );
  CLKBUF_X1 U19 ( .A(D3_i[4]), .Z(n70) );
  INV_X1 U20 ( .A(D2_i[1]), .ZN(n94) );
  OAI221_X1 U21 ( .B1(n97), .B2(rAdec_i[1]), .C1(n34), .C2(rAdec_i[3]), .A(n48), .ZN(n47) );
  NAND3_X1 U22 ( .A1(n92), .A2(n93), .A3(n49), .ZN(n46) );
  CLKBUF_X1 U23 ( .A(n30), .Z(n71) );
  INV_X1 U25 ( .A(D3_i[0]), .ZN(n22) );
  NOR3_X1 U26 ( .A1(n31), .A2(n32), .A3(n95), .ZN(S_FWB[0]) );
  NAND2_X1 U27 ( .A1(S_mem_W), .A2(S_mem_LOAD), .ZN(n30) );
  NOR4_X1 U28 ( .A1(n47), .A2(n46), .A3(n30), .A4(n45), .ZN(n101) );
  NOR4_X1 U29 ( .A1(n102), .A2(n50), .A3(n51), .A4(n52), .ZN(S_FWA[1]) );
  INV_X1 U30 ( .A(D3_i[1]), .ZN(n88) );
  INV_X1 U31 ( .A(D3_i[1]), .ZN(n24) );
  OR2_X1 U32 ( .A1(n41), .A2(n39), .ZN(n74) );
  INV_X1 U35 ( .A(S_wb_W), .ZN(n83) );
  INV_X1 U36 ( .A(D3_i[3]), .ZN(n82) );
  NOR3_X1 U41 ( .A1(n101), .A2(n40), .A3(n74), .ZN(S_FWAdec[1]) );
  INV_X1 U42 ( .A(n79), .ZN(n78) );
  NOR3_X1 U43 ( .A1(n31), .A2(n32), .A3(n95), .ZN(n103) );
  OR2_X1 U44 ( .A1(n29), .A2(n30), .ZN(n95) );
  INV_X1 U45 ( .A(D2_i[4]), .ZN(n36) );
  NOR4_X2 U46 ( .A1(n45), .A2(n71), .A3(n46), .A4(n47), .ZN(S_FWAdec[0]) );
  OAI221_X1 U47 ( .B1(n24), .B2(rAdec_i[1]), .C1(n25), .C2(rAdec_i[2]), .A(n43), .ZN(n40) );
  OAI22_X1 U48 ( .A1(rB_i[3]), .A2(n28), .B1(n69), .B2(rB_i[0]), .ZN(n90) );
  NOR2_X1 U49 ( .A1(n75), .A2(n103), .ZN(S_FWB[1]) );
  NAND3_X1 U50 ( .A1(n77), .A2(n76), .A3(n78), .ZN(n75) );
  NAND2_X1 U51 ( .A1(n88), .A2(rB_i[1]), .ZN(n87) );
  AOI21_X1 U52 ( .B1(n82), .B2(rB_i[3]), .A(n83), .ZN(n80) );
  OAI211_X1 U56 ( .C1(n24), .C2(rB_i[1]), .A(n81), .B(n80), .ZN(n79) );
  NAND2_X1 U57 ( .A1(n66), .A2(rB_i[4]), .ZN(n89) );
  OAI21_X1 U58 ( .B1(n73), .B2(rB_i[4]), .A(n89), .ZN(n84) );
  NAND2_X1 U59 ( .A1(n22), .A2(rB_i[0]), .ZN(n86) );
  OAI211_X1 U60 ( .C1(rB_i[2]), .C2(n25), .A(n86), .B(n87), .ZN(n85) );
  NAND2_X1 U61 ( .A1(n25), .A2(rB_i[2]), .ZN(n81) );
  NOR2_X1 U62 ( .A1(n84), .A2(n85), .ZN(n77) );
  AOI22_X1 U63 ( .A1(n66), .A2(rAdec_i[4]), .B1(n22), .B2(rAdec_i[0]), .ZN(n42) );
  OAI221_X1 U64 ( .B1(D3_i[3]), .B2(n44), .C1(n28), .C2(rAdec_i[3]), .A(S_wb_W), .ZN(n39) );
  OAI221_X1 U65 ( .B1(n73), .B2(rAdec_i[4]), .C1(n69), .C2(rAdec_i[0]), .A(n42), .ZN(n41) );
  AOI22_X1 U66 ( .A1(n24), .A2(rAdec_i[1]), .B1(rAdec_i[2]), .B2(n25), .ZN(n43) );
  INV_X1 U67 ( .A(D2_i[4]), .ZN(n96) );
  OAI221_X1 U68 ( .B1(n96), .B2(rA_i[4]), .C1(n37), .C2(rA_i[0]), .A(n64), 
        .ZN(n61) );
  OAI221_X1 U69 ( .B1(n94), .B2(rA_i[1]), .C1(n34), .C2(rA_i[3]), .A(n63), 
        .ZN(n62) );
  OAI221_X1 U70 ( .B1(n36), .B2(rB_i[4]), .C1(n37), .C2(rB_i[0]), .A(n38), 
        .ZN(n31) );
  AOI22_X1 U71 ( .A1(n56), .A2(n65), .B1(D3_i[2]), .B2(n57), .ZN(n58) );
  OAI221_X1 U72 ( .B1(n56), .B2(n65), .C1(n57), .C2(D3_i[2]), .A(n58), .ZN(n51) );
  OAI221_X1 U73 ( .B1(n53), .B2(n70), .C1(n54), .C2(n91), .A(n55), .ZN(n52) );
  AOI22_X1 U74 ( .A1(n53), .A2(n70), .B1(n91), .B2(n54), .ZN(n55) );
  NAND3_X1 U75 ( .A1(n99), .A2(n100), .A3(n35), .ZN(n32) );
  AOI22_X1 U76 ( .A1(n97), .A2(rAdec_i[1]), .B1(rAdec_i[3]), .B2(n34), .ZN(n48) );
  AOI22_X1 U77 ( .A1(n97), .A2(rA_i[1]), .B1(rA_i[3]), .B2(n34), .ZN(n63) );
  AOI22_X1 U78 ( .A1(n96), .A2(rA_i[4]), .B1(rA_i[0]), .B2(n37), .ZN(n64) );
  AOI22_X1 U79 ( .A1(n36), .A2(rB_i[4]), .B1(rB_i[0]), .B2(n37), .ZN(n38) );
  AOI22_X1 U80 ( .A1(n94), .A2(rB_i[1]), .B1(rB_i[3]), .B2(n34), .ZN(n35) );
  INV_X1 U81 ( .A(D2_i[0]), .ZN(n37) );
  INV_X1 U82 ( .A(D2_i[3]), .ZN(n34) );
endmodule


module mem_block ( X_i, LOAD_i, W_o, S_MUX_MEM_i_BAR );
  input [31:0] X_i;
  input [31:0] LOAD_i;
  output [31:0] W_o;
  input S_MUX_MEM_i_BAR;
  wire   S_MUX_MEM_i;
  assign S_MUX_MEM_i = S_MUX_MEM_i_BAR;

  mux21_3 MUXMEM ( .IN0(X_i), .IN1(LOAD_i), .OUT1(W_o), .CTRL_BAR(S_MUX_MEM_i)
         );
endmodule


module mem_regs ( W_i, D3_i, W_o, D3_o, clk, rst );
  input [31:0] W_i;
  input [4:0] D3_i;
  output [31:0] W_o;
  output [4:0] D3_o;
  input clk, rst;


  ff32_SIZE32 W ( .D(W_i), .clk(clk), .rst(rst), .Q(W_o) );
  ff32_SIZE5 D3 ( .D(D3_i), .clk(clk), .rst(rst), .Q(D3_o) );
endmodule


module execute_block ( IMM_i, A_i, rB_i, rC_i, MUXED_B_i, S_MUX_ALUIN_i, 
        FW_X_i, FW_W_i, S_FW_A_i, S_FW_B_i, muxed_dest, muxed_B, S_MUX_DEST_i, 
    .OP({\OP[4] , \OP[3] , \OP[2] , \OP[1] , \OP[0] }), ALUW_i, DOUT, stall_o, 
        Clock, Reset );
  input [31:0] IMM_i;
  input [31:0] A_i;
  input [4:0] rB_i;
  input [4:0] rC_i;
  input [31:0] MUXED_B_i;
  input [31:0] FW_X_i;
  input [31:0] FW_W_i;
  input [1:0] S_FW_A_i;
  input [1:0] S_FW_B_i;
  output [4:0] muxed_dest;
  output [31:0] muxed_B;
  input [1:0] S_MUX_DEST_i;
  input [12:0] ALUW_i;
  output [31:0] DOUT;
  input S_MUX_ALUIN_i, \OP[4] , \OP[3] , \OP[2] , \OP[1] , \OP[0] , Clock,
         Reset;
  output stall_o;
  wire   n6;
  wire   [31:0] FWB2alu;
  wire   [31:0] FWA2alu;

  mux21_0 ALUIN_MUX ( .IN0({muxed_B[31:10], n6, muxed_B[8:0]}), .IN1(IMM_i), 
        .CTRL(S_MUX_ALUIN_i), .OUT1(FWB2alu) );
  real_alu_DATA_SIZE32 ALU ( .IN1(FWA2alu), .IN2(FWB2alu), .ALUW_i(ALUW_i), 
        .DOUT(DOUT), .stall_o(stall_o), .Clock(Clock), .Reset(Reset) );
  mux41_MUX_SIZE5 MUXDEST ( .IN0({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .IN1(rC_i), 
        .IN2(rB_i), .IN3({1'b1, 1'b1, 1'b1, 1'b1, 1'b1}), .CTRL(S_MUX_DEST_i), 
        .OUT1(muxed_dest) );
  mux41_MUX_SIZE32_0 MUX_FWA ( .IN0(A_i), .IN1(FW_X_i), .IN2(FW_W_i), .IN3({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CTRL(S_FW_A_i), 
        .OUT1(FWA2alu) );
  mux41_MUX_SIZE32_1 MUX_FWB ( .IN0(MUXED_B_i), .IN1(FW_X_i), .IN2(FW_W_i), 
        .IN3({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CTRL(S_FW_B_i), .OUT1({muxed_B[31:10], n6, muxed_B[8:0]}) );
  CLKBUF_X1 U5 ( .A(n6), .Z(muxed_B[9]) );
endmodule


module execute_regs ( X_i, S_i, D2_i, X_o, S_o, D2_o, stall_i, clk, rst );
  input [31:0] X_i;
  input [31:0] S_i;
  input [4:0] D2_i;
  output [31:0] X_o;
  output [31:0] S_o;
  output [4:0] D2_o;
  input stall_i, clk, rst;


  ff32_en_SIZE32_3 X ( .D(X_i), .en(1'b1), .clk(clk), .rst(rst), .Q(X_o) );
  ff32_en_SIZE32_2 S ( .D(S_i), .en(1'b1), .clk(clk), .rst(rst), .Q(S_o) );
  ff32_en_SIZE5_1 D2 ( .D(D2_i), .en(1'b1), .clk(clk), .rst(rst), .Q(D2_o) );
endmodule


module decode_regs ( A_i, B_i, rA_i, rB_i, rC_i, IMM_i, ALUW_i, A_o, B_o, rA_o, 
        rB_o, rC_o, IMM_o, ALUW_o, stall_i, clk, rst );
  input [31:0] A_i;
  input [31:0] B_i;
  input [4:0] rA_i;
  input [4:0] rB_i;
  input [4:0] rC_i;
  input [31:0] IMM_i;
  input [12:0] ALUW_i;
  output [31:0] A_o;
  output [31:0] B_o;
  output [4:0] rA_o;
  output [4:0] rB_o;
  output [4:0] rC_o;
  output [31:0] IMM_o;
  output [12:0] ALUW_o;
  input stall_i, clk, rst;
  wire   enable;

  ff32_en_SIZE32_0 A ( .D(A_i), .en(enable), .clk(clk), .rst(rst), .Q(A_o) );
  ff32_en_SIZE32_5 B ( .D(B_i), .en(enable), .clk(clk), .rst(rst), .Q(B_o) );
  ff32_en_SIZE5_0 rA ( .D(rA_i), .en(enable), .clk(clk), .rst(rst), .Q(rA_o)
         );
  ff32_en_SIZE5_3 rB ( .D(rB_i), .en(enable), .clk(clk), .rst(rst), .Q(rB_o)
         );
  ff32_en_SIZE5_2 rC ( .D(rC_i), .en(enable), .clk(clk), .rst(rst), .Q(rC_o)
         );
  ff32_en_SIZE32_4 IMM ( .D(IMM_i), .en(enable), .clk(clk), .rst(rst), .Q(
        IMM_o) );
  ff32_en_SIZE13 ALUW ( .D(ALUW_i), .en(enable), .clk(clk), .rst(rst), .Q(
        ALUW_o) );
  INV_X8 U1 ( .A(stall_i), .ZN(enable) );
endmodule


module dlx_regfile ( Clk, Rst, ENABLE, RD1, RD2, WR, ADD_WR, ADD_RD1, ADD_RD2, 
        DATAIN, OUT1, OUT2 );
  input [4:0] ADD_WR;
  input [4:0] ADD_RD1;
  input [4:0] ADD_RD2;
  input [31:0] DATAIN;
  output [31:0] OUT1;
  output [31:0] OUT2;
  input Clk, Rst, ENABLE, RD1, RD2, WR;
  wire   N4487, n2152, n2184, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n222,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n2087, n2219, n2220,
         n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230,
         n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240,
         n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2601, n2634,
         n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644,
         n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654,
         n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664,
         n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763,
         n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773,
         n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783,
         n3784, net644357, net644358, net644359, net644360, net644361,
         net644362, net644363, net644364, net644365, net644366, net644367,
         net644368, net644369, net644370, net644371, net644372, net644373,
         net644374, net644375, net644376, net644377, net644378, net644379,
         net644380, net644381, net644382, net644383, net644384, net644385,
         net644386, net644387, net644388, net644389, net644390, net644391,
         net644392, net644393, net644394, net644395, net644396, net644397,
         net644398, net644399, net644400, net644401, net644402, net644403,
         net644404, net644405, net644406, net644407, net644408, net644409,
         net644410, net644411, net644412, net644413, net644414, net644415,
         net644416, net644417, net644418, net644419, net644420, net644421,
         net644422, net644423, net644424, net644425, net644426, net644427,
         net644428, net644429, net644430, net644431, net644432, net644433,
         net644434, net644435, net644436, net644437, net644438, net644439,
         net644440, net644441, net644442, net644443, net644444, net644445,
         net644446, net644447, net644448, net644449, net644450, net644451,
         net644452, net644453, net644454, net644455, net644456, net644457,
         net644458, net644459, net644460, net644461, net644462, net644463,
         net644464, net644465, net644466, net644467, net644468, net644469,
         net644470, net644471, net644472, net644473, net644474, net644475,
         net644476, net644477, net644478, net644479, net644480, net644481,
         net644482, net644483, net644484, net644485, net644486, net644487,
         net644488, net644489, net644490, net644491, net644492, net644493,
         net644494, net644495, net644496, net644497, net644498, net644499,
         net644500, net644501, net644502, net644503, net644504, net644505,
         net644506, net644507, net644508, net644509, net644510, net644511,
         net644512, net644513, net644514, net644515, net644516, net644517,
         net644518, net644519, net644520, net644521, net644522, net644523,
         net644524, net644525, net644526, net644527, net644528, net644529,
         net644530, net644531, net644532, net644533, net644534, net644535,
         net644536, net644537, net644538, net644539, net644540, net644541,
         net644542, net644543, net644544, net644545, net644546, net644547,
         net644548, net644549, net644550, net644551, net644552, net644553,
         net644554, net644555, net644556, net644557, net644558, net644559,
         net644560, net644561, net644562, net644563, net644564, net644565,
         net644566, net644567, net644568, net644569, net644570, net644571,
         net644572, net644573, net644574, net644575, net644576, net644577,
         net644578, net644579, net644580, net644581, net644582, net644583,
         net644584, net644585, net644586, net644587, net644588, net644589,
         net644590, net644591, net644592, net644593, net644594, net644595,
         net644596, net644597, net644598, net644599, net644600, net644601,
         net644602, net644603, net644604, net644605, net644606, net644607,
         net644608, net644609, net644610, net644611, net644612, net644613,
         net644614, net644615, net644616, net644617, net644618, net644619,
         net644620, net644621, net644622, net644623, net644624, net644625,
         net644626, net644627, net644628, net644629, net644630, net644631,
         net644632, net644633, net644634, net644635, net644636, net644637,
         net644638, net644639, net644640, net644641, net644642, net644643,
         net644644, net644645, net644646, net644647, net644648, net644649,
         net644650, net644651, net644652, net644653, net644654, net644655,
         net644656, net644657, net644658, net644659, net644660, net644661,
         net644662, net644663, net644664, net644665, net644666, net644667,
         net644668, net644669, net644670, net644671, net644672, net644673,
         net644674, net644675, net644676, net644677, net644678, net644679,
         net644680, net644681, net644682, net644683, net644684, net644685,
         net644686, net644687, net644688, net644689, net644690, net644691,
         net644692, net644693, net644694, net644695, net644696, net644697,
         net644698, net644699, net644700, net644701, net644702, net644703,
         net644704, net644705, net644706, net644707, net644708, net644709,
         net644710, net644711, net644712, net644713, net644714, net644715,
         net644716, net644717, net644718, net644719, net644720, net644721,
         net644722, net644723, net644724, net644725, net644726, net644727,
         net644728, net644729, net644730, net644731, net644732, net644733,
         net644734, net644735, net644736, net644737, net644738, net644739,
         net644740, net644741, net644742, net644743, net644744, net644745,
         net644746, net644747, net644748, net644749, net644750, net644751,
         net644752, net644753, net644754, net644755, net644756, net644757,
         net644758, net644759, net644760, net644761, net644762, net644763,
         net644764, net644765, net644766, net644767, net644768, net644769,
         net644770, net644771, net644772, net644773, net644774, net644775,
         net644776, net644777, net644778, net644779, net644780, net644781,
         net644782, net644783, net644784, net644785, net644786, net644787,
         net644788, net644789, net644790, net644791, net644792, net644793,
         net644794, net644795, net644796, net644797, net644798, net644799,
         net644800, net644801, net644802, net644803, net644804, net644805,
         net644806, net644807, net644808, net644809, net644810, net644811,
         net644812, net644813, net644814, net644815, net644816, net644817,
         net644818, net644819, net644820, net644821, net644822, net644823,
         net644824, net644825, net644826, net644827, net644828, net644829,
         net644830, net644831, net644832, net644833, net644834, net644835,
         net644836, net644837, net644838, net644839, net644840, net644841,
         net644842, net644843, net644844, net644845, net644846, net644847,
         net644848, net644849, net644850, net644851, net644852, net644853,
         net644854, net644855, net644856, net644857, net644858, net644859,
         net644860, net644861, net644862, net644863, net644864, net644865,
         net644866, net644867, net644868, net644869, net644870, net644871,
         net644872, net644873, net644874, net644875, net644876, net644877,
         net644878, net644879, net644880, net644881, net644882, net644883,
         net644884, net644885, net644886, net644887, net644888, net644889,
         net644890, net644891, net644892, net644893, net644894, net644895,
         net644896, net644897, net644898, net644899, net644900, net644901,
         net644902, net644903, net644904, net644905, net644906, net644907,
         net644908, net644909, net644910, net644911, net644912, net644913,
         net644914, net644915, net644916, net644917, net644918, net644919,
         net644920, net644921, net644922, net644923, net644924, net644925,
         net644926, net644927, net644928, net644929, net644930, net644931,
         net644932, net644933, n1662, n1663, n1664, n1666, n1668, n1670, n1672,
         n1674, n1676, n1678, n1680, n1682, n1684, n1686, n1688, n1690, n1692,
         n1694, n1696, n1698, n1700, n1702, n1704, n1706, n1708, n1710, n1712,
         n1714, n1716, n1718, n1720, n1722, n1724, n1726, n1728, n1729, n1730,
         n1731, n1733, n1735, n1736, n1768, n1769, n1770, n1772, n1773, n1805,
         n1806, n1807, n1808, n1811, n1812, n1843, n1844, n1846, n1847, n1848,
         n1850, n1852, n1853, n1885, n1886, n1917, n1918, n1919, n1921, n1922,
         n1954, n1956, n1957, n1990, n1991, n2023, n2024, n2025, n2027, n2028,
         n2060, n2062, n2063, n3888, n3889, n3892, n3893, n3924, n3926, n3927,
         n3959, n3961, n3962, n3994, n3995, n3996, n3997, n4000, n4001, n4033,
         n4035, n4036, n4068, n4069, n4073, n4074, n4106, n4107, n4108, n4110,
         n4111, n4143, n4145, n4146, n4178, n4180, n4181, n4182, n4183, n4184,
         n4185, n4186, n4187, n4188, n4189, n4190, n4192, n4194, n4195, n4196,
         n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4207,
         n4208, n4209, n4210, n4211, n4212, n4214, n4215, n4216, n4217, n4218,
         n4219, n4220, n4221, n4223, n4224, n4225, n4226, n4228, n4229, n4231,
         n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241,
         n4243, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4254, n4255,
         n4256, n4257, n4258, n4259, n4260, n4261, n4264, n4265, n4266, n4267,
         n4270, n4271, n4272, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4294, n4295,
         n4296, n4297, n4300, n4301, n4302, n4306, n4307, n4308, n4309, n4310,
         n4311, n4312, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321,
         n4324, n4325, n4326, n4327, n4330, n4331, n4332, n4336, n4337, n4338,
         n4339, n4340, n4341, n4342, n4344, n4345, n4346, n4347, n4348, n4349,
         n4350, n4351, n4354, n4355, n4356, n4357, n4360, n4361, n4362, n4366,
         n4367, n4368, n4369, n4370, n4371, n4372, n4374, n4375, n4376, n4377,
         n4378, n4379, n4380, n4381, n4384, n4385, n4386, n4387, n4390, n4391,
         n4392, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4404, n4405,
         n4406, n4407, n4408, n4409, n4410, n4411, n4414, n4415, n4416, n4417,
         n4420, n4421, n4422, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4444, n4445,
         n4446, n4447, n4450, n4451, n4452, n4456, n4457, n4458, n4459, n4460,
         n4461, n4462, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471,
         n4474, n4475, n4476, n4477, n4480, n4481, n4482, n4486, n4487, n4488,
         n4489, n4490, n4491, n4492, n4494, n4495, n4496, n4497, n4498, n4499,
         n4500, n4501, n4504, n4505, n4506, n4507, n4510, n4511, n4512, n4516,
         n4517, n4518, n4519, n4520, n4521, n4522, n4524, n4525, n4526, n4527,
         n4528, n4529, n4530, n4531, n4534, n4535, n4536, n4537, n4540, n4541,
         n4542, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4554, n4555,
         n4556, n4557, n4558, n4559, n4560, n4561, n4564, n4565, n4566, n4567,
         n4570, n4571, n4572, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4594, n4595,
         n4596, n4597, n4600, n4601, n4602, n4606, n4607, n4608, n4609, n4610,
         n4611, n4612, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621,
         n4624, n4625, n4626, n4627, n4630, n4631, n4632, n4636, n4637, n4638,
         n4639, n4640, n4641, n4642, n4644, n4645, n4646, n4647, n4648, n4649,
         n4650, n4651, n4654, n4655, n4656, n4657, n4660, n4661, n4662, n4666,
         n4667, n4668, n4669, n4670, n4671, n4672, n4674, n4675, n4676, n4677,
         n4678, n4679, n4680, n4681, n4684, n4685, n4686, n4687, n4690, n4691,
         n4692, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4704, n4705,
         n4706, n4707, n4708, n4709, n4710, n4711, n4714, n4715, n4716, n4717,
         n4720, n4721, n4722, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4744, n4745,
         n4746, n4747, n4750, n4751, n4752, n4756, n4757, n4758, n4759, n4760,
         n4761, n4762, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771,
         n4774, n4775, n4776, n4777, n4780, n4781, n4782, n4786, n4787, n4788,
         n4789, n4790, n4791, n4792, n4794, n4795, n4796, n4797, n4798, n4799,
         n4800, n4801, n4804, n4805, n4806, n4807, n4810, n4811, n4812, n4816,
         n4817, n4818, n4819, n4820, n4821, n4822, n4824, n4825, n4826, n4827,
         n4828, n4829, n4830, n4831, n4834, n4835, n4836, n4837, n4840, n4841,
         n4842, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4854, n4855,
         n4856, n4857, n4858, n4859, n4860, n4861, n4864, n4865, n4866, n4867,
         n4870, n4871, n4872, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4894, n4895,
         n4896, n4897, n4900, n4901, n4902, n4906, n4907, n4908, n4909, n4910,
         n4911, n4912, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921,
         n4924, n4925, n4926, n4927, n4930, n4931, n4932, n4936, n4937, n4938,
         n4939, n4940, n4941, n4942, n4944, n4945, n4946, n4947, n4948, n4949,
         n4950, n4951, n4954, n4955, n4956, n4957, n4960, n4961, n4962, n4966,
         n4967, n4968, n4969, n4970, n4971, n4972, n4974, n4975, n4976, n4977,
         n4978, n4979, n4980, n4981, n4984, n4985, n4986, n4987, n4990, n4991,
         n4992, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5004, n5005,
         n5006, n5007, n5008, n5009, n5010, n5011, n5014, n5015, n5016, n5017,
         n5020, n5021, n5022, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5044, n5045,
         n5046, n5047, n5050, n5051, n5052, n5056, n5057, n5058, n5059, n5060,
         n5061, n5062, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071,
         n5074, n5075, n5076, n5077, n5080, n5081, n5082, n5086, n5087, n5088,
         n5089, n5090, n5091, n5092, n5094, n5095, n5096, n5097, n5098, n5099,
         n5100, n5101, n5104, n5105, n5106, n5107, n5110, n5111, n5112, n5116,
         n5117, n5118, n5119, n5120, n5121, n5122, n5124, n5125, n5126, n5127,
         n5128, n5129, n5130, n5131, n5132, n5135, n5136, n5137, n5138, n5140,
         n5141, n5142, n5143, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163,
         n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173,
         n5175, n5176, n5177, n5178, n5179, n5181, n5182, n5184, n5185, n5186,
         n5187, n5189, n5190, n5191, n5192, n5194, n5195, n5196, n5197, n5198,
         n5199, n5200, n5201, n5202, n5205, n5206, n5207, n5208, n5209, n5210,
         n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5219, n5220, n5221,
         n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231,
         n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241,
         n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943,
         n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953,
         n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963,
         n5964, n5966, n5967, n5968, n5969, n5971, n5972, n5973, n5974, n5975,
         n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n3880,
         n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3890, n3891, n3894,
         n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904,
         n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914,
         n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3925,
         n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937,
         n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947,
         n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957,
         n3958, n3960, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970,
         n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980,
         n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990,
         n3991, n3992, n3993, n3998, n3999, n4002, n4003, n4004, n4005, n4006,
         n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016,
         n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026,
         n4027, n4028, n4029, n4030, n4031, n4032, n4034, n4037, n4038, n4039,
         n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049,
         n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059,
         n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4070, n4071,
         n4072, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083,
         n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093,
         n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103,
         n4104, n4105, n4109, n4112, n4113, n4114, n4115, n4116, n4117, n4118,
         n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128,
         n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138,
         n4139, n4140, n4141, n4142, n4144, n4147, n4148, n4149, n4150, n4151,
         n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161,
         n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171,
         n4172, n4173, n4174, n4175, n4176, n4177, n4179, n4191, n4193, n4206,
         n4213, n4222, n4227, n4230, n4242, n4244, n4245, n4253, n4262, n4263,
         n4268, n4269, n4273, n4274, n4275, n4283, n4292, n4293, n4298, n4299,
         n4303, n4304, n4305, n4313, n4322, n4323, n4328, n4329, n4333, n4334,
         n4335, n4343, n4352, n4353, n4358, n4359, n4363, n4364, n4365, n4373,
         n4382, n4383, n4388, n4389, n4393, n4394, n4395, n4403, n4412, n4413,
         n4418, n4419, n4423, n4424, n4425, n4433, n4442, n4443, n4448, n4449,
         n4453, n4454, n4455, n4463, n4472, n4473, n4478, n4479, n4483, n4484,
         n4485, n4493, n4502, n4503, n4508, n4509, n4513, n4514, n4515, n4523,
         n4532, n4533, n4538, n4539, n4543, n4544, n4545, n4553, n4562, n4563,
         n4568, n4569, n4573, n4574, n4575, n4583, n4592, n4593, n4598, n4599,
         n4603, n4604, n4605, n4613, n4622, n4623, n4628, n4629, n4633, n4634,
         n4635, n4643, n4652, n4653, n4658, n4659, n4663, n4664, n4665, n4673,
         n4682, n4683, n4688, n4689, n4693, n4694, n4695, n4703, n4712, n4713,
         n4718, n4719, n4723, n4724, n4725, n4733, n4742, n4743, n4748, n4749,
         n4753, n4754, n4755, n4763, n4772, n4773, n4778, n4779, n4783, n4784,
         n4785, n4793, n4802, n4803, n4808, n4809, n4813, n4814, n4815, n4823,
         n4832, n4833, n4838, n4839, n4843, n4844, n4845, n4853, n4862, n4863,
         n4868, n4869, n4873, n4874, n4875, n4883, n4892, n4893, n4898, n4899,
         n4903, n4904, n4905, n4913, n4922, n4923, n4928, n4929, n4933, n4934,
         n4935, n4943, n4952, n4953, n4958, n4959, n4963, n4964, n4965, n4973,
         n4982, n4983, n4988, n4989, n4993, n4994, n4995, n5003, n5012, n5013,
         n5018, n5019, n5023, n5024, n5025, n5033, n5042, n5043, n5048, n5049,
         n5053, n5054, n5055, n5063, n5072, n5073, n5078, n5079, n5083, n5084,
         n5085, n5093, n5102, n5103, n5108, n5109, n5113, n5114, n5115, n5123,
         n5133, n5134, n5139, n5144, n5145, n5153, n5174, n5180, n5183, n5188,
         n5193, n5203, n5204, n5218, n5252, n5933, n5965, n5970, n5985, n5986,
         n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996,
         n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006,
         n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016,
         n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026,
         n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036,
         n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046,
         n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056,
         n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066,
         n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076,
         n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086,
         n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096,
         n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106,
         n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116,
         n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126,
         n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136,
         n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146,
         n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156,
         n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166,
         n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176,
         n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186,
         n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196,
         n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206,
         n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216,
         n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226,
         n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236,
         n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246,
         n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256,
         n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266,
         n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276,
         n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286,
         n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296,
         n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306,
         n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316,
         n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326,
         n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336,
         n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346,
         n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356,
         n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366,
         n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376,
         n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386,
         n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396,
         n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406,
         n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416,
         n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426,
         n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436,
         n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446;
  assign N4487 = Rst;

  DFF_X1 \REGISTERS_reg[1][31]  ( .D(n3751), .CK(Clk), .Q(net644933), .QN(
        n6055) );
  DFF_X1 \REGISTERS_reg[1][30]  ( .D(n3750), .CK(Clk), .Q(net644932), .QN(
        n6054) );
  DFF_X1 \REGISTERS_reg[1][29]  ( .D(n3749), .CK(Clk), .Q(net644931), .QN(
        n6053) );
  DFF_X1 \REGISTERS_reg[1][28]  ( .D(n3748), .CK(Clk), .Q(net644930), .QN(
        n6052) );
  DFF_X1 \REGISTERS_reg[1][27]  ( .D(n3747), .CK(Clk), .Q(net644929), .QN(
        n6051) );
  DFF_X1 \REGISTERS_reg[1][26]  ( .D(n3746), .CK(Clk), .Q(net644928), .QN(
        n6050) );
  DFF_X1 \REGISTERS_reg[1][25]  ( .D(n3745), .CK(Clk), .Q(net644927), .QN(
        n6049) );
  DFF_X1 \REGISTERS_reg[1][24]  ( .D(n3744), .CK(Clk), .Q(net644926), .QN(
        n6048) );
  DFF_X1 \REGISTERS_reg[1][23]  ( .D(n3743), .CK(Clk), .Q(net644925), .QN(
        n6047) );
  DFF_X1 \REGISTERS_reg[1][22]  ( .D(n3742), .CK(Clk), .Q(net644924), .QN(
        n6046) );
  DFF_X1 \REGISTERS_reg[1][21]  ( .D(n3741), .CK(Clk), .Q(net644923), .QN(
        n6045) );
  DFF_X1 \REGISTERS_reg[1][20]  ( .D(n3740), .CK(Clk), .Q(net644922), .QN(
        n6044) );
  DFF_X1 \REGISTERS_reg[1][19]  ( .D(n3739), .CK(Clk), .Q(net644921), .QN(
        n6043) );
  DFF_X1 \REGISTERS_reg[1][18]  ( .D(n3738), .CK(Clk), .Q(net644920), .QN(
        n6042) );
  DFF_X1 \REGISTERS_reg[1][17]  ( .D(n3737), .CK(Clk), .Q(net644919), .QN(
        n6041) );
  DFF_X1 \REGISTERS_reg[1][16]  ( .D(n3736), .CK(Clk), .Q(net644918), .QN(
        n6040) );
  DFF_X1 \REGISTERS_reg[1][15]  ( .D(n3735), .CK(Clk), .Q(net644917), .QN(
        n6039) );
  DFF_X1 \REGISTERS_reg[1][14]  ( .D(n3734), .CK(Clk), .Q(net644916), .QN(
        n6038) );
  DFF_X1 \REGISTERS_reg[1][13]  ( .D(n3733), .CK(Clk), .Q(net644915), .QN(
        n6037) );
  DFF_X1 \REGISTERS_reg[1][12]  ( .D(n3732), .CK(Clk), .Q(net644914), .QN(
        n6036) );
  DFF_X1 \REGISTERS_reg[1][11]  ( .D(n3731), .CK(Clk), .Q(net644913), .QN(
        n6035) );
  DFF_X1 \REGISTERS_reg[1][10]  ( .D(n3730), .CK(Clk), .Q(net644912), .QN(
        n6034) );
  DFF_X1 \REGISTERS_reg[1][9]  ( .D(n3729), .CK(Clk), .Q(net644911), .QN(n6033) );
  DFF_X1 \REGISTERS_reg[1][8]  ( .D(n3728), .CK(Clk), .Q(net644910), .QN(n6032) );
  DFF_X1 \REGISTERS_reg[1][7]  ( .D(n3727), .CK(Clk), .Q(net644909), .QN(n6031) );
  DFF_X1 \REGISTERS_reg[1][6]  ( .D(n3726), .CK(Clk), .Q(net644908), .QN(n6030) );
  DFF_X1 \REGISTERS_reg[1][5]  ( .D(n3725), .CK(Clk), .Q(net644907), .QN(n6029) );
  DFF_X1 \REGISTERS_reg[1][4]  ( .D(n3724), .CK(Clk), .Q(net644906), .QN(n6028) );
  DFF_X1 \REGISTERS_reg[1][3]  ( .D(n3723), .CK(Clk), .Q(net644905), .QN(n6027) );
  DFF_X1 \REGISTERS_reg[1][2]  ( .D(n3722), .CK(Clk), .Q(net644904), .QN(n6026) );
  DFF_X1 \REGISTERS_reg[1][1]  ( .D(n3721), .CK(Clk), .Q(net644903), .QN(n6025) );
  DFF_X1 \REGISTERS_reg[1][0]  ( .D(n3720), .CK(Clk), .Q(net644902), .QN(n6346) );
  DFF_X1 \REGISTERS_reg[2][31]  ( .D(n3719), .CK(Clk), .Q(n3949), .QN(n577) );
  DFF_X1 \REGISTERS_reg[2][30]  ( .D(n3718), .CK(Clk), .Q(n3948), .QN(n578) );
  DFF_X1 \REGISTERS_reg[2][29]  ( .D(n3717), .CK(Clk), .Q(n3947), .QN(n579) );
  DFF_X1 \REGISTERS_reg[2][28]  ( .D(n3716), .CK(Clk), .Q(n3946), .QN(n580) );
  DFF_X1 \REGISTERS_reg[2][27]  ( .D(n3715), .CK(Clk), .Q(n3945), .QN(n581) );
  DFF_X1 \REGISTERS_reg[2][26]  ( .D(n3714), .CK(Clk), .Q(n3944), .QN(n582) );
  DFF_X1 \REGISTERS_reg[2][25]  ( .D(n3713), .CK(Clk), .Q(n3943), .QN(n583) );
  DFF_X1 \REGISTERS_reg[2][24]  ( .D(n3712), .CK(Clk), .Q(n3942), .QN(n584) );
  DFF_X1 \REGISTERS_reg[2][23]  ( .D(n3711), .CK(Clk), .Q(n3941), .QN(n585) );
  DFF_X1 \REGISTERS_reg[2][22]  ( .D(n3710), .CK(Clk), .Q(n3940), .QN(n586) );
  DFF_X1 \REGISTERS_reg[2][21]  ( .D(n3709), .CK(Clk), .Q(n3939), .QN(n587) );
  DFF_X1 \REGISTERS_reg[2][20]  ( .D(n3708), .CK(Clk), .Q(n3938), .QN(n588) );
  DFF_X1 \REGISTERS_reg[2][19]  ( .D(n3707), .CK(Clk), .Q(n3937), .QN(n589) );
  DFF_X1 \REGISTERS_reg[2][18]  ( .D(n3706), .CK(Clk), .Q(n3936), .QN(n590) );
  DFF_X1 \REGISTERS_reg[2][17]  ( .D(n3705), .CK(Clk), .Q(n3935), .QN(n591) );
  DFF_X1 \REGISTERS_reg[2][16]  ( .D(n3704), .CK(Clk), .Q(n3934), .QN(n592) );
  DFF_X1 \REGISTERS_reg[2][15]  ( .D(n3703), .CK(Clk), .Q(n3933), .QN(n593) );
  DFF_X1 \REGISTERS_reg[2][14]  ( .D(n3702), .CK(Clk), .Q(n3932), .QN(n594) );
  DFF_X1 \REGISTERS_reg[2][13]  ( .D(n3701), .CK(Clk), .Q(n3931), .QN(n595) );
  DFF_X1 \REGISTERS_reg[2][12]  ( .D(n3700), .CK(Clk), .Q(n3930), .QN(n596) );
  DFF_X1 \REGISTERS_reg[2][11]  ( .D(n3699), .CK(Clk), .Q(n3929), .QN(n597) );
  DFF_X1 \REGISTERS_reg[2][10]  ( .D(n3698), .CK(Clk), .Q(n3928), .QN(n598) );
  DFF_X1 \REGISTERS_reg[2][9]  ( .D(n3697), .CK(Clk), .Q(n3925), .QN(n599) );
  DFF_X1 \REGISTERS_reg[2][8]  ( .D(n3696), .CK(Clk), .Q(n3923), .QN(n600) );
  DFF_X1 \REGISTERS_reg[2][7]  ( .D(n3695), .CK(Clk), .Q(n3922), .QN(n601) );
  DFF_X1 \REGISTERS_reg[2][6]  ( .D(n3694), .CK(Clk), .Q(n3921), .QN(n602) );
  DFF_X1 \REGISTERS_reg[2][5]  ( .D(n3693), .CK(Clk), .Q(n3920), .QN(n603) );
  DFF_X1 \REGISTERS_reg[2][4]  ( .D(n3692), .CK(Clk), .Q(n3919), .QN(n604) );
  DFF_X1 \REGISTERS_reg[2][3]  ( .D(n3691), .CK(Clk), .Q(n3918), .QN(n605) );
  DFF_X1 \REGISTERS_reg[2][2]  ( .D(n3690), .CK(Clk), .Q(n3917), .QN(n606) );
  DFF_X1 \REGISTERS_reg[2][1]  ( .D(n3689), .CK(Clk), .Q(n3916), .QN(n607) );
  DFF_X1 \REGISTERS_reg[2][0]  ( .D(n3688), .CK(Clk), .Q(net644901), .QN(n6345) );
  DFF_X1 \REGISTERS_reg[3][31]  ( .D(n3687), .CK(Clk), .Q(net644900), .QN(
        n6024) );
  DFF_X1 \REGISTERS_reg[3][30]  ( .D(n3686), .CK(Clk), .Q(net644899), .QN(
        n6023) );
  DFF_X1 \REGISTERS_reg[3][29]  ( .D(n3685), .CK(Clk), .Q(net644898), .QN(
        n6022) );
  DFF_X1 \REGISTERS_reg[3][28]  ( .D(n3684), .CK(Clk), .Q(net644897), .QN(
        n6021) );
  DFF_X1 \REGISTERS_reg[3][27]  ( .D(n3683), .CK(Clk), .Q(net644896), .QN(
        n6020) );
  DFF_X1 \REGISTERS_reg[3][26]  ( .D(n3682), .CK(Clk), .Q(net644895), .QN(
        n6019) );
  DFF_X1 \REGISTERS_reg[3][25]  ( .D(n3681), .CK(Clk), .Q(net644894), .QN(
        n6018) );
  DFF_X1 \REGISTERS_reg[3][24]  ( .D(n3680), .CK(Clk), .Q(net644893), .QN(
        n6017) );
  DFF_X1 \REGISTERS_reg[3][23]  ( .D(n3679), .CK(Clk), .Q(net644892), .QN(
        n6016) );
  DFF_X1 \REGISTERS_reg[3][22]  ( .D(n3678), .CK(Clk), .Q(net644891), .QN(
        n6015) );
  DFF_X1 \REGISTERS_reg[3][21]  ( .D(n3677), .CK(Clk), .Q(net644890), .QN(
        n6014) );
  DFF_X1 \REGISTERS_reg[3][20]  ( .D(n3676), .CK(Clk), .Q(net644889), .QN(
        n6013) );
  DFF_X1 \REGISTERS_reg[3][19]  ( .D(n3675), .CK(Clk), .Q(net644888), .QN(
        n6012) );
  DFF_X1 \REGISTERS_reg[3][18]  ( .D(n3674), .CK(Clk), .Q(net644887), .QN(
        n6011) );
  DFF_X1 \REGISTERS_reg[3][17]  ( .D(n3673), .CK(Clk), .Q(net644886), .QN(
        n6010) );
  DFF_X1 \REGISTERS_reg[3][16]  ( .D(n3672), .CK(Clk), .Q(net644885), .QN(
        n6009) );
  DFF_X1 \REGISTERS_reg[3][15]  ( .D(n3671), .CK(Clk), .Q(net644884), .QN(
        n6008) );
  DFF_X1 \REGISTERS_reg[3][14]  ( .D(n3670), .CK(Clk), .Q(net644883), .QN(
        n6007) );
  DFF_X1 \REGISTERS_reg[3][13]  ( .D(n3669), .CK(Clk), .Q(net644882), .QN(
        n6006) );
  DFF_X1 \REGISTERS_reg[3][12]  ( .D(n3668), .CK(Clk), .Q(net644881), .QN(
        n6005) );
  DFF_X1 \REGISTERS_reg[3][11]  ( .D(n3667), .CK(Clk), .Q(net644880), .QN(
        n6004) );
  DFF_X1 \REGISTERS_reg[3][10]  ( .D(n3666), .CK(Clk), .Q(net644879), .QN(
        n6003) );
  DFF_X1 \REGISTERS_reg[3][9]  ( .D(n3665), .CK(Clk), .Q(net644878), .QN(n6002) );
  DFF_X1 \REGISTERS_reg[3][8]  ( .D(n3664), .CK(Clk), .Q(net644877), .QN(n6001) );
  DFF_X1 \REGISTERS_reg[3][7]  ( .D(n3663), .CK(Clk), .Q(net644876), .QN(n6000) );
  DFF_X1 \REGISTERS_reg[3][6]  ( .D(n3662), .CK(Clk), .Q(net644875), .QN(n5999) );
  DFF_X1 \REGISTERS_reg[3][5]  ( .D(n3661), .CK(Clk), .Q(net644874), .QN(n5998) );
  DFF_X1 \REGISTERS_reg[3][4]  ( .D(n3660), .CK(Clk), .Q(net644873), .QN(n5997) );
  DFF_X1 \REGISTERS_reg[3][3]  ( .D(n3659), .CK(Clk), .Q(net644872), .QN(n5996) );
  DFF_X1 \REGISTERS_reg[3][2]  ( .D(n3658), .CK(Clk), .Q(net644871), .QN(n5995) );
  DFF_X1 \REGISTERS_reg[3][1]  ( .D(n3657), .CK(Clk), .Q(net644870), .QN(n5994) );
  DFF_X1 \REGISTERS_reg[3][0]  ( .D(n3656), .CK(Clk), .Q(net644869), .QN(n6354) );
  DFF_X1 \REGISTERS_reg[4][31]  ( .D(n3655), .CK(Clk), .Q(n388), .QN(n4413) );
  DFF_X1 \REGISTERS_reg[4][30]  ( .D(n3654), .CK(Clk), .Q(n391), .QN(n4412) );
  DFF_X1 \REGISTERS_reg[4][29]  ( .D(n3653), .CK(Clk), .Q(n394), .QN(n4403) );
  DFF_X1 \REGISTERS_reg[4][28]  ( .D(n3652), .CK(Clk), .Q(n397), .QN(n4395) );
  DFF_X1 \REGISTERS_reg[4][27]  ( .D(n3651), .CK(Clk), .Q(n400), .QN(n4394) );
  DFF_X1 \REGISTERS_reg[4][26]  ( .D(n3650), .CK(Clk), .Q(n403), .QN(n4393) );
  DFF_X1 \REGISTERS_reg[4][25]  ( .D(n3649), .CK(Clk), .Q(n406), .QN(n4389) );
  DFF_X1 \REGISTERS_reg[4][24]  ( .D(n3648), .CK(Clk), .Q(n409), .QN(n4388) );
  DFF_X1 \REGISTERS_reg[4][23]  ( .D(n3647), .CK(Clk), .Q(n412), .QN(n4383) );
  DFF_X1 \REGISTERS_reg[4][22]  ( .D(n3646), .CK(Clk), .Q(n415), .QN(n4382) );
  DFF_X1 \REGISTERS_reg[4][21]  ( .D(n3645), .CK(Clk), .Q(n418), .QN(n4373) );
  DFF_X1 \REGISTERS_reg[4][20]  ( .D(n3644), .CK(Clk), .Q(n421), .QN(n4365) );
  DFF_X1 \REGISTERS_reg[4][19]  ( .D(n3643), .CK(Clk), .Q(n424), .QN(n4364) );
  DFF_X1 \REGISTERS_reg[4][18]  ( .D(n3642), .CK(Clk), .Q(n427), .QN(n4363) );
  DFF_X1 \REGISTERS_reg[4][17]  ( .D(n3641), .CK(Clk), .Q(n430), .QN(n4359) );
  DFF_X1 \REGISTERS_reg[4][16]  ( .D(n3640), .CK(Clk), .Q(n433), .QN(n4358) );
  DFF_X1 \REGISTERS_reg[4][15]  ( .D(n3639), .CK(Clk), .Q(n436), .QN(n4353) );
  DFF_X1 \REGISTERS_reg[4][14]  ( .D(n3638), .CK(Clk), .Q(n439), .QN(n4352) );
  DFF_X1 \REGISTERS_reg[4][13]  ( .D(n3637), .CK(Clk), .Q(n442), .QN(n4343) );
  DFF_X1 \REGISTERS_reg[4][12]  ( .D(n3636), .CK(Clk), .Q(n445), .QN(n4335) );
  DFF_X1 \REGISTERS_reg[4][11]  ( .D(n3635), .CK(Clk), .Q(n448), .QN(n4334) );
  DFF_X1 \REGISTERS_reg[4][10]  ( .D(n3634), .CK(Clk), .Q(n451), .QN(n4333) );
  DFF_X1 \REGISTERS_reg[4][9]  ( .D(n3633), .CK(Clk), .Q(n454), .QN(n4329) );
  DFF_X1 \REGISTERS_reg[4][8]  ( .D(n3632), .CK(Clk), .Q(n457), .QN(n4328) );
  DFF_X1 \REGISTERS_reg[4][7]  ( .D(n3631), .CK(Clk), .Q(n460), .QN(n4323) );
  DFF_X1 \REGISTERS_reg[4][6]  ( .D(n3630), .CK(Clk), .Q(n463), .QN(n4322) );
  DFF_X1 \REGISTERS_reg[4][5]  ( .D(n3629), .CK(Clk), .Q(n466), .QN(n4313) );
  DFF_X1 \REGISTERS_reg[4][4]  ( .D(n3628), .CK(Clk), .Q(n469), .QN(n4305) );
  DFF_X1 \REGISTERS_reg[4][3]  ( .D(n3627), .CK(Clk), .Q(n472), .QN(n4304) );
  DFF_X1 \REGISTERS_reg[4][2]  ( .D(n3626), .CK(Clk), .Q(n475), .QN(n4303) );
  DFF_X1 \REGISTERS_reg[4][1]  ( .D(n3625), .CK(Clk), .Q(n478), .QN(n4299) );
  DFF_X1 \REGISTERS_reg[4][0]  ( .D(n3624), .CK(Clk), .Q(net644868), .QN(n6353) );
  DFF_X1 \REGISTERS_reg[5][31]  ( .D(n3623), .CK(Clk), .Q(n4058), .QN(n3784)
         );
  DFF_X1 \REGISTERS_reg[5][30]  ( .D(n3622), .CK(Clk), .Q(n4055), .QN(n3783)
         );
  DFF_X1 \REGISTERS_reg[5][29]  ( .D(n3621), .CK(Clk), .Q(n4052), .QN(n3782)
         );
  DFF_X1 \REGISTERS_reg[5][28]  ( .D(n3620), .CK(Clk), .Q(n4049), .QN(n3781)
         );
  DFF_X1 \REGISTERS_reg[5][27]  ( .D(n3619), .CK(Clk), .Q(n4046), .QN(n3780)
         );
  DFF_X1 \REGISTERS_reg[5][26]  ( .D(n3618), .CK(Clk), .Q(n4043), .QN(n3779)
         );
  DFF_X1 \REGISTERS_reg[5][25]  ( .D(n3617), .CK(Clk), .Q(n4040), .QN(n3778)
         );
  DFF_X1 \REGISTERS_reg[5][24]  ( .D(n3616), .CK(Clk), .Q(n4037), .QN(n3777)
         );
  DFF_X1 \REGISTERS_reg[5][23]  ( .D(n3615), .CK(Clk), .Q(n4031), .QN(n3776)
         );
  DFF_X1 \REGISTERS_reg[5][22]  ( .D(n3614), .CK(Clk), .Q(n4028), .QN(n3775)
         );
  DFF_X1 \REGISTERS_reg[5][21]  ( .D(n3613), .CK(Clk), .Q(n4025), .QN(n3774)
         );
  DFF_X1 \REGISTERS_reg[5][20]  ( .D(n3612), .CK(Clk), .Q(n4022), .QN(n3773)
         );
  DFF_X1 \REGISTERS_reg[5][19]  ( .D(n3611), .CK(Clk), .Q(n4019), .QN(n3772)
         );
  DFF_X1 \REGISTERS_reg[5][18]  ( .D(n3610), .CK(Clk), .Q(n4016), .QN(n3771)
         );
  DFF_X1 \REGISTERS_reg[5][17]  ( .D(n3609), .CK(Clk), .Q(n4013), .QN(n3770)
         );
  DFF_X1 \REGISTERS_reg[5][16]  ( .D(n3608), .CK(Clk), .Q(n4010), .QN(n3769)
         );
  DFF_X1 \REGISTERS_reg[5][15]  ( .D(n3607), .CK(Clk), .Q(n4007), .QN(n3768)
         );
  DFF_X1 \REGISTERS_reg[5][14]  ( .D(n3606), .CK(Clk), .Q(n4004), .QN(n3767)
         );
  DFF_X1 \REGISTERS_reg[5][13]  ( .D(n3605), .CK(Clk), .Q(n3999), .QN(n3766)
         );
  DFF_X1 \REGISTERS_reg[5][12]  ( .D(n3604), .CK(Clk), .Q(n3992), .QN(n3765)
         );
  DFF_X1 \REGISTERS_reg[5][11]  ( .D(n3603), .CK(Clk), .Q(n3989), .QN(n3764)
         );
  DFF_X1 \REGISTERS_reg[5][10]  ( .D(n3602), .CK(Clk), .Q(n3986), .QN(n3763)
         );
  DFF_X1 \REGISTERS_reg[5][9]  ( .D(n3601), .CK(Clk), .Q(n3983), .QN(n3762) );
  DFF_X1 \REGISTERS_reg[5][8]  ( .D(n3600), .CK(Clk), .Q(n3980), .QN(n3761) );
  DFF_X1 \REGISTERS_reg[5][7]  ( .D(n3599), .CK(Clk), .Q(n3977), .QN(n3760) );
  DFF_X1 \REGISTERS_reg[5][6]  ( .D(n3598), .CK(Clk), .Q(n3974), .QN(n3759) );
  DFF_X1 \REGISTERS_reg[5][5]  ( .D(n3597), .CK(Clk), .Q(n3971), .QN(n3758) );
  DFF_X1 \REGISTERS_reg[5][4]  ( .D(n3596), .CK(Clk), .Q(n3968), .QN(n3757) );
  DFF_X1 \REGISTERS_reg[5][3]  ( .D(n3595), .CK(Clk), .Q(n3965), .QN(n3756) );
  DFF_X1 \REGISTERS_reg[5][2]  ( .D(n3594), .CK(Clk), .Q(n3960), .QN(n3755) );
  DFF_X1 \REGISTERS_reg[5][1]  ( .D(n3593), .CK(Clk), .Q(n3956), .QN(n3754) );
  DFF_X1 \REGISTERS_reg[5][0]  ( .D(n3592), .CK(Clk), .Q(net644867), .QN(n6344) );
  DFF_X1 \REGISTERS_reg[6][31]  ( .D(n3591), .CK(Clk), .Q(net644866), .QN(
        n6336) );
  DFF_X1 \REGISTERS_reg[6][30]  ( .D(n3590), .CK(Clk), .Q(net644865), .QN(
        n6335) );
  DFF_X1 \REGISTERS_reg[6][29]  ( .D(n3589), .CK(Clk), .Q(net644864), .QN(
        n6334) );
  DFF_X1 \REGISTERS_reg[6][28]  ( .D(n3588), .CK(Clk), .Q(net644863), .QN(
        n6333) );
  DFF_X1 \REGISTERS_reg[6][27]  ( .D(n3587), .CK(Clk), .Q(net644862), .QN(
        n6332) );
  DFF_X1 \REGISTERS_reg[6][26]  ( .D(n3586), .CK(Clk), .Q(net644861), .QN(
        n6331) );
  DFF_X1 \REGISTERS_reg[6][25]  ( .D(n3585), .CK(Clk), .Q(net644860), .QN(
        n6330) );
  DFF_X1 \REGISTERS_reg[6][24]  ( .D(n3584), .CK(Clk), .Q(net644859), .QN(
        n6329) );
  DFF_X1 \REGISTERS_reg[6][23]  ( .D(n3583), .CK(Clk), .Q(net644858), .QN(
        n6328) );
  DFF_X1 \REGISTERS_reg[6][22]  ( .D(n3582), .CK(Clk), .Q(net644857), .QN(
        n6327) );
  DFF_X1 \REGISTERS_reg[6][21]  ( .D(n3581), .CK(Clk), .Q(net644856), .QN(
        n6326) );
  DFF_X1 \REGISTERS_reg[6][20]  ( .D(n3580), .CK(Clk), .Q(net644855), .QN(
        n6325) );
  DFF_X1 \REGISTERS_reg[6][19]  ( .D(n3579), .CK(Clk), .Q(net644854), .QN(
        n6324) );
  DFF_X1 \REGISTERS_reg[6][18]  ( .D(n3578), .CK(Clk), .Q(net644853), .QN(
        n6323) );
  DFF_X1 \REGISTERS_reg[6][17]  ( .D(n3577), .CK(Clk), .Q(net644852), .QN(
        n6322) );
  DFF_X1 \REGISTERS_reg[6][16]  ( .D(n3576), .CK(Clk), .Q(net644851), .QN(
        n6321) );
  DFF_X1 \REGISTERS_reg[6][15]  ( .D(n3575), .CK(Clk), .Q(net644850), .QN(
        n6320) );
  DFF_X1 \REGISTERS_reg[6][14]  ( .D(n3574), .CK(Clk), .Q(net644849), .QN(
        n6319) );
  DFF_X1 \REGISTERS_reg[6][13]  ( .D(n3573), .CK(Clk), .Q(net644848), .QN(
        n6318) );
  DFF_X1 \REGISTERS_reg[6][12]  ( .D(n3572), .CK(Clk), .Q(net644847), .QN(
        n6317) );
  DFF_X1 \REGISTERS_reg[6][11]  ( .D(n3571), .CK(Clk), .Q(net644846), .QN(
        n6316) );
  DFF_X1 \REGISTERS_reg[6][10]  ( .D(n3570), .CK(Clk), .Q(net644845), .QN(
        n6315) );
  DFF_X1 \REGISTERS_reg[6][9]  ( .D(n3569), .CK(Clk), .Q(net644844), .QN(n6314) );
  DFF_X1 \REGISTERS_reg[6][8]  ( .D(n3568), .CK(Clk), .Q(net644843), .QN(n6313) );
  DFF_X1 \REGISTERS_reg[6][7]  ( .D(n3567), .CK(Clk), .Q(net644842), .QN(n6312) );
  DFF_X1 \REGISTERS_reg[6][6]  ( .D(n3566), .CK(Clk), .Q(net644841), .QN(n6311) );
  DFF_X1 \REGISTERS_reg[6][5]  ( .D(n3565), .CK(Clk), .Q(net644840), .QN(n6310) );
  DFF_X1 \REGISTERS_reg[6][4]  ( .D(n3564), .CK(Clk), .Q(net644839), .QN(n6309) );
  DFF_X1 \REGISTERS_reg[6][3]  ( .D(n3563), .CK(Clk), .Q(net644838), .QN(n6308) );
  DFF_X1 \REGISTERS_reg[6][2]  ( .D(n3562), .CK(Clk), .Q(net644837), .QN(n6307) );
  DFF_X1 \REGISTERS_reg[6][1]  ( .D(n3561), .CK(Clk), .Q(net644836), .QN(n6306) );
  DFF_X1 \REGISTERS_reg[6][0]  ( .D(n3560), .CK(Clk), .Q(n4059), .QN(n480) );
  DFF_X1 \REGISTERS_reg[7][31]  ( .D(n3559), .CK(Clk), .QN(n608) );
  DFF_X1 \REGISTERS_reg[7][30]  ( .D(n3558), .CK(Clk), .QN(n609) );
  DFF_X1 \REGISTERS_reg[7][29]  ( .D(n3557), .CK(Clk), .QN(n610) );
  DFF_X1 \REGISTERS_reg[7][28]  ( .D(n3556), .CK(Clk), .QN(n611) );
  DFF_X1 \REGISTERS_reg[7][27]  ( .D(n3555), .CK(Clk), .QN(n612) );
  DFF_X1 \REGISTERS_reg[7][26]  ( .D(n3554), .CK(Clk), .QN(n613) );
  DFF_X1 \REGISTERS_reg[7][25]  ( .D(n3553), .CK(Clk), .QN(n614) );
  DFF_X1 \REGISTERS_reg[7][24]  ( .D(n3552), .CK(Clk), .QN(n615) );
  DFF_X1 \REGISTERS_reg[7][23]  ( .D(n3551), .CK(Clk), .QN(n616) );
  DFF_X1 \REGISTERS_reg[7][22]  ( .D(n3550), .CK(Clk), .QN(n617) );
  DFF_X1 \REGISTERS_reg[7][21]  ( .D(n3549), .CK(Clk), .QN(n618) );
  DFF_X1 \REGISTERS_reg[7][20]  ( .D(n3548), .CK(Clk), .QN(n619) );
  DFF_X1 \REGISTERS_reg[7][19]  ( .D(n3547), .CK(Clk), .QN(n620) );
  DFF_X1 \REGISTERS_reg[7][18]  ( .D(n3546), .CK(Clk), .QN(n621) );
  DFF_X1 \REGISTERS_reg[7][17]  ( .D(n3545), .CK(Clk), .QN(n622) );
  DFF_X1 \REGISTERS_reg[7][16]  ( .D(n3544), .CK(Clk), .QN(n623) );
  DFF_X1 \REGISTERS_reg[7][15]  ( .D(n3543), .CK(Clk), .QN(n624) );
  DFF_X1 \REGISTERS_reg[7][14]  ( .D(n3542), .CK(Clk), .QN(n625) );
  DFF_X1 \REGISTERS_reg[7][13]  ( .D(n3541), .CK(Clk), .QN(n626) );
  DFF_X1 \REGISTERS_reg[7][12]  ( .D(n3540), .CK(Clk), .QN(n627) );
  DFF_X1 \REGISTERS_reg[7][11]  ( .D(n3539), .CK(Clk), .QN(n628) );
  DFF_X1 \REGISTERS_reg[7][10]  ( .D(n3538), .CK(Clk), .QN(n629) );
  DFF_X1 \REGISTERS_reg[7][9]  ( .D(n3537), .CK(Clk), .QN(n630) );
  DFF_X1 \REGISTERS_reg[7][8]  ( .D(n3536), .CK(Clk), .QN(n631) );
  DFF_X1 \REGISTERS_reg[7][7]  ( .D(n3535), .CK(Clk), .QN(n632) );
  DFF_X1 \REGISTERS_reg[7][6]  ( .D(n3534), .CK(Clk), .QN(n633) );
  DFF_X1 \REGISTERS_reg[7][5]  ( .D(n3533), .CK(Clk), .QN(n634) );
  DFF_X1 \REGISTERS_reg[7][4]  ( .D(n3532), .CK(Clk), .QN(n635) );
  DFF_X1 \REGISTERS_reg[7][3]  ( .D(n3531), .CK(Clk), .QN(n636) );
  DFF_X1 \REGISTERS_reg[7][2]  ( .D(n3530), .CK(Clk), .QN(n637) );
  DFF_X1 \REGISTERS_reg[7][1]  ( .D(n3529), .CK(Clk), .QN(n638) );
  DFF_X1 \REGISTERS_reg[7][0]  ( .D(n3528), .CK(Clk), .Q(net644835), .QN(n6343) );
  DFF_X1 \REGISTERS_reg[8][31]  ( .D(n3527), .CK(Clk), .Q(n4165), .QN(n2664)
         );
  DFF_X1 \REGISTERS_reg[8][30]  ( .D(n3526), .CK(Clk), .Q(n4162), .QN(n2663)
         );
  DFF_X1 \REGISTERS_reg[8][29]  ( .D(n3525), .CK(Clk), .Q(n4159), .QN(n2662)
         );
  DFF_X1 \REGISTERS_reg[8][28]  ( .D(n3524), .CK(Clk), .Q(n4156), .QN(n2661)
         );
  DFF_X1 \REGISTERS_reg[8][27]  ( .D(n3523), .CK(Clk), .Q(n4153), .QN(n2660)
         );
  DFF_X1 \REGISTERS_reg[8][26]  ( .D(n3522), .CK(Clk), .Q(n4150), .QN(n2659)
         );
  DFF_X1 \REGISTERS_reg[8][25]  ( .D(n3521), .CK(Clk), .Q(n4147), .QN(n2658)
         );
  DFF_X1 \REGISTERS_reg[8][24]  ( .D(n3520), .CK(Clk), .Q(n4141), .QN(n2657)
         );
  DFF_X1 \REGISTERS_reg[8][23]  ( .D(n3519), .CK(Clk), .Q(n4138), .QN(n2656)
         );
  DFF_X1 \REGISTERS_reg[8][22]  ( .D(n3518), .CK(Clk), .Q(n4135), .QN(n2655)
         );
  DFF_X1 \REGISTERS_reg[8][21]  ( .D(n3517), .CK(Clk), .Q(n4132), .QN(n2654)
         );
  DFF_X1 \REGISTERS_reg[8][20]  ( .D(n3516), .CK(Clk), .Q(n4129), .QN(n2653)
         );
  DFF_X1 \REGISTERS_reg[8][19]  ( .D(n3515), .CK(Clk), .Q(n4126), .QN(n2652)
         );
  DFF_X1 \REGISTERS_reg[8][18]  ( .D(n3514), .CK(Clk), .Q(n4123), .QN(n2651)
         );
  DFF_X1 \REGISTERS_reg[8][17]  ( .D(n3513), .CK(Clk), .Q(n4120), .QN(n2650)
         );
  DFF_X1 \REGISTERS_reg[8][16]  ( .D(n3512), .CK(Clk), .Q(n4117), .QN(n2649)
         );
  DFF_X1 \REGISTERS_reg[8][15]  ( .D(n3511), .CK(Clk), .Q(n4114), .QN(n2648)
         );
  DFF_X1 \REGISTERS_reg[8][14]  ( .D(n3510), .CK(Clk), .Q(n4109), .QN(n2647)
         );
  DFF_X1 \REGISTERS_reg[8][13]  ( .D(n3509), .CK(Clk), .Q(n4103), .QN(n2646)
         );
  DFF_X1 \REGISTERS_reg[8][12]  ( .D(n3508), .CK(Clk), .Q(n4100), .QN(n2645)
         );
  DFF_X1 \REGISTERS_reg[8][11]  ( .D(n3507), .CK(Clk), .Q(n4097), .QN(n2644)
         );
  DFF_X1 \REGISTERS_reg[8][10]  ( .D(n3506), .CK(Clk), .Q(n4094), .QN(n2643)
         );
  DFF_X1 \REGISTERS_reg[8][9]  ( .D(n3505), .CK(Clk), .Q(n4091), .QN(n2642) );
  DFF_X1 \REGISTERS_reg[8][8]  ( .D(n3504), .CK(Clk), .Q(n4088), .QN(n2641) );
  DFF_X1 \REGISTERS_reg[8][7]  ( .D(n3503), .CK(Clk), .Q(n4085), .QN(n2640) );
  DFF_X1 \REGISTERS_reg[8][6]  ( .D(n3502), .CK(Clk), .Q(n4082), .QN(n2639) );
  DFF_X1 \REGISTERS_reg[8][5]  ( .D(n3501), .CK(Clk), .Q(n4079), .QN(n2638) );
  DFF_X1 \REGISTERS_reg[8][4]  ( .D(n3500), .CK(Clk), .Q(n4076), .QN(n2637) );
  DFF_X1 \REGISTERS_reg[8][3]  ( .D(n3499), .CK(Clk), .Q(n4071), .QN(n2636) );
  DFF_X1 \REGISTERS_reg[8][2]  ( .D(n3498), .CK(Clk), .Q(n4066), .QN(n2635) );
  DFF_X1 \REGISTERS_reg[8][1]  ( .D(n3497), .CK(Clk), .Q(n4063), .QN(n2634) );
  DFF_X1 \REGISTERS_reg[8][0]  ( .D(n3496), .CK(Clk), .Q(n384), .QN(n4169) );
  DFF_X1 \REGISTERS_reg[9][31]  ( .D(n3495), .CK(Clk), .Q(n389), .QN(n5993) );
  DFF_X1 \REGISTERS_reg[9][30]  ( .D(n3494), .CK(Clk), .Q(n392), .QN(n5992) );
  DFF_X1 \REGISTERS_reg[9][29]  ( .D(n3493), .CK(Clk), .Q(n395), .QN(n5991) );
  DFF_X1 \REGISTERS_reg[9][28]  ( .D(n3492), .CK(Clk), .Q(n398), .QN(n5990) );
  DFF_X1 \REGISTERS_reg[9][27]  ( .D(n3491), .CK(Clk), .Q(n401), .QN(n5989) );
  DFF_X1 \REGISTERS_reg[9][26]  ( .D(n3490), .CK(Clk), .Q(n404), .QN(n5988) );
  DFF_X1 \REGISTERS_reg[9][25]  ( .D(n3489), .CK(Clk), .Q(n407), .QN(n5987) );
  DFF_X1 \REGISTERS_reg[9][24]  ( .D(n3488), .CK(Clk), .Q(n410), .QN(n5986) );
  DFF_X1 \REGISTERS_reg[9][23]  ( .D(n3487), .CK(Clk), .Q(n413), .QN(n5985) );
  DFF_X1 \REGISTERS_reg[9][22]  ( .D(n3486), .CK(Clk), .Q(n416), .QN(n5970) );
  DFF_X1 \REGISTERS_reg[9][21]  ( .D(n3485), .CK(Clk), .Q(n419), .QN(n5965) );
  DFF_X1 \REGISTERS_reg[9][20]  ( .D(n3484), .CK(Clk), .Q(n422), .QN(n5933) );
  DFF_X1 \REGISTERS_reg[9][19]  ( .D(n3483), .CK(Clk), .Q(n425), .QN(n5252) );
  DFF_X1 \REGISTERS_reg[9][18]  ( .D(n3482), .CK(Clk), .Q(n428), .QN(n5218) );
  DFF_X1 \REGISTERS_reg[9][17]  ( .D(n3481), .CK(Clk), .Q(n431), .QN(n5204) );
  DFF_X1 \REGISTERS_reg[9][16]  ( .D(n3480), .CK(Clk), .Q(n434), .QN(n5203) );
  DFF_X1 \REGISTERS_reg[9][15]  ( .D(n3479), .CK(Clk), .Q(n437), .QN(n5193) );
  DFF_X1 \REGISTERS_reg[9][14]  ( .D(n3478), .CK(Clk), .Q(n440), .QN(n5188) );
  DFF_X1 \REGISTERS_reg[9][13]  ( .D(n3477), .CK(Clk), .Q(n443), .QN(n5183) );
  DFF_X1 \REGISTERS_reg[9][12]  ( .D(n3476), .CK(Clk), .Q(n446), .QN(n5180) );
  DFF_X1 \REGISTERS_reg[9][11]  ( .D(n3475), .CK(Clk), .Q(n449), .QN(n5174) );
  DFF_X1 \REGISTERS_reg[9][10]  ( .D(n3474), .CK(Clk), .Q(n452), .QN(n5153) );
  DFF_X1 \REGISTERS_reg[9][9]  ( .D(n3473), .CK(Clk), .Q(n455), .QN(n5145) );
  DFF_X1 \REGISTERS_reg[9][8]  ( .D(n3472), .CK(Clk), .Q(n458), .QN(n5144) );
  DFF_X1 \REGISTERS_reg[9][7]  ( .D(n3471), .CK(Clk), .Q(n461), .QN(n5139) );
  DFF_X1 \REGISTERS_reg[9][6]  ( .D(n3470), .CK(Clk), .Q(n464), .QN(n5134) );
  DFF_X1 \REGISTERS_reg[9][5]  ( .D(n3469), .CK(Clk), .Q(n467), .QN(n5133) );
  DFF_X1 \REGISTERS_reg[9][4]  ( .D(n3468), .CK(Clk), .Q(n470), .QN(n5123) );
  DFF_X1 \REGISTERS_reg[9][3]  ( .D(n3467), .CK(Clk), .Q(n473), .QN(n5115) );
  DFF_X1 \REGISTERS_reg[9][2]  ( .D(n3466), .CK(Clk), .Q(n476), .QN(n5114) );
  DFF_X1 \REGISTERS_reg[9][1]  ( .D(n3465), .CK(Clk), .Q(n479), .QN(n5113) );
  DFF_X1 \REGISTERS_reg[9][0]  ( .D(n3464), .CK(Clk), .Q(n4062), .QN(n2601) );
  DFF_X1 \REGISTERS_reg[10][31]  ( .D(n3463), .CK(Clk), .Q(net644834), .QN(
        n5109) );
  DFF_X1 \REGISTERS_reg[10][30]  ( .D(n3462), .CK(Clk), .Q(net644833), .QN(
        n5108) );
  DFF_X1 \REGISTERS_reg[10][29]  ( .D(n3461), .CK(Clk), .Q(net644832), .QN(
        n5103) );
  DFF_X1 \REGISTERS_reg[10][28]  ( .D(n3460), .CK(Clk), .Q(net644831), .QN(
        n5102) );
  DFF_X1 \REGISTERS_reg[10][27]  ( .D(n3459), .CK(Clk), .Q(net644830), .QN(
        n5093) );
  DFF_X1 \REGISTERS_reg[10][26]  ( .D(n3458), .CK(Clk), .Q(net644829), .QN(
        n5085) );
  DFF_X1 \REGISTERS_reg[10][25]  ( .D(n3457), .CK(Clk), .Q(net644828), .QN(
        n5084) );
  DFF_X1 \REGISTERS_reg[10][24]  ( .D(n3456), .CK(Clk), .Q(net644827), .QN(
        n5083) );
  DFF_X1 \REGISTERS_reg[10][23]  ( .D(n3455), .CK(Clk), .Q(net644826), .QN(
        n5079) );
  DFF_X1 \REGISTERS_reg[10][22]  ( .D(n3454), .CK(Clk), .Q(net644825), .QN(
        n5078) );
  DFF_X1 \REGISTERS_reg[10][21]  ( .D(n3453), .CK(Clk), .Q(net644824), .QN(
        n5073) );
  DFF_X1 \REGISTERS_reg[10][20]  ( .D(n3452), .CK(Clk), .Q(net644823), .QN(
        n5072) );
  DFF_X1 \REGISTERS_reg[10][19]  ( .D(n3451), .CK(Clk), .Q(net644822), .QN(
        n5063) );
  DFF_X1 \REGISTERS_reg[10][18]  ( .D(n3450), .CK(Clk), .Q(net644821), .QN(
        n5055) );
  DFF_X1 \REGISTERS_reg[10][17]  ( .D(n3449), .CK(Clk), .Q(net644820), .QN(
        n5054) );
  DFF_X1 \REGISTERS_reg[10][16]  ( .D(n3448), .CK(Clk), .Q(net644819), .QN(
        n5053) );
  DFF_X1 \REGISTERS_reg[10][15]  ( .D(n3447), .CK(Clk), .Q(net644818), .QN(
        n5049) );
  DFF_X1 \REGISTERS_reg[10][14]  ( .D(n3446), .CK(Clk), .Q(net644817), .QN(
        n5048) );
  DFF_X1 \REGISTERS_reg[10][13]  ( .D(n3445), .CK(Clk), .Q(net644816), .QN(
        n5043) );
  DFF_X1 \REGISTERS_reg[10][12]  ( .D(n3444), .CK(Clk), .Q(net644815), .QN(
        n5042) );
  DFF_X1 \REGISTERS_reg[10][11]  ( .D(n3443), .CK(Clk), .Q(net644814), .QN(
        n5033) );
  DFF_X1 \REGISTERS_reg[10][10]  ( .D(n3442), .CK(Clk), .Q(net644813), .QN(
        n5025) );
  DFF_X1 \REGISTERS_reg[10][9]  ( .D(n3441), .CK(Clk), .Q(net644812), .QN(
        n5024) );
  DFF_X1 \REGISTERS_reg[10][8]  ( .D(n3440), .CK(Clk), .Q(net644811), .QN(
        n5023) );
  DFF_X1 \REGISTERS_reg[10][7]  ( .D(n3439), .CK(Clk), .Q(net644810), .QN(
        n5019) );
  DFF_X1 \REGISTERS_reg[10][6]  ( .D(n3438), .CK(Clk), .Q(net644809), .QN(
        n5018) );
  DFF_X1 \REGISTERS_reg[10][5]  ( .D(n3437), .CK(Clk), .Q(net644808), .QN(
        n5013) );
  DFF_X1 \REGISTERS_reg[10][4]  ( .D(n3436), .CK(Clk), .Q(net644807), .QN(
        n5012) );
  DFF_X1 \REGISTERS_reg[10][3]  ( .D(n3435), .CK(Clk), .Q(net644806), .QN(
        n5003) );
  DFF_X1 \REGISTERS_reg[10][2]  ( .D(n3434), .CK(Clk), .Q(net644805), .QN(
        n4995) );
  DFF_X1 \REGISTERS_reg[10][1]  ( .D(n3433), .CK(Clk), .Q(net644804), .QN(
        n4994) );
  DFF_X1 \REGISTERS_reg[10][0]  ( .D(n3432), .CK(Clk), .QN(n481) );
  DFF_X1 \REGISTERS_reg[11][31]  ( .D(n3431), .CK(Clk), .Q(n4056), .QN(n482)
         );
  DFF_X1 \REGISTERS_reg[11][30]  ( .D(n3430), .CK(Clk), .Q(n4053), .QN(n483)
         );
  DFF_X1 \REGISTERS_reg[11][29]  ( .D(n3429), .CK(Clk), .Q(n4050), .QN(n484)
         );
  DFF_X1 \REGISTERS_reg[11][28]  ( .D(n3428), .CK(Clk), .Q(n4047), .QN(n485)
         );
  DFF_X1 \REGISTERS_reg[11][27]  ( .D(n3427), .CK(Clk), .Q(n4044), .QN(n486)
         );
  DFF_X1 \REGISTERS_reg[11][26]  ( .D(n3426), .CK(Clk), .Q(n4041), .QN(n487)
         );
  DFF_X1 \REGISTERS_reg[11][25]  ( .D(n3425), .CK(Clk), .Q(n4038), .QN(n488)
         );
  DFF_X1 \REGISTERS_reg[11][24]  ( .D(n3424), .CK(Clk), .Q(n4032), .QN(n489)
         );
  DFF_X1 \REGISTERS_reg[11][23]  ( .D(n3423), .CK(Clk), .Q(n4029), .QN(n490)
         );
  DFF_X1 \REGISTERS_reg[11][22]  ( .D(n3422), .CK(Clk), .Q(n4026), .QN(n491)
         );
  DFF_X1 \REGISTERS_reg[11][21]  ( .D(n3421), .CK(Clk), .Q(n4023), .QN(n492)
         );
  DFF_X1 \REGISTERS_reg[11][20]  ( .D(n3420), .CK(Clk), .Q(n4020), .QN(n493)
         );
  DFF_X1 \REGISTERS_reg[11][19]  ( .D(n3419), .CK(Clk), .Q(n4017), .QN(n494)
         );
  DFF_X1 \REGISTERS_reg[11][18]  ( .D(n3418), .CK(Clk), .Q(n4014), .QN(n495)
         );
  DFF_X1 \REGISTERS_reg[11][17]  ( .D(n3417), .CK(Clk), .Q(n4011), .QN(n496)
         );
  DFF_X1 \REGISTERS_reg[11][16]  ( .D(n3416), .CK(Clk), .Q(n4008), .QN(n497)
         );
  DFF_X1 \REGISTERS_reg[11][15]  ( .D(n3415), .CK(Clk), .Q(n4005), .QN(n498)
         );
  DFF_X1 \REGISTERS_reg[11][14]  ( .D(n3414), .CK(Clk), .Q(n4002), .QN(n499)
         );
  DFF_X1 \REGISTERS_reg[11][13]  ( .D(n3413), .CK(Clk), .Q(n3993), .QN(n500)
         );
  DFF_X1 \REGISTERS_reg[11][12]  ( .D(n3412), .CK(Clk), .Q(n3990), .QN(n501)
         );
  DFF_X1 \REGISTERS_reg[11][11]  ( .D(n3411), .CK(Clk), .Q(n3987), .QN(n502)
         );
  DFF_X1 \REGISTERS_reg[11][10]  ( .D(n3410), .CK(Clk), .Q(n3984), .QN(n503)
         );
  DFF_X1 \REGISTERS_reg[11][9]  ( .D(n3409), .CK(Clk), .Q(n3981), .QN(n504) );
  DFF_X1 \REGISTERS_reg[11][8]  ( .D(n3408), .CK(Clk), .Q(n3978), .QN(n505) );
  DFF_X1 \REGISTERS_reg[11][7]  ( .D(n3407), .CK(Clk), .Q(n3975), .QN(n506) );
  DFF_X1 \REGISTERS_reg[11][6]  ( .D(n3406), .CK(Clk), .Q(n3972), .QN(n507) );
  DFF_X1 \REGISTERS_reg[11][5]  ( .D(n3405), .CK(Clk), .Q(n3969), .QN(n508) );
  DFF_X1 \REGISTERS_reg[11][4]  ( .D(n3404), .CK(Clk), .Q(n3966), .QN(n509) );
  DFF_X1 \REGISTERS_reg[11][3]  ( .D(n3403), .CK(Clk), .Q(n3963), .QN(n510) );
  DFF_X1 \REGISTERS_reg[11][2]  ( .D(n3402), .CK(Clk), .Q(n3957), .QN(n511) );
  DFF_X1 \REGISTERS_reg[11][1]  ( .D(n3401), .CK(Clk), .Q(n3954), .QN(n512) );
  DFF_X1 \REGISTERS_reg[11][0]  ( .D(n3400), .CK(Clk), .Q(n3915), .QN(n639) );
  DFF_X1 \REGISTERS_reg[12][31]  ( .D(n3399), .CK(Clk), .Q(net644803), .QN(
        n4993) );
  DFF_X1 \REGISTERS_reg[12][30]  ( .D(n3398), .CK(Clk), .Q(net644802), .QN(
        n4989) );
  DFF_X1 \REGISTERS_reg[12][29]  ( .D(n3397), .CK(Clk), .Q(net644801), .QN(
        n4988) );
  DFF_X1 \REGISTERS_reg[12][28]  ( .D(n3396), .CK(Clk), .Q(net644800), .QN(
        n4983) );
  DFF_X1 \REGISTERS_reg[12][27]  ( .D(n3395), .CK(Clk), .Q(net644799), .QN(
        n4982) );
  DFF_X1 \REGISTERS_reg[12][26]  ( .D(n3394), .CK(Clk), .Q(net644798), .QN(
        n4973) );
  DFF_X1 \REGISTERS_reg[12][25]  ( .D(n3393), .CK(Clk), .Q(net644797), .QN(
        n4965) );
  DFF_X1 \REGISTERS_reg[12][24]  ( .D(n3392), .CK(Clk), .Q(net644796), .QN(
        n4964) );
  DFF_X1 \REGISTERS_reg[12][23]  ( .D(n3391), .CK(Clk), .Q(net644795), .QN(
        n4963) );
  DFF_X1 \REGISTERS_reg[12][22]  ( .D(n3390), .CK(Clk), .Q(net644794), .QN(
        n4959) );
  DFF_X1 \REGISTERS_reg[12][21]  ( .D(n3389), .CK(Clk), .Q(net644793), .QN(
        n4958) );
  DFF_X1 \REGISTERS_reg[12][20]  ( .D(n3388), .CK(Clk), .Q(net644792), .QN(
        n4953) );
  DFF_X1 \REGISTERS_reg[12][19]  ( .D(n3387), .CK(Clk), .Q(net644791), .QN(
        n4952) );
  DFF_X1 \REGISTERS_reg[12][18]  ( .D(n3386), .CK(Clk), .Q(net644790), .QN(
        n4943) );
  DFF_X1 \REGISTERS_reg[12][17]  ( .D(n3385), .CK(Clk), .Q(net644789), .QN(
        n4935) );
  DFF_X1 \REGISTERS_reg[12][16]  ( .D(n3384), .CK(Clk), .Q(net644788), .QN(
        n4934) );
  DFF_X1 \REGISTERS_reg[12][15]  ( .D(n3383), .CK(Clk), .Q(net644787), .QN(
        n4933) );
  DFF_X1 \REGISTERS_reg[12][14]  ( .D(n3382), .CK(Clk), .Q(net644786), .QN(
        n4929) );
  DFF_X1 \REGISTERS_reg[12][13]  ( .D(n3381), .CK(Clk), .Q(net644785), .QN(
        n4928) );
  DFF_X1 \REGISTERS_reg[12][12]  ( .D(n3380), .CK(Clk), .Q(net644784), .QN(
        n4923) );
  DFF_X1 \REGISTERS_reg[12][11]  ( .D(n3379), .CK(Clk), .Q(net644783), .QN(
        n4922) );
  DFF_X1 \REGISTERS_reg[12][10]  ( .D(n3378), .CK(Clk), .Q(net644782), .QN(
        n4913) );
  DFF_X1 \REGISTERS_reg[12][9]  ( .D(n3377), .CK(Clk), .Q(net644781), .QN(
        n4905) );
  DFF_X1 \REGISTERS_reg[12][8]  ( .D(n3376), .CK(Clk), .Q(net644780), .QN(
        n4904) );
  DFF_X1 \REGISTERS_reg[12][7]  ( .D(n3375), .CK(Clk), .Q(net644779), .QN(
        n4903) );
  DFF_X1 \REGISTERS_reg[12][6]  ( .D(n3374), .CK(Clk), .Q(net644778), .QN(
        n4899) );
  DFF_X1 \REGISTERS_reg[12][5]  ( .D(n3373), .CK(Clk), .Q(net644777), .QN(
        n4898) );
  DFF_X1 \REGISTERS_reg[12][4]  ( .D(n3372), .CK(Clk), .Q(net644776), .QN(
        n4893) );
  DFF_X1 \REGISTERS_reg[12][3]  ( .D(n3371), .CK(Clk), .Q(net644775), .QN(
        n4892) );
  DFF_X1 \REGISTERS_reg[12][2]  ( .D(n3370), .CK(Clk), .Q(net644774), .QN(
        n4883) );
  DFF_X1 \REGISTERS_reg[12][1]  ( .D(n3369), .CK(Clk), .Q(net644773), .QN(
        n4875) );
  DFF_X1 \REGISTERS_reg[12][0]  ( .D(n3368), .CK(Clk), .Q(net644772), .QN(
        n6342) );
  DFF_X1 \REGISTERS_reg[13][31]  ( .D(n3367), .CK(Clk), .Q(net644771), .QN(
        n6305) );
  DFF_X1 \REGISTERS_reg[13][30]  ( .D(n3366), .CK(Clk), .Q(net644770), .QN(
        n6304) );
  DFF_X1 \REGISTERS_reg[13][29]  ( .D(n3365), .CK(Clk), .Q(net644769), .QN(
        n6303) );
  DFF_X1 \REGISTERS_reg[13][28]  ( .D(n3364), .CK(Clk), .Q(net644768), .QN(
        n6302) );
  DFF_X1 \REGISTERS_reg[13][27]  ( .D(n3363), .CK(Clk), .Q(net644767), .QN(
        n6301) );
  DFF_X1 \REGISTERS_reg[13][26]  ( .D(n3362), .CK(Clk), .Q(net644766), .QN(
        n6300) );
  DFF_X1 \REGISTERS_reg[13][25]  ( .D(n3361), .CK(Clk), .Q(net644765), .QN(
        n6299) );
  DFF_X1 \REGISTERS_reg[13][24]  ( .D(n3360), .CK(Clk), .Q(net644764), .QN(
        n6298) );
  DFF_X1 \REGISTERS_reg[13][23]  ( .D(n3359), .CK(Clk), .Q(net644763), .QN(
        n6297) );
  DFF_X1 \REGISTERS_reg[13][22]  ( .D(n3358), .CK(Clk), .Q(net644762), .QN(
        n6296) );
  DFF_X1 \REGISTERS_reg[13][21]  ( .D(n3357), .CK(Clk), .Q(net644761), .QN(
        n6295) );
  DFF_X1 \REGISTERS_reg[13][20]  ( .D(n3356), .CK(Clk), .Q(net644760), .QN(
        n6294) );
  DFF_X1 \REGISTERS_reg[13][19]  ( .D(n3355), .CK(Clk), .Q(net644759), .QN(
        n6293) );
  DFF_X1 \REGISTERS_reg[13][18]  ( .D(n3354), .CK(Clk), .Q(net644758), .QN(
        n6292) );
  DFF_X1 \REGISTERS_reg[13][17]  ( .D(n3353), .CK(Clk), .Q(net644757), .QN(
        n6291) );
  DFF_X1 \REGISTERS_reg[13][16]  ( .D(n3352), .CK(Clk), .Q(net644756), .QN(
        n6290) );
  DFF_X1 \REGISTERS_reg[13][15]  ( .D(n3351), .CK(Clk), .Q(net644755), .QN(
        n6289) );
  DFF_X1 \REGISTERS_reg[13][14]  ( .D(n3350), .CK(Clk), .Q(net644754), .QN(
        n6288) );
  DFF_X1 \REGISTERS_reg[13][13]  ( .D(n3349), .CK(Clk), .Q(net644753), .QN(
        n6287) );
  DFF_X1 \REGISTERS_reg[13][12]  ( .D(n3348), .CK(Clk), .Q(net644752), .QN(
        n6286) );
  DFF_X1 \REGISTERS_reg[13][11]  ( .D(n3347), .CK(Clk), .Q(net644751), .QN(
        n6285) );
  DFF_X1 \REGISTERS_reg[13][10]  ( .D(n3346), .CK(Clk), .Q(net644750), .QN(
        n6284) );
  DFF_X1 \REGISTERS_reg[13][9]  ( .D(n3345), .CK(Clk), .Q(net644749), .QN(
        n6283) );
  DFF_X1 \REGISTERS_reg[13][8]  ( .D(n3344), .CK(Clk), .Q(net644748), .QN(
        n6282) );
  DFF_X1 \REGISTERS_reg[13][7]  ( .D(n3343), .CK(Clk), .Q(net644747), .QN(
        n6281) );
  DFF_X1 \REGISTERS_reg[13][6]  ( .D(n3342), .CK(Clk), .Q(net644746), .QN(
        n6280) );
  DFF_X1 \REGISTERS_reg[13][5]  ( .D(n3341), .CK(Clk), .Q(net644745), .QN(
        n6279) );
  DFF_X1 \REGISTERS_reg[13][4]  ( .D(n3340), .CK(Clk), .Q(net644744), .QN(
        n6278) );
  DFF_X1 \REGISTERS_reg[13][3]  ( .D(n3339), .CK(Clk), .Q(net644743), .QN(
        n6277) );
  DFF_X1 \REGISTERS_reg[13][2]  ( .D(n3338), .CK(Clk), .Q(net644742), .QN(
        n6276) );
  DFF_X1 \REGISTERS_reg[13][1]  ( .D(n3337), .CK(Clk), .Q(net644741), .QN(
        n6275) );
  DFF_X1 \REGISTERS_reg[13][0]  ( .D(n3336), .CK(Clk), .Q(net644740), .QN(
        n6352) );
  DFF_X1 \REGISTERS_reg[14][31]  ( .D(n3335), .CK(Clk), .Q(net644739), .QN(
        n6118) );
  DFF_X1 \REGISTERS_reg[14][30]  ( .D(n3334), .CK(Clk), .Q(net644738), .QN(
        n6117) );
  DFF_X1 \REGISTERS_reg[14][29]  ( .D(n3333), .CK(Clk), .Q(net644737), .QN(
        n6116) );
  DFF_X1 \REGISTERS_reg[14][28]  ( .D(n3332), .CK(Clk), .Q(net644736), .QN(
        n6115) );
  DFF_X1 \REGISTERS_reg[14][27]  ( .D(n3331), .CK(Clk), .Q(net644735), .QN(
        n6114) );
  DFF_X1 \REGISTERS_reg[14][26]  ( .D(n3330), .CK(Clk), .Q(net644734), .QN(
        n6113) );
  DFF_X1 \REGISTERS_reg[14][25]  ( .D(n3329), .CK(Clk), .Q(net644733), .QN(
        n6112) );
  DFF_X1 \REGISTERS_reg[14][24]  ( .D(n3328), .CK(Clk), .Q(net644732), .QN(
        n6111) );
  DFF_X1 \REGISTERS_reg[14][23]  ( .D(n3327), .CK(Clk), .Q(net644731), .QN(
        n6110) );
  DFF_X1 \REGISTERS_reg[14][22]  ( .D(n3326), .CK(Clk), .Q(net644730), .QN(
        n6109) );
  DFF_X1 \REGISTERS_reg[14][21]  ( .D(n3325), .CK(Clk), .Q(net644729), .QN(
        n6108) );
  DFF_X1 \REGISTERS_reg[14][20]  ( .D(n3324), .CK(Clk), .Q(net644728), .QN(
        n6107) );
  DFF_X1 \REGISTERS_reg[14][19]  ( .D(n3323), .CK(Clk), .Q(net644727), .QN(
        n6106) );
  DFF_X1 \REGISTERS_reg[14][18]  ( .D(n3322), .CK(Clk), .Q(net644726), .QN(
        n6105) );
  DFF_X1 \REGISTERS_reg[14][17]  ( .D(n3321), .CK(Clk), .Q(net644725), .QN(
        n6104) );
  DFF_X1 \REGISTERS_reg[14][16]  ( .D(n3320), .CK(Clk), .Q(net644724), .QN(
        n6103) );
  DFF_X1 \REGISTERS_reg[14][15]  ( .D(n3319), .CK(Clk), .Q(net644723), .QN(
        n6102) );
  DFF_X1 \REGISTERS_reg[14][14]  ( .D(n3318), .CK(Clk), .Q(net644722), .QN(
        n6101) );
  DFF_X1 \REGISTERS_reg[14][13]  ( .D(n3317), .CK(Clk), .Q(net644721), .QN(
        n6100) );
  DFF_X1 \REGISTERS_reg[14][12]  ( .D(n3316), .CK(Clk), .Q(net644720), .QN(
        n6099) );
  DFF_X1 \REGISTERS_reg[14][11]  ( .D(n3315), .CK(Clk), .Q(net644719), .QN(
        n6098) );
  DFF_X1 \REGISTERS_reg[14][10]  ( .D(n3314), .CK(Clk), .Q(net644718), .QN(
        n6097) );
  DFF_X1 \REGISTERS_reg[14][9]  ( .D(n3313), .CK(Clk), .Q(net644717), .QN(
        n6096) );
  DFF_X1 \REGISTERS_reg[14][8]  ( .D(n3312), .CK(Clk), .Q(net644716), .QN(
        n6095) );
  DFF_X1 \REGISTERS_reg[14][7]  ( .D(n3311), .CK(Clk), .Q(net644715), .QN(
        n6094) );
  DFF_X1 \REGISTERS_reg[14][6]  ( .D(n3310), .CK(Clk), .Q(net644714), .QN(
        n6093) );
  DFF_X1 \REGISTERS_reg[14][5]  ( .D(n3309), .CK(Clk), .Q(net644713), .QN(
        n6092) );
  DFF_X1 \REGISTERS_reg[14][4]  ( .D(n3308), .CK(Clk), .Q(net644712), .QN(
        n6091) );
  DFF_X1 \REGISTERS_reg[14][3]  ( .D(n3307), .CK(Clk), .Q(net644711), .QN(
        n6090) );
  DFF_X1 \REGISTERS_reg[14][2]  ( .D(n3306), .CK(Clk), .Q(net644710), .QN(
        n6089) );
  DFF_X1 \REGISTERS_reg[14][1]  ( .D(n3305), .CK(Clk), .Q(net644709), .QN(
        n6088) );
  DFF_X1 \REGISTERS_reg[14][0]  ( .D(n3304), .CK(Clk), .Q(net644708), .QN(
        n6087) );
  DFF_X1 \REGISTERS_reg[15][31]  ( .D(n3303), .CK(Clk), .Q(n4057), .QN(n704)
         );
  DFF_X1 \REGISTERS_reg[15][30]  ( .D(n3302), .CK(Clk), .Q(n4054), .QN(n705)
         );
  DFF_X1 \REGISTERS_reg[15][29]  ( .D(n3301), .CK(Clk), .Q(n4051), .QN(n706)
         );
  DFF_X1 \REGISTERS_reg[15][28]  ( .D(n3300), .CK(Clk), .Q(n4048), .QN(n707)
         );
  DFF_X1 \REGISTERS_reg[15][27]  ( .D(n3299), .CK(Clk), .Q(n4045), .QN(n708)
         );
  DFF_X1 \REGISTERS_reg[15][26]  ( .D(n3298), .CK(Clk), .Q(n4042), .QN(n709)
         );
  DFF_X1 \REGISTERS_reg[15][25]  ( .D(n3297), .CK(Clk), .Q(n4039), .QN(n710)
         );
  DFF_X1 \REGISTERS_reg[15][24]  ( .D(n3296), .CK(Clk), .Q(n4034), .QN(n711)
         );
  DFF_X1 \REGISTERS_reg[15][23]  ( .D(n3295), .CK(Clk), .Q(n4030), .QN(n712)
         );
  DFF_X1 \REGISTERS_reg[15][22]  ( .D(n3294), .CK(Clk), .Q(n4027), .QN(n713)
         );
  DFF_X1 \REGISTERS_reg[15][21]  ( .D(n3293), .CK(Clk), .Q(n4024), .QN(n714)
         );
  DFF_X1 \REGISTERS_reg[15][20]  ( .D(n3292), .CK(Clk), .Q(n4021), .QN(n715)
         );
  DFF_X1 \REGISTERS_reg[15][19]  ( .D(n3291), .CK(Clk), .Q(n4018), .QN(n716)
         );
  DFF_X1 \REGISTERS_reg[15][18]  ( .D(n3290), .CK(Clk), .Q(n4015), .QN(n717)
         );
  DFF_X1 \REGISTERS_reg[15][17]  ( .D(n3289), .CK(Clk), .Q(n4012), .QN(n718)
         );
  DFF_X1 \REGISTERS_reg[15][16]  ( .D(n3288), .CK(Clk), .Q(n4009), .QN(n719)
         );
  DFF_X1 \REGISTERS_reg[15][15]  ( .D(n3287), .CK(Clk), .Q(n4006), .QN(n720)
         );
  DFF_X1 \REGISTERS_reg[15][14]  ( .D(n3286), .CK(Clk), .Q(n4003), .QN(n721)
         );
  DFF_X1 \REGISTERS_reg[15][13]  ( .D(n3285), .CK(Clk), .Q(n3998), .QN(n722)
         );
  DFF_X1 \REGISTERS_reg[15][12]  ( .D(n3284), .CK(Clk), .Q(n3991), .QN(n723)
         );
  DFF_X1 \REGISTERS_reg[15][11]  ( .D(n3283), .CK(Clk), .Q(n3988), .QN(n724)
         );
  DFF_X1 \REGISTERS_reg[15][10]  ( .D(n3282), .CK(Clk), .Q(n3985), .QN(n725)
         );
  DFF_X1 \REGISTERS_reg[15][9]  ( .D(n3281), .CK(Clk), .Q(n3982), .QN(n726) );
  DFF_X1 \REGISTERS_reg[15][8]  ( .D(n3280), .CK(Clk), .Q(n3979), .QN(n727) );
  DFF_X1 \REGISTERS_reg[15][7]  ( .D(n3279), .CK(Clk), .Q(n3976), .QN(n728) );
  DFF_X1 \REGISTERS_reg[15][6]  ( .D(n3278), .CK(Clk), .Q(n3973), .QN(n729) );
  DFF_X1 \REGISTERS_reg[15][5]  ( .D(n3277), .CK(Clk), .Q(n3970), .QN(n730) );
  DFF_X1 \REGISTERS_reg[15][4]  ( .D(n3276), .CK(Clk), .Q(n3967), .QN(n731) );
  DFF_X1 \REGISTERS_reg[15][3]  ( .D(n3275), .CK(Clk), .Q(n3964), .QN(n732) );
  DFF_X1 \REGISTERS_reg[15][2]  ( .D(n3274), .CK(Clk), .Q(n3958), .QN(n733) );
  DFF_X1 \REGISTERS_reg[15][1]  ( .D(n3273), .CK(Clk), .Q(n3955), .QN(n734) );
  DFF_X1 \REGISTERS_reg[15][0]  ( .D(n3272), .CK(Clk), .Q(n4061), .QN(n513) );
  DFF_X1 \REGISTERS_reg[16][31]  ( .D(n3271), .CK(Clk), .Q(net644707), .QN(
        n6274) );
  DFF_X1 \REGISTERS_reg[16][30]  ( .D(n3270), .CK(Clk), .Q(net644706), .QN(
        n6273) );
  DFF_X1 \REGISTERS_reg[16][29]  ( .D(n3269), .CK(Clk), .Q(net644705), .QN(
        n6272) );
  DFF_X1 \REGISTERS_reg[16][28]  ( .D(n3268), .CK(Clk), .Q(net644704), .QN(
        n6271) );
  DFF_X1 \REGISTERS_reg[16][27]  ( .D(n3267), .CK(Clk), .Q(net644703), .QN(
        n6270) );
  DFF_X1 \REGISTERS_reg[16][26]  ( .D(n3266), .CK(Clk), .Q(net644702), .QN(
        n6269) );
  DFF_X1 \REGISTERS_reg[16][25]  ( .D(n3265), .CK(Clk), .Q(net644701), .QN(
        n6268) );
  DFF_X1 \REGISTERS_reg[16][24]  ( .D(n3264), .CK(Clk), .Q(net644700), .QN(
        n6267) );
  DFF_X1 \REGISTERS_reg[16][23]  ( .D(n3263), .CK(Clk), .Q(net644699), .QN(
        n6266) );
  DFF_X1 \REGISTERS_reg[16][22]  ( .D(n3262), .CK(Clk), .Q(net644698), .QN(
        n6265) );
  DFF_X1 \REGISTERS_reg[16][21]  ( .D(n3261), .CK(Clk), .Q(net644697), .QN(
        n6264) );
  DFF_X1 \REGISTERS_reg[16][20]  ( .D(n3260), .CK(Clk), .Q(net644696), .QN(
        n6263) );
  DFF_X1 \REGISTERS_reg[16][19]  ( .D(n3259), .CK(Clk), .Q(net644695), .QN(
        n6262) );
  DFF_X1 \REGISTERS_reg[16][18]  ( .D(n3258), .CK(Clk), .Q(net644694), .QN(
        n6261) );
  DFF_X1 \REGISTERS_reg[16][17]  ( .D(n3257), .CK(Clk), .Q(net644693), .QN(
        n6260) );
  DFF_X1 \REGISTERS_reg[16][16]  ( .D(n3256), .CK(Clk), .Q(net644692), .QN(
        n6259) );
  DFF_X1 \REGISTERS_reg[16][15]  ( .D(n3255), .CK(Clk), .Q(net644691), .QN(
        n6258) );
  DFF_X1 \REGISTERS_reg[16][14]  ( .D(n3254), .CK(Clk), .Q(net644690), .QN(
        n6257) );
  DFF_X1 \REGISTERS_reg[16][13]  ( .D(n3253), .CK(Clk), .Q(net644689), .QN(
        n6256) );
  DFF_X1 \REGISTERS_reg[16][12]  ( .D(n3252), .CK(Clk), .Q(net644688), .QN(
        n6255) );
  DFF_X1 \REGISTERS_reg[16][11]  ( .D(n3251), .CK(Clk), .Q(net644687), .QN(
        n6254) );
  DFF_X1 \REGISTERS_reg[16][10]  ( .D(n3250), .CK(Clk), .Q(net644686), .QN(
        n6253) );
  DFF_X1 \REGISTERS_reg[16][9]  ( .D(n3249), .CK(Clk), .Q(net644685), .QN(
        n6252) );
  DFF_X1 \REGISTERS_reg[16][8]  ( .D(n3248), .CK(Clk), .Q(net644684), .QN(
        n6251) );
  DFF_X1 \REGISTERS_reg[16][7]  ( .D(n3247), .CK(Clk), .Q(net644683), .QN(
        n6250) );
  DFF_X1 \REGISTERS_reg[16][6]  ( .D(n3246), .CK(Clk), .Q(net644682), .QN(
        n6249) );
  DFF_X1 \REGISTERS_reg[16][5]  ( .D(n3245), .CK(Clk), .Q(net644681), .QN(
        n6248) );
  DFF_X1 \REGISTERS_reg[16][4]  ( .D(n3244), .CK(Clk), .Q(net644680), .QN(
        n6247) );
  DFF_X1 \REGISTERS_reg[16][3]  ( .D(n3243), .CK(Clk), .Q(net644679), .QN(
        n6246) );
  DFF_X1 \REGISTERS_reg[16][2]  ( .D(n3242), .CK(Clk), .Q(net644678), .QN(
        n6245) );
  DFF_X1 \REGISTERS_reg[16][1]  ( .D(n3241), .CK(Clk), .Q(net644677), .QN(
        n6244) );
  DFF_X1 \REGISTERS_reg[16][0]  ( .D(n3240), .CK(Clk), .Q(net644676), .QN(
        n6351) );
  DFF_X1 \REGISTERS_reg[17][31]  ( .D(n3239), .CK(Clk), .Q(n353), .QN(n4298)
         );
  DFF_X1 \REGISTERS_reg[17][30]  ( .D(n3238), .CK(Clk), .Q(n354), .QN(n4293)
         );
  DFF_X1 \REGISTERS_reg[17][29]  ( .D(n3237), .CK(Clk), .Q(n355), .QN(n4292)
         );
  DFF_X1 \REGISTERS_reg[17][28]  ( .D(n3236), .CK(Clk), .Q(n356), .QN(n4283)
         );
  DFF_X1 \REGISTERS_reg[17][27]  ( .D(n3235), .CK(Clk), .Q(n357), .QN(n4275)
         );
  DFF_X1 \REGISTERS_reg[17][26]  ( .D(n3234), .CK(Clk), .Q(n358), .QN(n4274)
         );
  DFF_X1 \REGISTERS_reg[17][25]  ( .D(n3233), .CK(Clk), .Q(n359), .QN(n4273)
         );
  DFF_X1 \REGISTERS_reg[17][24]  ( .D(n3232), .CK(Clk), .Q(n360), .QN(n4269)
         );
  DFF_X1 \REGISTERS_reg[17][23]  ( .D(n3231), .CK(Clk), .Q(n361), .QN(n4268)
         );
  DFF_X1 \REGISTERS_reg[17][22]  ( .D(n3230), .CK(Clk), .Q(n362), .QN(n4263)
         );
  DFF_X1 \REGISTERS_reg[17][21]  ( .D(n3229), .CK(Clk), .Q(n363), .QN(n4262)
         );
  DFF_X1 \REGISTERS_reg[17][20]  ( .D(n3228), .CK(Clk), .Q(n364), .QN(n4253)
         );
  DFF_X1 \REGISTERS_reg[17][19]  ( .D(n3227), .CK(Clk), .Q(n365), .QN(n4245)
         );
  DFF_X1 \REGISTERS_reg[17][18]  ( .D(n3226), .CK(Clk), .Q(n366), .QN(n4244)
         );
  DFF_X1 \REGISTERS_reg[17][17]  ( .D(n3225), .CK(Clk), .Q(n367), .QN(n4242)
         );
  DFF_X1 \REGISTERS_reg[17][16]  ( .D(n3224), .CK(Clk), .Q(n368), .QN(n4230)
         );
  DFF_X1 \REGISTERS_reg[17][15]  ( .D(n3223), .CK(Clk), .Q(n369), .QN(n4227)
         );
  DFF_X1 \REGISTERS_reg[17][14]  ( .D(n3222), .CK(Clk), .Q(n370), .QN(n4222)
         );
  DFF_X1 \REGISTERS_reg[17][13]  ( .D(n3221), .CK(Clk), .Q(n371), .QN(n4213)
         );
  DFF_X1 \REGISTERS_reg[17][12]  ( .D(n3220), .CK(Clk), .Q(n372), .QN(n4206)
         );
  DFF_X1 \REGISTERS_reg[17][11]  ( .D(n3219), .CK(Clk), .Q(n373), .QN(n4193)
         );
  DFF_X1 \REGISTERS_reg[17][10]  ( .D(n3218), .CK(Clk), .Q(n374), .QN(n4191)
         );
  DFF_X1 \REGISTERS_reg[17][9]  ( .D(n3217), .CK(Clk), .Q(n375), .QN(n4179) );
  DFF_X1 \REGISTERS_reg[17][8]  ( .D(n3216), .CK(Clk), .Q(n376), .QN(n4177) );
  DFF_X1 \REGISTERS_reg[17][7]  ( .D(n3215), .CK(Clk), .Q(n377), .QN(n4176) );
  DFF_X1 \REGISTERS_reg[17][6]  ( .D(n3214), .CK(Clk), .Q(n378), .QN(n4175) );
  DFF_X1 \REGISTERS_reg[17][5]  ( .D(n3213), .CK(Clk), .Q(n379), .QN(n4174) );
  DFF_X1 \REGISTERS_reg[17][4]  ( .D(n3212), .CK(Clk), .Q(n380), .QN(n4173) );
  DFF_X1 \REGISTERS_reg[17][3]  ( .D(n3211), .CK(Clk), .Q(n381), .QN(n4172) );
  DFF_X1 \REGISTERS_reg[17][2]  ( .D(n3210), .CK(Clk), .Q(n382), .QN(n4171) );
  DFF_X1 \REGISTERS_reg[17][1]  ( .D(n3209), .CK(Clk), .Q(n383), .QN(n4170) );
  DFF_X1 \REGISTERS_reg[17][0]  ( .D(n3208), .CK(Clk), .Q(n386), .QN(n4168) );
  DFF_X1 \REGISTERS_reg[18][31]  ( .D(n3207), .CK(Clk), .QN(n640) );
  DFF_X1 \REGISTERS_reg[18][30]  ( .D(n3206), .CK(Clk), .QN(n641) );
  DFF_X1 \REGISTERS_reg[18][29]  ( .D(n3205), .CK(Clk), .QN(n642) );
  DFF_X1 \REGISTERS_reg[18][28]  ( .D(n3204), .CK(Clk), .QN(n643) );
  DFF_X1 \REGISTERS_reg[18][27]  ( .D(n3203), .CK(Clk), .QN(n644) );
  DFF_X1 \REGISTERS_reg[18][26]  ( .D(n3202), .CK(Clk), .QN(n645) );
  DFF_X1 \REGISTERS_reg[18][25]  ( .D(n3201), .CK(Clk), .QN(n646) );
  DFF_X1 \REGISTERS_reg[18][24]  ( .D(n3200), .CK(Clk), .QN(n647) );
  DFF_X1 \REGISTERS_reg[18][23]  ( .D(n3199), .CK(Clk), .QN(n648) );
  DFF_X1 \REGISTERS_reg[18][22]  ( .D(n3198), .CK(Clk), .QN(n649) );
  DFF_X1 \REGISTERS_reg[18][21]  ( .D(n3197), .CK(Clk), .QN(n650) );
  DFF_X1 \REGISTERS_reg[18][20]  ( .D(n3196), .CK(Clk), .QN(n651) );
  DFF_X1 \REGISTERS_reg[18][19]  ( .D(n3195), .CK(Clk), .QN(n652) );
  DFF_X1 \REGISTERS_reg[18][18]  ( .D(n3194), .CK(Clk), .QN(n653) );
  DFF_X1 \REGISTERS_reg[18][17]  ( .D(n3193), .CK(Clk), .QN(n654) );
  DFF_X1 \REGISTERS_reg[18][16]  ( .D(n3192), .CK(Clk), .QN(n655) );
  DFF_X1 \REGISTERS_reg[18][15]  ( .D(n3191), .CK(Clk), .QN(n656) );
  DFF_X1 \REGISTERS_reg[18][14]  ( .D(n3190), .CK(Clk), .QN(n657) );
  DFF_X1 \REGISTERS_reg[18][13]  ( .D(n3189), .CK(Clk), .QN(n658) );
  DFF_X1 \REGISTERS_reg[18][12]  ( .D(n3188), .CK(Clk), .QN(n659) );
  DFF_X1 \REGISTERS_reg[18][11]  ( .D(n3187), .CK(Clk), .QN(n660) );
  DFF_X1 \REGISTERS_reg[18][10]  ( .D(n3186), .CK(Clk), .QN(n661) );
  DFF_X1 \REGISTERS_reg[18][9]  ( .D(n3185), .CK(Clk), .QN(n662) );
  DFF_X1 \REGISTERS_reg[18][8]  ( .D(n3184), .CK(Clk), .QN(n663) );
  DFF_X1 \REGISTERS_reg[18][7]  ( .D(n3183), .CK(Clk), .QN(n664) );
  DFF_X1 \REGISTERS_reg[18][6]  ( .D(n3182), .CK(Clk), .QN(n665) );
  DFF_X1 \REGISTERS_reg[18][5]  ( .D(n3181), .CK(Clk), .QN(n666) );
  DFF_X1 \REGISTERS_reg[18][4]  ( .D(n3180), .CK(Clk), .QN(n667) );
  DFF_X1 \REGISTERS_reg[18][3]  ( .D(n3179), .CK(Clk), .QN(n668) );
  DFF_X1 \REGISTERS_reg[18][2]  ( .D(n3178), .CK(Clk), .QN(n669) );
  DFF_X1 \REGISTERS_reg[18][1]  ( .D(n3177), .CK(Clk), .QN(n670) );
  DFF_X1 \REGISTERS_reg[18][0]  ( .D(n3176), .CK(Clk), .Q(net644675), .QN(
        n6337) );
  DFF_X1 \REGISTERS_reg[19][31]  ( .D(n3175), .CK(Clk), .Q(net644674), .QN(
        n6086) );
  DFF_X1 \REGISTERS_reg[19][30]  ( .D(n3174), .CK(Clk), .Q(net644673), .QN(
        n6085) );
  DFF_X1 \REGISTERS_reg[19][29]  ( .D(n3173), .CK(Clk), .Q(net644672), .QN(
        n6084) );
  DFF_X1 \REGISTERS_reg[19][28]  ( .D(n3172), .CK(Clk), .Q(net644671), .QN(
        n6083) );
  DFF_X1 \REGISTERS_reg[19][27]  ( .D(n3171), .CK(Clk), .Q(net644670), .QN(
        n6082) );
  DFF_X1 \REGISTERS_reg[19][26]  ( .D(n3170), .CK(Clk), .Q(net644669), .QN(
        n6081) );
  DFF_X1 \REGISTERS_reg[19][25]  ( .D(n3169), .CK(Clk), .Q(net644668), .QN(
        n6080) );
  DFF_X1 \REGISTERS_reg[19][24]  ( .D(n3168), .CK(Clk), .Q(net644667), .QN(
        n6079) );
  DFF_X1 \REGISTERS_reg[19][23]  ( .D(n3167), .CK(Clk), .Q(net644666), .QN(
        n6078) );
  DFF_X1 \REGISTERS_reg[19][22]  ( .D(n3166), .CK(Clk), .Q(net644665), .QN(
        n6077) );
  DFF_X1 \REGISTERS_reg[19][21]  ( .D(n3165), .CK(Clk), .Q(net644664), .QN(
        n6076) );
  DFF_X1 \REGISTERS_reg[19][20]  ( .D(n3164), .CK(Clk), .Q(net644663), .QN(
        n6075) );
  DFF_X1 \REGISTERS_reg[19][19]  ( .D(n3163), .CK(Clk), .Q(net644662), .QN(
        n6074) );
  DFF_X1 \REGISTERS_reg[19][18]  ( .D(n3162), .CK(Clk), .Q(net644661), .QN(
        n6073) );
  DFF_X1 \REGISTERS_reg[19][17]  ( .D(n3161), .CK(Clk), .Q(net644660), .QN(
        n6072) );
  DFF_X1 \REGISTERS_reg[19][16]  ( .D(n3160), .CK(Clk), .Q(net644659), .QN(
        n6071) );
  DFF_X1 \REGISTERS_reg[19][15]  ( .D(n3159), .CK(Clk), .Q(net644658), .QN(
        n6070) );
  DFF_X1 \REGISTERS_reg[19][14]  ( .D(n3158), .CK(Clk), .Q(net644657), .QN(
        n6069) );
  DFF_X1 \REGISTERS_reg[19][13]  ( .D(n3157), .CK(Clk), .Q(net644656), .QN(
        n6068) );
  DFF_X1 \REGISTERS_reg[19][12]  ( .D(n3156), .CK(Clk), .Q(net644655), .QN(
        n6067) );
  DFF_X1 \REGISTERS_reg[19][11]  ( .D(n3155), .CK(Clk), .Q(net644654), .QN(
        n6066) );
  DFF_X1 \REGISTERS_reg[19][10]  ( .D(n3154), .CK(Clk), .Q(net644653), .QN(
        n6065) );
  DFF_X1 \REGISTERS_reg[19][9]  ( .D(n3153), .CK(Clk), .Q(net644652), .QN(
        n6064) );
  DFF_X1 \REGISTERS_reg[19][8]  ( .D(n3152), .CK(Clk), .Q(net644651), .QN(
        n6063) );
  DFF_X1 \REGISTERS_reg[19][7]  ( .D(n3151), .CK(Clk), .Q(net644650), .QN(
        n6062) );
  DFF_X1 \REGISTERS_reg[19][6]  ( .D(n3150), .CK(Clk), .Q(net644649), .QN(
        n6061) );
  DFF_X1 \REGISTERS_reg[19][5]  ( .D(n3149), .CK(Clk), .Q(net644648), .QN(
        n6060) );
  DFF_X1 \REGISTERS_reg[19][4]  ( .D(n3148), .CK(Clk), .Q(net644647), .QN(
        n6059) );
  DFF_X1 \REGISTERS_reg[19][3]  ( .D(n3147), .CK(Clk), .Q(net644646), .QN(
        n6058) );
  DFF_X1 \REGISTERS_reg[19][2]  ( .D(n3146), .CK(Clk), .Q(net644645), .QN(
        n6057) );
  DFF_X1 \REGISTERS_reg[19][1]  ( .D(n3145), .CK(Clk), .Q(net644644), .QN(
        n6056) );
  DFF_X1 \REGISTERS_reg[19][0]  ( .D(n3144), .CK(Clk), .QN(n514) );
  DFF_X1 \REGISTERS_reg[20][31]  ( .D(n3143), .CK(Clk), .Q(net644643), .QN(
        n4874) );
  DFF_X1 \REGISTERS_reg[20][30]  ( .D(n3142), .CK(Clk), .Q(net644642), .QN(
        n4873) );
  DFF_X1 \REGISTERS_reg[20][29]  ( .D(n3141), .CK(Clk), .Q(net644641), .QN(
        n4869) );
  DFF_X1 \REGISTERS_reg[20][28]  ( .D(n3140), .CK(Clk), .Q(net644640), .QN(
        n4868) );
  DFF_X1 \REGISTERS_reg[20][27]  ( .D(n3139), .CK(Clk), .Q(net644639), .QN(
        n4863) );
  DFF_X1 \REGISTERS_reg[20][26]  ( .D(n3138), .CK(Clk), .Q(net644638), .QN(
        n4862) );
  DFF_X1 \REGISTERS_reg[20][25]  ( .D(n3137), .CK(Clk), .Q(net644637), .QN(
        n4853) );
  DFF_X1 \REGISTERS_reg[20][24]  ( .D(n3136), .CK(Clk), .Q(net644636), .QN(
        n4845) );
  DFF_X1 \REGISTERS_reg[20][23]  ( .D(n3135), .CK(Clk), .Q(net644635), .QN(
        n4844) );
  DFF_X1 \REGISTERS_reg[20][22]  ( .D(n3134), .CK(Clk), .Q(net644634), .QN(
        n4843) );
  DFF_X1 \REGISTERS_reg[20][21]  ( .D(n3133), .CK(Clk), .Q(net644633), .QN(
        n4839) );
  DFF_X1 \REGISTERS_reg[20][20]  ( .D(n3132), .CK(Clk), .Q(net644632), .QN(
        n4838) );
  DFF_X1 \REGISTERS_reg[20][19]  ( .D(n3131), .CK(Clk), .Q(net644631), .QN(
        n4833) );
  DFF_X1 \REGISTERS_reg[20][18]  ( .D(n3130), .CK(Clk), .Q(net644630), .QN(
        n4832) );
  DFF_X1 \REGISTERS_reg[20][17]  ( .D(n3129), .CK(Clk), .Q(net644629), .QN(
        n4823) );
  DFF_X1 \REGISTERS_reg[20][16]  ( .D(n3128), .CK(Clk), .Q(net644628), .QN(
        n4815) );
  DFF_X1 \REGISTERS_reg[20][15]  ( .D(n3127), .CK(Clk), .Q(net644627), .QN(
        n4814) );
  DFF_X1 \REGISTERS_reg[20][14]  ( .D(n3126), .CK(Clk), .Q(net644626), .QN(
        n4813) );
  DFF_X1 \REGISTERS_reg[20][13]  ( .D(n3125), .CK(Clk), .Q(net644625), .QN(
        n4809) );
  DFF_X1 \REGISTERS_reg[20][12]  ( .D(n3124), .CK(Clk), .Q(net644624), .QN(
        n4808) );
  DFF_X1 \REGISTERS_reg[20][11]  ( .D(n3123), .CK(Clk), .Q(net644623), .QN(
        n4803) );
  DFF_X1 \REGISTERS_reg[20][10]  ( .D(n3122), .CK(Clk), .Q(net644622), .QN(
        n4802) );
  DFF_X1 \REGISTERS_reg[20][9]  ( .D(n3121), .CK(Clk), .Q(net644621), .QN(
        n4793) );
  DFF_X1 \REGISTERS_reg[20][8]  ( .D(n3120), .CK(Clk), .Q(net644620), .QN(
        n4785) );
  DFF_X1 \REGISTERS_reg[20][7]  ( .D(n3119), .CK(Clk), .Q(net644619), .QN(
        n4784) );
  DFF_X1 \REGISTERS_reg[20][6]  ( .D(n3118), .CK(Clk), .Q(net644618), .QN(
        n4783) );
  DFF_X1 \REGISTERS_reg[20][5]  ( .D(n3117), .CK(Clk), .Q(net644617), .QN(
        n4779) );
  DFF_X1 \REGISTERS_reg[20][4]  ( .D(n3116), .CK(Clk), .Q(net644616), .QN(
        n4778) );
  DFF_X1 \REGISTERS_reg[20][3]  ( .D(n3115), .CK(Clk), .Q(net644615), .QN(
        n4773) );
  DFF_X1 \REGISTERS_reg[20][2]  ( .D(n3114), .CK(Clk), .Q(net644614), .QN(
        n4772) );
  DFF_X1 \REGISTERS_reg[20][1]  ( .D(n3113), .CK(Clk), .Q(net644613), .QN(
        n4763) );
  DFF_X1 \REGISTERS_reg[20][0]  ( .D(n3112), .CK(Clk), .Q(net644612), .QN(
        n6341) );
  DFF_X1 \REGISTERS_reg[21][31]  ( .D(n3111), .CK(Clk), .Q(net644611), .QN(
        n4755) );
  DFF_X1 \REGISTERS_reg[21][30]  ( .D(n3110), .CK(Clk), .Q(net644610), .QN(
        n4754) );
  DFF_X1 \REGISTERS_reg[21][29]  ( .D(n3109), .CK(Clk), .Q(net644609), .QN(
        n4753) );
  DFF_X1 \REGISTERS_reg[21][28]  ( .D(n3108), .CK(Clk), .Q(net644608), .QN(
        n4749) );
  DFF_X1 \REGISTERS_reg[21][27]  ( .D(n3107), .CK(Clk), .Q(net644607), .QN(
        n4748) );
  DFF_X1 \REGISTERS_reg[21][26]  ( .D(n3106), .CK(Clk), .Q(net644606), .QN(
        n4743) );
  DFF_X1 \REGISTERS_reg[21][25]  ( .D(n3105), .CK(Clk), .Q(net644605), .QN(
        n4742) );
  DFF_X1 \REGISTERS_reg[21][24]  ( .D(n3104), .CK(Clk), .Q(net644604), .QN(
        n4733) );
  DFF_X1 \REGISTERS_reg[21][23]  ( .D(n3103), .CK(Clk), .Q(net644603), .QN(
        n4725) );
  DFF_X1 \REGISTERS_reg[21][22]  ( .D(n3102), .CK(Clk), .Q(net644602), .QN(
        n4724) );
  DFF_X1 \REGISTERS_reg[21][21]  ( .D(n3101), .CK(Clk), .Q(net644601), .QN(
        n4723) );
  DFF_X1 \REGISTERS_reg[21][20]  ( .D(n3100), .CK(Clk), .Q(net644600), .QN(
        n4719) );
  DFF_X1 \REGISTERS_reg[21][19]  ( .D(n3099), .CK(Clk), .Q(net644599), .QN(
        n4718) );
  DFF_X1 \REGISTERS_reg[21][18]  ( .D(n3098), .CK(Clk), .Q(net644598), .QN(
        n4713) );
  DFF_X1 \REGISTERS_reg[21][17]  ( .D(n3097), .CK(Clk), .Q(net644597), .QN(
        n4712) );
  DFF_X1 \REGISTERS_reg[21][16]  ( .D(n3096), .CK(Clk), .Q(net644596), .QN(
        n4703) );
  DFF_X1 \REGISTERS_reg[21][15]  ( .D(n3095), .CK(Clk), .Q(net644595), .QN(
        n4695) );
  DFF_X1 \REGISTERS_reg[21][14]  ( .D(n3094), .CK(Clk), .Q(net644594), .QN(
        n4694) );
  DFF_X1 \REGISTERS_reg[21][13]  ( .D(n3093), .CK(Clk), .Q(net644593), .QN(
        n4693) );
  DFF_X1 \REGISTERS_reg[21][12]  ( .D(n3092), .CK(Clk), .Q(net644592), .QN(
        n4689) );
  DFF_X1 \REGISTERS_reg[21][11]  ( .D(n3091), .CK(Clk), .Q(net644591), .QN(
        n4688) );
  DFF_X1 \REGISTERS_reg[21][10]  ( .D(n3090), .CK(Clk), .Q(net644590), .QN(
        n4683) );
  DFF_X1 \REGISTERS_reg[21][9]  ( .D(n3089), .CK(Clk), .Q(net644589), .QN(
        n4682) );
  DFF_X1 \REGISTERS_reg[21][8]  ( .D(n3088), .CK(Clk), .Q(net644588), .QN(
        n4673) );
  DFF_X1 \REGISTERS_reg[21][7]  ( .D(n3087), .CK(Clk), .Q(net644587), .QN(
        n4665) );
  DFF_X1 \REGISTERS_reg[21][6]  ( .D(n3086), .CK(Clk), .Q(net644586), .QN(
        n4664) );
  DFF_X1 \REGISTERS_reg[21][5]  ( .D(n3085), .CK(Clk), .Q(net644585), .QN(
        n4663) );
  DFF_X1 \REGISTERS_reg[21][4]  ( .D(n3084), .CK(Clk), .Q(net644584), .QN(
        n4659) );
  DFF_X1 \REGISTERS_reg[21][3]  ( .D(n3083), .CK(Clk), .Q(net644583), .QN(
        n4658) );
  DFF_X1 \REGISTERS_reg[21][2]  ( .D(n3082), .CK(Clk), .Q(net644582), .QN(
        n4653) );
  DFF_X1 \REGISTERS_reg[21][1]  ( .D(n3081), .CK(Clk), .Q(net644581), .QN(
        n4652) );
  DFF_X1 \REGISTERS_reg[21][0]  ( .D(n3080), .CK(Clk), .Q(net644580), .QN(
        n6340) );
  DFF_X1 \REGISTERS_reg[22][31]  ( .D(n3079), .CK(Clk), .QN(n515) );
  DFF_X1 \REGISTERS_reg[22][30]  ( .D(n3078), .CK(Clk), .QN(n516) );
  DFF_X1 \REGISTERS_reg[22][29]  ( .D(n3077), .CK(Clk), .QN(n517) );
  DFF_X1 \REGISTERS_reg[22][28]  ( .D(n3076), .CK(Clk), .QN(n518) );
  DFF_X1 \REGISTERS_reg[22][27]  ( .D(n3075), .CK(Clk), .QN(n519) );
  DFF_X1 \REGISTERS_reg[22][26]  ( .D(n3074), .CK(Clk), .QN(n520) );
  DFF_X1 \REGISTERS_reg[22][25]  ( .D(n3073), .CK(Clk), .QN(n521) );
  DFF_X1 \REGISTERS_reg[22][24]  ( .D(n3072), .CK(Clk), .QN(n522) );
  DFF_X1 \REGISTERS_reg[22][23]  ( .D(n3071), .CK(Clk), .QN(n523) );
  DFF_X1 \REGISTERS_reg[22][22]  ( .D(n3070), .CK(Clk), .QN(n524) );
  DFF_X1 \REGISTERS_reg[22][21]  ( .D(n3069), .CK(Clk), .QN(n525) );
  DFF_X1 \REGISTERS_reg[22][20]  ( .D(n3068), .CK(Clk), .QN(n526) );
  DFF_X1 \REGISTERS_reg[22][19]  ( .D(n3067), .CK(Clk), .QN(n527) );
  DFF_X1 \REGISTERS_reg[22][18]  ( .D(n3066), .CK(Clk), .QN(n528) );
  DFF_X1 \REGISTERS_reg[22][17]  ( .D(n3065), .CK(Clk), .QN(n529) );
  DFF_X1 \REGISTERS_reg[22][16]  ( .D(n3064), .CK(Clk), .QN(n530) );
  DFF_X1 \REGISTERS_reg[22][15]  ( .D(n3063), .CK(Clk), .QN(n531) );
  DFF_X1 \REGISTERS_reg[22][14]  ( .D(n3062), .CK(Clk), .QN(n532) );
  DFF_X1 \REGISTERS_reg[22][13]  ( .D(n3061), .CK(Clk), .QN(n533) );
  DFF_X1 \REGISTERS_reg[22][12]  ( .D(n3060), .CK(Clk), .QN(n534) );
  DFF_X1 \REGISTERS_reg[22][11]  ( .D(n3059), .CK(Clk), .QN(n535) );
  DFF_X1 \REGISTERS_reg[22][10]  ( .D(n3058), .CK(Clk), .QN(n536) );
  DFF_X1 \REGISTERS_reg[22][9]  ( .D(n3057), .CK(Clk), .QN(n537) );
  DFF_X1 \REGISTERS_reg[22][8]  ( .D(n3056), .CK(Clk), .QN(n538) );
  DFF_X1 \REGISTERS_reg[22][7]  ( .D(n3055), .CK(Clk), .QN(n539) );
  DFF_X1 \REGISTERS_reg[22][6]  ( .D(n3054), .CK(Clk), .QN(n540) );
  DFF_X1 \REGISTERS_reg[22][5]  ( .D(n3053), .CK(Clk), .QN(n541) );
  DFF_X1 \REGISTERS_reg[22][4]  ( .D(n3052), .CK(Clk), .QN(n542) );
  DFF_X1 \REGISTERS_reg[22][3]  ( .D(n3051), .CK(Clk), .QN(n543) );
  DFF_X1 \REGISTERS_reg[22][2]  ( .D(n3050), .CK(Clk), .QN(n544) );
  DFF_X1 \REGISTERS_reg[22][1]  ( .D(n3049), .CK(Clk), .QN(n545) );
  DFF_X1 \REGISTERS_reg[22][0]  ( .D(n3048), .CK(Clk), .QN(n671) );
  DFF_X1 \REGISTERS_reg[23][31]  ( .D(n3047), .CK(Clk), .Q(n4166), .QN(n672)
         );
  DFF_X1 \REGISTERS_reg[23][30]  ( .D(n3046), .CK(Clk), .Q(n4163), .QN(n673)
         );
  DFF_X1 \REGISTERS_reg[23][29]  ( .D(n3045), .CK(Clk), .Q(n4160), .QN(n674)
         );
  DFF_X1 \REGISTERS_reg[23][28]  ( .D(n3044), .CK(Clk), .Q(n4157), .QN(n675)
         );
  DFF_X1 \REGISTERS_reg[23][27]  ( .D(n3043), .CK(Clk), .Q(n4154), .QN(n676)
         );
  DFF_X1 \REGISTERS_reg[23][26]  ( .D(n3042), .CK(Clk), .Q(n4151), .QN(n677)
         );
  DFF_X1 \REGISTERS_reg[23][25]  ( .D(n3041), .CK(Clk), .Q(n4148), .QN(n678)
         );
  DFF_X1 \REGISTERS_reg[23][24]  ( .D(n3040), .CK(Clk), .Q(n4142), .QN(n679)
         );
  DFF_X1 \REGISTERS_reg[23][23]  ( .D(n3039), .CK(Clk), .Q(n4139), .QN(n680)
         );
  DFF_X1 \REGISTERS_reg[23][22]  ( .D(n3038), .CK(Clk), .Q(n4136), .QN(n681)
         );
  DFF_X1 \REGISTERS_reg[23][21]  ( .D(n3037), .CK(Clk), .Q(n4133), .QN(n682)
         );
  DFF_X1 \REGISTERS_reg[23][20]  ( .D(n3036), .CK(Clk), .Q(n4130), .QN(n683)
         );
  DFF_X1 \REGISTERS_reg[23][19]  ( .D(n3035), .CK(Clk), .Q(n4127), .QN(n684)
         );
  DFF_X1 \REGISTERS_reg[23][18]  ( .D(n3034), .CK(Clk), .Q(n4124), .QN(n685)
         );
  DFF_X1 \REGISTERS_reg[23][17]  ( .D(n3033), .CK(Clk), .Q(n4121), .QN(n686)
         );
  DFF_X1 \REGISTERS_reg[23][16]  ( .D(n3032), .CK(Clk), .Q(n4118), .QN(n687)
         );
  DFF_X1 \REGISTERS_reg[23][15]  ( .D(n3031), .CK(Clk), .Q(n4115), .QN(n688)
         );
  DFF_X1 \REGISTERS_reg[23][14]  ( .D(n3030), .CK(Clk), .Q(n4112), .QN(n689)
         );
  DFF_X1 \REGISTERS_reg[23][13]  ( .D(n3029), .CK(Clk), .Q(n4104), .QN(n690)
         );
  DFF_X1 \REGISTERS_reg[23][12]  ( .D(n3028), .CK(Clk), .Q(n4101), .QN(n691)
         );
  DFF_X1 \REGISTERS_reg[23][11]  ( .D(n3027), .CK(Clk), .Q(n4098), .QN(n692)
         );
  DFF_X1 \REGISTERS_reg[23][10]  ( .D(n3026), .CK(Clk), .Q(n4095), .QN(n693)
         );
  DFF_X1 \REGISTERS_reg[23][9]  ( .D(n3025), .CK(Clk), .Q(n4092), .QN(n694) );
  DFF_X1 \REGISTERS_reg[23][8]  ( .D(n3024), .CK(Clk), .Q(n4089), .QN(n695) );
  DFF_X1 \REGISTERS_reg[23][7]  ( .D(n3023), .CK(Clk), .Q(n4086), .QN(n696) );
  DFF_X1 \REGISTERS_reg[23][6]  ( .D(n3022), .CK(Clk), .Q(n4083), .QN(n697) );
  DFF_X1 \REGISTERS_reg[23][5]  ( .D(n3021), .CK(Clk), .Q(n4080), .QN(n698) );
  DFF_X1 \REGISTERS_reg[23][4]  ( .D(n3020), .CK(Clk), .Q(n4077), .QN(n699) );
  DFF_X1 \REGISTERS_reg[23][3]  ( .D(n3019), .CK(Clk), .Q(n4072), .QN(n700) );
  DFF_X1 \REGISTERS_reg[23][2]  ( .D(n3018), .CK(Clk), .Q(n4067), .QN(n701) );
  DFF_X1 \REGISTERS_reg[23][1]  ( .D(n3017), .CK(Clk), .Q(n4064), .QN(n702) );
  DFF_X1 \REGISTERS_reg[23][0]  ( .D(n3016), .CK(Clk), .Q(net644579), .QN(
        n6350) );
  DFF_X1 \REGISTERS_reg[24][31]  ( .D(n3015), .CK(Clk), .Q(net644578), .QN(
        n6149) );
  DFF_X1 \REGISTERS_reg[24][30]  ( .D(n3014), .CK(Clk), .Q(net644577), .QN(
        n6148) );
  DFF_X1 \REGISTERS_reg[24][29]  ( .D(n3013), .CK(Clk), .Q(net644576), .QN(
        n6147) );
  DFF_X1 \REGISTERS_reg[24][28]  ( .D(n3012), .CK(Clk), .Q(net644575), .QN(
        n6146) );
  DFF_X1 \REGISTERS_reg[24][27]  ( .D(n3011), .CK(Clk), .Q(net644574), .QN(
        n6145) );
  DFF_X1 \REGISTERS_reg[24][26]  ( .D(n3010), .CK(Clk), .Q(net644573), .QN(
        n6144) );
  DFF_X1 \REGISTERS_reg[24][25]  ( .D(n3009), .CK(Clk), .Q(net644572), .QN(
        n6143) );
  DFF_X1 \REGISTERS_reg[24][24]  ( .D(n3008), .CK(Clk), .Q(net644571), .QN(
        n6142) );
  DFF_X1 \REGISTERS_reg[24][23]  ( .D(n3007), .CK(Clk), .Q(net644570), .QN(
        n6141) );
  DFF_X1 \REGISTERS_reg[24][22]  ( .D(n3006), .CK(Clk), .Q(net644569), .QN(
        n6140) );
  DFF_X1 \REGISTERS_reg[24][21]  ( .D(n3005), .CK(Clk), .Q(net644568), .QN(
        n6139) );
  DFF_X1 \REGISTERS_reg[24][20]  ( .D(n3004), .CK(Clk), .Q(net644567), .QN(
        n6138) );
  DFF_X1 \REGISTERS_reg[24][19]  ( .D(n3003), .CK(Clk), .Q(net644566), .QN(
        n6137) );
  DFF_X1 \REGISTERS_reg[24][18]  ( .D(n3002), .CK(Clk), .Q(net644565), .QN(
        n6136) );
  DFF_X1 \REGISTERS_reg[24][17]  ( .D(n3001), .CK(Clk), .Q(net644564), .QN(
        n6135) );
  DFF_X1 \REGISTERS_reg[24][16]  ( .D(n3000), .CK(Clk), .Q(net644563), .QN(
        n6134) );
  DFF_X1 \REGISTERS_reg[24][15]  ( .D(n2999), .CK(Clk), .Q(net644562), .QN(
        n6133) );
  DFF_X1 \REGISTERS_reg[24][14]  ( .D(n2998), .CK(Clk), .Q(net644561), .QN(
        n6132) );
  DFF_X1 \REGISTERS_reg[24][13]  ( .D(n2997), .CK(Clk), .Q(net644560), .QN(
        n6131) );
  DFF_X1 \REGISTERS_reg[24][12]  ( .D(n2996), .CK(Clk), .Q(net644559), .QN(
        n6130) );
  DFF_X1 \REGISTERS_reg[24][11]  ( .D(n2995), .CK(Clk), .Q(net644558), .QN(
        n6129) );
  DFF_X1 \REGISTERS_reg[24][10]  ( .D(n2994), .CK(Clk), .Q(net644557), .QN(
        n6128) );
  DFF_X1 \REGISTERS_reg[24][9]  ( .D(n2993), .CK(Clk), .Q(net644556), .QN(
        n6127) );
  DFF_X1 \REGISTERS_reg[24][8]  ( .D(n2992), .CK(Clk), .Q(net644555), .QN(
        n6126) );
  DFF_X1 \REGISTERS_reg[24][7]  ( .D(n2991), .CK(Clk), .Q(net644554), .QN(
        n6125) );
  DFF_X1 \REGISTERS_reg[24][6]  ( .D(n2990), .CK(Clk), .Q(net644553), .QN(
        n6124) );
  DFF_X1 \REGISTERS_reg[24][5]  ( .D(n2989), .CK(Clk), .Q(net644552), .QN(
        n6123) );
  DFF_X1 \REGISTERS_reg[24][4]  ( .D(n2988), .CK(Clk), .Q(net644551), .QN(
        n6122) );
  DFF_X1 \REGISTERS_reg[24][3]  ( .D(n2987), .CK(Clk), .Q(net644550), .QN(
        n6121) );
  DFF_X1 \REGISTERS_reg[24][2]  ( .D(n2986), .CK(Clk), .Q(net644549), .QN(
        n6120) );
  DFF_X1 \REGISTERS_reg[24][1]  ( .D(n2985), .CK(Clk), .Q(net644548), .QN(
        n6119) );
  DFF_X1 \REGISTERS_reg[24][0]  ( .D(n2984), .CK(Clk), .Q(net644547), .QN(
        n6349) );
  DFF_X1 \REGISTERS_reg[25][31]  ( .D(n2983), .CK(Clk), .Q(net644546), .QN(
        n6180) );
  DFF_X1 \REGISTERS_reg[25][30]  ( .D(n2982), .CK(Clk), .Q(net644545), .QN(
        n6179) );
  DFF_X1 \REGISTERS_reg[25][29]  ( .D(n2981), .CK(Clk), .Q(net644544), .QN(
        n6178) );
  DFF_X1 \REGISTERS_reg[25][28]  ( .D(n2980), .CK(Clk), .Q(net644543), .QN(
        n6177) );
  DFF_X1 \REGISTERS_reg[25][27]  ( .D(n2979), .CK(Clk), .Q(net644542), .QN(
        n6176) );
  DFF_X1 \REGISTERS_reg[25][26]  ( .D(n2978), .CK(Clk), .Q(net644541), .QN(
        n6175) );
  DFF_X1 \REGISTERS_reg[25][25]  ( .D(n2977), .CK(Clk), .Q(net644540), .QN(
        n6174) );
  DFF_X1 \REGISTERS_reg[25][24]  ( .D(n2976), .CK(Clk), .Q(net644539), .QN(
        n6173) );
  DFF_X1 \REGISTERS_reg[25][23]  ( .D(n2975), .CK(Clk), .Q(net644538), .QN(
        n6172) );
  DFF_X1 \REGISTERS_reg[25][22]  ( .D(n2974), .CK(Clk), .Q(net644537), .QN(
        n6171) );
  DFF_X1 \REGISTERS_reg[25][21]  ( .D(n2973), .CK(Clk), .Q(net644536), .QN(
        n6170) );
  DFF_X1 \REGISTERS_reg[25][20]  ( .D(n2972), .CK(Clk), .Q(net644535), .QN(
        n6169) );
  DFF_X1 \REGISTERS_reg[25][19]  ( .D(n2971), .CK(Clk), .Q(net644534), .QN(
        n6168) );
  DFF_X1 \REGISTERS_reg[25][18]  ( .D(n2970), .CK(Clk), .Q(net644533), .QN(
        n6167) );
  DFF_X1 \REGISTERS_reg[25][17]  ( .D(n2969), .CK(Clk), .Q(net644532), .QN(
        n6166) );
  DFF_X1 \REGISTERS_reg[25][16]  ( .D(n2968), .CK(Clk), .Q(net644531), .QN(
        n6165) );
  DFF_X1 \REGISTERS_reg[25][15]  ( .D(n2967), .CK(Clk), .Q(net644530), .QN(
        n6164) );
  DFF_X1 \REGISTERS_reg[25][14]  ( .D(n2966), .CK(Clk), .Q(net644529), .QN(
        n6163) );
  DFF_X1 \REGISTERS_reg[25][13]  ( .D(n2965), .CK(Clk), .Q(net644528), .QN(
        n6162) );
  DFF_X1 \REGISTERS_reg[25][12]  ( .D(n2964), .CK(Clk), .Q(net644527), .QN(
        n6161) );
  DFF_X1 \REGISTERS_reg[25][11]  ( .D(n2963), .CK(Clk), .Q(net644526), .QN(
        n6160) );
  DFF_X1 \REGISTERS_reg[25][10]  ( .D(n2962), .CK(Clk), .Q(net644525), .QN(
        n6159) );
  DFF_X1 \REGISTERS_reg[25][9]  ( .D(n2961), .CK(Clk), .Q(net644524), .QN(
        n6158) );
  DFF_X1 \REGISTERS_reg[25][8]  ( .D(n2960), .CK(Clk), .Q(net644523), .QN(
        n6157) );
  DFF_X1 \REGISTERS_reg[25][7]  ( .D(n2959), .CK(Clk), .Q(net644522), .QN(
        n6156) );
  DFF_X1 \REGISTERS_reg[25][6]  ( .D(n2958), .CK(Clk), .Q(net644521), .QN(
        n6155) );
  DFF_X1 \REGISTERS_reg[25][5]  ( .D(n2957), .CK(Clk), .Q(net644520), .QN(
        n6154) );
  DFF_X1 \REGISTERS_reg[25][4]  ( .D(n2956), .CK(Clk), .Q(net644519), .QN(
        n6153) );
  DFF_X1 \REGISTERS_reg[25][3]  ( .D(n2955), .CK(Clk), .Q(net644518), .QN(
        n6152) );
  DFF_X1 \REGISTERS_reg[25][2]  ( .D(n2954), .CK(Clk), .Q(net644517), .QN(
        n6151) );
  DFF_X1 \REGISTERS_reg[25][1]  ( .D(n2953), .CK(Clk), .Q(net644516), .QN(
        n6150) );
  DFF_X1 \REGISTERS_reg[25][0]  ( .D(n2952), .CK(Clk), .Q(net644515), .QN(
        n6339) );
  DFF_X1 \REGISTERS_reg[26][31]  ( .D(n2951), .CK(Clk), .Q(n4164), .QN(n2248)
         );
  DFF_X1 \REGISTERS_reg[26][30]  ( .D(n2950), .CK(Clk), .Q(n4161), .QN(n2247)
         );
  DFF_X1 \REGISTERS_reg[26][29]  ( .D(n2949), .CK(Clk), .Q(n4158), .QN(n2246)
         );
  DFF_X1 \REGISTERS_reg[26][28]  ( .D(n2948), .CK(Clk), .Q(n4155), .QN(n2245)
         );
  DFF_X1 \REGISTERS_reg[26][27]  ( .D(n2947), .CK(Clk), .Q(n4152), .QN(n2244)
         );
  DFF_X1 \REGISTERS_reg[26][26]  ( .D(n2946), .CK(Clk), .Q(n4149), .QN(n2243)
         );
  DFF_X1 \REGISTERS_reg[26][25]  ( .D(n2945), .CK(Clk), .Q(n4144), .QN(n2242)
         );
  DFF_X1 \REGISTERS_reg[26][24]  ( .D(n2944), .CK(Clk), .Q(n4140), .QN(n2241)
         );
  DFF_X1 \REGISTERS_reg[26][23]  ( .D(n2943), .CK(Clk), .Q(n4137), .QN(n2240)
         );
  DFF_X1 \REGISTERS_reg[26][22]  ( .D(n2942), .CK(Clk), .Q(n4134), .QN(n2239)
         );
  DFF_X1 \REGISTERS_reg[26][21]  ( .D(n2941), .CK(Clk), .Q(n4131), .QN(n2238)
         );
  DFF_X1 \REGISTERS_reg[26][20]  ( .D(n2940), .CK(Clk), .Q(n4128), .QN(n2237)
         );
  DFF_X1 \REGISTERS_reg[26][19]  ( .D(n2939), .CK(Clk), .Q(n4125), .QN(n2236)
         );
  DFF_X1 \REGISTERS_reg[26][18]  ( .D(n2938), .CK(Clk), .Q(n4122), .QN(n2235)
         );
  DFF_X1 \REGISTERS_reg[26][17]  ( .D(n2937), .CK(Clk), .Q(n4119), .QN(n2234)
         );
  DFF_X1 \REGISTERS_reg[26][16]  ( .D(n2936), .CK(Clk), .Q(n4116), .QN(n2233)
         );
  DFF_X1 \REGISTERS_reg[26][15]  ( .D(n2935), .CK(Clk), .Q(n4113), .QN(n2232)
         );
  DFF_X1 \REGISTERS_reg[26][14]  ( .D(n2934), .CK(Clk), .Q(n4105), .QN(n2231)
         );
  DFF_X1 \REGISTERS_reg[26][13]  ( .D(n2933), .CK(Clk), .Q(n4102), .QN(n2230)
         );
  DFF_X1 \REGISTERS_reg[26][12]  ( .D(n2932), .CK(Clk), .Q(n4099), .QN(n2229)
         );
  DFF_X1 \REGISTERS_reg[26][11]  ( .D(n2931), .CK(Clk), .Q(n4096), .QN(n2228)
         );
  DFF_X1 \REGISTERS_reg[26][10]  ( .D(n2930), .CK(Clk), .Q(n4093), .QN(n2227)
         );
  DFF_X1 \REGISTERS_reg[26][9]  ( .D(n2929), .CK(Clk), .Q(n4090), .QN(n2226)
         );
  DFF_X1 \REGISTERS_reg[26][8]  ( .D(n2928), .CK(Clk), .Q(n4087), .QN(n2225)
         );
  DFF_X1 \REGISTERS_reg[26][7]  ( .D(n2927), .CK(Clk), .Q(n4084), .QN(n2224)
         );
  DFF_X1 \REGISTERS_reg[26][6]  ( .D(n2926), .CK(Clk), .Q(n4081), .QN(n2223)
         );
  DFF_X1 \REGISTERS_reg[26][5]  ( .D(n2925), .CK(Clk), .Q(n4078), .QN(n2222)
         );
  DFF_X1 \REGISTERS_reg[26][4]  ( .D(n2924), .CK(Clk), .Q(n4075), .QN(n2221)
         );
  DFF_X1 \REGISTERS_reg[26][3]  ( .D(n2923), .CK(Clk), .Q(n4070), .QN(n2220)
         );
  DFF_X1 \REGISTERS_reg[26][2]  ( .D(n2922), .CK(Clk), .Q(n4065), .QN(n2219)
         );
  DFF_X1 \REGISTERS_reg[26][1]  ( .D(n2921), .CK(Clk), .Q(n222), .QN(n6243) );
  DFF_X1 \REGISTERS_reg[26][0]  ( .D(n2920), .CK(Clk), .Q(n385), .QN(n4167) );
  DFF_X1 \REGISTERS_reg[27][31]  ( .D(n2919), .CK(Clk), .Q(net644514), .QN(
        n6242) );
  DFF_X1 \REGISTERS_reg[27][30]  ( .D(n2918), .CK(Clk), .Q(net644513), .QN(
        n6241) );
  DFF_X1 \REGISTERS_reg[27][29]  ( .D(n2917), .CK(Clk), .Q(net644512), .QN(
        n6240) );
  DFF_X1 \REGISTERS_reg[27][28]  ( .D(n2916), .CK(Clk), .Q(net644511), .QN(
        n6239) );
  DFF_X1 \REGISTERS_reg[27][27]  ( .D(n2915), .CK(Clk), .Q(net644510), .QN(
        n6238) );
  DFF_X1 \REGISTERS_reg[27][26]  ( .D(n2914), .CK(Clk), .Q(net644509), .QN(
        n6237) );
  DFF_X1 \REGISTERS_reg[27][25]  ( .D(n2913), .CK(Clk), .Q(net644508), .QN(
        n6236) );
  DFF_X1 \REGISTERS_reg[27][24]  ( .D(n2912), .CK(Clk), .Q(net644507), .QN(
        n6235) );
  DFF_X1 \REGISTERS_reg[27][23]  ( .D(n2911), .CK(Clk), .Q(net644506), .QN(
        n6234) );
  DFF_X1 \REGISTERS_reg[27][22]  ( .D(n2910), .CK(Clk), .Q(net644505), .QN(
        n6233) );
  DFF_X1 \REGISTERS_reg[27][21]  ( .D(n2909), .CK(Clk), .Q(net644504), .QN(
        n6232) );
  DFF_X1 \REGISTERS_reg[27][20]  ( .D(n2908), .CK(Clk), .Q(net644503), .QN(
        n6231) );
  DFF_X1 \REGISTERS_reg[27][19]  ( .D(n2907), .CK(Clk), .Q(net644502), .QN(
        n6230) );
  DFF_X1 \REGISTERS_reg[27][18]  ( .D(n2906), .CK(Clk), .Q(net644501), .QN(
        n6229) );
  DFF_X1 \REGISTERS_reg[27][17]  ( .D(n2905), .CK(Clk), .Q(net644500), .QN(
        n6228) );
  DFF_X1 \REGISTERS_reg[27][16]  ( .D(n2904), .CK(Clk), .Q(net644499), .QN(
        n6227) );
  DFF_X1 \REGISTERS_reg[27][15]  ( .D(n2903), .CK(Clk), .Q(net644498), .QN(
        n6226) );
  DFF_X1 \REGISTERS_reg[27][14]  ( .D(n2902), .CK(Clk), .Q(net644497), .QN(
        n6225) );
  DFF_X1 \REGISTERS_reg[27][13]  ( .D(n2901), .CK(Clk), .Q(net644496), .QN(
        n6224) );
  DFF_X1 \REGISTERS_reg[27][12]  ( .D(n2900), .CK(Clk), .Q(net644495), .QN(
        n6223) );
  DFF_X1 \REGISTERS_reg[27][11]  ( .D(n2899), .CK(Clk), .Q(net644494), .QN(
        n6222) );
  DFF_X1 \REGISTERS_reg[27][10]  ( .D(n2898), .CK(Clk), .Q(net644493), .QN(
        n6221) );
  DFF_X1 \REGISTERS_reg[27][9]  ( .D(n2897), .CK(Clk), .Q(net644492), .QN(
        n6220) );
  DFF_X1 \REGISTERS_reg[27][8]  ( .D(n2896), .CK(Clk), .Q(net644491), .QN(
        n6219) );
  DFF_X1 \REGISTERS_reg[27][7]  ( .D(n2895), .CK(Clk), .Q(net644490), .QN(
        n6218) );
  DFF_X1 \REGISTERS_reg[27][6]  ( .D(n2894), .CK(Clk), .Q(net644489), .QN(
        n6217) );
  DFF_X1 \REGISTERS_reg[27][5]  ( .D(n2893), .CK(Clk), .Q(net644488), .QN(
        n6216) );
  DFF_X1 \REGISTERS_reg[27][4]  ( .D(n2892), .CK(Clk), .Q(net644487), .QN(
        n6215) );
  DFF_X1 \REGISTERS_reg[27][3]  ( .D(n2891), .CK(Clk), .Q(net644486), .QN(
        n6214) );
  DFF_X1 \REGISTERS_reg[27][2]  ( .D(n2890), .CK(Clk), .Q(net644485), .QN(
        n6213) );
  DFF_X1 \REGISTERS_reg[27][1]  ( .D(n2889), .CK(Clk), .Q(net644484), .QN(
        n6212) );
  DFF_X1 \REGISTERS_reg[27][0]  ( .D(n2888), .CK(Clk), .Q(net644483), .QN(
        n6348) );
  DFF_X1 \REGISTERS_reg[28][31]  ( .D(n2887), .CK(Clk), .QN(n546) );
  DFF_X1 \REGISTERS_reg[28][30]  ( .D(n2886), .CK(Clk), .QN(n547) );
  DFF_X1 \REGISTERS_reg[28][29]  ( .D(n2885), .CK(Clk), .QN(n548) );
  DFF_X1 \REGISTERS_reg[28][28]  ( .D(n2884), .CK(Clk), .QN(n549) );
  DFF_X1 \REGISTERS_reg[28][27]  ( .D(n2883), .CK(Clk), .QN(n550) );
  DFF_X1 \REGISTERS_reg[28][26]  ( .D(n2882), .CK(Clk), .QN(n551) );
  DFF_X1 \REGISTERS_reg[28][25]  ( .D(n2881), .CK(Clk), .QN(n552) );
  DFF_X1 \REGISTERS_reg[28][24]  ( .D(n2880), .CK(Clk), .QN(n553) );
  DFF_X1 \REGISTERS_reg[28][23]  ( .D(n2879), .CK(Clk), .QN(n554) );
  DFF_X1 \REGISTERS_reg[28][22]  ( .D(n2878), .CK(Clk), .QN(n555) );
  DFF_X1 \REGISTERS_reg[28][21]  ( .D(n2877), .CK(Clk), .QN(n556) );
  DFF_X1 \REGISTERS_reg[28][20]  ( .D(n2876), .CK(Clk), .QN(n557) );
  DFF_X1 \REGISTERS_reg[28][19]  ( .D(n2875), .CK(Clk), .QN(n558) );
  DFF_X1 \REGISTERS_reg[28][18]  ( .D(n2874), .CK(Clk), .QN(n559) );
  DFF_X1 \REGISTERS_reg[28][17]  ( .D(n2873), .CK(Clk), .QN(n560) );
  DFF_X1 \REGISTERS_reg[28][16]  ( .D(n2872), .CK(Clk), .QN(n561) );
  DFF_X1 \REGISTERS_reg[28][15]  ( .D(n2871), .CK(Clk), .QN(n562) );
  DFF_X1 \REGISTERS_reg[28][14]  ( .D(n2870), .CK(Clk), .QN(n563) );
  DFF_X1 \REGISTERS_reg[28][13]  ( .D(n2869), .CK(Clk), .QN(n564) );
  DFF_X1 \REGISTERS_reg[28][12]  ( .D(n2868), .CK(Clk), .QN(n565) );
  DFF_X1 \REGISTERS_reg[28][11]  ( .D(n2867), .CK(Clk), .QN(n566) );
  DFF_X1 \REGISTERS_reg[28][10]  ( .D(n2866), .CK(Clk), .QN(n567) );
  DFF_X1 \REGISTERS_reg[28][9]  ( .D(n2865), .CK(Clk), .QN(n568) );
  DFF_X1 \REGISTERS_reg[28][8]  ( .D(n2864), .CK(Clk), .QN(n569) );
  DFF_X1 \REGISTERS_reg[28][7]  ( .D(n2863), .CK(Clk), .QN(n570) );
  DFF_X1 \REGISTERS_reg[28][6]  ( .D(n2862), .CK(Clk), .QN(n571) );
  DFF_X1 \REGISTERS_reg[28][5]  ( .D(n2861), .CK(Clk), .QN(n572) );
  DFF_X1 \REGISTERS_reg[28][4]  ( .D(n2860), .CK(Clk), .QN(n573) );
  DFF_X1 \REGISTERS_reg[28][3]  ( .D(n2859), .CK(Clk), .QN(n574) );
  DFF_X1 \REGISTERS_reg[28][2]  ( .D(n2858), .CK(Clk), .QN(n575) );
  DFF_X1 \REGISTERS_reg[28][1]  ( .D(n2857), .CK(Clk), .QN(n576) );
  DFF_X1 \REGISTERS_reg[28][0]  ( .D(n2856), .CK(Clk), .QN(n703) );
  DFF_X1 \REGISTERS_reg[29][31]  ( .D(n2855), .CK(Clk), .Q(net644482), .QN(
        n4643) );
  DFF_X1 \REGISTERS_reg[29][30]  ( .D(n2854), .CK(Clk), .Q(net644481), .QN(
        n4635) );
  DFF_X1 \REGISTERS_reg[29][29]  ( .D(n2853), .CK(Clk), .Q(net644480), .QN(
        n4634) );
  DFF_X1 \REGISTERS_reg[29][28]  ( .D(n2852), .CK(Clk), .Q(net644479), .QN(
        n4633) );
  DFF_X1 \REGISTERS_reg[29][27]  ( .D(n2851), .CK(Clk), .Q(net644478), .QN(
        n4629) );
  DFF_X1 \REGISTERS_reg[29][26]  ( .D(n2850), .CK(Clk), .Q(net644477), .QN(
        n4628) );
  DFF_X1 \REGISTERS_reg[29][25]  ( .D(n2849), .CK(Clk), .Q(net644476), .QN(
        n4623) );
  DFF_X1 \REGISTERS_reg[29][24]  ( .D(n2848), .CK(Clk), .Q(net644475), .QN(
        n4622) );
  DFF_X1 \REGISTERS_reg[29][23]  ( .D(n2847), .CK(Clk), .Q(net644474), .QN(
        n4613) );
  DFF_X1 \REGISTERS_reg[29][22]  ( .D(n2846), .CK(Clk), .Q(net644473), .QN(
        n4605) );
  DFF_X1 \REGISTERS_reg[29][21]  ( .D(n2845), .CK(Clk), .Q(net644472), .QN(
        n4604) );
  DFF_X1 \REGISTERS_reg[29][20]  ( .D(n2844), .CK(Clk), .Q(net644471), .QN(
        n4603) );
  DFF_X1 \REGISTERS_reg[29][19]  ( .D(n2843), .CK(Clk), .Q(net644470), .QN(
        n4599) );
  DFF_X1 \REGISTERS_reg[29][18]  ( .D(n2842), .CK(Clk), .Q(net644469), .QN(
        n4598) );
  DFF_X1 \REGISTERS_reg[29][17]  ( .D(n2841), .CK(Clk), .Q(net644468), .QN(
        n4593) );
  DFF_X1 \REGISTERS_reg[29][16]  ( .D(n2840), .CK(Clk), .Q(net644467), .QN(
        n4592) );
  DFF_X1 \REGISTERS_reg[29][15]  ( .D(n2839), .CK(Clk), .Q(net644466), .QN(
        n4583) );
  DFF_X1 \REGISTERS_reg[29][14]  ( .D(n2838), .CK(Clk), .Q(net644465), .QN(
        n4575) );
  DFF_X1 \REGISTERS_reg[29][13]  ( .D(n2837), .CK(Clk), .Q(net644464), .QN(
        n4574) );
  DFF_X1 \REGISTERS_reg[29][12]  ( .D(n2836), .CK(Clk), .Q(net644463), .QN(
        n4573) );
  DFF_X1 \REGISTERS_reg[29][11]  ( .D(n2835), .CK(Clk), .Q(net644462), .QN(
        n4569) );
  DFF_X1 \REGISTERS_reg[29][10]  ( .D(n2834), .CK(Clk), .Q(net644461), .QN(
        n4568) );
  DFF_X1 \REGISTERS_reg[29][9]  ( .D(n2833), .CK(Clk), .Q(net644460), .QN(
        n4563) );
  DFF_X1 \REGISTERS_reg[29][8]  ( .D(n2832), .CK(Clk), .Q(net644459), .QN(
        n4562) );
  DFF_X1 \REGISTERS_reg[29][7]  ( .D(n2831), .CK(Clk), .Q(net644458), .QN(
        n4553) );
  DFF_X1 \REGISTERS_reg[29][6]  ( .D(n2830), .CK(Clk), .Q(net644457), .QN(
        n4545) );
  DFF_X1 \REGISTERS_reg[29][5]  ( .D(n2829), .CK(Clk), .Q(net644456), .QN(
        n4544) );
  DFF_X1 \REGISTERS_reg[29][4]  ( .D(n2828), .CK(Clk), .Q(net644455), .QN(
        n4543) );
  DFF_X1 \REGISTERS_reg[29][3]  ( .D(n2827), .CK(Clk), .Q(net644454), .QN(
        n4539) );
  DFF_X1 \REGISTERS_reg[29][2]  ( .D(n2826), .CK(Clk), .Q(net644453), .QN(
        n4538) );
  DFF_X1 \REGISTERS_reg[29][1]  ( .D(n2825), .CK(Clk), .Q(net644452), .QN(
        n4533) );
  DFF_X1 \REGISTERS_reg[29][0]  ( .D(n2824), .CK(Clk), .Q(net644451), .QN(
        n6338) );
  DFF_X1 \REGISTERS_reg[30][31]  ( .D(n2823), .CK(Clk), .Q(net644450), .QN(
        n6211) );
  DFF_X1 \REGISTERS_reg[30][30]  ( .D(n2822), .CK(Clk), .Q(net644449), .QN(
        n6210) );
  DFF_X1 \REGISTERS_reg[30][29]  ( .D(n2821), .CK(Clk), .Q(net644448), .QN(
        n6209) );
  DFF_X1 \REGISTERS_reg[30][28]  ( .D(n2820), .CK(Clk), .Q(net644447), .QN(
        n6208) );
  DFF_X1 \REGISTERS_reg[30][27]  ( .D(n2819), .CK(Clk), .Q(net644446), .QN(
        n6207) );
  DFF_X1 \REGISTERS_reg[30][26]  ( .D(n2818), .CK(Clk), .Q(net644445), .QN(
        n6206) );
  DFF_X1 \REGISTERS_reg[30][25]  ( .D(n2817), .CK(Clk), .Q(net644444), .QN(
        n6205) );
  DFF_X1 \REGISTERS_reg[30][24]  ( .D(n2816), .CK(Clk), .Q(net644443), .QN(
        n6204) );
  DFF_X1 \REGISTERS_reg[30][23]  ( .D(n2815), .CK(Clk), .Q(net644442), .QN(
        n6203) );
  DFF_X1 \REGISTERS_reg[30][22]  ( .D(n2814), .CK(Clk), .Q(net644441), .QN(
        n6202) );
  DFF_X1 \REGISTERS_reg[30][21]  ( .D(n2813), .CK(Clk), .Q(net644440), .QN(
        n6201) );
  DFF_X1 \REGISTERS_reg[30][20]  ( .D(n2812), .CK(Clk), .Q(net644439), .QN(
        n6200) );
  DFF_X1 \REGISTERS_reg[30][19]  ( .D(n2811), .CK(Clk), .Q(net644438), .QN(
        n6199) );
  DFF_X1 \REGISTERS_reg[30][18]  ( .D(n2810), .CK(Clk), .Q(net644437), .QN(
        n6198) );
  DFF_X1 \REGISTERS_reg[30][17]  ( .D(n2809), .CK(Clk), .Q(net644436), .QN(
        n6197) );
  DFF_X1 \REGISTERS_reg[30][16]  ( .D(n2808), .CK(Clk), .Q(net644435), .QN(
        n6196) );
  DFF_X1 \REGISTERS_reg[30][15]  ( .D(n2807), .CK(Clk), .Q(net644434), .QN(
        n6195) );
  DFF_X1 \REGISTERS_reg[30][14]  ( .D(n2806), .CK(Clk), .Q(net644433), .QN(
        n6194) );
  DFF_X1 \REGISTERS_reg[30][13]  ( .D(n2805), .CK(Clk), .Q(net644432), .QN(
        n6193) );
  DFF_X1 \REGISTERS_reg[30][12]  ( .D(n2804), .CK(Clk), .Q(net644431), .QN(
        n6192) );
  DFF_X1 \REGISTERS_reg[30][11]  ( .D(n2803), .CK(Clk), .Q(net644430), .QN(
        n6191) );
  DFF_X1 \REGISTERS_reg[30][10]  ( .D(n2802), .CK(Clk), .Q(net644429), .QN(
        n6190) );
  DFF_X1 \REGISTERS_reg[30][9]  ( .D(n2801), .CK(Clk), .Q(net644428), .QN(
        n6189) );
  DFF_X1 \REGISTERS_reg[30][8]  ( .D(n2800), .CK(Clk), .Q(net644427), .QN(
        n6188) );
  DFF_X1 \REGISTERS_reg[30][7]  ( .D(n2799), .CK(Clk), .Q(net644426), .QN(
        n6187) );
  DFF_X1 \REGISTERS_reg[30][6]  ( .D(n2798), .CK(Clk), .Q(net644425), .QN(
        n6186) );
  DFF_X1 \REGISTERS_reg[30][5]  ( .D(n2797), .CK(Clk), .Q(net644424), .QN(
        n6185) );
  DFF_X1 \REGISTERS_reg[30][4]  ( .D(n2796), .CK(Clk), .Q(net644423), .QN(
        n6184) );
  DFF_X1 \REGISTERS_reg[30][3]  ( .D(n2795), .CK(Clk), .Q(net644422), .QN(
        n6183) );
  DFF_X1 \REGISTERS_reg[30][2]  ( .D(n2794), .CK(Clk), .Q(net644421), .QN(
        n6182) );
  DFF_X1 \REGISTERS_reg[30][1]  ( .D(n2793), .CK(Clk), .Q(net644420), .QN(
        n6181) );
  DFF_X1 \REGISTERS_reg[30][0]  ( .D(n2792), .CK(Clk), .Q(net644419), .QN(
        n6347) );
  DFF_X1 \REGISTERS_reg[31][31]  ( .D(n2791), .CK(Clk), .Q(n387), .QN(n4532)
         );
  DFF_X1 \OUT2_reg[31]  ( .D(n2790), .CK(Clk), .Q(OUT2[31]), .QN(net644418) );
  DFF_X1 \REGISTERS_reg[31][30]  ( .D(n2789), .CK(Clk), .Q(n390), .QN(n4523)
         );
  DFF_X1 \OUT2_reg[30]  ( .D(n2788), .CK(Clk), .Q(OUT2[30]), .QN(net644417) );
  DFF_X1 \REGISTERS_reg[31][29]  ( .D(n2787), .CK(Clk), .Q(n393), .QN(n4515)
         );
  DFF_X1 \OUT2_reg[29]  ( .D(n2786), .CK(Clk), .Q(OUT2[29]), .QN(net644416) );
  DFF_X1 \REGISTERS_reg[31][28]  ( .D(n2785), .CK(Clk), .Q(n396), .QN(n4514)
         );
  DFF_X1 \OUT2_reg[28]  ( .D(n2784), .CK(Clk), .Q(OUT2[28]), .QN(net644415) );
  DFF_X1 \REGISTERS_reg[31][27]  ( .D(n2783), .CK(Clk), .Q(n399), .QN(n4513)
         );
  DFF_X1 \OUT2_reg[27]  ( .D(n2782), .CK(Clk), .Q(OUT2[27]), .QN(net644414) );
  DFF_X1 \REGISTERS_reg[31][26]  ( .D(n2781), .CK(Clk), .Q(n402), .QN(n4509)
         );
  DFF_X1 \OUT2_reg[26]  ( .D(n2780), .CK(Clk), .Q(OUT2[26]), .QN(net644413) );
  DFF_X1 \REGISTERS_reg[31][25]  ( .D(n2779), .CK(Clk), .Q(n405), .QN(n4508)
         );
  DFF_X1 \OUT2_reg[25]  ( .D(n2778), .CK(Clk), .Q(OUT2[25]), .QN(net644412) );
  DFF_X1 \REGISTERS_reg[31][24]  ( .D(n2777), .CK(Clk), .Q(n408), .QN(n4503)
         );
  DFF_X1 \OUT2_reg[24]  ( .D(n2776), .CK(Clk), .Q(OUT2[24]), .QN(net644411) );
  DFF_X1 \REGISTERS_reg[31][23]  ( .D(n2775), .CK(Clk), .Q(n411), .QN(n4502)
         );
  DFF_X1 \OUT2_reg[23]  ( .D(n2774), .CK(Clk), .Q(OUT2[23]), .QN(net644410) );
  DFF_X1 \REGISTERS_reg[31][22]  ( .D(n2773), .CK(Clk), .Q(n414), .QN(n4493)
         );
  DFF_X1 \OUT2_reg[22]  ( .D(n2772), .CK(Clk), .Q(OUT2[22]), .QN(net644409) );
  DFF_X1 \REGISTERS_reg[31][21]  ( .D(n2771), .CK(Clk), .Q(n417), .QN(n4485)
         );
  DFF_X1 \OUT2_reg[21]  ( .D(n2770), .CK(Clk), .Q(OUT2[21]), .QN(net644408) );
  DFF_X1 \REGISTERS_reg[31][20]  ( .D(n2769), .CK(Clk), .Q(n420), .QN(n4484)
         );
  DFF_X1 \OUT2_reg[20]  ( .D(n2768), .CK(Clk), .Q(OUT2[20]), .QN(net644407) );
  DFF_X1 \REGISTERS_reg[31][19]  ( .D(n2767), .CK(Clk), .Q(n423), .QN(n4483)
         );
  DFF_X1 \OUT2_reg[19]  ( .D(n2766), .CK(Clk), .Q(OUT2[19]), .QN(net644406) );
  DFF_X1 \REGISTERS_reg[31][18]  ( .D(n2765), .CK(Clk), .Q(n426), .QN(n4479)
         );
  DFF_X1 \OUT2_reg[18]  ( .D(n2764), .CK(Clk), .Q(OUT2[18]), .QN(net644405) );
  DFF_X1 \REGISTERS_reg[31][17]  ( .D(n2763), .CK(Clk), .Q(n429), .QN(n4478)
         );
  DFF_X1 \OUT2_reg[17]  ( .D(n2762), .CK(Clk), .Q(OUT2[17]), .QN(net644404) );
  DFF_X1 \REGISTERS_reg[31][16]  ( .D(n2761), .CK(Clk), .Q(n432), .QN(n4473)
         );
  DFF_X1 \OUT2_reg[16]  ( .D(n2760), .CK(Clk), .Q(OUT2[16]), .QN(net644403) );
  DFF_X1 \REGISTERS_reg[31][15]  ( .D(n2759), .CK(Clk), .Q(n435), .QN(n4472)
         );
  DFF_X1 \OUT2_reg[15]  ( .D(n2758), .CK(Clk), .Q(OUT2[15]), .QN(net644402) );
  DFF_X1 \REGISTERS_reg[31][14]  ( .D(n2757), .CK(Clk), .Q(n438), .QN(n4463)
         );
  DFF_X1 \OUT2_reg[14]  ( .D(n2756), .CK(Clk), .Q(OUT2[14]), .QN(net644401) );
  DFF_X1 \REGISTERS_reg[31][13]  ( .D(n2755), .CK(Clk), .Q(n441), .QN(n4455)
         );
  DFF_X1 \OUT2_reg[13]  ( .D(n2754), .CK(Clk), .Q(OUT2[13]), .QN(net644400) );
  DFF_X1 \REGISTERS_reg[31][12]  ( .D(n2753), .CK(Clk), .Q(n444), .QN(n4454)
         );
  DFF_X1 \OUT2_reg[12]  ( .D(n2752), .CK(Clk), .Q(OUT2[12]), .QN(net644399) );
  DFF_X1 \REGISTERS_reg[31][11]  ( .D(n2751), .CK(Clk), .Q(n447), .QN(n4453)
         );
  DFF_X1 \OUT2_reg[11]  ( .D(n2750), .CK(Clk), .Q(OUT2[11]), .QN(net644398) );
  DFF_X1 \REGISTERS_reg[31][10]  ( .D(n2749), .CK(Clk), .Q(n450), .QN(n4449)
         );
  DFF_X1 \OUT2_reg[10]  ( .D(n2748), .CK(Clk), .Q(OUT2[10]), .QN(net644397) );
  DFF_X1 \REGISTERS_reg[31][9]  ( .D(n2747), .CK(Clk), .Q(n453), .QN(n4448) );
  DFF_X1 \OUT2_reg[9]  ( .D(n2746), .CK(Clk), .Q(OUT2[9]), .QN(net644396) );
  DFF_X1 \REGISTERS_reg[31][8]  ( .D(n2745), .CK(Clk), .Q(n456), .QN(n4443) );
  DFF_X1 \OUT2_reg[8]  ( .D(n2744), .CK(Clk), .Q(OUT2[8]), .QN(net644395) );
  DFF_X1 \REGISTERS_reg[31][7]  ( .D(n2743), .CK(Clk), .Q(n459), .QN(n4442) );
  DFF_X1 \OUT2_reg[7]  ( .D(n2742), .CK(Clk), .Q(OUT2[7]), .QN(net644394) );
  DFF_X1 \REGISTERS_reg[31][6]  ( .D(n2741), .CK(Clk), .Q(n462), .QN(n4433) );
  DFF_X1 \OUT2_reg[6]  ( .D(n2740), .CK(Clk), .Q(OUT2[6]), .QN(net644393) );
  DFF_X1 \REGISTERS_reg[31][5]  ( .D(n2739), .CK(Clk), .Q(n465), .QN(n4425) );
  DFF_X1 \OUT2_reg[5]  ( .D(n2738), .CK(Clk), .Q(OUT2[5]), .QN(net644392) );
  DFF_X1 \REGISTERS_reg[31][4]  ( .D(n2737), .CK(Clk), .Q(n468), .QN(n4424) );
  DFF_X1 \OUT2_reg[4]  ( .D(n2736), .CK(Clk), .Q(OUT2[4]), .QN(net644391) );
  DFF_X1 \REGISTERS_reg[31][3]  ( .D(n2735), .CK(Clk), .Q(n471), .QN(n4423) );
  DFF_X1 \OUT2_reg[3]  ( .D(n2734), .CK(Clk), .Q(OUT2[3]), .QN(net644390) );
  DFF_X1 \REGISTERS_reg[31][2]  ( .D(n2733), .CK(Clk), .Q(n474), .QN(n4419) );
  DFF_X1 \OUT2_reg[2]  ( .D(n2732), .CK(Clk), .Q(OUT2[2]), .QN(net644389) );
  DFF_X1 \REGISTERS_reg[31][1]  ( .D(n2731), .CK(Clk), .Q(n477), .QN(n4418) );
  DFF_X1 \OUT2_reg[1]  ( .D(n2730), .CK(Clk), .Q(OUT2[1]), .QN(net644388) );
  DFF_X1 \REGISTERS_reg[31][0]  ( .D(n2729), .CK(Clk), .Q(n4060), .QN(n2087)
         );
  DFF_X1 \OUT2_reg[0]  ( .D(n2728), .CK(Clk), .Q(OUT2[0]), .QN(n2184) );
  DFF_X1 \OUT1_reg[31]  ( .D(n2727), .CK(Clk), .Q(OUT1[31]), .QN(net644387) );
  DFF_X1 \OUT1_reg[30]  ( .D(n2726), .CK(Clk), .Q(OUT1[30]), .QN(net644386) );
  DFF_X1 \OUT1_reg[29]  ( .D(n2725), .CK(Clk), .Q(OUT1[29]), .QN(net644385) );
  DFF_X1 \OUT1_reg[28]  ( .D(n2724), .CK(Clk), .Q(OUT1[28]), .QN(net644384) );
  DFF_X1 \OUT1_reg[27]  ( .D(n2723), .CK(Clk), .Q(OUT1[27]), .QN(net644383) );
  DFF_X1 \OUT1_reg[26]  ( .D(n2722), .CK(Clk), .Q(OUT1[26]), .QN(net644382) );
  DFF_X1 \OUT1_reg[25]  ( .D(n2721), .CK(Clk), .Q(OUT1[25]), .QN(net644381) );
  DFF_X1 \OUT1_reg[24]  ( .D(n2720), .CK(Clk), .Q(OUT1[24]), .QN(net644380) );
  DFF_X1 \OUT1_reg[23]  ( .D(n2719), .CK(Clk), .Q(OUT1[23]), .QN(net644379) );
  DFF_X1 \OUT1_reg[22]  ( .D(n2718), .CK(Clk), .Q(OUT1[22]), .QN(net644378) );
  DFF_X1 \OUT1_reg[21]  ( .D(n2717), .CK(Clk), .Q(OUT1[21]), .QN(net644377) );
  DFF_X1 \OUT1_reg[20]  ( .D(n2716), .CK(Clk), .Q(OUT1[20]), .QN(net644376) );
  DFF_X1 \OUT1_reg[19]  ( .D(n2715), .CK(Clk), .Q(OUT1[19]), .QN(net644375) );
  DFF_X1 \OUT1_reg[18]  ( .D(n2714), .CK(Clk), .Q(OUT1[18]), .QN(net644374) );
  DFF_X1 \OUT1_reg[17]  ( .D(n2713), .CK(Clk), .Q(OUT1[17]), .QN(net644373) );
  DFF_X1 \OUT1_reg[16]  ( .D(n2712), .CK(Clk), .Q(OUT1[16]), .QN(net644372) );
  DFF_X1 \OUT1_reg[15]  ( .D(n2711), .CK(Clk), .Q(OUT1[15]), .QN(net644371) );
  DFF_X1 \OUT1_reg[14]  ( .D(n2710), .CK(Clk), .Q(OUT1[14]), .QN(net644370) );
  DFF_X1 \OUT1_reg[13]  ( .D(n2709), .CK(Clk), .Q(OUT1[13]), .QN(net644369) );
  DFF_X1 \OUT1_reg[12]  ( .D(n2708), .CK(Clk), .Q(OUT1[12]), .QN(net644368) );
  DFF_X1 \OUT1_reg[11]  ( .D(n2707), .CK(Clk), .Q(OUT1[11]), .QN(net644367) );
  DFF_X1 \OUT1_reg[10]  ( .D(n2706), .CK(Clk), .Q(OUT1[10]), .QN(net644366) );
  DFF_X1 \OUT1_reg[9]  ( .D(n2705), .CK(Clk), .Q(OUT1[9]), .QN(net644365) );
  DFF_X1 \OUT1_reg[8]  ( .D(n2704), .CK(Clk), .Q(OUT1[8]), .QN(net644364) );
  DFF_X1 \OUT1_reg[7]  ( .D(n2703), .CK(Clk), .Q(OUT1[7]), .QN(net644363) );
  DFF_X1 \OUT1_reg[6]  ( .D(n2702), .CK(Clk), .Q(OUT1[6]), .QN(net644362) );
  DFF_X1 \OUT1_reg[5]  ( .D(n2701), .CK(Clk), .Q(OUT1[5]), .QN(net644361) );
  DFF_X1 \OUT1_reg[4]  ( .D(n2700), .CK(Clk), .Q(OUT1[4]), .QN(net644360) );
  DFF_X1 \OUT1_reg[3]  ( .D(n2699), .CK(Clk), .Q(OUT1[3]), .QN(net644359) );
  DFF_X1 \OUT1_reg[2]  ( .D(n2698), .CK(Clk), .Q(OUT1[2]), .QN(net644358) );
  DFF_X1 \OUT1_reg[1]  ( .D(n2697), .CK(Clk), .Q(OUT1[1]), .QN(net644357) );
  DFF_X1 \OUT1_reg[0]  ( .D(n2696), .CK(Clk), .Q(OUT1[0]), .QN(n2152) );
  NAND3_X1 U3574 ( .A1(ADD_RD2[4]), .A2(ADD_RD2[3]), .A3(n5189), .ZN(n5170) );
  NAND3_X1 U3575 ( .A1(ADD_RD2[3]), .A2(n5189), .A3(n5190), .ZN(n5158) );
  NAND3_X1 U3576 ( .A1(n5194), .A2(ADD_RD2[4]), .A3(ADD_RD2[0]), .ZN(n5155) );
  NAND3_X1 U3577 ( .A1(ADD_RD2[0]), .A2(ADD_RD2[4]), .A3(ADD_RD2[3]), .ZN(
        n5181) );
  NAND3_X1 U3578 ( .A1(ADD_RD2[4]), .A2(n5189), .A3(n5194), .ZN(n5179) );
  NAND3_X1 U3579 ( .A1(ADD_RD2[0]), .A2(n5190), .A3(n5194), .ZN(n5157) );
  NAND3_X1 U3580 ( .A1(n5189), .A2(n5190), .A3(n5194), .ZN(n5169) );
  NAND3_X1 U3581 ( .A1(ADD_RD2[0]), .A2(ADD_RD2[3]), .A3(n5190), .ZN(n5173) );
  NAND3_X1 U3582 ( .A1(ADD_RD1[3]), .A2(ADD_RD1[4]), .A3(n5966), .ZN(n5950) );
  NAND3_X1 U3583 ( .A1(ADD_RD1[3]), .A2(n5967), .A3(n5966), .ZN(n5938) );
  NAND3_X1 U3584 ( .A1(n5971), .A2(ADD_RD1[4]), .A3(ADD_RD1[0]), .ZN(n5935) );
  NAND3_X1 U3585 ( .A1(ADD_RD1[4]), .A2(ADD_RD1[3]), .A3(ADD_RD1[0]), .ZN(
        n5959) );
  NAND3_X1 U3586 ( .A1(ADD_RD1[4]), .A2(n5971), .A3(n5966), .ZN(n5958) );
  NAND3_X1 U3587 ( .A1(ADD_RD1[0]), .A2(n5967), .A3(n5971), .ZN(n5937) );
  NAND3_X1 U3588 ( .A1(n5967), .A2(n5971), .A3(n5966), .ZN(n5949) );
  NAND3_X1 U3589 ( .A1(ADD_RD1[3]), .A2(ADD_RD1[0]), .A3(n5967), .ZN(n5953) );
  NOR3_X1 U3557 ( .A1(n5979), .A2(n5973), .A3(n5978), .ZN(n5980) );
  NAND2_X1 U3553 ( .A1(n5984), .A2(n1769), .ZN(n5983) );
  AOI22_X1 U3549 ( .A1(n1919), .A2(ADD_RD1[2]), .B1(n5146), .B2(ADD_RD1[4]), 
        .ZN(n5982) );
  OAI221_X1 U3548 ( .B1(n1919), .B2(ADD_RD1[2]), .C1(n5146), .C2(ADD_RD1[4]), 
        .A(n5982), .ZN(n5981) );
  AOI22_X1 U3534 ( .A1(n6355), .A2(n3915), .B1(n6357), .B2(n4059), .ZN(n5927)
         );
  AOI22_X1 U3531 ( .A1(net644901), .A2(n6356), .B1(net644869), .B2(n6358), 
        .ZN(n5928) );
  NOR2_X1 U3530 ( .A1(n5958), .A2(n5939), .ZN(n5925) );
  NOR2_X1 U3525 ( .A1(n5978), .A2(n5979), .ZN(n5976) );
  NAND2_X1 U3524 ( .A1(n5976), .A2(n5977), .ZN(n5975) );
  NOR4_X1 U3523 ( .A1(N4487), .A2(n5973), .A3(n5974), .A4(n5975), .ZN(n5260)
         );
  AOI22_X1 U3522 ( .A1(net644451), .A2(n6360), .B1(DATAIN[0]), .B2(n6359), 
        .ZN(n5972) );
  OAI21_X1 U3521 ( .B1(n5257), .B2(n2152), .A(n5972), .ZN(n5968) );
  OAI22_X1 U3517 ( .A1(n671), .A2(n5255), .B1(n514), .B2(n3952), .ZN(n5969) );
  AOI211_X1 U3516 ( .C1(net644675), .C2(n5925), .A(n5968), .B(n5969), .ZN(
        n5929) );
  NAND2_X1 U3512 ( .A1(n5963), .A2(n5964), .ZN(n5952) );
  AOI22_X1 U3509 ( .A1(net644515), .A2(n6363), .B1(net644547), .B2(n6362), 
        .ZN(n5940) );
  AOI22_X1 U3505 ( .A1(n6364), .A2(n385), .B1(n5248), .B2(n4060), .ZN(n5954)
         );
  AOI22_X1 U3502 ( .A1(net644612), .A2(n3911), .B1(net644483), .B2(n3912), 
        .ZN(n5955) );
  AOI22_X1 U3498 ( .A1(n6366), .A2(n386), .B1(n5244), .B2(n4061), .ZN(n5956)
         );
  AOI22_X1 U3495 ( .A1(net644580), .A2(n3913), .B1(net644676), .B2(n3914), 
        .ZN(n5957) );
  NAND4_X1 U3494 ( .A1(n5954), .A2(n5955), .A3(n5956), .A4(n5957), .ZN(n5942)
         );
  AOI22_X1 U3490 ( .A1(n6368), .A2(n384), .B1(n5236), .B2(n4062), .ZN(n5944)
         );
  AOI22_X1 U3487 ( .A1(net644772), .A2(n3910), .B1(net644740), .B2(n3909), 
        .ZN(n5945) );
  AOI22_X1 U3484 ( .A1(net644902), .A2(n3908), .B1(net644419), .B2(n3907), 
        .ZN(n5946) );
  AOI22_X1 U3481 ( .A1(net644867), .A2(n3906), .B1(net644868), .B2(n3905), 
        .ZN(n5947) );
  NAND4_X1 U3480 ( .A1(n5944), .A2(n5945), .A3(n5946), .A4(n5947), .ZN(n5943)
         );
  OAI21_X1 U3479 ( .B1(n5942), .B2(n5943), .A(n6370), .ZN(n5941) );
  OAI211_X1 U3478 ( .C1(n703), .C2(n5220), .A(n5940), .B(n5941), .ZN(n5931) );
  NOR2_X1 U3475 ( .A1(n5937), .A2(n5936), .ZN(n5910) );
  AOI22_X1 U3473 ( .A1(net644835), .A2(n5910), .B1(net644579), .B2(n5219), 
        .ZN(n5934) );
  OAI21_X1 U3472 ( .B1(n481), .B2(n3953), .A(n5934), .ZN(n5932) );
  AOI211_X1 U3471 ( .C1(n6374), .C2(net644708), .A(n5931), .B(n5932), .ZN(
        n5930) );
  NAND4_X1 U3470 ( .A1(n5927), .A2(n5928), .A3(n5929), .A4(n5930), .ZN(n2696)
         );
  AOI22_X1 U2534 ( .A1(ADD_WR[2]), .A2(ADD_RD2[2]), .B1(n5186), .B2(n1919), 
        .ZN(n5196) );
  NOR3_X1 U2531 ( .A1(n5202), .A2(n5196), .A3(n5201), .ZN(n5205) );
  AOI22_X1 U2530 ( .A1(n5146), .A2(ADD_RD2[4]), .B1(ADD_RD2[3]), .B2(n1846), 
        .ZN(n5208) );
  OAI221_X1 U2529 ( .B1(n5146), .B2(ADD_RD2[4]), .C1(n1846), .C2(ADD_RD2[3]), 
        .A(n5208), .ZN(n5207) );
  NOR2_X1 U2528 ( .A1(n5206), .A2(n5207), .ZN(n5200) );
  AOI22_X1 U2517 ( .A1(n4241), .A2(n3915), .B1(n6377), .B2(n4059), .ZN(n5147)
         );
  AOI22_X1 U2514 ( .A1(net644901), .A2(n6375), .B1(net644869), .B2(n6378), 
        .ZN(n5148) );
  NOR2_X1 U2513 ( .A1(n5179), .A2(n5159), .ZN(n5142) );
  NOR2_X1 U2508 ( .A1(n5201), .A2(n5202), .ZN(n5199) );
  NAND2_X1 U2507 ( .A1(n5199), .A2(n5200), .ZN(n5198) );
  NOR4_X1 U2506 ( .A1(N4487), .A2(n5196), .A3(n5197), .A4(n5198), .ZN(n4238)
         );
  AOI22_X1 U2505 ( .A1(net644451), .A2(n4237), .B1(DATAIN[0]), .B2(n6379), 
        .ZN(n5195) );
  OAI21_X1 U2504 ( .B1(n4235), .B2(n2184), .A(n5195), .ZN(n5191) );
  OAI22_X1 U2500 ( .A1(n671), .A2(n4234), .B1(n514), .B2(n3950), .ZN(n5192) );
  AOI211_X1 U2499 ( .C1(net644675), .C2(n5142), .A(n5191), .B(n5192), .ZN(
        n5149) );
  NAND2_X1 U2495 ( .A1(n5186), .A2(n5187), .ZN(n5172) );
  AOI22_X1 U2492 ( .A1(net644515), .A2(n3880), .B1(net644547), .B2(n4228), 
        .ZN(n5160) );
  AOI22_X1 U2489 ( .A1(n3896), .A2(n385), .B1(n4225), .B2(n4060), .ZN(n5175)
         );
  AOI22_X1 U2486 ( .A1(net644612), .A2(n4223), .B1(net644483), .B2(n3894), 
        .ZN(n5176) );
  AOI22_X1 U2483 ( .A1(n6384), .A2(n386), .B1(n3891), .B2(n4061), .ZN(n5177)
         );
  AOI22_X1 U2480 ( .A1(net644580), .A2(n3890), .B1(net644676), .B2(n4219), 
        .ZN(n5178) );
  NAND4_X1 U2479 ( .A1(n5175), .A2(n5176), .A3(n5177), .A4(n5178), .ZN(n5162)
         );
  AOI22_X1 U2476 ( .A1(n3903), .A2(n384), .B1(n3904), .B2(n4062), .ZN(n5164)
         );
  AOI22_X1 U2473 ( .A1(net644772), .A2(n4209), .B1(net644740), .B2(n3901), 
        .ZN(n5165) );
  AOI22_X1 U2470 ( .A1(net644902), .A2(n4207), .B1(net644419), .B2(n3899), 
        .ZN(n5166) );
  NOR2_X1 U2468 ( .A1(n5168), .A2(n5169), .ZN(n4204) );
  AOI22_X1 U2467 ( .A1(net644867), .A2(n3898), .B1(net644868), .B2(n6385), 
        .ZN(n5167) );
  NAND4_X1 U2466 ( .A1(n5164), .A2(n5165), .A3(n5166), .A4(n5167), .ZN(n5163)
         );
  OAI21_X1 U2465 ( .B1(n5162), .B2(n5163), .A(n6386), .ZN(n5161) );
  OAI211_X1 U2464 ( .C1(n703), .C2(n4194), .A(n5160), .B(n5161), .ZN(n5151) );
  NOR2_X1 U2461 ( .A1(n5157), .A2(n5156), .ZN(n5124) );
  AOI22_X1 U2459 ( .A1(net644835), .A2(n5124), .B1(net644579), .B2(n6388), 
        .ZN(n5154) );
  OAI21_X1 U2458 ( .B1(n481), .B2(n3951), .A(n5154), .ZN(n5152) );
  AOI211_X1 U2457 ( .C1(net644708), .C2(n4186), .A(n5151), .B(n5152), .ZN(
        n5150) );
  NAND4_X1 U2456 ( .A1(n5147), .A2(n5148), .A3(n5149), .A4(n5150), .ZN(n2728)
         );
  AOI22_X1 U2596 ( .A1(n5263), .A2(n3948), .B1(n5264), .B2(n4053), .ZN(n5265)
         );
  AOI22_X1 U2595 ( .A1(n5261), .A2(net644899), .B1(n5262), .B2(net644865), 
        .ZN(n5266) );
  AOI22_X1 U2594 ( .A1(n6360), .A2(net644481), .B1(n6359), .B2(DATAIN[30]), 
        .ZN(n5286) );
  OAI21_X1 U2593 ( .B1(n5257), .B2(net644386), .A(n5286), .ZN(n5284) );
  OAI22_X1 U2592 ( .A1(n516), .A2(n5255), .B1(n641), .B2(n5256), .ZN(n5285) );
  AOI211_X1 U2591 ( .C1(n6361), .C2(net644673), .A(n5284), .B(n5285), .ZN(
        n5267) );
  AOI22_X1 U2590 ( .A1(n6363), .A2(net644545), .B1(n6362), .B2(net644577), 
        .ZN(n5272) );
  AOI22_X1 U2588 ( .A1(n5248), .A2(n390), .B1(n5249), .B2(n4161), .ZN(n5280)
         );
  AOI22_X1 U2587 ( .A1(n3911), .A2(net644642), .B1(n3912), .B2(net644513), 
        .ZN(n5281) );
  AOI22_X1 U2585 ( .A1(n5244), .A2(n4054), .B1(n5245), .B2(n354), .ZN(n5282)
         );
  AOI22_X1 U2584 ( .A1(n3913), .A2(net644610), .B1(n3914), .B2(net644706), 
        .ZN(n5283) );
  NAND4_X1 U2583 ( .A1(n5280), .A2(n5281), .A3(n5282), .A4(n5283), .ZN(n5274)
         );
  AOI22_X1 U2581 ( .A1(n5236), .A2(n392), .B1(n5237), .B2(n4162), .ZN(n5276)
         );
  AOI22_X1 U2580 ( .A1(n3910), .A2(net644802), .B1(n3909), .B2(net644770), 
        .ZN(n5277) );
  AOI22_X1 U2579 ( .A1(n3908), .A2(net644932), .B1(n3907), .B2(net644449), 
        .ZN(n5278) );
  AOI22_X1 U2577 ( .A1(n3906), .A2(n4055), .B1(n3905), .B2(n391), .ZN(n5279)
         );
  NAND4_X1 U2576 ( .A1(n5276), .A2(n5277), .A3(n5278), .A4(n5279), .ZN(n5275)
         );
  OAI21_X1 U2575 ( .B1(n5274), .B2(n5275), .A(n6370), .ZN(n5273) );
  OAI211_X1 U2574 ( .C1(n547), .C2(n5220), .A(n5272), .B(n5273), .ZN(n5269) );
  AOI22_X1 U2572 ( .A1(n6373), .A2(net644833), .B1(n6372), .B2(n4163), .ZN(
        n5271) );
  OAI21_X1 U2571 ( .B1(n609), .B2(n5216), .A(n5271), .ZN(n5270) );
  AOI211_X1 U2570 ( .C1(n5213), .C2(net644738), .A(n5269), .B(n5270), .ZN(
        n5268) );
  NAND4_X1 U2569 ( .A1(n5265), .A2(n5266), .A3(n5267), .A4(n5268), .ZN(n2726)
         );
  AOI22_X1 U2626 ( .A1(n5263), .A2(n3947), .B1(n5264), .B2(n4050), .ZN(n5287)
         );
  AOI22_X1 U2625 ( .A1(n5261), .A2(net644898), .B1(n5262), .B2(net644864), 
        .ZN(n5288) );
  AOI22_X1 U2624 ( .A1(n5259), .A2(net644480), .B1(n5260), .B2(DATAIN[29]), 
        .ZN(n5308) );
  OAI21_X1 U2623 ( .B1(n5257), .B2(net644385), .A(n5308), .ZN(n5306) );
  OAI22_X1 U2622 ( .A1(n517), .A2(n5255), .B1(n642), .B2(n5256), .ZN(n5307) );
  AOI211_X1 U2621 ( .C1(n6361), .C2(net644672), .A(n5306), .B(n5307), .ZN(
        n5289) );
  AOI22_X1 U2620 ( .A1(n5250), .A2(net644544), .B1(n5251), .B2(net644576), 
        .ZN(n5294) );
  AOI22_X1 U2618 ( .A1(n5248), .A2(n393), .B1(n5249), .B2(n4158), .ZN(n5302)
         );
  AOI22_X1 U2617 ( .A1(n3911), .A2(net644641), .B1(n3912), .B2(net644512), 
        .ZN(n5303) );
  AOI22_X1 U2615 ( .A1(n5244), .A2(n4051), .B1(n5245), .B2(n355), .ZN(n5304)
         );
  AOI22_X1 U2614 ( .A1(n3913), .A2(net644609), .B1(n3914), .B2(net644705), 
        .ZN(n5305) );
  NAND4_X1 U2613 ( .A1(n5302), .A2(n5303), .A3(n5304), .A4(n5305), .ZN(n5296)
         );
  AOI22_X1 U2611 ( .A1(n5236), .A2(n395), .B1(n5237), .B2(n4159), .ZN(n5298)
         );
  AOI22_X1 U2610 ( .A1(n3910), .A2(net644801), .B1(n3909), .B2(net644769), 
        .ZN(n5299) );
  AOI22_X1 U2609 ( .A1(n3908), .A2(net644931), .B1(n3907), .B2(net644448), 
        .ZN(n5300) );
  AOI22_X1 U2607 ( .A1(n3906), .A2(n4052), .B1(n3905), .B2(n394), .ZN(n5301)
         );
  NAND4_X1 U2606 ( .A1(n5298), .A2(n5299), .A3(n5300), .A4(n5301), .ZN(n5297)
         );
  OAI21_X1 U2605 ( .B1(n5296), .B2(n5297), .A(n6370), .ZN(n5295) );
  OAI211_X1 U2604 ( .C1(n548), .C2(n5220), .A(n5294), .B(n5295), .ZN(n5291) );
  AOI22_X1 U2602 ( .A1(n6373), .A2(net644832), .B1(n6372), .B2(n4160), .ZN(
        n5293) );
  OAI21_X1 U2601 ( .B1(n610), .B2(n5216), .A(n5293), .ZN(n5292) );
  AOI211_X1 U2600 ( .C1(n5213), .C2(net644737), .A(n5291), .B(n5292), .ZN(
        n5290) );
  NAND4_X1 U2599 ( .A1(n5287), .A2(n5288), .A3(n5289), .A4(n5290), .ZN(n2725)
         );
  AOI22_X1 U2656 ( .A1(n5263), .A2(n3946), .B1(n5264), .B2(n4047), .ZN(n5309)
         );
  AOI22_X1 U2655 ( .A1(n5261), .A2(net644897), .B1(n5262), .B2(net644863), 
        .ZN(n5310) );
  AOI22_X1 U2654 ( .A1(n6360), .A2(net644479), .B1(n5260), .B2(DATAIN[28]), 
        .ZN(n5330) );
  OAI21_X1 U2653 ( .B1(n5257), .B2(net644384), .A(n5330), .ZN(n5328) );
  OAI22_X1 U2652 ( .A1(n518), .A2(n5255), .B1(n643), .B2(n5256), .ZN(n5329) );
  AOI211_X1 U2651 ( .C1(n6361), .C2(net644671), .A(n5328), .B(n5329), .ZN(
        n5311) );
  AOI22_X1 U2650 ( .A1(n6363), .A2(net644543), .B1(n5251), .B2(net644575), 
        .ZN(n5316) );
  AOI22_X1 U2648 ( .A1(n5248), .A2(n396), .B1(n5249), .B2(n4155), .ZN(n5324)
         );
  AOI22_X1 U2647 ( .A1(n3911), .A2(net644640), .B1(n3912), .B2(net644511), 
        .ZN(n5325) );
  AOI22_X1 U2645 ( .A1(n5244), .A2(n4048), .B1(n5245), .B2(n356), .ZN(n5326)
         );
  AOI22_X1 U2644 ( .A1(n3913), .A2(net644608), .B1(n3914), .B2(net644704), 
        .ZN(n5327) );
  NAND4_X1 U2643 ( .A1(n5324), .A2(n5325), .A3(n5326), .A4(n5327), .ZN(n5318)
         );
  AOI22_X1 U2641 ( .A1(n5236), .A2(n398), .B1(n5237), .B2(n4156), .ZN(n5320)
         );
  AOI22_X1 U2640 ( .A1(n3910), .A2(net644800), .B1(n3909), .B2(net644768), 
        .ZN(n5321) );
  AOI22_X1 U2639 ( .A1(n3908), .A2(net644930), .B1(n3907), .B2(net644447), 
        .ZN(n5322) );
  AOI22_X1 U2637 ( .A1(n3906), .A2(n4049), .B1(n3905), .B2(n397), .ZN(n5323)
         );
  NAND4_X1 U2636 ( .A1(n5320), .A2(n5321), .A3(n5322), .A4(n5323), .ZN(n5319)
         );
  OAI21_X1 U2635 ( .B1(n5318), .B2(n5319), .A(n6370), .ZN(n5317) );
  OAI211_X1 U2634 ( .C1(n549), .C2(n5220), .A(n5316), .B(n5317), .ZN(n5313) );
  AOI22_X1 U2632 ( .A1(n6373), .A2(net644831), .B1(n6372), .B2(n4157), .ZN(
        n5315) );
  OAI21_X1 U2631 ( .B1(n611), .B2(n5216), .A(n5315), .ZN(n5314) );
  AOI211_X1 U2630 ( .C1(n5213), .C2(net644736), .A(n5313), .B(n5314), .ZN(
        n5312) );
  NAND4_X1 U2629 ( .A1(n5309), .A2(n5310), .A3(n5311), .A4(n5312), .ZN(n2724)
         );
  AOI22_X1 U2566 ( .A1(n5263), .A2(n3949), .B1(n5264), .B2(n4056), .ZN(n5209)
         );
  AOI22_X1 U2565 ( .A1(n6358), .A2(net644900), .B1(n5262), .B2(net644866), 
        .ZN(n5210) );
  AOI22_X1 U2564 ( .A1(n5259), .A2(net644482), .B1(n6359), .B2(DATAIN[31]), 
        .ZN(n5258) );
  OAI21_X1 U2563 ( .B1(n5257), .B2(net644387), .A(n5258), .ZN(n5253) );
  OAI22_X1 U2562 ( .A1(n515), .A2(n5255), .B1(n640), .B2(n5256), .ZN(n5254) );
  AOI211_X1 U2561 ( .C1(n6361), .C2(net644674), .A(n5253), .B(n5254), .ZN(
        n5211) );
  AOI22_X1 U2560 ( .A1(n5250), .A2(net644546), .B1(n6362), .B2(net644578), 
        .ZN(n5221) );
  AOI22_X1 U2558 ( .A1(n6365), .A2(n387), .B1(n5249), .B2(n4164), .ZN(n5238)
         );
  AOI22_X1 U2557 ( .A1(n3911), .A2(net644643), .B1(n3912), .B2(net644514), 
        .ZN(n5239) );
  AOI22_X1 U2555 ( .A1(n6367), .A2(n4057), .B1(n5245), .B2(n353), .ZN(n5240)
         );
  AOI22_X1 U2554 ( .A1(n3913), .A2(net644611), .B1(n3914), .B2(net644707), 
        .ZN(n5241) );
  NAND4_X1 U2553 ( .A1(n5238), .A2(n5239), .A3(n5240), .A4(n5241), .ZN(n5223)
         );
  AOI22_X1 U2551 ( .A1(n6369), .A2(n389), .B1(n5237), .B2(n4165), .ZN(n5226)
         );
  AOI22_X1 U2550 ( .A1(n3910), .A2(net644803), .B1(n3909), .B2(net644771), 
        .ZN(n5227) );
  AOI22_X1 U2549 ( .A1(n3908), .A2(net644933), .B1(n3907), .B2(net644450), 
        .ZN(n5228) );
  AOI22_X1 U2547 ( .A1(n3906), .A2(n4058), .B1(n3905), .B2(n388), .ZN(n5229)
         );
  NAND4_X1 U2546 ( .A1(n5226), .A2(n5227), .A3(n5228), .A4(n5229), .ZN(n5224)
         );
  OAI21_X1 U2545 ( .B1(n5223), .B2(n5224), .A(n6370), .ZN(n5222) );
  OAI211_X1 U2544 ( .C1(n546), .C2(n5220), .A(n5221), .B(n5222), .ZN(n5214) );
  AOI22_X1 U2542 ( .A1(n6373), .A2(net644834), .B1(n6372), .B2(n4166), .ZN(
        n5217) );
  OAI21_X1 U2541 ( .B1(n608), .B2(n5216), .A(n5217), .ZN(n5215) );
  AOI211_X1 U2540 ( .C1(n5213), .C2(net644739), .A(n5214), .B(n5215), .ZN(
        n5212) );
  NAND4_X1 U2539 ( .A1(n5209), .A2(n5210), .A3(n5211), .A4(n5212), .ZN(n2727)
         );
  AOI22_X1 U2746 ( .A1(n6356), .A2(n3943), .B1(n5264), .B2(n4038), .ZN(n5375)
         );
  AOI22_X1 U2745 ( .A1(n6358), .A2(net644894), .B1(n5262), .B2(net644860), 
        .ZN(n5376) );
  AOI22_X1 U2744 ( .A1(n6360), .A2(net644476), .B1(n6359), .B2(DATAIN[25]), 
        .ZN(n5396) );
  OAI21_X1 U2743 ( .B1(n5257), .B2(net644381), .A(n5396), .ZN(n5394) );
  OAI22_X1 U2742 ( .A1(n521), .A2(n5255), .B1(n646), .B2(n5256), .ZN(n5395) );
  AOI211_X1 U2741 ( .C1(n6361), .C2(net644668), .A(n5394), .B(n5395), .ZN(
        n5377) );
  AOI22_X1 U2740 ( .A1(n6363), .A2(net644540), .B1(n6362), .B2(net644572), 
        .ZN(n5382) );
  AOI22_X1 U2738 ( .A1(n6365), .A2(n405), .B1(n5249), .B2(n4144), .ZN(n5390)
         );
  AOI22_X1 U2737 ( .A1(n3911), .A2(net644637), .B1(n3912), .B2(net644508), 
        .ZN(n5391) );
  AOI22_X1 U2735 ( .A1(n5244), .A2(n4039), .B1(n5245), .B2(n359), .ZN(n5392)
         );
  AOI22_X1 U2734 ( .A1(n3913), .A2(net644605), .B1(n3914), .B2(net644701), 
        .ZN(n5393) );
  NAND4_X1 U2733 ( .A1(n5390), .A2(n5391), .A3(n5392), .A4(n5393), .ZN(n5384)
         );
  AOI22_X1 U2731 ( .A1(n5236), .A2(n407), .B1(n5237), .B2(n4147), .ZN(n5386)
         );
  AOI22_X1 U2730 ( .A1(n3910), .A2(net644797), .B1(n3909), .B2(net644765), 
        .ZN(n5387) );
  AOI22_X1 U2729 ( .A1(n3908), .A2(net644927), .B1(n3907), .B2(net644444), 
        .ZN(n5388) );
  AOI22_X1 U2727 ( .A1(n3906), .A2(n4040), .B1(n3905), .B2(n406), .ZN(n5389)
         );
  NAND4_X1 U2726 ( .A1(n5386), .A2(n5387), .A3(n5388), .A4(n5389), .ZN(n5385)
         );
  OAI21_X1 U2725 ( .B1(n5384), .B2(n5385), .A(n6370), .ZN(n5383) );
  OAI211_X1 U2724 ( .C1(n552), .C2(n5220), .A(n5382), .B(n5383), .ZN(n5379) );
  AOI22_X1 U2722 ( .A1(n6373), .A2(net644828), .B1(n6372), .B2(n4148), .ZN(
        n5381) );
  OAI21_X1 U2721 ( .B1(n614), .B2(n5216), .A(n5381), .ZN(n5380) );
  AOI211_X1 U2720 ( .C1(n5213), .C2(net644733), .A(n5379), .B(n5380), .ZN(
        n5378) );
  NAND4_X1 U2719 ( .A1(n5375), .A2(n5376), .A3(n5377), .A4(n5378), .ZN(n2721)
         );
  AOI22_X1 U3046 ( .A1(n6356), .A2(n3933), .B1(n5264), .B2(n4005), .ZN(n5595)
         );
  AOI22_X1 U3045 ( .A1(n6358), .A2(net644884), .B1(n6357), .B2(net644850), 
        .ZN(n5596) );
  AOI22_X1 U3044 ( .A1(n6360), .A2(net644466), .B1(n6359), .B2(DATAIN[15]), 
        .ZN(n5616) );
  OAI21_X1 U3043 ( .B1(n5257), .B2(net644371), .A(n5616), .ZN(n5614) );
  OAI22_X1 U3042 ( .A1(n531), .A2(n5255), .B1(n656), .B2(n5256), .ZN(n5615) );
  AOI211_X1 U3041 ( .C1(n6361), .C2(net644658), .A(n5614), .B(n5615), .ZN(
        n5597) );
  AOI22_X1 U3040 ( .A1(n6363), .A2(net644530), .B1(n6362), .B2(net644562), 
        .ZN(n5602) );
  AOI22_X1 U3038 ( .A1(n6365), .A2(n435), .B1(n5249), .B2(n4113), .ZN(n5610)
         );
  AOI22_X1 U3037 ( .A1(n3911), .A2(net644627), .B1(n3912), .B2(net644498), 
        .ZN(n5611) );
  AOI22_X1 U3035 ( .A1(n6367), .A2(n4006), .B1(n5245), .B2(n369), .ZN(n5612)
         );
  AOI22_X1 U3034 ( .A1(n3913), .A2(net644595), .B1(n3914), .B2(net644691), 
        .ZN(n5613) );
  NAND4_X1 U3033 ( .A1(n5610), .A2(n5611), .A3(n5612), .A4(n5613), .ZN(n5604)
         );
  AOI22_X1 U3031 ( .A1(n6369), .A2(n437), .B1(n5237), .B2(n4114), .ZN(n5606)
         );
  AOI22_X1 U3030 ( .A1(n3910), .A2(net644787), .B1(n3909), .B2(net644755), 
        .ZN(n5607) );
  AOI22_X1 U3029 ( .A1(n3908), .A2(net644917), .B1(n3907), .B2(net644434), 
        .ZN(n5608) );
  AOI22_X1 U3027 ( .A1(n3906), .A2(n4007), .B1(n3905), .B2(n436), .ZN(n5609)
         );
  NAND4_X1 U3026 ( .A1(n5606), .A2(n5607), .A3(n5608), .A4(n5609), .ZN(n5605)
         );
  OAI21_X1 U3025 ( .B1(n5604), .B2(n5605), .A(n6370), .ZN(n5603) );
  OAI211_X1 U3024 ( .C1(n562), .C2(n5220), .A(n5602), .B(n5603), .ZN(n5599) );
  AOI22_X1 U3022 ( .A1(n6373), .A2(net644818), .B1(n6372), .B2(n4115), .ZN(
        n5601) );
  OAI21_X1 U3021 ( .B1(n624), .B2(n5216), .A(n5601), .ZN(n5600) );
  AOI211_X1 U3020 ( .C1(n5213), .C2(net644723), .A(n5599), .B(n5600), .ZN(
        n5598) );
  NAND4_X1 U3019 ( .A1(n5595), .A2(n5596), .A3(n5597), .A4(n5598), .ZN(n2711)
         );
  AOI22_X1 U3076 ( .A1(n6356), .A2(n3932), .B1(n5264), .B2(n4002), .ZN(n5617)
         );
  AOI22_X1 U3075 ( .A1(n6358), .A2(net644883), .B1(n6357), .B2(net644849), 
        .ZN(n5618) );
  AOI22_X1 U3074 ( .A1(n6360), .A2(net644465), .B1(n6359), .B2(DATAIN[14]), 
        .ZN(n5638) );
  OAI21_X1 U3073 ( .B1(n5257), .B2(net644370), .A(n5638), .ZN(n5636) );
  OAI22_X1 U3072 ( .A1(n532), .A2(n5255), .B1(n657), .B2(n5256), .ZN(n5637) );
  AOI211_X1 U3071 ( .C1(n6361), .C2(net644657), .A(n5636), .B(n5637), .ZN(
        n5619) );
  AOI22_X1 U3070 ( .A1(n6363), .A2(net644529), .B1(n6362), .B2(net644561), 
        .ZN(n5624) );
  AOI22_X1 U3068 ( .A1(n6365), .A2(n438), .B1(n5249), .B2(n4105), .ZN(n5632)
         );
  AOI22_X1 U3067 ( .A1(n3911), .A2(net644626), .B1(n3912), .B2(net644497), 
        .ZN(n5633) );
  AOI22_X1 U3065 ( .A1(n6367), .A2(n4003), .B1(n5245), .B2(n370), .ZN(n5634)
         );
  AOI22_X1 U3064 ( .A1(n3913), .A2(net644594), .B1(n3914), .B2(net644690), 
        .ZN(n5635) );
  NAND4_X1 U3063 ( .A1(n5632), .A2(n5633), .A3(n5634), .A4(n5635), .ZN(n5626)
         );
  AOI22_X1 U3061 ( .A1(n6369), .A2(n440), .B1(n5237), .B2(n4109), .ZN(n5628)
         );
  AOI22_X1 U3060 ( .A1(n3910), .A2(net644786), .B1(n3909), .B2(net644754), 
        .ZN(n5629) );
  AOI22_X1 U3059 ( .A1(n3908), .A2(net644916), .B1(n3907), .B2(net644433), 
        .ZN(n5630) );
  AOI22_X1 U3057 ( .A1(n3906), .A2(n4004), .B1(n3905), .B2(n439), .ZN(n5631)
         );
  NAND4_X1 U3056 ( .A1(n5628), .A2(n5629), .A3(n5630), .A4(n5631), .ZN(n5627)
         );
  OAI21_X1 U3055 ( .B1(n5626), .B2(n5627), .A(n6370), .ZN(n5625) );
  OAI211_X1 U3054 ( .C1(n563), .C2(n5220), .A(n5624), .B(n5625), .ZN(n5621) );
  AOI22_X1 U3052 ( .A1(n6373), .A2(net644817), .B1(n6372), .B2(n4112), .ZN(
        n5623) );
  OAI21_X1 U3051 ( .B1(n625), .B2(n5216), .A(n5623), .ZN(n5622) );
  AOI211_X1 U3050 ( .C1(n5213), .C2(net644722), .A(n5621), .B(n5622), .ZN(
        n5620) );
  NAND4_X1 U3049 ( .A1(n5617), .A2(n5618), .A3(n5619), .A4(n5620), .ZN(n2710)
         );
  AOI22_X1 U3226 ( .A1(n6356), .A2(n3925), .B1(n6355), .B2(n3981), .ZN(n5727)
         );
  AOI22_X1 U3225 ( .A1(n6358), .A2(net644878), .B1(n6357), .B2(net644844), 
        .ZN(n5728) );
  AOI22_X1 U3224 ( .A1(n6360), .A2(net644460), .B1(n6359), .B2(DATAIN[9]), 
        .ZN(n5748) );
  OAI21_X1 U3223 ( .B1(n5257), .B2(net644365), .A(n5748), .ZN(n5746) );
  OAI22_X1 U3222 ( .A1(n537), .A2(n5255), .B1(n662), .B2(n5256), .ZN(n5747) );
  AOI211_X1 U3221 ( .C1(n6361), .C2(net644652), .A(n5746), .B(n5747), .ZN(
        n5729) );
  AOI22_X1 U3220 ( .A1(n6363), .A2(net644524), .B1(n6362), .B2(net644556), 
        .ZN(n5734) );
  AOI22_X1 U3218 ( .A1(n6365), .A2(n453), .B1(n6364), .B2(n4090), .ZN(n5742)
         );
  AOI22_X1 U3217 ( .A1(n3911), .A2(net644621), .B1(n3912), .B2(net644492), 
        .ZN(n5743) );
  AOI22_X1 U3215 ( .A1(n6367), .A2(n3982), .B1(n6366), .B2(n375), .ZN(n5744)
         );
  AOI22_X1 U3214 ( .A1(n3913), .A2(net644589), .B1(n3914), .B2(net644685), 
        .ZN(n5745) );
  NAND4_X1 U3213 ( .A1(n5742), .A2(n5743), .A3(n5744), .A4(n5745), .ZN(n5736)
         );
  AOI22_X1 U3211 ( .A1(n6369), .A2(n455), .B1(n6368), .B2(n4091), .ZN(n5738)
         );
  AOI22_X1 U3210 ( .A1(n3910), .A2(net644781), .B1(n3909), .B2(net644749), 
        .ZN(n5739) );
  AOI22_X1 U3209 ( .A1(n3908), .A2(net644911), .B1(n3907), .B2(net644428), 
        .ZN(n5740) );
  AOI22_X1 U3207 ( .A1(n3906), .A2(n3983), .B1(n3905), .B2(n454), .ZN(n5741)
         );
  NAND4_X1 U3206 ( .A1(n5738), .A2(n5739), .A3(n5740), .A4(n5741), .ZN(n5737)
         );
  OAI21_X1 U3205 ( .B1(n5736), .B2(n5737), .A(n6370), .ZN(n5735) );
  OAI211_X1 U3204 ( .C1(n568), .C2(n5220), .A(n5734), .B(n5735), .ZN(n5731) );
  AOI22_X1 U3202 ( .A1(n6373), .A2(net644812), .B1(n6372), .B2(n4092), .ZN(
        n5733) );
  OAI21_X1 U3201 ( .B1(n630), .B2(n5216), .A(n5733), .ZN(n5732) );
  AOI211_X1 U3200 ( .C1(n6374), .C2(net644717), .A(n5731), .B(n5732), .ZN(
        n5730) );
  NAND4_X1 U3199 ( .A1(n5727), .A2(n5728), .A3(n5729), .A4(n5730), .ZN(n2705)
         );
  AOI22_X1 U3106 ( .A1(n6356), .A2(n3931), .B1(n5264), .B2(n3993), .ZN(n5639)
         );
  AOI22_X1 U3105 ( .A1(n6358), .A2(net644882), .B1(n6357), .B2(net644848), 
        .ZN(n5640) );
  AOI22_X1 U3104 ( .A1(n6360), .A2(net644464), .B1(n6359), .B2(DATAIN[13]), 
        .ZN(n5660) );
  OAI21_X1 U3103 ( .B1(n5257), .B2(net644369), .A(n5660), .ZN(n5658) );
  OAI22_X1 U3102 ( .A1(n533), .A2(n5255), .B1(n658), .B2(n5256), .ZN(n5659) );
  AOI211_X1 U3101 ( .C1(n6361), .C2(net644656), .A(n5658), .B(n5659), .ZN(
        n5641) );
  AOI22_X1 U3100 ( .A1(n6363), .A2(net644528), .B1(n6362), .B2(net644560), 
        .ZN(n5646) );
  AOI22_X1 U3098 ( .A1(n6365), .A2(n441), .B1(n5249), .B2(n4102), .ZN(n5654)
         );
  AOI22_X1 U3097 ( .A1(n3911), .A2(net644625), .B1(n3912), .B2(net644496), 
        .ZN(n5655) );
  AOI22_X1 U3095 ( .A1(n6367), .A2(n3998), .B1(n5245), .B2(n371), .ZN(n5656)
         );
  AOI22_X1 U3094 ( .A1(n3913), .A2(net644593), .B1(n3914), .B2(net644689), 
        .ZN(n5657) );
  NAND4_X1 U3093 ( .A1(n5654), .A2(n5655), .A3(n5656), .A4(n5657), .ZN(n5648)
         );
  AOI22_X1 U3091 ( .A1(n6369), .A2(n443), .B1(n5237), .B2(n4103), .ZN(n5650)
         );
  AOI22_X1 U3090 ( .A1(n3910), .A2(net644785), .B1(n3909), .B2(net644753), 
        .ZN(n5651) );
  AOI22_X1 U3089 ( .A1(n3908), .A2(net644915), .B1(n3907), .B2(net644432), 
        .ZN(n5652) );
  AOI22_X1 U3087 ( .A1(n3906), .A2(n3999), .B1(n3905), .B2(n442), .ZN(n5653)
         );
  NAND4_X1 U3086 ( .A1(n5650), .A2(n5651), .A3(n5652), .A4(n5653), .ZN(n5649)
         );
  OAI21_X1 U3085 ( .B1(n5648), .B2(n5649), .A(n6370), .ZN(n5647) );
  OAI211_X1 U3084 ( .C1(n564), .C2(n5220), .A(n5646), .B(n5647), .ZN(n5643) );
  AOI22_X1 U3082 ( .A1(n6373), .A2(net644816), .B1(n6372), .B2(n4104), .ZN(
        n5645) );
  OAI21_X1 U3081 ( .B1(n626), .B2(n5216), .A(n5645), .ZN(n5644) );
  AOI211_X1 U3080 ( .C1(n5213), .C2(net644721), .A(n5643), .B(n5644), .ZN(
        n5642) );
  NAND4_X1 U3079 ( .A1(n5639), .A2(n5640), .A3(n5641), .A4(n5642), .ZN(n2709)
         );
  AOI22_X1 U2986 ( .A1(n5263), .A2(n3935), .B1(n5264), .B2(n4011), .ZN(n5551)
         );
  AOI22_X1 U2985 ( .A1(n6358), .A2(net644886), .B1(n6357), .B2(net644852), 
        .ZN(n5552) );
  AOI22_X1 U2984 ( .A1(n5259), .A2(net644468), .B1(n6359), .B2(DATAIN[17]), 
        .ZN(n5572) );
  OAI21_X1 U2983 ( .B1(n5257), .B2(net644373), .A(n5572), .ZN(n5570) );
  OAI22_X1 U2982 ( .A1(n529), .A2(n5255), .B1(n654), .B2(n5256), .ZN(n5571) );
  AOI211_X1 U2981 ( .C1(n6361), .C2(net644660), .A(n5570), .B(n5571), .ZN(
        n5553) );
  AOI22_X1 U2980 ( .A1(n5250), .A2(net644532), .B1(n6362), .B2(net644564), 
        .ZN(n5558) );
  AOI22_X1 U2978 ( .A1(n6365), .A2(n429), .B1(n5249), .B2(n4119), .ZN(n5566)
         );
  AOI22_X1 U2977 ( .A1(n3911), .A2(net644629), .B1(n3912), .B2(net644500), 
        .ZN(n5567) );
  AOI22_X1 U2975 ( .A1(n6367), .A2(n4012), .B1(n5245), .B2(n367), .ZN(n5568)
         );
  AOI22_X1 U2974 ( .A1(n3913), .A2(net644597), .B1(n3914), .B2(net644693), 
        .ZN(n5569) );
  NAND4_X1 U2973 ( .A1(n5566), .A2(n5567), .A3(n5568), .A4(n5569), .ZN(n5560)
         );
  AOI22_X1 U2971 ( .A1(n6369), .A2(n431), .B1(n5237), .B2(n4120), .ZN(n5562)
         );
  AOI22_X1 U2970 ( .A1(n3910), .A2(net644789), .B1(n3909), .B2(net644757), 
        .ZN(n5563) );
  AOI22_X1 U2969 ( .A1(n3908), .A2(net644919), .B1(n3907), .B2(net644436), 
        .ZN(n5564) );
  AOI22_X1 U2967 ( .A1(n3906), .A2(n4013), .B1(n3905), .B2(n430), .ZN(n5565)
         );
  NAND4_X1 U2966 ( .A1(n5562), .A2(n5563), .A3(n5564), .A4(n5565), .ZN(n5561)
         );
  OAI21_X1 U2965 ( .B1(n5560), .B2(n5561), .A(n6370), .ZN(n5559) );
  OAI211_X1 U2964 ( .C1(n560), .C2(n5220), .A(n5558), .B(n5559), .ZN(n5555) );
  AOI22_X1 U2962 ( .A1(n6373), .A2(net644820), .B1(n6372), .B2(n4121), .ZN(
        n5557) );
  OAI21_X1 U2961 ( .B1(n622), .B2(n5216), .A(n5557), .ZN(n5556) );
  AOI211_X1 U2960 ( .C1(n5213), .C2(net644725), .A(n5555), .B(n5556), .ZN(
        n5554) );
  NAND4_X1 U2959 ( .A1(n5551), .A2(n5552), .A3(n5553), .A4(n5554), .ZN(n2713)
         );
  AOI22_X1 U3436 ( .A1(n6356), .A2(n3917), .B1(n6355), .B2(n3957), .ZN(n5881)
         );
  AOI22_X1 U3435 ( .A1(n6358), .A2(net644871), .B1(n5262), .B2(net644837), 
        .ZN(n5882) );
  AOI22_X1 U3434 ( .A1(n6360), .A2(net644453), .B1(n6359), .B2(DATAIN[2]), 
        .ZN(n5902) );
  OAI21_X1 U3433 ( .B1(n5257), .B2(net644358), .A(n5902), .ZN(n5900) );
  OAI22_X1 U3432 ( .A1(n544), .A2(n5255), .B1(n669), .B2(n5256), .ZN(n5901) );
  AOI211_X1 U3431 ( .C1(n6361), .C2(net644645), .A(n5900), .B(n5901), .ZN(
        n5883) );
  AOI22_X1 U3430 ( .A1(n6363), .A2(net644517), .B1(n6362), .B2(net644549), 
        .ZN(n5888) );
  AOI22_X1 U3428 ( .A1(n5248), .A2(n474), .B1(n6364), .B2(n4065), .ZN(n5896)
         );
  AOI22_X1 U3427 ( .A1(n3911), .A2(net644614), .B1(n3912), .B2(net644485), 
        .ZN(n5897) );
  AOI22_X1 U3425 ( .A1(n5244), .A2(n3958), .B1(n6366), .B2(n382), .ZN(n5898)
         );
  AOI22_X1 U3424 ( .A1(n3913), .A2(net644582), .B1(n3914), .B2(net644678), 
        .ZN(n5899) );
  NAND4_X1 U3423 ( .A1(n5896), .A2(n5897), .A3(n5898), .A4(n5899), .ZN(n5890)
         );
  AOI22_X1 U3421 ( .A1(n5236), .A2(n476), .B1(n6368), .B2(n4066), .ZN(n5892)
         );
  AOI22_X1 U3420 ( .A1(n3910), .A2(net644774), .B1(n3909), .B2(net644742), 
        .ZN(n5893) );
  AOI22_X1 U3419 ( .A1(n3908), .A2(net644904), .B1(n3907), .B2(net644421), 
        .ZN(n5894) );
  AOI22_X1 U3417 ( .A1(n3906), .A2(n3960), .B1(n3905), .B2(n475), .ZN(n5895)
         );
  NAND4_X1 U3416 ( .A1(n5892), .A2(n5893), .A3(n5894), .A4(n5895), .ZN(n5891)
         );
  OAI21_X1 U3415 ( .B1(n5890), .B2(n5891), .A(n6370), .ZN(n5889) );
  OAI211_X1 U3414 ( .C1(n575), .C2(n5220), .A(n5888), .B(n5889), .ZN(n5885) );
  AOI22_X1 U3412 ( .A1(n6373), .A2(net644805), .B1(n6372), .B2(n4067), .ZN(
        n5887) );
  OAI21_X1 U3411 ( .B1(n637), .B2(n5216), .A(n5887), .ZN(n5886) );
  AOI211_X1 U3410 ( .C1(n6374), .C2(net644710), .A(n5885), .B(n5886), .ZN(
        n5884) );
  NAND4_X1 U3409 ( .A1(n5881), .A2(n5882), .A3(n5883), .A4(n5884), .ZN(n2698)
         );
  AOI22_X1 U3136 ( .A1(n6356), .A2(n3930), .B1(n6355), .B2(n3990), .ZN(n5661)
         );
  AOI22_X1 U3135 ( .A1(n6358), .A2(net644881), .B1(n6357), .B2(net644847), 
        .ZN(n5662) );
  AOI22_X1 U3134 ( .A1(n6360), .A2(net644463), .B1(n6359), .B2(DATAIN[12]), 
        .ZN(n5682) );
  OAI21_X1 U3133 ( .B1(n5257), .B2(net644368), .A(n5682), .ZN(n5680) );
  OAI22_X1 U3132 ( .A1(n534), .A2(n5255), .B1(n659), .B2(n5256), .ZN(n5681) );
  AOI211_X1 U3131 ( .C1(n6361), .C2(net644655), .A(n5680), .B(n5681), .ZN(
        n5663) );
  AOI22_X1 U3130 ( .A1(n6363), .A2(net644527), .B1(n6362), .B2(net644559), 
        .ZN(n5668) );
  AOI22_X1 U3128 ( .A1(n6365), .A2(n444), .B1(n6364), .B2(n4099), .ZN(n5676)
         );
  AOI22_X1 U3127 ( .A1(n3911), .A2(net644624), .B1(n3912), .B2(net644495), 
        .ZN(n5677) );
  AOI22_X1 U3125 ( .A1(n6367), .A2(n3991), .B1(n6366), .B2(n372), .ZN(n5678)
         );
  AOI22_X1 U3124 ( .A1(n3913), .A2(net644592), .B1(n3914), .B2(net644688), 
        .ZN(n5679) );
  NAND4_X1 U3123 ( .A1(n5676), .A2(n5677), .A3(n5678), .A4(n5679), .ZN(n5670)
         );
  AOI22_X1 U3121 ( .A1(n6369), .A2(n446), .B1(n6368), .B2(n4100), .ZN(n5672)
         );
  AOI22_X1 U3120 ( .A1(n3910), .A2(net644784), .B1(n3909), .B2(net644752), 
        .ZN(n5673) );
  AOI22_X1 U3119 ( .A1(n3908), .A2(net644914), .B1(n3907), .B2(net644431), 
        .ZN(n5674) );
  AOI22_X1 U3117 ( .A1(n3906), .A2(n3992), .B1(n3905), .B2(n445), .ZN(n5675)
         );
  NAND4_X1 U3116 ( .A1(n5672), .A2(n5673), .A3(n5674), .A4(n5675), .ZN(n5671)
         );
  OAI21_X1 U3115 ( .B1(n5670), .B2(n5671), .A(n5225), .ZN(n5669) );
  OAI211_X1 U3114 ( .C1(n565), .C2(n5220), .A(n5668), .B(n5669), .ZN(n5665) );
  AOI22_X1 U3112 ( .A1(n6373), .A2(net644815), .B1(n6372), .B2(n4101), .ZN(
        n5667) );
  OAI21_X1 U3111 ( .B1(n627), .B2(n5216), .A(n5667), .ZN(n5666) );
  AOI211_X1 U3110 ( .C1(n6374), .C2(net644720), .A(n5665), .B(n5666), .ZN(
        n5664) );
  NAND4_X1 U3109 ( .A1(n5661), .A2(n5662), .A3(n5663), .A4(n5664), .ZN(n2708)
         );
  AOI22_X1 U3196 ( .A1(n6356), .A2(n3928), .B1(n6355), .B2(n3984), .ZN(n5705)
         );
  AOI22_X1 U3195 ( .A1(n6358), .A2(net644879), .B1(n6357), .B2(net644845), 
        .ZN(n5706) );
  AOI22_X1 U3194 ( .A1(n6360), .A2(net644461), .B1(n6359), .B2(DATAIN[10]), 
        .ZN(n5726) );
  OAI21_X1 U3193 ( .B1(n5257), .B2(net644366), .A(n5726), .ZN(n5724) );
  OAI22_X1 U3192 ( .A1(n536), .A2(n5255), .B1(n661), .B2(n5256), .ZN(n5725) );
  AOI211_X1 U3191 ( .C1(n6361), .C2(net644653), .A(n5724), .B(n5725), .ZN(
        n5707) );
  AOI22_X1 U3190 ( .A1(n6363), .A2(net644525), .B1(n6362), .B2(net644557), 
        .ZN(n5712) );
  AOI22_X1 U3188 ( .A1(n6365), .A2(n450), .B1(n6364), .B2(n4093), .ZN(n5720)
         );
  AOI22_X1 U3187 ( .A1(n3911), .A2(net644622), .B1(n3912), .B2(net644493), 
        .ZN(n5721) );
  AOI22_X1 U3185 ( .A1(n6367), .A2(n3985), .B1(n6366), .B2(n374), .ZN(n5722)
         );
  AOI22_X1 U3184 ( .A1(n3913), .A2(net644590), .B1(n3914), .B2(net644686), 
        .ZN(n5723) );
  NAND4_X1 U3183 ( .A1(n5720), .A2(n5721), .A3(n5722), .A4(n5723), .ZN(n5714)
         );
  AOI22_X1 U3181 ( .A1(n6369), .A2(n452), .B1(n6368), .B2(n4094), .ZN(n5716)
         );
  AOI22_X1 U3180 ( .A1(n3910), .A2(net644782), .B1(n3909), .B2(net644750), 
        .ZN(n5717) );
  AOI22_X1 U3179 ( .A1(n3908), .A2(net644912), .B1(n3907), .B2(net644429), 
        .ZN(n5718) );
  AOI22_X1 U3177 ( .A1(n3906), .A2(n3986), .B1(n3905), .B2(n451), .ZN(n5719)
         );
  NAND4_X1 U3176 ( .A1(n5716), .A2(n5717), .A3(n5718), .A4(n5719), .ZN(n5715)
         );
  OAI21_X1 U3175 ( .B1(n5714), .B2(n5715), .A(n6370), .ZN(n5713) );
  OAI211_X1 U3174 ( .C1(n567), .C2(n5220), .A(n5712), .B(n5713), .ZN(n5709) );
  AOI22_X1 U3172 ( .A1(n6373), .A2(net644813), .B1(n6372), .B2(n4095), .ZN(
        n5711) );
  OAI21_X1 U3171 ( .B1(n629), .B2(n5216), .A(n5711), .ZN(n5710) );
  AOI211_X1 U3170 ( .C1(n6374), .C2(net644718), .A(n5709), .B(n5710), .ZN(
        n5708) );
  NAND4_X1 U3169 ( .A1(n5705), .A2(n5706), .A3(n5707), .A4(n5708), .ZN(n2706)
         );
  AOI22_X1 U3166 ( .A1(n6356), .A2(n3929), .B1(n6355), .B2(n3987), .ZN(n5683)
         );
  AOI22_X1 U3165 ( .A1(n6358), .A2(net644880), .B1(n6357), .B2(net644846), 
        .ZN(n5684) );
  AOI22_X1 U3164 ( .A1(n6360), .A2(net644462), .B1(n6359), .B2(DATAIN[11]), 
        .ZN(n5704) );
  OAI21_X1 U3163 ( .B1(n5257), .B2(net644367), .A(n5704), .ZN(n5702) );
  OAI22_X1 U3162 ( .A1(n535), .A2(n5255), .B1(n660), .B2(n5256), .ZN(n5703) );
  AOI211_X1 U3161 ( .C1(n6361), .C2(net644654), .A(n5702), .B(n5703), .ZN(
        n5685) );
  AOI22_X1 U3160 ( .A1(n6363), .A2(net644526), .B1(n6362), .B2(net644558), 
        .ZN(n5690) );
  AOI22_X1 U3158 ( .A1(n6365), .A2(n447), .B1(n6364), .B2(n4096), .ZN(n5698)
         );
  AOI22_X1 U3157 ( .A1(n3911), .A2(net644623), .B1(n3912), .B2(net644494), 
        .ZN(n5699) );
  AOI22_X1 U3155 ( .A1(n6367), .A2(n3988), .B1(n6366), .B2(n373), .ZN(n5700)
         );
  AOI22_X1 U3154 ( .A1(n3913), .A2(net644591), .B1(n3914), .B2(net644687), 
        .ZN(n5701) );
  NAND4_X1 U3153 ( .A1(n5698), .A2(n5699), .A3(n5700), .A4(n5701), .ZN(n5692)
         );
  AOI22_X1 U3151 ( .A1(n6369), .A2(n449), .B1(n6368), .B2(n4097), .ZN(n5694)
         );
  AOI22_X1 U3150 ( .A1(n3910), .A2(net644783), .B1(n3909), .B2(net644751), 
        .ZN(n5695) );
  AOI22_X1 U3149 ( .A1(n3908), .A2(net644913), .B1(n3907), .B2(net644430), 
        .ZN(n5696) );
  AOI22_X1 U3147 ( .A1(n3906), .A2(n3989), .B1(n3905), .B2(n448), .ZN(n5697)
         );
  NAND4_X1 U3146 ( .A1(n5694), .A2(n5695), .A3(n5696), .A4(n5697), .ZN(n5693)
         );
  OAI21_X1 U3145 ( .B1(n5692), .B2(n5693), .A(n6370), .ZN(n5691) );
  OAI211_X1 U3144 ( .C1(n566), .C2(n5220), .A(n5690), .B(n5691), .ZN(n5687) );
  AOI22_X1 U3142 ( .A1(n6373), .A2(net644814), .B1(n6372), .B2(n4098), .ZN(
        n5689) );
  OAI21_X1 U3141 ( .B1(n628), .B2(n5216), .A(n5689), .ZN(n5688) );
  AOI211_X1 U3140 ( .C1(n6374), .C2(net644719), .A(n5687), .B(n5688), .ZN(
        n5686) );
  NAND4_X1 U3139 ( .A1(n5683), .A2(n5684), .A3(n5685), .A4(n5686), .ZN(n2707)
         );
  AOI22_X1 U3406 ( .A1(n6356), .A2(n3918), .B1(n6355), .B2(n3963), .ZN(n5859)
         );
  AOI22_X1 U3405 ( .A1(n6358), .A2(net644872), .B1(n5262), .B2(net644838), 
        .ZN(n5860) );
  AOI22_X1 U3404 ( .A1(n6360), .A2(net644454), .B1(n6359), .B2(DATAIN[3]), 
        .ZN(n5880) );
  OAI21_X1 U3403 ( .B1(n5257), .B2(net644359), .A(n5880), .ZN(n5878) );
  OAI22_X1 U3402 ( .A1(n543), .A2(n5255), .B1(n668), .B2(n5256), .ZN(n5879) );
  AOI211_X1 U3401 ( .C1(n6361), .C2(net644646), .A(n5878), .B(n5879), .ZN(
        n5861) );
  AOI22_X1 U3400 ( .A1(n6363), .A2(net644518), .B1(n6362), .B2(net644550), 
        .ZN(n5866) );
  AOI22_X1 U3398 ( .A1(n5248), .A2(n471), .B1(n6364), .B2(n4070), .ZN(n5874)
         );
  AOI22_X1 U3397 ( .A1(n3911), .A2(net644615), .B1(n3912), .B2(net644486), 
        .ZN(n5875) );
  AOI22_X1 U3395 ( .A1(n5244), .A2(n3964), .B1(n6366), .B2(n381), .ZN(n5876)
         );
  AOI22_X1 U3394 ( .A1(n3913), .A2(net644583), .B1(n3914), .B2(net644679), 
        .ZN(n5877) );
  NAND4_X1 U3393 ( .A1(n5874), .A2(n5875), .A3(n5876), .A4(n5877), .ZN(n5868)
         );
  AOI22_X1 U3391 ( .A1(n5236), .A2(n473), .B1(n6368), .B2(n4071), .ZN(n5870)
         );
  AOI22_X1 U3390 ( .A1(n3910), .A2(net644775), .B1(n3909), .B2(net644743), 
        .ZN(n5871) );
  AOI22_X1 U3389 ( .A1(n3908), .A2(net644905), .B1(n3907), .B2(net644422), 
        .ZN(n5872) );
  AOI22_X1 U3387 ( .A1(n3906), .A2(n3965), .B1(n3905), .B2(n472), .ZN(n5873)
         );
  NAND4_X1 U3386 ( .A1(n5870), .A2(n5871), .A3(n5872), .A4(n5873), .ZN(n5869)
         );
  OAI21_X1 U3385 ( .B1(n5868), .B2(n5869), .A(n6370), .ZN(n5867) );
  OAI211_X1 U3384 ( .C1(n574), .C2(n5220), .A(n5866), .B(n5867), .ZN(n5863) );
  AOI22_X1 U3382 ( .A1(n6373), .A2(net644806), .B1(n6372), .B2(n4072), .ZN(
        n5865) );
  OAI21_X1 U3381 ( .B1(n636), .B2(n5216), .A(n5865), .ZN(n5864) );
  AOI211_X1 U3380 ( .C1(n6374), .C2(net644711), .A(n5863), .B(n5864), .ZN(
        n5862) );
  NAND4_X1 U3379 ( .A1(n5859), .A2(n5860), .A3(n5861), .A4(n5862), .ZN(n2699)
         );
  AOI22_X1 U2926 ( .A1(n5263), .A2(n3937), .B1(n6355), .B2(n4017), .ZN(n5507)
         );
  AOI22_X1 U2925 ( .A1(n5261), .A2(net644888), .B1(n6357), .B2(net644854), 
        .ZN(n5508) );
  AOI22_X1 U2924 ( .A1(n6360), .A2(net644470), .B1(n6359), .B2(DATAIN[19]), 
        .ZN(n5528) );
  OAI21_X1 U2923 ( .B1(n5257), .B2(net644375), .A(n5528), .ZN(n5526) );
  OAI22_X1 U2922 ( .A1(n527), .A2(n5255), .B1(n652), .B2(n5256), .ZN(n5527) );
  AOI211_X1 U2921 ( .C1(n6361), .C2(net644662), .A(n5526), .B(n5527), .ZN(
        n5509) );
  AOI22_X1 U2920 ( .A1(n6363), .A2(net644534), .B1(n6362), .B2(net644566), 
        .ZN(n5514) );
  AOI22_X1 U2918 ( .A1(n6365), .A2(n423), .B1(n6364), .B2(n4125), .ZN(n5522)
         );
  AOI22_X1 U2917 ( .A1(n3911), .A2(net644631), .B1(n3912), .B2(net644502), 
        .ZN(n5523) );
  AOI22_X1 U2915 ( .A1(n6367), .A2(n4018), .B1(n6366), .B2(n365), .ZN(n5524)
         );
  AOI22_X1 U2914 ( .A1(n3913), .A2(net644599), .B1(n3914), .B2(net644695), 
        .ZN(n5525) );
  NAND4_X1 U2913 ( .A1(n5522), .A2(n5523), .A3(n5524), .A4(n5525), .ZN(n5516)
         );
  AOI22_X1 U2911 ( .A1(n6369), .A2(n425), .B1(n6368), .B2(n4126), .ZN(n5518)
         );
  AOI22_X1 U2910 ( .A1(n3910), .A2(net644791), .B1(n3909), .B2(net644759), 
        .ZN(n5519) );
  AOI22_X1 U2909 ( .A1(n3908), .A2(net644921), .B1(n3907), .B2(net644438), 
        .ZN(n5520) );
  AOI22_X1 U2907 ( .A1(n3906), .A2(n4019), .B1(n3905), .B2(n424), .ZN(n5521)
         );
  NAND4_X1 U2906 ( .A1(n5518), .A2(n5519), .A3(n5520), .A4(n5521), .ZN(n5517)
         );
  OAI21_X1 U2905 ( .B1(n5516), .B2(n5517), .A(n6370), .ZN(n5515) );
  OAI211_X1 U2904 ( .C1(n558), .C2(n5220), .A(n5514), .B(n5515), .ZN(n5511) );
  AOI22_X1 U2902 ( .A1(n6373), .A2(net644822), .B1(n6372), .B2(n4127), .ZN(
        n5513) );
  OAI21_X1 U2901 ( .B1(n620), .B2(n5216), .A(n5513), .ZN(n5512) );
  AOI211_X1 U2900 ( .C1(n6374), .C2(net644727), .A(n5511), .B(n5512), .ZN(
        n5510) );
  NAND4_X1 U2899 ( .A1(n5507), .A2(n5508), .A3(n5509), .A4(n5510), .ZN(n2715)
         );
  AOI22_X1 U2896 ( .A1(n6356), .A2(n3938), .B1(n6355), .B2(n4020), .ZN(n5485)
         );
  AOI22_X1 U2895 ( .A1(n6358), .A2(net644889), .B1(n6357), .B2(net644855), 
        .ZN(n5486) );
  AOI22_X1 U2894 ( .A1(n6360), .A2(net644471), .B1(n6359), .B2(DATAIN[20]), 
        .ZN(n5506) );
  OAI21_X1 U2893 ( .B1(n5257), .B2(net644376), .A(n5506), .ZN(n5504) );
  OAI22_X1 U2892 ( .A1(n526), .A2(n5255), .B1(n651), .B2(n5256), .ZN(n5505) );
  AOI211_X1 U2891 ( .C1(n6361), .C2(net644663), .A(n5504), .B(n5505), .ZN(
        n5487) );
  AOI22_X1 U2890 ( .A1(n6363), .A2(net644535), .B1(n6362), .B2(net644567), 
        .ZN(n5492) );
  AOI22_X1 U2888 ( .A1(n6365), .A2(n420), .B1(n6364), .B2(n4128), .ZN(n5500)
         );
  AOI22_X1 U2887 ( .A1(n3911), .A2(net644632), .B1(n3912), .B2(net644503), 
        .ZN(n5501) );
  AOI22_X1 U2885 ( .A1(n6367), .A2(n4021), .B1(n6366), .B2(n364), .ZN(n5502)
         );
  AOI22_X1 U2884 ( .A1(n3913), .A2(net644600), .B1(n3914), .B2(net644696), 
        .ZN(n5503) );
  NAND4_X1 U2883 ( .A1(n5500), .A2(n5501), .A3(n5502), .A4(n5503), .ZN(n5494)
         );
  AOI22_X1 U2881 ( .A1(n6369), .A2(n422), .B1(n6368), .B2(n4129), .ZN(n5496)
         );
  AOI22_X1 U2880 ( .A1(n3910), .A2(net644792), .B1(n3909), .B2(net644760), 
        .ZN(n5497) );
  AOI22_X1 U2879 ( .A1(n3908), .A2(net644922), .B1(n3907), .B2(net644439), 
        .ZN(n5498) );
  AOI22_X1 U2877 ( .A1(n3906), .A2(n4022), .B1(n3905), .B2(n421), .ZN(n5499)
         );
  NAND4_X1 U2876 ( .A1(n5496), .A2(n5497), .A3(n5498), .A4(n5499), .ZN(n5495)
         );
  OAI21_X1 U2875 ( .B1(n5494), .B2(n5495), .A(n6370), .ZN(n5493) );
  OAI211_X1 U2874 ( .C1(n557), .C2(n5220), .A(n5492), .B(n5493), .ZN(n5489) );
  AOI22_X1 U2872 ( .A1(n6373), .A2(net644823), .B1(n6372), .B2(n4130), .ZN(
        n5491) );
  OAI21_X1 U2871 ( .B1(n619), .B2(n5216), .A(n5491), .ZN(n5490) );
  AOI211_X1 U2870 ( .C1(n6374), .C2(net644728), .A(n5489), .B(n5490), .ZN(
        n5488) );
  NAND4_X1 U2869 ( .A1(n5485), .A2(n5486), .A3(n5487), .A4(n5488), .ZN(n2716)
         );
  AOI22_X1 U2956 ( .A1(n6356), .A2(n3936), .B1(n5264), .B2(n4014), .ZN(n5529)
         );
  AOI22_X1 U2955 ( .A1(n5261), .A2(net644887), .B1(n6357), .B2(net644853), 
        .ZN(n5530) );
  AOI22_X1 U2954 ( .A1(n6360), .A2(net644469), .B1(n6359), .B2(DATAIN[18]), 
        .ZN(n5550) );
  OAI21_X1 U2953 ( .B1(n5257), .B2(net644374), .A(n5550), .ZN(n5548) );
  OAI22_X1 U2952 ( .A1(n528), .A2(n5255), .B1(n653), .B2(n5256), .ZN(n5549) );
  AOI211_X1 U2951 ( .C1(n6361), .C2(net644661), .A(n5548), .B(n5549), .ZN(
        n5531) );
  AOI22_X1 U2950 ( .A1(n6363), .A2(net644533), .B1(n5251), .B2(net644565), 
        .ZN(n5536) );
  AOI22_X1 U2948 ( .A1(n6365), .A2(n426), .B1(n5249), .B2(n4122), .ZN(n5544)
         );
  AOI22_X1 U2947 ( .A1(n3911), .A2(net644630), .B1(n3912), .B2(net644501), 
        .ZN(n5545) );
  AOI22_X1 U2945 ( .A1(n6367), .A2(n4015), .B1(n5245), .B2(n366), .ZN(n5546)
         );
  AOI22_X1 U2944 ( .A1(n3913), .A2(net644598), .B1(n3914), .B2(net644694), 
        .ZN(n5547) );
  NAND4_X1 U2943 ( .A1(n5544), .A2(n5545), .A3(n5546), .A4(n5547), .ZN(n5538)
         );
  AOI22_X1 U2941 ( .A1(n6369), .A2(n428), .B1(n5237), .B2(n4123), .ZN(n5540)
         );
  AOI22_X1 U2940 ( .A1(n3910), .A2(net644790), .B1(n3909), .B2(net644758), 
        .ZN(n5541) );
  AOI22_X1 U2939 ( .A1(n3908), .A2(net644920), .B1(n3907), .B2(net644437), 
        .ZN(n5542) );
  AOI22_X1 U2937 ( .A1(n3906), .A2(n4016), .B1(n3905), .B2(n427), .ZN(n5543)
         );
  NAND4_X1 U2936 ( .A1(n5540), .A2(n5541), .A3(n5542), .A4(n5543), .ZN(n5539)
         );
  OAI21_X1 U2935 ( .B1(n5538), .B2(n5539), .A(n6370), .ZN(n5537) );
  OAI211_X1 U2934 ( .C1(n559), .C2(n5220), .A(n5536), .B(n5537), .ZN(n5533) );
  AOI22_X1 U2932 ( .A1(n6373), .A2(net644821), .B1(n6372), .B2(n4124), .ZN(
        n5535) );
  OAI21_X1 U2931 ( .B1(n621), .B2(n5216), .A(n5535), .ZN(n5534) );
  AOI211_X1 U2930 ( .C1(n6374), .C2(net644726), .A(n5533), .B(n5534), .ZN(
        n5532) );
  NAND4_X1 U2929 ( .A1(n5529), .A2(n5530), .A3(n5531), .A4(n5532), .ZN(n2714)
         );
  AOI22_X1 U2776 ( .A1(n6356), .A2(n3942), .B1(n5264), .B2(n4032), .ZN(n5397)
         );
  AOI22_X1 U2775 ( .A1(n6358), .A2(net644893), .B1(n5262), .B2(net644859), 
        .ZN(n5398) );
  AOI22_X1 U2774 ( .A1(n6360), .A2(net644475), .B1(n6359), .B2(DATAIN[24]), 
        .ZN(n5418) );
  OAI21_X1 U2773 ( .B1(n5257), .B2(net644380), .A(n5418), .ZN(n5416) );
  OAI22_X1 U2772 ( .A1(n522), .A2(n5255), .B1(n647), .B2(n5256), .ZN(n5417) );
  AOI211_X1 U2771 ( .C1(n6361), .C2(net644667), .A(n5416), .B(n5417), .ZN(
        n5399) );
  AOI22_X1 U2770 ( .A1(n6363), .A2(net644539), .B1(n6362), .B2(net644571), 
        .ZN(n5404) );
  AOI22_X1 U2768 ( .A1(n6365), .A2(n408), .B1(n5249), .B2(n4140), .ZN(n5412)
         );
  AOI22_X1 U2767 ( .A1(n3911), .A2(net644636), .B1(n3912), .B2(net644507), 
        .ZN(n5413) );
  AOI22_X1 U2765 ( .A1(n6367), .A2(n4034), .B1(n5245), .B2(n360), .ZN(n5414)
         );
  AOI22_X1 U2764 ( .A1(n3913), .A2(net644604), .B1(n3914), .B2(net644700), 
        .ZN(n5415) );
  NAND4_X1 U2763 ( .A1(n5412), .A2(n5413), .A3(n5414), .A4(n5415), .ZN(n5406)
         );
  AOI22_X1 U2761 ( .A1(n6369), .A2(n410), .B1(n5237), .B2(n4141), .ZN(n5408)
         );
  AOI22_X1 U2760 ( .A1(n3910), .A2(net644796), .B1(n3909), .B2(net644764), 
        .ZN(n5409) );
  AOI22_X1 U2759 ( .A1(n3908), .A2(net644926), .B1(n3907), .B2(net644443), 
        .ZN(n5410) );
  AOI22_X1 U2757 ( .A1(n3906), .A2(n4037), .B1(n3905), .B2(n409), .ZN(n5411)
         );
  NAND4_X1 U2756 ( .A1(n5408), .A2(n5409), .A3(n5410), .A4(n5411), .ZN(n5407)
         );
  OAI21_X1 U2755 ( .B1(n5406), .B2(n5407), .A(n6370), .ZN(n5405) );
  OAI211_X1 U2754 ( .C1(n553), .C2(n5220), .A(n5404), .B(n5405), .ZN(n5401) );
  AOI22_X1 U2752 ( .A1(n6373), .A2(net644827), .B1(n6372), .B2(n4142), .ZN(
        n5403) );
  OAI21_X1 U2751 ( .B1(n615), .B2(n5216), .A(n5403), .ZN(n5402) );
  AOI211_X1 U2750 ( .C1(n5213), .C2(net644732), .A(n5401), .B(n5402), .ZN(
        n5400) );
  NAND4_X1 U2749 ( .A1(n5397), .A2(n5398), .A3(n5399), .A4(n5400), .ZN(n2720)
         );
  AOI22_X1 U2866 ( .A1(n6356), .A2(n3939), .B1(n6355), .B2(n4023), .ZN(n5463)
         );
  AOI22_X1 U2865 ( .A1(n6358), .A2(net644890), .B1(n6357), .B2(net644856), 
        .ZN(n5464) );
  AOI22_X1 U2864 ( .A1(n6360), .A2(net644472), .B1(n6359), .B2(DATAIN[21]), 
        .ZN(n5484) );
  OAI21_X1 U2863 ( .B1(n5257), .B2(net644377), .A(n5484), .ZN(n5482) );
  OAI22_X1 U2862 ( .A1(n525), .A2(n5255), .B1(n650), .B2(n5256), .ZN(n5483) );
  AOI211_X1 U2861 ( .C1(n6361), .C2(net644664), .A(n5482), .B(n5483), .ZN(
        n5465) );
  AOI22_X1 U2860 ( .A1(n6363), .A2(net644536), .B1(n6362), .B2(net644568), 
        .ZN(n5470) );
  AOI22_X1 U2858 ( .A1(n6365), .A2(n417), .B1(n6364), .B2(n4131), .ZN(n5478)
         );
  AOI22_X1 U2857 ( .A1(n3911), .A2(net644633), .B1(n3912), .B2(net644504), 
        .ZN(n5479) );
  AOI22_X1 U2855 ( .A1(n6367), .A2(n4024), .B1(n6366), .B2(n363), .ZN(n5480)
         );
  AOI22_X1 U2854 ( .A1(n3913), .A2(net644601), .B1(n3914), .B2(net644697), 
        .ZN(n5481) );
  NAND4_X1 U2853 ( .A1(n5478), .A2(n5479), .A3(n5480), .A4(n5481), .ZN(n5472)
         );
  AOI22_X1 U2851 ( .A1(n6369), .A2(n419), .B1(n6368), .B2(n4132), .ZN(n5474)
         );
  AOI22_X1 U2850 ( .A1(n3910), .A2(net644793), .B1(n3909), .B2(net644761), 
        .ZN(n5475) );
  AOI22_X1 U2849 ( .A1(n3908), .A2(net644923), .B1(n3907), .B2(net644440), 
        .ZN(n5476) );
  AOI22_X1 U2847 ( .A1(n3906), .A2(n4025), .B1(n3905), .B2(n418), .ZN(n5477)
         );
  NAND4_X1 U2846 ( .A1(n5474), .A2(n5475), .A3(n5476), .A4(n5477), .ZN(n5473)
         );
  OAI21_X1 U2845 ( .B1(n5472), .B2(n5473), .A(n6370), .ZN(n5471) );
  OAI211_X1 U2844 ( .C1(n556), .C2(n5220), .A(n5470), .B(n5471), .ZN(n5467) );
  AOI22_X1 U2842 ( .A1(n6373), .A2(net644824), .B1(n6372), .B2(n4133), .ZN(
        n5469) );
  OAI21_X1 U2841 ( .B1(n618), .B2(n5216), .A(n5469), .ZN(n5468) );
  AOI211_X1 U2840 ( .C1(n6374), .C2(net644729), .A(n5467), .B(n5468), .ZN(
        n5466) );
  NAND4_X1 U2839 ( .A1(n5463), .A2(n5464), .A3(n5465), .A4(n5466), .ZN(n2717)
         );
  AOI22_X1 U3016 ( .A1(n6356), .A2(n3934), .B1(n5264), .B2(n4008), .ZN(n5573)
         );
  AOI22_X1 U3015 ( .A1(n6358), .A2(net644885), .B1(n6357), .B2(net644851), 
        .ZN(n5574) );
  AOI22_X1 U3014 ( .A1(n6360), .A2(net644467), .B1(n6359), .B2(DATAIN[16]), 
        .ZN(n5594) );
  OAI21_X1 U3013 ( .B1(n5257), .B2(net644372), .A(n5594), .ZN(n5592) );
  OAI22_X1 U3012 ( .A1(n530), .A2(n5255), .B1(n655), .B2(n5256), .ZN(n5593) );
  AOI211_X1 U3011 ( .C1(n6361), .C2(net644659), .A(n5592), .B(n5593), .ZN(
        n5575) );
  AOI22_X1 U3010 ( .A1(n6363), .A2(net644531), .B1(n6362), .B2(net644563), 
        .ZN(n5580) );
  AOI22_X1 U3008 ( .A1(n6365), .A2(n432), .B1(n5249), .B2(n4116), .ZN(n5588)
         );
  AOI22_X1 U3007 ( .A1(n3911), .A2(net644628), .B1(n3912), .B2(net644499), 
        .ZN(n5589) );
  AOI22_X1 U3005 ( .A1(n6367), .A2(n4009), .B1(n5245), .B2(n368), .ZN(n5590)
         );
  AOI22_X1 U3004 ( .A1(n3913), .A2(net644596), .B1(n3914), .B2(net644692), 
        .ZN(n5591) );
  NAND4_X1 U3003 ( .A1(n5588), .A2(n5589), .A3(n5590), .A4(n5591), .ZN(n5582)
         );
  AOI22_X1 U3001 ( .A1(n6369), .A2(n434), .B1(n5237), .B2(n4117), .ZN(n5584)
         );
  AOI22_X1 U3000 ( .A1(n3910), .A2(net644788), .B1(n3909), .B2(net644756), 
        .ZN(n5585) );
  AOI22_X1 U2999 ( .A1(n3908), .A2(net644918), .B1(n3907), .B2(net644435), 
        .ZN(n5586) );
  AOI22_X1 U2997 ( .A1(n3906), .A2(n4010), .B1(n3905), .B2(n433), .ZN(n5587)
         );
  NAND4_X1 U2996 ( .A1(n5584), .A2(n5585), .A3(n5586), .A4(n5587), .ZN(n5583)
         );
  OAI21_X1 U2995 ( .B1(n5582), .B2(n5583), .A(n6370), .ZN(n5581) );
  OAI211_X1 U2994 ( .C1(n561), .C2(n5220), .A(n5580), .B(n5581), .ZN(n5577) );
  AOI22_X1 U2992 ( .A1(n6373), .A2(net644819), .B1(n6372), .B2(n4118), .ZN(
        n5579) );
  OAI21_X1 U2991 ( .B1(n623), .B2(n5216), .A(n5579), .ZN(n5578) );
  AOI211_X1 U2990 ( .C1(n5213), .C2(net644724), .A(n5577), .B(n5578), .ZN(
        n5576) );
  NAND4_X1 U2989 ( .A1(n5573), .A2(n5574), .A3(n5575), .A4(n5576), .ZN(n2712)
         );
  AOI22_X1 U3256 ( .A1(n6356), .A2(n3923), .B1(n6355), .B2(n3978), .ZN(n5749)
         );
  AOI22_X1 U3255 ( .A1(n6358), .A2(net644877), .B1(n6357), .B2(net644843), 
        .ZN(n5750) );
  AOI22_X1 U3254 ( .A1(n6360), .A2(net644459), .B1(n6359), .B2(DATAIN[8]), 
        .ZN(n5770) );
  OAI21_X1 U3253 ( .B1(n5257), .B2(net644364), .A(n5770), .ZN(n5768) );
  OAI22_X1 U3252 ( .A1(n538), .A2(n5255), .B1(n663), .B2(n5256), .ZN(n5769) );
  AOI211_X1 U3251 ( .C1(n6361), .C2(net644651), .A(n5768), .B(n5769), .ZN(
        n5751) );
  AOI22_X1 U3250 ( .A1(n6363), .A2(net644523), .B1(n6362), .B2(net644555), 
        .ZN(n5756) );
  AOI22_X1 U3248 ( .A1(n6365), .A2(n456), .B1(n6364), .B2(n4087), .ZN(n5764)
         );
  AOI22_X1 U3247 ( .A1(n3911), .A2(net644620), .B1(n3912), .B2(net644491), 
        .ZN(n5765) );
  AOI22_X1 U3245 ( .A1(n6367), .A2(n3979), .B1(n6366), .B2(n376), .ZN(n5766)
         );
  AOI22_X1 U3244 ( .A1(n3913), .A2(net644588), .B1(n3914), .B2(net644684), 
        .ZN(n5767) );
  NAND4_X1 U3243 ( .A1(n5764), .A2(n5765), .A3(n5766), .A4(n5767), .ZN(n5758)
         );
  AOI22_X1 U3241 ( .A1(n6369), .A2(n458), .B1(n6368), .B2(n4088), .ZN(n5760)
         );
  AOI22_X1 U3240 ( .A1(n3910), .A2(net644780), .B1(n3909), .B2(net644748), 
        .ZN(n5761) );
  AOI22_X1 U3239 ( .A1(n3908), .A2(net644910), .B1(n3907), .B2(net644427), 
        .ZN(n5762) );
  AOI22_X1 U3237 ( .A1(n3906), .A2(n3980), .B1(n3905), .B2(n457), .ZN(n5763)
         );
  NAND4_X1 U3236 ( .A1(n5760), .A2(n5761), .A3(n5762), .A4(n5763), .ZN(n5759)
         );
  OAI21_X1 U3235 ( .B1(n5758), .B2(n5759), .A(n6370), .ZN(n5757) );
  OAI211_X1 U3234 ( .C1(n569), .C2(n5220), .A(n5756), .B(n5757), .ZN(n5753) );
  AOI22_X1 U3232 ( .A1(n6373), .A2(net644811), .B1(n6372), .B2(n4089), .ZN(
        n5755) );
  OAI21_X1 U3231 ( .B1(n631), .B2(n5216), .A(n5755), .ZN(n5754) );
  AOI211_X1 U3230 ( .C1(n6374), .C2(net644716), .A(n5753), .B(n5754), .ZN(
        n5752) );
  NAND4_X1 U3229 ( .A1(n5749), .A2(n5750), .A3(n5751), .A4(n5752), .ZN(n2704)
         );
  AOI22_X1 U3316 ( .A1(n6356), .A2(n3921), .B1(n6355), .B2(n3972), .ZN(n5793)
         );
  AOI22_X1 U3315 ( .A1(n6358), .A2(net644875), .B1(n5262), .B2(net644841), 
        .ZN(n5794) );
  AOI22_X1 U3314 ( .A1(n6360), .A2(net644457), .B1(n6359), .B2(DATAIN[6]), 
        .ZN(n5814) );
  OAI21_X1 U3313 ( .B1(n5257), .B2(net644362), .A(n5814), .ZN(n5812) );
  OAI22_X1 U3312 ( .A1(n540), .A2(n5255), .B1(n665), .B2(n5256), .ZN(n5813) );
  AOI211_X1 U3311 ( .C1(n6361), .C2(net644649), .A(n5812), .B(n5813), .ZN(
        n5795) );
  AOI22_X1 U3310 ( .A1(n6363), .A2(net644521), .B1(n6362), .B2(net644553), 
        .ZN(n5800) );
  AOI22_X1 U3308 ( .A1(n5248), .A2(n462), .B1(n6364), .B2(n4081), .ZN(n5808)
         );
  AOI22_X1 U3307 ( .A1(n3911), .A2(net644618), .B1(n3912), .B2(net644489), 
        .ZN(n5809) );
  AOI22_X1 U3305 ( .A1(n5244), .A2(n3973), .B1(n6366), .B2(n378), .ZN(n5810)
         );
  AOI22_X1 U3304 ( .A1(n3913), .A2(net644586), .B1(n3914), .B2(net644682), 
        .ZN(n5811) );
  NAND4_X1 U3303 ( .A1(n5808), .A2(n5809), .A3(n5810), .A4(n5811), .ZN(n5802)
         );
  AOI22_X1 U3301 ( .A1(n5236), .A2(n464), .B1(n6368), .B2(n4082), .ZN(n5804)
         );
  AOI22_X1 U3300 ( .A1(n3910), .A2(net644778), .B1(n3909), .B2(net644746), 
        .ZN(n5805) );
  AOI22_X1 U3299 ( .A1(n3908), .A2(net644908), .B1(n3907), .B2(net644425), 
        .ZN(n5806) );
  AOI22_X1 U3297 ( .A1(n3906), .A2(n3974), .B1(n3905), .B2(n463), .ZN(n5807)
         );
  NAND4_X1 U3296 ( .A1(n5804), .A2(n5805), .A3(n5806), .A4(n5807), .ZN(n5803)
         );
  OAI21_X1 U3295 ( .B1(n5802), .B2(n5803), .A(n6370), .ZN(n5801) );
  OAI211_X1 U3294 ( .C1(n571), .C2(n5220), .A(n5800), .B(n5801), .ZN(n5797) );
  AOI22_X1 U3292 ( .A1(n6373), .A2(net644809), .B1(n6372), .B2(n4083), .ZN(
        n5799) );
  OAI21_X1 U3291 ( .B1(n633), .B2(n5216), .A(n5799), .ZN(n5798) );
  AOI211_X1 U3290 ( .C1(n6374), .C2(net644714), .A(n5797), .B(n5798), .ZN(
        n5796) );
  NAND4_X1 U3289 ( .A1(n5793), .A2(n5794), .A3(n5795), .A4(n5796), .ZN(n2702)
         );
  AOI22_X1 U2836 ( .A1(n6356), .A2(n3940), .B1(n6355), .B2(n4026), .ZN(n5441)
         );
  AOI22_X1 U2835 ( .A1(n6358), .A2(net644891), .B1(n6357), .B2(net644857), 
        .ZN(n5442) );
  AOI22_X1 U2834 ( .A1(n6360), .A2(net644473), .B1(n6359), .B2(DATAIN[22]), 
        .ZN(n5462) );
  OAI21_X1 U2833 ( .B1(n5257), .B2(net644378), .A(n5462), .ZN(n5460) );
  OAI22_X1 U2832 ( .A1(n524), .A2(n5255), .B1(n649), .B2(n5256), .ZN(n5461) );
  AOI211_X1 U2831 ( .C1(n6361), .C2(net644665), .A(n5460), .B(n5461), .ZN(
        n5443) );
  AOI22_X1 U2830 ( .A1(n6363), .A2(net644537), .B1(n6362), .B2(net644569), 
        .ZN(n5448) );
  AOI22_X1 U2828 ( .A1(n6365), .A2(n414), .B1(n6364), .B2(n4134), .ZN(n5456)
         );
  AOI22_X1 U2827 ( .A1(n3911), .A2(net644634), .B1(n3912), .B2(net644505), 
        .ZN(n5457) );
  AOI22_X1 U2825 ( .A1(n6367), .A2(n4027), .B1(n6366), .B2(n362), .ZN(n5458)
         );
  AOI22_X1 U2824 ( .A1(n3913), .A2(net644602), .B1(n3914), .B2(net644698), 
        .ZN(n5459) );
  NAND4_X1 U2823 ( .A1(n5456), .A2(n5457), .A3(n5458), .A4(n5459), .ZN(n5450)
         );
  AOI22_X1 U2821 ( .A1(n6369), .A2(n416), .B1(n6368), .B2(n4135), .ZN(n5452)
         );
  AOI22_X1 U2820 ( .A1(n3910), .A2(net644794), .B1(n3909), .B2(net644762), 
        .ZN(n5453) );
  AOI22_X1 U2819 ( .A1(n3908), .A2(net644924), .B1(n3907), .B2(net644441), 
        .ZN(n5454) );
  AOI22_X1 U2817 ( .A1(n3906), .A2(n4028), .B1(n3905), .B2(n415), .ZN(n5455)
         );
  NAND4_X1 U2816 ( .A1(n5452), .A2(n5453), .A3(n5454), .A4(n5455), .ZN(n5451)
         );
  OAI21_X1 U2815 ( .B1(n5450), .B2(n5451), .A(n6370), .ZN(n5449) );
  OAI211_X1 U2814 ( .C1(n555), .C2(n5220), .A(n5448), .B(n5449), .ZN(n5445) );
  AOI22_X1 U2812 ( .A1(n6373), .A2(net644825), .B1(n6372), .B2(n4136), .ZN(
        n5447) );
  OAI21_X1 U2811 ( .B1(n617), .B2(n5216), .A(n5447), .ZN(n5446) );
  AOI211_X1 U2810 ( .C1(n6374), .C2(net644730), .A(n5445), .B(n5446), .ZN(
        n5444) );
  NAND4_X1 U2809 ( .A1(n5441), .A2(n5442), .A3(n5443), .A4(n5444), .ZN(n2718)
         );
  AOI22_X1 U2686 ( .A1(n6356), .A2(n3945), .B1(n5264), .B2(n4044), .ZN(n5331)
         );
  AOI22_X1 U2685 ( .A1(n5261), .A2(net644896), .B1(n5262), .B2(net644862), 
        .ZN(n5332) );
  AOI22_X1 U2684 ( .A1(n5259), .A2(net644478), .B1(n5260), .B2(DATAIN[27]), 
        .ZN(n5352) );
  OAI21_X1 U2683 ( .B1(n5257), .B2(net644383), .A(n5352), .ZN(n5350) );
  OAI22_X1 U2682 ( .A1(n519), .A2(n5255), .B1(n644), .B2(n5256), .ZN(n5351) );
  AOI211_X1 U2681 ( .C1(n6361), .C2(net644670), .A(n5350), .B(n5351), .ZN(
        n5333) );
  AOI22_X1 U2680 ( .A1(n5250), .A2(net644542), .B1(n5251), .B2(net644574), 
        .ZN(n5338) );
  AOI22_X1 U2678 ( .A1(n5248), .A2(n399), .B1(n5249), .B2(n4152), .ZN(n5346)
         );
  AOI22_X1 U2677 ( .A1(n3911), .A2(net644639), .B1(n3912), .B2(net644510), 
        .ZN(n5347) );
  AOI22_X1 U2675 ( .A1(n6367), .A2(n4045), .B1(n5245), .B2(n357), .ZN(n5348)
         );
  AOI22_X1 U2674 ( .A1(n3913), .A2(net644607), .B1(n3914), .B2(net644703), 
        .ZN(n5349) );
  NAND4_X1 U2673 ( .A1(n5346), .A2(n5347), .A3(n5348), .A4(n5349), .ZN(n5340)
         );
  AOI22_X1 U2671 ( .A1(n6369), .A2(n401), .B1(n5237), .B2(n4153), .ZN(n5342)
         );
  AOI22_X1 U2670 ( .A1(n3910), .A2(net644799), .B1(n3909), .B2(net644767), 
        .ZN(n5343) );
  AOI22_X1 U2669 ( .A1(n3908), .A2(net644929), .B1(n3907), .B2(net644446), 
        .ZN(n5344) );
  AOI22_X1 U2667 ( .A1(n3906), .A2(n4046), .B1(n3905), .B2(n400), .ZN(n5345)
         );
  NAND4_X1 U2666 ( .A1(n5342), .A2(n5343), .A3(n5344), .A4(n5345), .ZN(n5341)
         );
  OAI21_X1 U2665 ( .B1(n5340), .B2(n5341), .A(n6370), .ZN(n5339) );
  OAI211_X1 U2664 ( .C1(n550), .C2(n5220), .A(n5338), .B(n5339), .ZN(n5335) );
  AOI22_X1 U2662 ( .A1(n6373), .A2(net644830), .B1(n6372), .B2(n4154), .ZN(
        n5337) );
  OAI21_X1 U2661 ( .B1(n612), .B2(n5216), .A(n5337), .ZN(n5336) );
  AOI211_X1 U2660 ( .C1(n5213), .C2(net644735), .A(n5335), .B(n5336), .ZN(
        n5334) );
  NAND4_X1 U2659 ( .A1(n5331), .A2(n5332), .A3(n5333), .A4(n5334), .ZN(n2723)
         );
  AOI22_X1 U2806 ( .A1(n6356), .A2(n3941), .B1(n6355), .B2(n4029), .ZN(n5419)
         );
  AOI22_X1 U2805 ( .A1(n6358), .A2(net644892), .B1(n6357), .B2(net644858), 
        .ZN(n5420) );
  AOI22_X1 U2804 ( .A1(n5259), .A2(net644474), .B1(n6359), .B2(DATAIN[23]), 
        .ZN(n5440) );
  OAI21_X1 U2803 ( .B1(n5257), .B2(net644379), .A(n5440), .ZN(n5438) );
  OAI22_X1 U2802 ( .A1(n523), .A2(n5255), .B1(n648), .B2(n5256), .ZN(n5439) );
  AOI211_X1 U2801 ( .C1(n6361), .C2(net644666), .A(n5438), .B(n5439), .ZN(
        n5421) );
  AOI22_X1 U2800 ( .A1(n5250), .A2(net644538), .B1(n5251), .B2(net644570), 
        .ZN(n5426) );
  AOI22_X1 U2798 ( .A1(n6365), .A2(n411), .B1(n6364), .B2(n4137), .ZN(n5434)
         );
  AOI22_X1 U2797 ( .A1(n3911), .A2(net644635), .B1(n3912), .B2(net644506), 
        .ZN(n5435) );
  AOI22_X1 U2795 ( .A1(n6367), .A2(n4030), .B1(n6366), .B2(n361), .ZN(n5436)
         );
  AOI22_X1 U2794 ( .A1(n3913), .A2(net644603), .B1(n3914), .B2(net644699), 
        .ZN(n5437) );
  NAND4_X1 U2793 ( .A1(n5434), .A2(n5435), .A3(n5436), .A4(n5437), .ZN(n5428)
         );
  AOI22_X1 U2791 ( .A1(n6369), .A2(n413), .B1(n6368), .B2(n4138), .ZN(n5430)
         );
  AOI22_X1 U2790 ( .A1(n3910), .A2(net644795), .B1(n3909), .B2(net644763), 
        .ZN(n5431) );
  AOI22_X1 U2789 ( .A1(n3908), .A2(net644925), .B1(n3907), .B2(net644442), 
        .ZN(n5432) );
  AOI22_X1 U2787 ( .A1(n3906), .A2(n4031), .B1(n3905), .B2(n412), .ZN(n5433)
         );
  NAND4_X1 U2786 ( .A1(n5430), .A2(n5431), .A3(n5432), .A4(n5433), .ZN(n5429)
         );
  OAI21_X1 U2785 ( .B1(n5428), .B2(n5429), .A(n6370), .ZN(n5427) );
  OAI211_X1 U2784 ( .C1(n554), .C2(n5220), .A(n5426), .B(n5427), .ZN(n5423) );
  AOI22_X1 U2782 ( .A1(n6373), .A2(net644826), .B1(n6372), .B2(n4139), .ZN(
        n5425) );
  OAI21_X1 U2781 ( .B1(n616), .B2(n5216), .A(n5425), .ZN(n5424) );
  AOI211_X1 U2780 ( .C1(n6374), .C2(net644731), .A(n5423), .B(n5424), .ZN(
        n5422) );
  NAND4_X1 U2779 ( .A1(n5419), .A2(n5420), .A3(n5421), .A4(n5422), .ZN(n2719)
         );
  AOI22_X1 U1691 ( .A1(n4241), .A2(n4053), .B1(n6375), .B2(n3948), .ZN(n4246)
         );
  AOI22_X1 U1690 ( .A1(net644899), .A2(n4239), .B1(net644865), .B2(n4240), 
        .ZN(n4247) );
  AOI22_X1 U1689 ( .A1(net644481), .A2(n6380), .B1(DATAIN[30]), .B2(n6379), 
        .ZN(n4272) );
  OAI21_X1 U1688 ( .B1(n4235), .B2(net644417), .A(n4272), .ZN(n4270) );
  OAI22_X1 U1687 ( .A1(n641), .A2(n4233), .B1(n516), .B2(n4234), .ZN(n4271) );
  AOI211_X1 U1686 ( .C1(net644673), .C2(n6381), .A(n4270), .B(n4271), .ZN(
        n4248) );
  AOI22_X1 U1685 ( .A1(net644577), .A2(n6382), .B1(net644545), .B2(n3880), 
        .ZN(n4254) );
  AOI22_X1 U1684 ( .A1(n390), .A2(n6383), .B1(n3896), .B2(n4161), .ZN(n4264)
         );
  AOI22_X1 U1683 ( .A1(net644642), .A2(n3895), .B1(net644513), .B2(n3894), 
        .ZN(n4265) );
  AOI22_X1 U1682 ( .A1(n4220), .A2(n354), .B1(n3891), .B2(n4054), .ZN(n4266)
         );
  AOI22_X1 U1681 ( .A1(net644610), .A2(n3890), .B1(net644706), .B2(n3897), 
        .ZN(n4267) );
  NAND4_X1 U1680 ( .A1(n4264), .A2(n4265), .A3(n4266), .A4(n4267), .ZN(n4256)
         );
  AOI22_X1 U1679 ( .A1(n392), .A2(n3904), .B1(n3903), .B2(n4162), .ZN(n4258)
         );
  AOI22_X1 U1678 ( .A1(net644802), .A2(n3902), .B1(net644770), .B2(n3901), 
        .ZN(n4259) );
  AOI22_X1 U1677 ( .A1(net644932), .A2(n3900), .B1(net644449), .B2(n3899), 
        .ZN(n4260) );
  AOI22_X1 U1676 ( .A1(n4204), .A2(n391), .B1(n3898), .B2(n4055), .ZN(n4261)
         );
  NAND4_X1 U1675 ( .A1(n4258), .A2(n4259), .A3(n4260), .A4(n4261), .ZN(n4257)
         );
  OAI21_X1 U1674 ( .B1(n4256), .B2(n4257), .A(n6386), .ZN(n4255) );
  OAI211_X1 U1673 ( .C1(n547), .C2(n4194), .A(n4254), .B(n4255), .ZN(n4250) );
  AOI22_X1 U1672 ( .A1(net644833), .A2(n6389), .B1(n6388), .B2(n4163), .ZN(
        n4252) );
  OAI21_X1 U1671 ( .B1(n609), .B2(n4189), .A(n4252), .ZN(n4251) );
  AOI211_X1 U1670 ( .C1(net644738), .C2(n6390), .A(n4250), .B(n4251), .ZN(
        n4249) );
  NAND4_X1 U1669 ( .A1(n4246), .A2(n4247), .A3(n4248), .A4(n4249), .ZN(n2788)
         );
  AOI22_X1 U1743 ( .A1(n4241), .A2(n4047), .B1(n4243), .B2(n3946), .ZN(n4306)
         );
  AOI22_X1 U1742 ( .A1(net644897), .A2(n6378), .B1(net644863), .B2(n4240), 
        .ZN(n4307) );
  AOI22_X1 U1741 ( .A1(net644479), .A2(n6380), .B1(DATAIN[28]), .B2(n6379), 
        .ZN(n4332) );
  OAI21_X1 U1740 ( .B1(n4235), .B2(net644415), .A(n4332), .ZN(n4330) );
  OAI22_X1 U1739 ( .A1(n643), .A2(n4233), .B1(n518), .B2(n4234), .ZN(n4331) );
  AOI211_X1 U1738 ( .C1(net644671), .C2(n6381), .A(n4330), .B(n4331), .ZN(
        n4308) );
  AOI22_X1 U1737 ( .A1(net644575), .A2(n6382), .B1(net644543), .B2(n3880), 
        .ZN(n4314) );
  AOI22_X1 U1736 ( .A1(n396), .A2(n6383), .B1(n3896), .B2(n4155), .ZN(n4324)
         );
  AOI22_X1 U1735 ( .A1(net644640), .A2(n3895), .B1(net644511), .B2(n3894), 
        .ZN(n4325) );
  AOI22_X1 U1734 ( .A1(n4220), .A2(n356), .B1(n4221), .B2(n4048), .ZN(n4326)
         );
  AOI22_X1 U1733 ( .A1(net644608), .A2(n3890), .B1(net644704), .B2(n3897), 
        .ZN(n4327) );
  NAND4_X1 U1732 ( .A1(n4324), .A2(n4325), .A3(n4326), .A4(n4327), .ZN(n4316)
         );
  AOI22_X1 U1731 ( .A1(n398), .A2(n3904), .B1(n4212), .B2(n4156), .ZN(n4318)
         );
  AOI22_X1 U1730 ( .A1(net644800), .A2(n3902), .B1(net644768), .B2(n3901), 
        .ZN(n4319) );
  AOI22_X1 U1729 ( .A1(net644930), .A2(n3900), .B1(net644447), .B2(n3899), 
        .ZN(n4320) );
  AOI22_X1 U1728 ( .A1(n4204), .A2(n397), .B1(n3898), .B2(n4049), .ZN(n4321)
         );
  NAND4_X1 U1727 ( .A1(n4318), .A2(n4319), .A3(n4320), .A4(n4321), .ZN(n4317)
         );
  OAI21_X1 U1726 ( .B1(n4316), .B2(n4317), .A(n6386), .ZN(n4315) );
  OAI211_X1 U1725 ( .C1(n549), .C2(n4194), .A(n4314), .B(n4315), .ZN(n4310) );
  AOI22_X1 U1724 ( .A1(net644831), .A2(n6389), .B1(n4192), .B2(n4157), .ZN(
        n4312) );
  OAI21_X1 U1723 ( .B1(n611), .B2(n4189), .A(n4312), .ZN(n4311) );
  AOI211_X1 U1722 ( .C1(net644736), .C2(n6390), .A(n4310), .B(n4311), .ZN(
        n4309) );
  NAND4_X1 U1721 ( .A1(n4306), .A2(n4307), .A3(n4308), .A4(n4309), .ZN(n2784)
         );
  AOI22_X1 U1665 ( .A1(n4241), .A2(n4056), .B1(n4243), .B2(n3949), .ZN(n4182)
         );
  AOI22_X1 U1664 ( .A1(net644900), .A2(n4239), .B1(net644866), .B2(n4240), 
        .ZN(n4183) );
  AOI22_X1 U1663 ( .A1(net644482), .A2(n6380), .B1(DATAIN[31]), .B2(n6379), 
        .ZN(n4236) );
  OAI21_X1 U1662 ( .B1(n4235), .B2(net644418), .A(n4236), .ZN(n4231) );
  OAI22_X1 U1661 ( .A1(n640), .A2(n4233), .B1(n515), .B2(n4234), .ZN(n4232) );
  AOI211_X1 U1660 ( .C1(net644674), .C2(n6381), .A(n4231), .B(n4232), .ZN(
        n4184) );
  AOI22_X1 U1659 ( .A1(net644578), .A2(n4228), .B1(net644546), .B2(n3880), 
        .ZN(n4195) );
  AOI22_X1 U1658 ( .A1(n387), .A2(n6383), .B1(n3896), .B2(n4164), .ZN(n4214)
         );
  AOI22_X1 U1657 ( .A1(net644643), .A2(n3895), .B1(net644514), .B2(n3894), 
        .ZN(n4215) );
  AOI22_X1 U1656 ( .A1(n4220), .A2(n353), .B1(n3891), .B2(n4057), .ZN(n4216)
         );
  AOI22_X1 U1655 ( .A1(net644611), .A2(n3890), .B1(net644707), .B2(n3897), 
        .ZN(n4217) );
  NAND4_X1 U1654 ( .A1(n4214), .A2(n4215), .A3(n4216), .A4(n4217), .ZN(n4197)
         );
  AOI22_X1 U1653 ( .A1(n389), .A2(n3904), .B1(n3903), .B2(n4165), .ZN(n4200)
         );
  AOI22_X1 U1652 ( .A1(net644803), .A2(n3902), .B1(net644771), .B2(n3901), 
        .ZN(n4201) );
  AOI22_X1 U1651 ( .A1(net644933), .A2(n3900), .B1(net644450), .B2(n3899), 
        .ZN(n4202) );
  AOI22_X1 U1650 ( .A1(n6385), .A2(n388), .B1(n3898), .B2(n4058), .ZN(n4203)
         );
  NAND4_X1 U1649 ( .A1(n4200), .A2(n4201), .A3(n4202), .A4(n4203), .ZN(n4198)
         );
  OAI21_X1 U1648 ( .B1(n4197), .B2(n4198), .A(n6386), .ZN(n4196) );
  OAI211_X1 U1647 ( .C1(n546), .C2(n4194), .A(n4195), .B(n4196), .ZN(n4187) );
  AOI22_X1 U1646 ( .A1(net644834), .A2(n6389), .B1(n4192), .B2(n4166), .ZN(
        n4190) );
  OAI21_X1 U1645 ( .B1(n608), .B2(n4189), .A(n4190), .ZN(n4188) );
  AOI211_X1 U1644 ( .C1(net644739), .C2(n6390), .A(n4187), .B(n4188), .ZN(
        n4185) );
  NAND4_X1 U1643 ( .A1(n4182), .A2(n4183), .A3(n4184), .A4(n4185), .ZN(n2790)
         );
  AOI22_X1 U1717 ( .A1(n4241), .A2(n4050), .B1(n6375), .B2(n3947), .ZN(n4276)
         );
  AOI22_X1 U1716 ( .A1(net644898), .A2(n6378), .B1(net644864), .B2(n4240), 
        .ZN(n4277) );
  AOI22_X1 U1715 ( .A1(net644480), .A2(n6380), .B1(DATAIN[29]), .B2(n6379), 
        .ZN(n4302) );
  OAI21_X1 U1714 ( .B1(n4235), .B2(net644416), .A(n4302), .ZN(n4300) );
  OAI22_X1 U1713 ( .A1(n642), .A2(n4233), .B1(n517), .B2(n4234), .ZN(n4301) );
  AOI211_X1 U1712 ( .C1(net644672), .C2(n6381), .A(n4300), .B(n4301), .ZN(
        n4278) );
  AOI22_X1 U1711 ( .A1(net644576), .A2(n6382), .B1(net644544), .B2(n3880), 
        .ZN(n4284) );
  AOI22_X1 U1710 ( .A1(n393), .A2(n6383), .B1(n3896), .B2(n4158), .ZN(n4294)
         );
  AOI22_X1 U1709 ( .A1(net644641), .A2(n3895), .B1(net644512), .B2(n3894), 
        .ZN(n4295) );
  AOI22_X1 U1708 ( .A1(n4220), .A2(n355), .B1(n4221), .B2(n4051), .ZN(n4296)
         );
  AOI22_X1 U1707 ( .A1(net644609), .A2(n3890), .B1(net644705), .B2(n3897), 
        .ZN(n4297) );
  NAND4_X1 U1706 ( .A1(n4294), .A2(n4295), .A3(n4296), .A4(n4297), .ZN(n4286)
         );
  AOI22_X1 U1705 ( .A1(n395), .A2(n3904), .B1(n4212), .B2(n4159), .ZN(n4288)
         );
  AOI22_X1 U1704 ( .A1(net644801), .A2(n3902), .B1(net644769), .B2(n3901), 
        .ZN(n4289) );
  AOI22_X1 U1703 ( .A1(net644931), .A2(n3900), .B1(net644448), .B2(n3899), 
        .ZN(n4290) );
  AOI22_X1 U1702 ( .A1(n6385), .A2(n394), .B1(n3898), .B2(n4052), .ZN(n4291)
         );
  NAND4_X1 U1701 ( .A1(n4288), .A2(n4289), .A3(n4290), .A4(n4291), .ZN(n4287)
         );
  OAI21_X1 U1700 ( .B1(n4286), .B2(n4287), .A(n6386), .ZN(n4285) );
  OAI211_X1 U1699 ( .C1(n548), .C2(n4194), .A(n4284), .B(n4285), .ZN(n4280) );
  AOI22_X1 U1698 ( .A1(net644832), .A2(n6389), .B1(n6388), .B2(n4160), .ZN(
        n4282) );
  OAI21_X1 U1697 ( .B1(n610), .B2(n4189), .A(n4282), .ZN(n4281) );
  AOI211_X1 U1696 ( .C1(net644737), .C2(n6390), .A(n4280), .B(n4281), .ZN(
        n4279) );
  NAND4_X1 U1695 ( .A1(n4276), .A2(n4277), .A3(n4278), .A4(n4279), .ZN(n2786)
         );
  AOI22_X1 U1821 ( .A1(n4241), .A2(n4038), .B1(n6375), .B2(n3943), .ZN(n4396)
         );
  AOI22_X1 U1820 ( .A1(net644894), .A2(n4239), .B1(net644860), .B2(n4240), 
        .ZN(n4397) );
  AOI22_X1 U1819 ( .A1(net644476), .A2(n6380), .B1(DATAIN[25]), .B2(n6379), 
        .ZN(n4422) );
  OAI21_X1 U1818 ( .B1(n4235), .B2(net644412), .A(n4422), .ZN(n4420) );
  OAI22_X1 U1817 ( .A1(n646), .A2(n4233), .B1(n521), .B2(n4234), .ZN(n4421) );
  AOI211_X1 U1816 ( .C1(net644668), .C2(n6381), .A(n4420), .B(n4421), .ZN(
        n4398) );
  AOI22_X1 U1815 ( .A1(net644572), .A2(n6382), .B1(net644540), .B2(n3880), 
        .ZN(n4404) );
  AOI22_X1 U1814 ( .A1(n405), .A2(n6383), .B1(n3896), .B2(n4144), .ZN(n4414)
         );
  AOI22_X1 U1813 ( .A1(net644637), .A2(n3895), .B1(net644508), .B2(n3894), 
        .ZN(n4415) );
  AOI22_X1 U1812 ( .A1(n4220), .A2(n359), .B1(n4221), .B2(n4039), .ZN(n4416)
         );
  AOI22_X1 U1811 ( .A1(net644605), .A2(n3890), .B1(net644701), .B2(n3897), 
        .ZN(n4417) );
  NAND4_X1 U1810 ( .A1(n4414), .A2(n4415), .A3(n4416), .A4(n4417), .ZN(n4406)
         );
  AOI22_X1 U1809 ( .A1(n407), .A2(n3904), .B1(n4212), .B2(n4147), .ZN(n4408)
         );
  AOI22_X1 U1808 ( .A1(net644797), .A2(n3902), .B1(net644765), .B2(n3901), 
        .ZN(n4409) );
  AOI22_X1 U1807 ( .A1(net644927), .A2(n3900), .B1(net644444), .B2(n3899), 
        .ZN(n4410) );
  AOI22_X1 U1806 ( .A1(n6385), .A2(n406), .B1(n3898), .B2(n4040), .ZN(n4411)
         );
  NAND4_X1 U1805 ( .A1(n4408), .A2(n4409), .A3(n4410), .A4(n4411), .ZN(n4407)
         );
  OAI21_X1 U1804 ( .B1(n4406), .B2(n4407), .A(n6386), .ZN(n4405) );
  OAI211_X1 U1803 ( .C1(n552), .C2(n4194), .A(n4404), .B(n4405), .ZN(n4400) );
  AOI22_X1 U1802 ( .A1(net644828), .A2(n6389), .B1(n4192), .B2(n4148), .ZN(
        n4402) );
  OAI21_X1 U1801 ( .B1(n614), .B2(n4189), .A(n4402), .ZN(n4401) );
  AOI211_X1 U1800 ( .C1(net644733), .C2(n6390), .A(n4400), .B(n4401), .ZN(
        n4399) );
  NAND4_X1 U1799 ( .A1(n4396), .A2(n4397), .A3(n4398), .A4(n4399), .ZN(n2778)
         );
  AOI22_X1 U2341 ( .A1(n6376), .A2(n3969), .B1(n6375), .B2(n3920), .ZN(n4996)
         );
  AOI22_X1 U2340 ( .A1(net644874), .A2(n6378), .B1(net644840), .B2(n6377), 
        .ZN(n4997) );
  AOI22_X1 U2339 ( .A1(net644456), .A2(n6380), .B1(DATAIN[5]), .B2(n6379), 
        .ZN(n5022) );
  OAI21_X1 U2338 ( .B1(n4235), .B2(net644392), .A(n5022), .ZN(n5020) );
  OAI22_X1 U2337 ( .A1(n666), .A2(n4233), .B1(n541), .B2(n4234), .ZN(n5021) );
  AOI211_X1 U2336 ( .C1(net644648), .C2(n6381), .A(n5020), .B(n5021), .ZN(
        n4998) );
  AOI22_X1 U2335 ( .A1(net644552), .A2(n6382), .B1(net644520), .B2(n3880), 
        .ZN(n5004) );
  AOI22_X1 U2334 ( .A1(n465), .A2(n4225), .B1(n3896), .B2(n4078), .ZN(n5014)
         );
  AOI22_X1 U2333 ( .A1(net644617), .A2(n3895), .B1(net644488), .B2(n3894), 
        .ZN(n5015) );
  AOI22_X1 U2332 ( .A1(n6384), .A2(n379), .B1(n3891), .B2(n3970), .ZN(n5016)
         );
  AOI22_X1 U2331 ( .A1(net644585), .A2(n3890), .B1(net644681), .B2(n3897), 
        .ZN(n5017) );
  NAND4_X1 U2330 ( .A1(n5014), .A2(n5015), .A3(n5016), .A4(n5017), .ZN(n5006)
         );
  AOI22_X1 U2329 ( .A1(n467), .A2(n3904), .B1(n3903), .B2(n4079), .ZN(n5008)
         );
  AOI22_X1 U2328 ( .A1(net644777), .A2(n3902), .B1(net644745), .B2(n3901), 
        .ZN(n5009) );
  AOI22_X1 U2327 ( .A1(net644907), .A2(n3900), .B1(net644424), .B2(n3899), 
        .ZN(n5010) );
  AOI22_X1 U2326 ( .A1(n6385), .A2(n466), .B1(n3898), .B2(n3971), .ZN(n5011)
         );
  NAND4_X1 U2325 ( .A1(n5008), .A2(n5009), .A3(n5010), .A4(n5011), .ZN(n5007)
         );
  OAI21_X1 U2324 ( .B1(n5006), .B2(n5007), .A(n6386), .ZN(n5005) );
  OAI211_X1 U2323 ( .C1(n572), .C2(n4194), .A(n5004), .B(n5005), .ZN(n5000) );
  AOI22_X1 U2322 ( .A1(net644808), .A2(n6389), .B1(n6388), .B2(n4080), .ZN(
        n5002) );
  OAI21_X1 U2321 ( .B1(n634), .B2(n4189), .A(n5002), .ZN(n5001) );
  AOI211_X1 U2320 ( .C1(net644713), .C2(n6390), .A(n5000), .B(n5001), .ZN(
        n4999) );
  NAND4_X1 U2319 ( .A1(n4996), .A2(n4997), .A3(n4998), .A4(n4999), .ZN(n2738)
         );
  AOI22_X1 U2185 ( .A1(n6376), .A2(n3987), .B1(n6375), .B2(n3929), .ZN(n4816)
         );
  AOI22_X1 U2184 ( .A1(net644880), .A2(n6378), .B1(net644846), .B2(n6377), 
        .ZN(n4817) );
  AOI22_X1 U2183 ( .A1(net644462), .A2(n4237), .B1(DATAIN[11]), .B2(n4238), 
        .ZN(n4842) );
  OAI21_X1 U2182 ( .B1(n4235), .B2(net644398), .A(n4842), .ZN(n4840) );
  OAI22_X1 U2181 ( .A1(n660), .A2(n4233), .B1(n535), .B2(n4234), .ZN(n4841) );
  AOI211_X1 U2180 ( .C1(net644654), .C2(n6381), .A(n4840), .B(n4841), .ZN(
        n4818) );
  AOI22_X1 U2179 ( .A1(net644558), .A2(n6382), .B1(net644526), .B2(n3880), 
        .ZN(n4824) );
  AOI22_X1 U2178 ( .A1(n447), .A2(n6383), .B1(n3896), .B2(n4096), .ZN(n4834)
         );
  AOI22_X1 U2177 ( .A1(net644623), .A2(n3895), .B1(net644494), .B2(n3894), 
        .ZN(n4835) );
  AOI22_X1 U2176 ( .A1(n6384), .A2(n373), .B1(n3891), .B2(n3988), .ZN(n4836)
         );
  AOI22_X1 U2175 ( .A1(net644591), .A2(n3890), .B1(net644687), .B2(n4219), 
        .ZN(n4837) );
  NAND4_X1 U2174 ( .A1(n4834), .A2(n4835), .A3(n4836), .A4(n4837), .ZN(n4826)
         );
  AOI22_X1 U2173 ( .A1(n449), .A2(n3904), .B1(n3903), .B2(n4097), .ZN(n4828)
         );
  AOI22_X1 U2172 ( .A1(net644783), .A2(n3902), .B1(net644751), .B2(n3901), 
        .ZN(n4829) );
  AOI22_X1 U2171 ( .A1(net644913), .A2(n3900), .B1(net644430), .B2(n3899), 
        .ZN(n4830) );
  AOI22_X1 U2170 ( .A1(n6385), .A2(n448), .B1(n3898), .B2(n3989), .ZN(n4831)
         );
  NAND4_X1 U2169 ( .A1(n4828), .A2(n4829), .A3(n4830), .A4(n4831), .ZN(n4827)
         );
  OAI21_X1 U2168 ( .B1(n4826), .B2(n4827), .A(n6386), .ZN(n4825) );
  OAI211_X1 U2167 ( .C1(n566), .C2(n4194), .A(n4824), .B(n4825), .ZN(n4820) );
  AOI22_X1 U2166 ( .A1(net644814), .A2(n6389), .B1(n6388), .B2(n4098), .ZN(
        n4822) );
  OAI21_X1 U2165 ( .B1(n628), .B2(n4189), .A(n4822), .ZN(n4821) );
  AOI211_X1 U2164 ( .C1(net644719), .C2(n4186), .A(n4820), .B(n4821), .ZN(
        n4819) );
  NAND4_X1 U2163 ( .A1(n4816), .A2(n4817), .A3(n4818), .A4(n4819), .ZN(n2750)
         );
  AOI22_X1 U2159 ( .A1(n6376), .A2(n3990), .B1(n6375), .B2(n3930), .ZN(n4786)
         );
  AOI22_X1 U2158 ( .A1(net644881), .A2(n6378), .B1(net644847), .B2(n6377), 
        .ZN(n4787) );
  AOI22_X1 U2157 ( .A1(net644463), .A2(n6380), .B1(DATAIN[12]), .B2(n6379), 
        .ZN(n4812) );
  OAI21_X1 U2156 ( .B1(n4235), .B2(net644399), .A(n4812), .ZN(n4810) );
  OAI22_X1 U2155 ( .A1(n659), .A2(n4233), .B1(n534), .B2(n4234), .ZN(n4811) );
  AOI211_X1 U2154 ( .C1(net644655), .C2(n6381), .A(n4810), .B(n4811), .ZN(
        n4788) );
  AOI22_X1 U2153 ( .A1(net644559), .A2(n6382), .B1(net644527), .B2(n4229), 
        .ZN(n4794) );
  AOI22_X1 U2152 ( .A1(n444), .A2(n4225), .B1(n3896), .B2(n4099), .ZN(n4804)
         );
  AOI22_X1 U2151 ( .A1(net644624), .A2(n3895), .B1(net644495), .B2(n4224), 
        .ZN(n4805) );
  AOI22_X1 U2150 ( .A1(n6384), .A2(n372), .B1(n3891), .B2(n3991), .ZN(n4806)
         );
  AOI22_X1 U2149 ( .A1(net644592), .A2(n4218), .B1(net644688), .B2(n3897), 
        .ZN(n4807) );
  NAND4_X1 U2148 ( .A1(n4804), .A2(n4805), .A3(n4806), .A4(n4807), .ZN(n4796)
         );
  AOI22_X1 U2147 ( .A1(n446), .A2(n3904), .B1(n3903), .B2(n4100), .ZN(n4798)
         );
  AOI22_X1 U2146 ( .A1(net644784), .A2(n3902), .B1(net644752), .B2(n4210), 
        .ZN(n4799) );
  AOI22_X1 U2145 ( .A1(net644914), .A2(n3900), .B1(net644431), .B2(n4208), 
        .ZN(n4800) );
  AOI22_X1 U2144 ( .A1(n6385), .A2(n445), .B1(n3898), .B2(n3992), .ZN(n4801)
         );
  NAND4_X1 U2143 ( .A1(n4798), .A2(n4799), .A3(n4800), .A4(n4801), .ZN(n4797)
         );
  OAI21_X1 U2142 ( .B1(n4796), .B2(n4797), .A(n4199), .ZN(n4795) );
  OAI211_X1 U2141 ( .C1(n565), .C2(n4194), .A(n4794), .B(n4795), .ZN(n4790) );
  AOI22_X1 U2140 ( .A1(net644815), .A2(n6389), .B1(n6388), .B2(n4101), .ZN(
        n4792) );
  OAI21_X1 U2139 ( .B1(n627), .B2(n4189), .A(n4792), .ZN(n4791) );
  AOI211_X1 U2138 ( .C1(net644720), .C2(n6390), .A(n4790), .B(n4791), .ZN(
        n4789) );
  NAND4_X1 U2137 ( .A1(n4786), .A2(n4787), .A3(n4788), .A4(n4789), .ZN(n2752)
         );
  AOI22_X1 U2447 ( .A1(n4241), .A2(n3954), .B1(n6375), .B2(n3916), .ZN(n5116)
         );
  AOI22_X1 U2446 ( .A1(net644870), .A2(n6378), .B1(net644836), .B2(n6377), 
        .ZN(n5117) );
  AOI22_X1 U2445 ( .A1(net644452), .A2(n4237), .B1(DATAIN[1]), .B2(n6379), 
        .ZN(n5143) );
  OAI21_X1 U2444 ( .B1(n4235), .B2(net644388), .A(n5143), .ZN(n5140) );
  OAI22_X1 U2442 ( .A1(n670), .A2(n4233), .B1(n545), .B2(n4234), .ZN(n5141) );
  AOI211_X1 U2441 ( .C1(net644644), .C2(n6381), .A(n5140), .B(n5141), .ZN(
        n5118) );
  AOI22_X1 U2440 ( .A1(net644548), .A2(n6382), .B1(net644516), .B2(n3880), 
        .ZN(n5125) );
  AOI22_X1 U2439 ( .A1(n477), .A2(n4225), .B1(n222), .B2(n3896), .ZN(n5135) );
  AOI22_X1 U2438 ( .A1(net644613), .A2(n3895), .B1(net644484), .B2(n3894), 
        .ZN(n5136) );
  AOI22_X1 U2437 ( .A1(n6384), .A2(n383), .B1(n3891), .B2(n3955), .ZN(n5137)
         );
  AOI22_X1 U2436 ( .A1(net644581), .A2(n3890), .B1(net644677), .B2(n3897), 
        .ZN(n5138) );
  NAND4_X1 U2435 ( .A1(n5135), .A2(n5136), .A3(n5137), .A4(n5138), .ZN(n5127)
         );
  AOI22_X1 U2434 ( .A1(n479), .A2(n3904), .B1(n3903), .B2(n4063), .ZN(n5129)
         );
  AOI22_X1 U2433 ( .A1(net644773), .A2(n3902), .B1(net644741), .B2(n3901), 
        .ZN(n5130) );
  AOI22_X1 U2432 ( .A1(net644903), .A2(n3900), .B1(net644420), .B2(n3899), 
        .ZN(n5131) );
  AOI22_X1 U2431 ( .A1(n6385), .A2(n478), .B1(n3898), .B2(n3956), .ZN(n5132)
         );
  NAND4_X1 U2430 ( .A1(n5129), .A2(n5130), .A3(n5131), .A4(n5132), .ZN(n5128)
         );
  OAI21_X1 U2429 ( .B1(n5127), .B2(n5128), .A(n6386), .ZN(n5126) );
  OAI211_X1 U2428 ( .C1(n576), .C2(n4194), .A(n5125), .B(n5126), .ZN(n5120) );
  AOI22_X1 U2426 ( .A1(net644804), .A2(n6389), .B1(n6388), .B2(n4064), .ZN(
        n5122) );
  OAI21_X1 U2425 ( .B1(n638), .B2(n4189), .A(n5122), .ZN(n5121) );
  AOI211_X1 U2424 ( .C1(net644709), .C2(n4186), .A(n5120), .B(n5121), .ZN(
        n5119) );
  NAND4_X1 U2423 ( .A1(n5116), .A2(n5117), .A3(n5118), .A4(n5119), .ZN(n2730)
         );
  AOI22_X1 U2419 ( .A1(n4241), .A2(n3957), .B1(n6375), .B2(n3917), .ZN(n5086)
         );
  AOI22_X1 U2418 ( .A1(net644871), .A2(n6378), .B1(net644837), .B2(n6377), 
        .ZN(n5087) );
  AOI22_X1 U2417 ( .A1(net644453), .A2(n4237), .B1(DATAIN[2]), .B2(n6379), 
        .ZN(n5112) );
  OAI21_X1 U2416 ( .B1(n4235), .B2(net644389), .A(n5112), .ZN(n5110) );
  OAI22_X1 U2415 ( .A1(n669), .A2(n4233), .B1(n544), .B2(n4234), .ZN(n5111) );
  AOI211_X1 U2414 ( .C1(net644645), .C2(n6381), .A(n5110), .B(n5111), .ZN(
        n5088) );
  AOI22_X1 U2413 ( .A1(net644549), .A2(n4228), .B1(net644517), .B2(n3880), 
        .ZN(n5094) );
  AOI22_X1 U2412 ( .A1(n474), .A2(n4225), .B1(n3896), .B2(n4065), .ZN(n5104)
         );
  AOI22_X1 U2411 ( .A1(net644614), .A2(n3895), .B1(net644485), .B2(n3894), 
        .ZN(n5105) );
  AOI22_X1 U2410 ( .A1(n6384), .A2(n382), .B1(n3891), .B2(n3958), .ZN(n5106)
         );
  AOI22_X1 U2409 ( .A1(net644582), .A2(n3890), .B1(net644678), .B2(n3897), 
        .ZN(n5107) );
  NAND4_X1 U2408 ( .A1(n5104), .A2(n5105), .A3(n5106), .A4(n5107), .ZN(n5096)
         );
  AOI22_X1 U2407 ( .A1(n476), .A2(n3904), .B1(n3903), .B2(n4066), .ZN(n5098)
         );
  AOI22_X1 U2406 ( .A1(net644774), .A2(n3902), .B1(net644742), .B2(n3901), 
        .ZN(n5099) );
  AOI22_X1 U2405 ( .A1(net644904), .A2(n3900), .B1(net644421), .B2(n3899), 
        .ZN(n5100) );
  AOI22_X1 U2404 ( .A1(n6385), .A2(n475), .B1(n3898), .B2(n3960), .ZN(n5101)
         );
  NAND4_X1 U2403 ( .A1(n5098), .A2(n5099), .A3(n5100), .A4(n5101), .ZN(n5097)
         );
  OAI21_X1 U2402 ( .B1(n5096), .B2(n5097), .A(n6386), .ZN(n5095) );
  OAI211_X1 U2401 ( .C1(n575), .C2(n4194), .A(n5094), .B(n5095), .ZN(n5090) );
  AOI22_X1 U2400 ( .A1(net644805), .A2(n6389), .B1(n6388), .B2(n4067), .ZN(
        n5092) );
  OAI21_X1 U2399 ( .B1(n637), .B2(n4189), .A(n5092), .ZN(n5091) );
  AOI211_X1 U2398 ( .C1(net644710), .C2(n4186), .A(n5090), .B(n5091), .ZN(
        n5089) );
  NAND4_X1 U2397 ( .A1(n5086), .A2(n5087), .A3(n5088), .A4(n5089), .ZN(n2732)
         );
  AOI22_X1 U2393 ( .A1(n6376), .A2(n3963), .B1(n6375), .B2(n3918), .ZN(n5056)
         );
  AOI22_X1 U2392 ( .A1(net644872), .A2(n6378), .B1(net644838), .B2(n6377), 
        .ZN(n5057) );
  AOI22_X1 U2391 ( .A1(net644454), .A2(n4237), .B1(DATAIN[3]), .B2(n4238), 
        .ZN(n5082) );
  OAI21_X1 U2390 ( .B1(n4235), .B2(net644390), .A(n5082), .ZN(n5080) );
  OAI22_X1 U2389 ( .A1(n668), .A2(n4233), .B1(n543), .B2(n4234), .ZN(n5081) );
  AOI211_X1 U2388 ( .C1(net644646), .C2(n6381), .A(n5080), .B(n5081), .ZN(
        n5058) );
  AOI22_X1 U2387 ( .A1(net644550), .A2(n6382), .B1(net644518), .B2(n3880), 
        .ZN(n5064) );
  AOI22_X1 U2386 ( .A1(n471), .A2(n6383), .B1(n3896), .B2(n4070), .ZN(n5074)
         );
  AOI22_X1 U2385 ( .A1(net644615), .A2(n3895), .B1(net644486), .B2(n3894), 
        .ZN(n5075) );
  AOI22_X1 U2384 ( .A1(n6384), .A2(n381), .B1(n3891), .B2(n3964), .ZN(n5076)
         );
  AOI22_X1 U2383 ( .A1(net644583), .A2(n3890), .B1(net644679), .B2(n3897), 
        .ZN(n5077) );
  NAND4_X1 U2382 ( .A1(n5074), .A2(n5075), .A3(n5076), .A4(n5077), .ZN(n5066)
         );
  AOI22_X1 U2381 ( .A1(n473), .A2(n3904), .B1(n3903), .B2(n4071), .ZN(n5068)
         );
  AOI22_X1 U2380 ( .A1(net644775), .A2(n3902), .B1(net644743), .B2(n3901), 
        .ZN(n5069) );
  AOI22_X1 U2379 ( .A1(net644905), .A2(n3900), .B1(net644422), .B2(n3899), 
        .ZN(n5070) );
  AOI22_X1 U2378 ( .A1(n6385), .A2(n472), .B1(n3898), .B2(n3965), .ZN(n5071)
         );
  NAND4_X1 U2377 ( .A1(n5068), .A2(n5069), .A3(n5070), .A4(n5071), .ZN(n5067)
         );
  OAI21_X1 U2376 ( .B1(n5066), .B2(n5067), .A(n6386), .ZN(n5065) );
  OAI211_X1 U2375 ( .C1(n574), .C2(n4194), .A(n5064), .B(n5065), .ZN(n5060) );
  AOI22_X1 U2374 ( .A1(net644806), .A2(n6389), .B1(n6388), .B2(n4072), .ZN(
        n5062) );
  OAI21_X1 U2373 ( .B1(n636), .B2(n4189), .A(n5062), .ZN(n5061) );
  AOI211_X1 U2372 ( .C1(net644711), .C2(n6390), .A(n5060), .B(n5061), .ZN(
        n5059) );
  NAND4_X1 U2371 ( .A1(n5056), .A2(n5057), .A3(n5058), .A4(n5059), .ZN(n2734)
         );
  AOI22_X1 U2055 ( .A1(n6376), .A2(n4008), .B1(n6375), .B2(n3934), .ZN(n4666)
         );
  AOI22_X1 U2054 ( .A1(net644885), .A2(n6378), .B1(net644851), .B2(n6377), 
        .ZN(n4667) );
  AOI22_X1 U2053 ( .A1(net644467), .A2(n4237), .B1(DATAIN[16]), .B2(n6379), 
        .ZN(n4692) );
  OAI21_X1 U2052 ( .B1(n4235), .B2(net644403), .A(n4692), .ZN(n4690) );
  OAI22_X1 U2051 ( .A1(n655), .A2(n4233), .B1(n530), .B2(n4234), .ZN(n4691) );
  AOI211_X1 U2050 ( .C1(net644659), .C2(n6381), .A(n4690), .B(n4691), .ZN(
        n4668) );
  AOI22_X1 U2049 ( .A1(net644563), .A2(n6382), .B1(net644531), .B2(n3880), 
        .ZN(n4674) );
  AOI22_X1 U2048 ( .A1(n432), .A2(n6383), .B1(n3896), .B2(n4116), .ZN(n4684)
         );
  AOI22_X1 U2047 ( .A1(net644628), .A2(n3895), .B1(net644499), .B2(n3894), 
        .ZN(n4685) );
  AOI22_X1 U2046 ( .A1(n6384), .A2(n368), .B1(n3891), .B2(n4009), .ZN(n4686)
         );
  AOI22_X1 U2045 ( .A1(net644596), .A2(n3890), .B1(net644692), .B2(n3897), 
        .ZN(n4687) );
  NAND4_X1 U2044 ( .A1(n4684), .A2(n4685), .A3(n4686), .A4(n4687), .ZN(n4676)
         );
  AOI22_X1 U2043 ( .A1(n434), .A2(n3904), .B1(n3903), .B2(n4117), .ZN(n4678)
         );
  AOI22_X1 U2042 ( .A1(net644788), .A2(n3902), .B1(net644756), .B2(n3901), 
        .ZN(n4679) );
  AOI22_X1 U2041 ( .A1(net644918), .A2(n3900), .B1(net644435), .B2(n3899), 
        .ZN(n4680) );
  AOI22_X1 U2040 ( .A1(n6385), .A2(n433), .B1(n3898), .B2(n4010), .ZN(n4681)
         );
  NAND4_X1 U2039 ( .A1(n4678), .A2(n4679), .A3(n4680), .A4(n4681), .ZN(n4677)
         );
  OAI21_X1 U2038 ( .B1(n4676), .B2(n4677), .A(n6386), .ZN(n4675) );
  OAI211_X1 U2037 ( .C1(n561), .C2(n4194), .A(n4674), .B(n4675), .ZN(n4670) );
  AOI22_X1 U2036 ( .A1(net644819), .A2(n6389), .B1(n4192), .B2(n4118), .ZN(
        n4672) );
  OAI21_X1 U2035 ( .B1(n623), .B2(n4189), .A(n4672), .ZN(n4671) );
  AOI211_X1 U2034 ( .C1(net644724), .C2(n4186), .A(n4670), .B(n4671), .ZN(
        n4669) );
  NAND4_X1 U2033 ( .A1(n4666), .A2(n4667), .A3(n4668), .A4(n4669), .ZN(n2760)
         );
  AOI22_X1 U2367 ( .A1(n4241), .A2(n3966), .B1(n6375), .B2(n3919), .ZN(n5026)
         );
  AOI22_X1 U2366 ( .A1(net644873), .A2(n6378), .B1(net644839), .B2(n6377), 
        .ZN(n5027) );
  AOI22_X1 U2365 ( .A1(net644455), .A2(n4237), .B1(DATAIN[4]), .B2(n6379), 
        .ZN(n5052) );
  OAI21_X1 U2364 ( .B1(n4235), .B2(net644391), .A(n5052), .ZN(n5050) );
  OAI22_X1 U2363 ( .A1(n667), .A2(n4233), .B1(n542), .B2(n4234), .ZN(n5051) );
  AOI211_X1 U2362 ( .C1(net644647), .C2(n6381), .A(n5050), .B(n5051), .ZN(
        n5028) );
  AOI22_X1 U2361 ( .A1(net644551), .A2(n6382), .B1(net644519), .B2(n3880), 
        .ZN(n5034) );
  AOI22_X1 U2360 ( .A1(n468), .A2(n4225), .B1(n3896), .B2(n4075), .ZN(n5044)
         );
  AOI22_X1 U2359 ( .A1(net644616), .A2(n3895), .B1(net644487), .B2(n3894), 
        .ZN(n5045) );
  AOI22_X1 U2358 ( .A1(n6384), .A2(n380), .B1(n3891), .B2(n3967), .ZN(n5046)
         );
  AOI22_X1 U2357 ( .A1(net644584), .A2(n3890), .B1(net644680), .B2(n3897), 
        .ZN(n5047) );
  NAND4_X1 U2356 ( .A1(n5044), .A2(n5045), .A3(n5046), .A4(n5047), .ZN(n5036)
         );
  AOI22_X1 U2355 ( .A1(n470), .A2(n3904), .B1(n3903), .B2(n4076), .ZN(n5038)
         );
  AOI22_X1 U2354 ( .A1(net644776), .A2(n3902), .B1(net644744), .B2(n3901), 
        .ZN(n5039) );
  AOI22_X1 U2353 ( .A1(net644906), .A2(n3900), .B1(net644423), .B2(n3899), 
        .ZN(n5040) );
  AOI22_X1 U2352 ( .A1(n6385), .A2(n469), .B1(n3898), .B2(n3968), .ZN(n5041)
         );
  NAND4_X1 U2351 ( .A1(n5038), .A2(n5039), .A3(n5040), .A4(n5041), .ZN(n5037)
         );
  OAI21_X1 U2350 ( .B1(n5036), .B2(n5037), .A(n6386), .ZN(n5035) );
  OAI211_X1 U2349 ( .C1(n573), .C2(n4194), .A(n5034), .B(n5035), .ZN(n5030) );
  AOI22_X1 U2348 ( .A1(net644807), .A2(n6389), .B1(n6388), .B2(n4077), .ZN(
        n5032) );
  OAI21_X1 U2347 ( .B1(n635), .B2(n4189), .A(n5032), .ZN(n5031) );
  AOI211_X1 U2346 ( .C1(net644712), .C2(n4186), .A(n5030), .B(n5031), .ZN(
        n5029) );
  NAND4_X1 U2345 ( .A1(n5026), .A2(n5027), .A3(n5028), .A4(n5029), .ZN(n2736)
         );
  AOI22_X1 U2315 ( .A1(n6376), .A2(n3972), .B1(n6375), .B2(n3921), .ZN(n4966)
         );
  AOI22_X1 U2314 ( .A1(net644875), .A2(n6378), .B1(net644841), .B2(n6377), 
        .ZN(n4967) );
  AOI22_X1 U2313 ( .A1(net644457), .A2(n6380), .B1(DATAIN[6]), .B2(n6379), 
        .ZN(n4992) );
  OAI21_X1 U2312 ( .B1(n4235), .B2(net644393), .A(n4992), .ZN(n4990) );
  OAI22_X1 U2311 ( .A1(n665), .A2(n4233), .B1(n540), .B2(n4234), .ZN(n4991) );
  AOI211_X1 U2310 ( .C1(net644649), .C2(n6381), .A(n4990), .B(n4991), .ZN(
        n4968) );
  AOI22_X1 U2309 ( .A1(net644553), .A2(n4228), .B1(net644521), .B2(n3880), 
        .ZN(n4974) );
  AOI22_X1 U2308 ( .A1(n462), .A2(n4225), .B1(n3896), .B2(n4081), .ZN(n4984)
         );
  AOI22_X1 U2307 ( .A1(net644618), .A2(n3895), .B1(net644489), .B2(n3894), 
        .ZN(n4985) );
  AOI22_X1 U2306 ( .A1(n6384), .A2(n378), .B1(n3891), .B2(n3973), .ZN(n4986)
         );
  AOI22_X1 U2305 ( .A1(net644586), .A2(n3890), .B1(net644682), .B2(n3897), 
        .ZN(n4987) );
  NAND4_X1 U2304 ( .A1(n4984), .A2(n4985), .A3(n4986), .A4(n4987), .ZN(n4976)
         );
  AOI22_X1 U2303 ( .A1(n464), .A2(n3904), .B1(n3903), .B2(n4082), .ZN(n4978)
         );
  AOI22_X1 U2302 ( .A1(net644778), .A2(n3902), .B1(net644746), .B2(n3901), 
        .ZN(n4979) );
  AOI22_X1 U2301 ( .A1(net644908), .A2(n3900), .B1(net644425), .B2(n3899), 
        .ZN(n4980) );
  AOI22_X1 U2300 ( .A1(n6385), .A2(n463), .B1(n3898), .B2(n3974), .ZN(n4981)
         );
  NAND4_X1 U2299 ( .A1(n4978), .A2(n4979), .A3(n4980), .A4(n4981), .ZN(n4977)
         );
  OAI21_X1 U2298 ( .B1(n4976), .B2(n4977), .A(n6386), .ZN(n4975) );
  OAI211_X1 U2297 ( .C1(n571), .C2(n4194), .A(n4974), .B(n4975), .ZN(n4970) );
  AOI22_X1 U2296 ( .A1(net644809), .A2(n6389), .B1(n6388), .B2(n4083), .ZN(
        n4972) );
  OAI21_X1 U2295 ( .B1(n633), .B2(n4189), .A(n4972), .ZN(n4971) );
  AOI211_X1 U2294 ( .C1(net644714), .C2(n6390), .A(n4970), .B(n4971), .ZN(
        n4969) );
  NAND4_X1 U2293 ( .A1(n4966), .A2(n4967), .A3(n4968), .A4(n4969), .ZN(n2740)
         );
  AOI22_X1 U2289 ( .A1(n6376), .A2(n3975), .B1(n6375), .B2(n3922), .ZN(n4936)
         );
  AOI22_X1 U2288 ( .A1(net644876), .A2(n6378), .B1(net644842), .B2(n6377), 
        .ZN(n4937) );
  AOI22_X1 U2287 ( .A1(net644458), .A2(n6380), .B1(DATAIN[7]), .B2(n4238), 
        .ZN(n4962) );
  OAI21_X1 U2286 ( .B1(n4235), .B2(net644394), .A(n4962), .ZN(n4960) );
  OAI22_X1 U2285 ( .A1(n664), .A2(n4233), .B1(n539), .B2(n4234), .ZN(n4961) );
  AOI211_X1 U2284 ( .C1(net644650), .C2(n6381), .A(n4960), .B(n4961), .ZN(
        n4938) );
  AOI22_X1 U2283 ( .A1(net644554), .A2(n4228), .B1(net644522), .B2(n3880), 
        .ZN(n4944) );
  AOI22_X1 U2282 ( .A1(n459), .A2(n6383), .B1(n3896), .B2(n4084), .ZN(n4954)
         );
  AOI22_X1 U2281 ( .A1(net644619), .A2(n3895), .B1(net644490), .B2(n3894), 
        .ZN(n4955) );
  AOI22_X1 U2280 ( .A1(n6384), .A2(n377), .B1(n3891), .B2(n3976), .ZN(n4956)
         );
  AOI22_X1 U2279 ( .A1(net644587), .A2(n3890), .B1(net644683), .B2(n3897), 
        .ZN(n4957) );
  NAND4_X1 U2278 ( .A1(n4954), .A2(n4955), .A3(n4956), .A4(n4957), .ZN(n4946)
         );
  AOI22_X1 U2277 ( .A1(n461), .A2(n3904), .B1(n3903), .B2(n4085), .ZN(n4948)
         );
  AOI22_X1 U2276 ( .A1(net644779), .A2(n3902), .B1(net644747), .B2(n3901), 
        .ZN(n4949) );
  AOI22_X1 U2275 ( .A1(net644909), .A2(n3900), .B1(net644426), .B2(n3899), 
        .ZN(n4950) );
  AOI22_X1 U2274 ( .A1(n6385), .A2(n460), .B1(n3898), .B2(n3977), .ZN(n4951)
         );
  NAND4_X1 U2273 ( .A1(n4948), .A2(n4949), .A3(n4950), .A4(n4951), .ZN(n4947)
         );
  OAI21_X1 U2272 ( .B1(n4946), .B2(n4947), .A(n6386), .ZN(n4945) );
  OAI211_X1 U2271 ( .C1(n570), .C2(n4194), .A(n4944), .B(n4945), .ZN(n4940) );
  AOI22_X1 U2270 ( .A1(net644810), .A2(n6389), .B1(n6388), .B2(n4086), .ZN(
        n4942) );
  OAI21_X1 U2269 ( .B1(n632), .B2(n4189), .A(n4942), .ZN(n4941) );
  AOI211_X1 U2268 ( .C1(net644715), .C2(n4186), .A(n4940), .B(n4941), .ZN(
        n4939) );
  NAND4_X1 U2267 ( .A1(n4936), .A2(n4937), .A3(n4938), .A4(n4939), .ZN(n2742)
         );
  AOI22_X1 U2263 ( .A1(n6376), .A2(n3978), .B1(n6375), .B2(n3923), .ZN(n4906)
         );
  AOI22_X1 U2262 ( .A1(net644877), .A2(n6378), .B1(net644843), .B2(n6377), 
        .ZN(n4907) );
  AOI22_X1 U2261 ( .A1(net644459), .A2(n4237), .B1(DATAIN[8]), .B2(n4238), 
        .ZN(n4932) );
  OAI21_X1 U2260 ( .B1(n4235), .B2(net644395), .A(n4932), .ZN(n4930) );
  OAI22_X1 U2259 ( .A1(n663), .A2(n4233), .B1(n538), .B2(n4234), .ZN(n4931) );
  AOI211_X1 U2258 ( .C1(net644651), .C2(n6381), .A(n4930), .B(n4931), .ZN(
        n4908) );
  AOI22_X1 U2257 ( .A1(net644555), .A2(n6382), .B1(net644523), .B2(n3880), 
        .ZN(n4914) );
  AOI22_X1 U2256 ( .A1(n456), .A2(n6383), .B1(n4226), .B2(n4087), .ZN(n4924)
         );
  AOI22_X1 U2255 ( .A1(net644620), .A2(n4223), .B1(net644491), .B2(n3894), 
        .ZN(n4925) );
  AOI22_X1 U2254 ( .A1(n6384), .A2(n376), .B1(n3891), .B2(n3979), .ZN(n4926)
         );
  AOI22_X1 U2253 ( .A1(net644588), .A2(n3890), .B1(net644684), .B2(n4219), 
        .ZN(n4927) );
  NAND4_X1 U2252 ( .A1(n4924), .A2(n4925), .A3(n4926), .A4(n4927), .ZN(n4916)
         );
  AOI22_X1 U2251 ( .A1(n458), .A2(n3904), .B1(n3903), .B2(n4088), .ZN(n4918)
         );
  AOI22_X1 U2250 ( .A1(net644780), .A2(n4209), .B1(net644748), .B2(n3901), 
        .ZN(n4919) );
  AOI22_X1 U2249 ( .A1(net644910), .A2(n4207), .B1(net644427), .B2(n3899), 
        .ZN(n4920) );
  AOI22_X1 U2248 ( .A1(n6385), .A2(n457), .B1(n3898), .B2(n3980), .ZN(n4921)
         );
  NAND4_X1 U2247 ( .A1(n4918), .A2(n4919), .A3(n4920), .A4(n4921), .ZN(n4917)
         );
  OAI21_X1 U2246 ( .B1(n4916), .B2(n4917), .A(n6386), .ZN(n4915) );
  OAI211_X1 U2245 ( .C1(n569), .C2(n4194), .A(n4914), .B(n4915), .ZN(n4910) );
  AOI22_X1 U2244 ( .A1(net644811), .A2(n6389), .B1(n6388), .B2(n4089), .ZN(
        n4912) );
  OAI21_X1 U2243 ( .B1(n631), .B2(n4189), .A(n4912), .ZN(n4911) );
  AOI211_X1 U2242 ( .C1(net644716), .C2(n4186), .A(n4910), .B(n4911), .ZN(
        n4909) );
  NAND4_X1 U2241 ( .A1(n4906), .A2(n4907), .A3(n4908), .A4(n4909), .ZN(n2744)
         );
  AOI22_X1 U2237 ( .A1(n6376), .A2(n3981), .B1(n6375), .B2(n3925), .ZN(n4876)
         );
  AOI22_X1 U2236 ( .A1(net644878), .A2(n6378), .B1(net644844), .B2(n4240), 
        .ZN(n4877) );
  AOI22_X1 U2235 ( .A1(net644460), .A2(n4237), .B1(DATAIN[9]), .B2(n6379), 
        .ZN(n4902) );
  OAI21_X1 U2234 ( .B1(n4235), .B2(net644396), .A(n4902), .ZN(n4900) );
  OAI22_X1 U2233 ( .A1(n662), .A2(n4233), .B1(n537), .B2(n4234), .ZN(n4901) );
  AOI211_X1 U2232 ( .C1(net644652), .C2(n6381), .A(n4900), .B(n4901), .ZN(
        n4878) );
  AOI22_X1 U2231 ( .A1(net644556), .A2(n6382), .B1(net644524), .B2(n3880), 
        .ZN(n4884) );
  AOI22_X1 U2230 ( .A1(n453), .A2(n6383), .B1(n3896), .B2(n4090), .ZN(n4894)
         );
  AOI22_X1 U2229 ( .A1(net644621), .A2(n4223), .B1(net644492), .B2(n3894), 
        .ZN(n4895) );
  AOI22_X1 U2228 ( .A1(n6384), .A2(n375), .B1(n3891), .B2(n3982), .ZN(n4896)
         );
  AOI22_X1 U2227 ( .A1(net644589), .A2(n3890), .B1(net644685), .B2(n4219), 
        .ZN(n4897) );
  NAND4_X1 U2226 ( .A1(n4894), .A2(n4895), .A3(n4896), .A4(n4897), .ZN(n4886)
         );
  AOI22_X1 U2225 ( .A1(n455), .A2(n3904), .B1(n3903), .B2(n4091), .ZN(n4888)
         );
  AOI22_X1 U2224 ( .A1(net644781), .A2(n4209), .B1(net644749), .B2(n3901), 
        .ZN(n4889) );
  AOI22_X1 U2223 ( .A1(net644911), .A2(n4207), .B1(net644428), .B2(n3899), 
        .ZN(n4890) );
  AOI22_X1 U2222 ( .A1(n6385), .A2(n454), .B1(n3898), .B2(n3983), .ZN(n4891)
         );
  NAND4_X1 U2221 ( .A1(n4888), .A2(n4889), .A3(n4890), .A4(n4891), .ZN(n4887)
         );
  OAI21_X1 U2220 ( .B1(n4886), .B2(n4887), .A(n6386), .ZN(n4885) );
  OAI211_X1 U2219 ( .C1(n568), .C2(n4194), .A(n4884), .B(n4885), .ZN(n4880) );
  AOI22_X1 U2218 ( .A1(net644812), .A2(n6389), .B1(n6388), .B2(n4092), .ZN(
        n4882) );
  OAI21_X1 U2217 ( .B1(n630), .B2(n4189), .A(n4882), .ZN(n4881) );
  AOI211_X1 U2216 ( .C1(net644717), .C2(n4186), .A(n4880), .B(n4881), .ZN(
        n4879) );
  NAND4_X1 U2215 ( .A1(n4876), .A2(n4877), .A3(n4878), .A4(n4879), .ZN(n2746)
         );
  AOI22_X1 U2211 ( .A1(n4241), .A2(n3984), .B1(n6375), .B2(n3928), .ZN(n4846)
         );
  AOI22_X1 U2210 ( .A1(net644879), .A2(n6378), .B1(net644845), .B2(n4240), 
        .ZN(n4847) );
  AOI22_X1 U2209 ( .A1(net644461), .A2(n4237), .B1(DATAIN[10]), .B2(n6379), 
        .ZN(n4872) );
  OAI21_X1 U2208 ( .B1(n4235), .B2(net644397), .A(n4872), .ZN(n4870) );
  OAI22_X1 U2207 ( .A1(n661), .A2(n4233), .B1(n536), .B2(n4234), .ZN(n4871) );
  AOI211_X1 U2206 ( .C1(net644653), .C2(n6381), .A(n4870), .B(n4871), .ZN(
        n4848) );
  AOI22_X1 U2205 ( .A1(net644557), .A2(n6382), .B1(net644525), .B2(n3880), 
        .ZN(n4854) );
  AOI22_X1 U2204 ( .A1(n450), .A2(n6383), .B1(n3896), .B2(n4093), .ZN(n4864)
         );
  AOI22_X1 U2203 ( .A1(net644622), .A2(n4223), .B1(net644493), .B2(n3894), 
        .ZN(n4865) );
  AOI22_X1 U2202 ( .A1(n6384), .A2(n374), .B1(n3891), .B2(n3985), .ZN(n4866)
         );
  AOI22_X1 U2201 ( .A1(net644590), .A2(n3890), .B1(net644686), .B2(n4219), 
        .ZN(n4867) );
  NAND4_X1 U2200 ( .A1(n4864), .A2(n4865), .A3(n4866), .A4(n4867), .ZN(n4856)
         );
  AOI22_X1 U2199 ( .A1(n452), .A2(n3904), .B1(n3903), .B2(n4094), .ZN(n4858)
         );
  AOI22_X1 U2198 ( .A1(net644782), .A2(n4209), .B1(net644750), .B2(n3901), 
        .ZN(n4859) );
  AOI22_X1 U2197 ( .A1(net644912), .A2(n4207), .B1(net644429), .B2(n3899), 
        .ZN(n4860) );
  AOI22_X1 U2196 ( .A1(n6385), .A2(n451), .B1(n3898), .B2(n3986), .ZN(n4861)
         );
  NAND4_X1 U2195 ( .A1(n4858), .A2(n4859), .A3(n4860), .A4(n4861), .ZN(n4857)
         );
  OAI21_X1 U2194 ( .B1(n4856), .B2(n4857), .A(n6386), .ZN(n4855) );
  OAI211_X1 U2193 ( .C1(n567), .C2(n4194), .A(n4854), .B(n4855), .ZN(n4850) );
  AOI22_X1 U2192 ( .A1(net644813), .A2(n6389), .B1(n6388), .B2(n4095), .ZN(
        n4852) );
  OAI21_X1 U2191 ( .B1(n629), .B2(n4189), .A(n4852), .ZN(n4851) );
  AOI211_X1 U2190 ( .C1(net644718), .C2(n4186), .A(n4850), .B(n4851), .ZN(
        n4849) );
  NAND4_X1 U2189 ( .A1(n4846), .A2(n4847), .A3(n4848), .A4(n4849), .ZN(n2748)
         );
  AOI22_X1 U1873 ( .A1(n6376), .A2(n4029), .B1(n4243), .B2(n3941), .ZN(n4456)
         );
  AOI22_X1 U1872 ( .A1(net644892), .A2(n6378), .B1(net644858), .B2(n4240), 
        .ZN(n4457) );
  AOI22_X1 U1871 ( .A1(net644474), .A2(n6380), .B1(DATAIN[23]), .B2(n6379), 
        .ZN(n4482) );
  OAI21_X1 U1870 ( .B1(n4235), .B2(net644410), .A(n4482), .ZN(n4480) );
  OAI22_X1 U1869 ( .A1(n648), .A2(n4233), .B1(n523), .B2(n4234), .ZN(n4481) );
  AOI211_X1 U1868 ( .C1(net644666), .C2(n6381), .A(n4480), .B(n4481), .ZN(
        n4458) );
  AOI22_X1 U1867 ( .A1(net644570), .A2(n6382), .B1(net644538), .B2(n4229), 
        .ZN(n4464) );
  AOI22_X1 U1866 ( .A1(n411), .A2(n6383), .B1(n3896), .B2(n4137), .ZN(n4474)
         );
  AOI22_X1 U1865 ( .A1(net644635), .A2(n3895), .B1(net644506), .B2(n4224), 
        .ZN(n4475) );
  AOI22_X1 U1864 ( .A1(n4220), .A2(n361), .B1(n3891), .B2(n4030), .ZN(n4476)
         );
  AOI22_X1 U1863 ( .A1(net644603), .A2(n4218), .B1(net644699), .B2(n3897), 
        .ZN(n4477) );
  NAND4_X1 U1862 ( .A1(n4474), .A2(n4475), .A3(n4476), .A4(n4477), .ZN(n4466)
         );
  AOI22_X1 U1861 ( .A1(n413), .A2(n4211), .B1(n3903), .B2(n4138), .ZN(n4468)
         );
  AOI22_X1 U1860 ( .A1(net644795), .A2(n3902), .B1(net644763), .B2(n4210), 
        .ZN(n4469) );
  AOI22_X1 U1859 ( .A1(net644925), .A2(n3900), .B1(net644442), .B2(n4208), 
        .ZN(n4470) );
  AOI22_X1 U1858 ( .A1(n6385), .A2(n412), .B1(n3898), .B2(n4031), .ZN(n4471)
         );
  NAND4_X1 U1857 ( .A1(n4468), .A2(n4469), .A3(n4470), .A4(n4471), .ZN(n4467)
         );
  OAI21_X1 U1856 ( .B1(n4466), .B2(n4467), .A(n6386), .ZN(n4465) );
  OAI211_X1 U1855 ( .C1(n554), .C2(n4194), .A(n4464), .B(n4465), .ZN(n4460) );
  AOI22_X1 U1854 ( .A1(net644826), .A2(n6389), .B1(n6388), .B2(n4139), .ZN(
        n4462) );
  OAI21_X1 U1853 ( .B1(n616), .B2(n4189), .A(n4462), .ZN(n4461) );
  AOI211_X1 U1852 ( .C1(net644731), .C2(n6390), .A(n4460), .B(n4461), .ZN(
        n4459) );
  NAND4_X1 U1851 ( .A1(n4456), .A2(n4457), .A3(n4458), .A4(n4459), .ZN(n2774)
         );
  AOI22_X1 U1847 ( .A1(n4241), .A2(n4032), .B1(n6375), .B2(n3942), .ZN(n4426)
         );
  AOI22_X1 U1846 ( .A1(net644893), .A2(n6378), .B1(net644859), .B2(n6377), 
        .ZN(n4427) );
  AOI22_X1 U1845 ( .A1(net644475), .A2(n6380), .B1(DATAIN[24]), .B2(n6379), 
        .ZN(n4452) );
  OAI21_X1 U1844 ( .B1(n4235), .B2(net644411), .A(n4452), .ZN(n4450) );
  OAI22_X1 U1843 ( .A1(n647), .A2(n4233), .B1(n522), .B2(n4234), .ZN(n4451) );
  AOI211_X1 U1842 ( .C1(net644667), .C2(n6381), .A(n4450), .B(n4451), .ZN(
        n4428) );
  AOI22_X1 U1841 ( .A1(net644571), .A2(n6382), .B1(net644539), .B2(n3880), 
        .ZN(n4434) );
  AOI22_X1 U1840 ( .A1(n408), .A2(n6383), .B1(n3896), .B2(n4140), .ZN(n4444)
         );
  AOI22_X1 U1839 ( .A1(net644636), .A2(n3895), .B1(net644507), .B2(n3894), 
        .ZN(n4445) );
  AOI22_X1 U1838 ( .A1(n4220), .A2(n360), .B1(n4221), .B2(n4034), .ZN(n4446)
         );
  AOI22_X1 U1837 ( .A1(net644604), .A2(n3890), .B1(net644700), .B2(n3897), 
        .ZN(n4447) );
  NAND4_X1 U1836 ( .A1(n4444), .A2(n4445), .A3(n4446), .A4(n4447), .ZN(n4436)
         );
  AOI22_X1 U1835 ( .A1(n410), .A2(n4211), .B1(n4212), .B2(n4141), .ZN(n4438)
         );
  AOI22_X1 U1834 ( .A1(net644796), .A2(n3902), .B1(net644764), .B2(n3901), 
        .ZN(n4439) );
  AOI22_X1 U1833 ( .A1(net644926), .A2(n3900), .B1(net644443), .B2(n3899), 
        .ZN(n4440) );
  AOI22_X1 U1832 ( .A1(n6385), .A2(n409), .B1(n3898), .B2(n4037), .ZN(n4441)
         );
  NAND4_X1 U1831 ( .A1(n4438), .A2(n4439), .A3(n4440), .A4(n4441), .ZN(n4437)
         );
  OAI21_X1 U1830 ( .B1(n4436), .B2(n4437), .A(n6386), .ZN(n4435) );
  OAI211_X1 U1829 ( .C1(n553), .C2(n4194), .A(n4434), .B(n4435), .ZN(n4430) );
  AOI22_X1 U1828 ( .A1(net644827), .A2(n6389), .B1(n6388), .B2(n4142), .ZN(
        n4432) );
  OAI21_X1 U1827 ( .B1(n615), .B2(n4189), .A(n4432), .ZN(n4431) );
  AOI211_X1 U1826 ( .C1(net644732), .C2(n6390), .A(n4430), .B(n4431), .ZN(
        n4429) );
  NAND4_X1 U1825 ( .A1(n4426), .A2(n4427), .A3(n4428), .A4(n4429), .ZN(n2776)
         );
  AOI22_X1 U2133 ( .A1(n6376), .A2(n3993), .B1(n6375), .B2(n3931), .ZN(n4756)
         );
  AOI22_X1 U2132 ( .A1(net644882), .A2(n6378), .B1(net644848), .B2(n6377), 
        .ZN(n4757) );
  AOI22_X1 U2131 ( .A1(net644464), .A2(n6380), .B1(DATAIN[13]), .B2(n6379), 
        .ZN(n4782) );
  OAI21_X1 U2130 ( .B1(n4235), .B2(net644400), .A(n4782), .ZN(n4780) );
  OAI22_X1 U2129 ( .A1(n658), .A2(n4233), .B1(n533), .B2(n4234), .ZN(n4781) );
  AOI211_X1 U2128 ( .C1(net644656), .C2(n6381), .A(n4780), .B(n4781), .ZN(
        n4758) );
  AOI22_X1 U2127 ( .A1(net644560), .A2(n6382), .B1(net644528), .B2(n3880), 
        .ZN(n4764) );
  AOI22_X1 U2126 ( .A1(n441), .A2(n4225), .B1(n3896), .B2(n4102), .ZN(n4774)
         );
  AOI22_X1 U2125 ( .A1(net644625), .A2(n3895), .B1(net644496), .B2(n3894), 
        .ZN(n4775) );
  AOI22_X1 U2124 ( .A1(n6384), .A2(n371), .B1(n3891), .B2(n3998), .ZN(n4776)
         );
  AOI22_X1 U2123 ( .A1(net644593), .A2(n3890), .B1(net644689), .B2(n3897), 
        .ZN(n4777) );
  NAND4_X1 U2122 ( .A1(n4774), .A2(n4775), .A3(n4776), .A4(n4777), .ZN(n4766)
         );
  AOI22_X1 U2121 ( .A1(n443), .A2(n3904), .B1(n3903), .B2(n4103), .ZN(n4768)
         );
  AOI22_X1 U2120 ( .A1(net644785), .A2(n3902), .B1(net644753), .B2(n3901), 
        .ZN(n4769) );
  AOI22_X1 U2119 ( .A1(net644915), .A2(n3900), .B1(net644432), .B2(n3899), 
        .ZN(n4770) );
  AOI22_X1 U2118 ( .A1(n6385), .A2(n442), .B1(n3898), .B2(n3999), .ZN(n4771)
         );
  NAND4_X1 U2117 ( .A1(n4768), .A2(n4769), .A3(n4770), .A4(n4771), .ZN(n4767)
         );
  OAI21_X1 U2116 ( .B1(n4766), .B2(n4767), .A(n6386), .ZN(n4765) );
  OAI211_X1 U2115 ( .C1(n564), .C2(n4194), .A(n4764), .B(n4765), .ZN(n4760) );
  AOI22_X1 U2114 ( .A1(net644816), .A2(n6389), .B1(n6388), .B2(n4104), .ZN(
        n4762) );
  OAI21_X1 U2113 ( .B1(n626), .B2(n4189), .A(n4762), .ZN(n4761) );
  AOI211_X1 U2112 ( .C1(net644721), .C2(n6390), .A(n4760), .B(n4761), .ZN(
        n4759) );
  NAND4_X1 U2111 ( .A1(n4756), .A2(n4757), .A3(n4758), .A4(n4759), .ZN(n2754)
         );
  AOI22_X1 U2107 ( .A1(n6376), .A2(n4002), .B1(n6375), .B2(n3932), .ZN(n4726)
         );
  AOI22_X1 U2106 ( .A1(net644883), .A2(n6378), .B1(net644849), .B2(n6377), 
        .ZN(n4727) );
  AOI22_X1 U2105 ( .A1(net644465), .A2(n6380), .B1(DATAIN[14]), .B2(n6379), 
        .ZN(n4752) );
  OAI21_X1 U2104 ( .B1(n4235), .B2(net644401), .A(n4752), .ZN(n4750) );
  OAI22_X1 U2103 ( .A1(n657), .A2(n4233), .B1(n532), .B2(n4234), .ZN(n4751) );
  AOI211_X1 U2102 ( .C1(net644657), .C2(n6381), .A(n4750), .B(n4751), .ZN(
        n4728) );
  AOI22_X1 U2101 ( .A1(net644561), .A2(n6382), .B1(net644529), .B2(n3880), 
        .ZN(n4734) );
  AOI22_X1 U2100 ( .A1(n438), .A2(n4225), .B1(n3896), .B2(n4105), .ZN(n4744)
         );
  AOI22_X1 U2099 ( .A1(net644626), .A2(n3895), .B1(net644497), .B2(n3894), 
        .ZN(n4745) );
  AOI22_X1 U2098 ( .A1(n6384), .A2(n370), .B1(n3891), .B2(n4003), .ZN(n4746)
         );
  AOI22_X1 U2097 ( .A1(net644594), .A2(n3890), .B1(net644690), .B2(n3897), 
        .ZN(n4747) );
  NAND4_X1 U2096 ( .A1(n4744), .A2(n4745), .A3(n4746), .A4(n4747), .ZN(n4736)
         );
  AOI22_X1 U2095 ( .A1(n440), .A2(n3904), .B1(n3903), .B2(n4109), .ZN(n4738)
         );
  AOI22_X1 U2094 ( .A1(net644786), .A2(n3902), .B1(net644754), .B2(n3901), 
        .ZN(n4739) );
  AOI22_X1 U2093 ( .A1(net644916), .A2(n3900), .B1(net644433), .B2(n3899), 
        .ZN(n4740) );
  AOI22_X1 U2092 ( .A1(n6385), .A2(n439), .B1(n3898), .B2(n4004), .ZN(n4741)
         );
  NAND4_X1 U2091 ( .A1(n4738), .A2(n4739), .A3(n4740), .A4(n4741), .ZN(n4737)
         );
  OAI21_X1 U2090 ( .B1(n4736), .B2(n4737), .A(n6386), .ZN(n4735) );
  OAI211_X1 U2089 ( .C1(n563), .C2(n4194), .A(n4734), .B(n4735), .ZN(n4730) );
  AOI22_X1 U2088 ( .A1(net644817), .A2(n6389), .B1(n6388), .B2(n4112), .ZN(
        n4732) );
  OAI21_X1 U2087 ( .B1(n625), .B2(n4189), .A(n4732), .ZN(n4731) );
  AOI211_X1 U2086 ( .C1(net644722), .C2(n6390), .A(n4730), .B(n4731), .ZN(
        n4729) );
  NAND4_X1 U2085 ( .A1(n4726), .A2(n4727), .A3(n4728), .A4(n4729), .ZN(n2756)
         );
  AOI22_X1 U2081 ( .A1(n6376), .A2(n4005), .B1(n4243), .B2(n3933), .ZN(n4696)
         );
  AOI22_X1 U2080 ( .A1(net644884), .A2(n6378), .B1(net644850), .B2(n4240), 
        .ZN(n4697) );
  AOI22_X1 U2079 ( .A1(net644466), .A2(n6380), .B1(DATAIN[15]), .B2(n6379), 
        .ZN(n4722) );
  OAI21_X1 U2078 ( .B1(n4235), .B2(net644402), .A(n4722), .ZN(n4720) );
  OAI22_X1 U2077 ( .A1(n656), .A2(n4233), .B1(n531), .B2(n4234), .ZN(n4721) );
  AOI211_X1 U2076 ( .C1(net644658), .C2(n6381), .A(n4720), .B(n4721), .ZN(
        n4698) );
  AOI22_X1 U2075 ( .A1(net644562), .A2(n6382), .B1(net644530), .B2(n3880), 
        .ZN(n4704) );
  AOI22_X1 U2074 ( .A1(n435), .A2(n6383), .B1(n3896), .B2(n4113), .ZN(n4714)
         );
  AOI22_X1 U2073 ( .A1(net644627), .A2(n3895), .B1(net644498), .B2(n3894), 
        .ZN(n4715) );
  AOI22_X1 U2072 ( .A1(n4220), .A2(n369), .B1(n3891), .B2(n4006), .ZN(n4716)
         );
  AOI22_X1 U2071 ( .A1(net644595), .A2(n3890), .B1(net644691), .B2(n3897), 
        .ZN(n4717) );
  NAND4_X1 U2070 ( .A1(n4714), .A2(n4715), .A3(n4716), .A4(n4717), .ZN(n4706)
         );
  AOI22_X1 U2069 ( .A1(n437), .A2(n3904), .B1(n3903), .B2(n4114), .ZN(n4708)
         );
  AOI22_X1 U2068 ( .A1(net644787), .A2(n3902), .B1(net644755), .B2(n3901), 
        .ZN(n4709) );
  AOI22_X1 U2067 ( .A1(net644917), .A2(n3900), .B1(net644434), .B2(n3899), 
        .ZN(n4710) );
  AOI22_X1 U2066 ( .A1(n6385), .A2(n436), .B1(n3898), .B2(n4007), .ZN(n4711)
         );
  NAND4_X1 U2065 ( .A1(n4708), .A2(n4709), .A3(n4710), .A4(n4711), .ZN(n4707)
         );
  OAI21_X1 U2064 ( .B1(n4706), .B2(n4707), .A(n6386), .ZN(n4705) );
  OAI211_X1 U2063 ( .C1(n562), .C2(n4194), .A(n4704), .B(n4705), .ZN(n4700) );
  AOI22_X1 U2062 ( .A1(net644818), .A2(n6389), .B1(n6388), .B2(n4115), .ZN(
        n4702) );
  OAI21_X1 U2061 ( .B1(n624), .B2(n4189), .A(n4702), .ZN(n4701) );
  AOI211_X1 U2060 ( .C1(net644723), .C2(n6390), .A(n4700), .B(n4701), .ZN(
        n4699) );
  NAND4_X1 U2059 ( .A1(n4696), .A2(n4697), .A3(n4698), .A4(n4699), .ZN(n2758)
         );
  AOI22_X1 U1925 ( .A1(n6376), .A2(n4023), .B1(n6375), .B2(n3939), .ZN(n4516)
         );
  AOI22_X1 U1924 ( .A1(net644890), .A2(n4239), .B1(net644856), .B2(n4240), 
        .ZN(n4517) );
  AOI22_X1 U1923 ( .A1(net644472), .A2(n4237), .B1(DATAIN[21]), .B2(n6379), 
        .ZN(n4542) );
  OAI21_X1 U1922 ( .B1(n4235), .B2(net644408), .A(n4542), .ZN(n4540) );
  OAI22_X1 U1921 ( .A1(n650), .A2(n4233), .B1(n525), .B2(n4234), .ZN(n4541) );
  AOI211_X1 U1920 ( .C1(net644664), .C2(n6381), .A(n4540), .B(n4541), .ZN(
        n4518) );
  AOI22_X1 U1919 ( .A1(net644568), .A2(n6382), .B1(net644536), .B2(n4229), 
        .ZN(n4524) );
  AOI22_X1 U1918 ( .A1(n417), .A2(n6383), .B1(n3896), .B2(n4131), .ZN(n4534)
         );
  AOI22_X1 U1917 ( .A1(net644633), .A2(n3895), .B1(net644504), .B2(n4224), 
        .ZN(n4535) );
  AOI22_X1 U1916 ( .A1(n4220), .A2(n363), .B1(n3891), .B2(n4024), .ZN(n4536)
         );
  AOI22_X1 U1915 ( .A1(net644601), .A2(n4218), .B1(net644697), .B2(n3897), 
        .ZN(n4537) );
  NAND4_X1 U1914 ( .A1(n4534), .A2(n4535), .A3(n4536), .A4(n4537), .ZN(n4526)
         );
  AOI22_X1 U1913 ( .A1(n419), .A2(n3904), .B1(n3903), .B2(n4132), .ZN(n4528)
         );
  AOI22_X1 U1912 ( .A1(net644793), .A2(n3902), .B1(net644761), .B2(n4210), 
        .ZN(n4529) );
  AOI22_X1 U1911 ( .A1(net644923), .A2(n3900), .B1(net644440), .B2(n4208), 
        .ZN(n4530) );
  AOI22_X1 U1910 ( .A1(n6385), .A2(n418), .B1(n3898), .B2(n4025), .ZN(n4531)
         );
  NAND4_X1 U1909 ( .A1(n4528), .A2(n4529), .A3(n4530), .A4(n4531), .ZN(n4527)
         );
  OAI21_X1 U1908 ( .B1(n4526), .B2(n4527), .A(n6386), .ZN(n4525) );
  OAI211_X1 U1907 ( .C1(n556), .C2(n4194), .A(n4524), .B(n4525), .ZN(n4520) );
  AOI22_X1 U1906 ( .A1(net644824), .A2(n6389), .B1(n6388), .B2(n4133), .ZN(
        n4522) );
  OAI21_X1 U1905 ( .B1(n618), .B2(n4189), .A(n4522), .ZN(n4521) );
  AOI211_X1 U1904 ( .C1(net644729), .C2(n4186), .A(n4520), .B(n4521), .ZN(
        n4519) );
  NAND4_X1 U1903 ( .A1(n4516), .A2(n4517), .A3(n4518), .A4(n4519), .ZN(n2770)
         );
  AOI22_X1 U2029 ( .A1(n6376), .A2(n4011), .B1(n6375), .B2(n3935), .ZN(n4636)
         );
  AOI22_X1 U2028 ( .A1(net644886), .A2(n6378), .B1(net644852), .B2(n6377), 
        .ZN(n4637) );
  AOI22_X1 U2027 ( .A1(net644468), .A2(n6380), .B1(DATAIN[17]), .B2(n6379), 
        .ZN(n4662) );
  OAI21_X1 U2026 ( .B1(n4235), .B2(net644404), .A(n4662), .ZN(n4660) );
  OAI22_X1 U2025 ( .A1(n654), .A2(n4233), .B1(n529), .B2(n4234), .ZN(n4661) );
  AOI211_X1 U2024 ( .C1(net644660), .C2(n6381), .A(n4660), .B(n4661), .ZN(
        n4638) );
  AOI22_X1 U2023 ( .A1(net644564), .A2(n6382), .B1(net644532), .B2(n3880), 
        .ZN(n4644) );
  AOI22_X1 U2022 ( .A1(n429), .A2(n4225), .B1(n3896), .B2(n4119), .ZN(n4654)
         );
  AOI22_X1 U2021 ( .A1(net644629), .A2(n3895), .B1(net644500), .B2(n3894), 
        .ZN(n4655) );
  AOI22_X1 U2020 ( .A1(n6384), .A2(n367), .B1(n3891), .B2(n4012), .ZN(n4656)
         );
  AOI22_X1 U2019 ( .A1(net644597), .A2(n3890), .B1(net644693), .B2(n3897), 
        .ZN(n4657) );
  NAND4_X1 U2018 ( .A1(n4654), .A2(n4655), .A3(n4656), .A4(n4657), .ZN(n4646)
         );
  AOI22_X1 U2017 ( .A1(n431), .A2(n3904), .B1(n3903), .B2(n4120), .ZN(n4648)
         );
  AOI22_X1 U2016 ( .A1(net644789), .A2(n3902), .B1(net644757), .B2(n3901), 
        .ZN(n4649) );
  AOI22_X1 U2015 ( .A1(net644919), .A2(n3900), .B1(net644436), .B2(n3899), 
        .ZN(n4650) );
  AOI22_X1 U2014 ( .A1(n6385), .A2(n430), .B1(n3898), .B2(n4013), .ZN(n4651)
         );
  NAND4_X1 U2013 ( .A1(n4648), .A2(n4649), .A3(n4650), .A4(n4651), .ZN(n4647)
         );
  OAI21_X1 U2012 ( .B1(n4646), .B2(n4647), .A(n6386), .ZN(n4645) );
  OAI211_X1 U2011 ( .C1(n560), .C2(n4194), .A(n4644), .B(n4645), .ZN(n4640) );
  AOI22_X1 U2010 ( .A1(net644820), .A2(n6389), .B1(n6388), .B2(n4121), .ZN(
        n4642) );
  OAI21_X1 U2009 ( .B1(n622), .B2(n4189), .A(n4642), .ZN(n4641) );
  AOI211_X1 U2008 ( .C1(net644725), .C2(n6390), .A(n4640), .B(n4641), .ZN(
        n4639) );
  NAND4_X1 U2007 ( .A1(n4636), .A2(n4637), .A3(n4638), .A4(n4639), .ZN(n2762)
         );
  AOI22_X1 U2003 ( .A1(n6376), .A2(n4014), .B1(n6375), .B2(n3936), .ZN(n4606)
         );
  AOI22_X1 U2002 ( .A1(net644887), .A2(n6378), .B1(net644853), .B2(n6377), 
        .ZN(n4607) );
  AOI22_X1 U2001 ( .A1(net644469), .A2(n6380), .B1(DATAIN[18]), .B2(n6379), 
        .ZN(n4632) );
  OAI21_X1 U2000 ( .B1(n4235), .B2(net644405), .A(n4632), .ZN(n4630) );
  OAI22_X1 U1999 ( .A1(n653), .A2(n4233), .B1(n528), .B2(n4234), .ZN(n4631) );
  AOI211_X1 U1998 ( .C1(net644661), .C2(n6381), .A(n4630), .B(n4631), .ZN(
        n4608) );
  AOI22_X1 U1997 ( .A1(net644565), .A2(n6382), .B1(net644533), .B2(n3880), 
        .ZN(n4614) );
  AOI22_X1 U1996 ( .A1(n426), .A2(n4225), .B1(n3896), .B2(n4122), .ZN(n4624)
         );
  AOI22_X1 U1995 ( .A1(net644630), .A2(n3895), .B1(net644501), .B2(n3894), 
        .ZN(n4625) );
  AOI22_X1 U1994 ( .A1(n6384), .A2(n366), .B1(n3891), .B2(n4015), .ZN(n4626)
         );
  AOI22_X1 U1993 ( .A1(net644598), .A2(n3890), .B1(net644694), .B2(n3897), 
        .ZN(n4627) );
  NAND4_X1 U1992 ( .A1(n4624), .A2(n4625), .A3(n4626), .A4(n4627), .ZN(n4616)
         );
  AOI22_X1 U1991 ( .A1(n428), .A2(n3904), .B1(n3903), .B2(n4123), .ZN(n4618)
         );
  AOI22_X1 U1990 ( .A1(net644790), .A2(n3902), .B1(net644758), .B2(n3901), 
        .ZN(n4619) );
  AOI22_X1 U1989 ( .A1(net644920), .A2(n3900), .B1(net644437), .B2(n3899), 
        .ZN(n4620) );
  AOI22_X1 U1988 ( .A1(n6385), .A2(n427), .B1(n3898), .B2(n4016), .ZN(n4621)
         );
  NAND4_X1 U1987 ( .A1(n4618), .A2(n4619), .A3(n4620), .A4(n4621), .ZN(n4617)
         );
  OAI21_X1 U1986 ( .B1(n4616), .B2(n4617), .A(n6386), .ZN(n4615) );
  OAI211_X1 U1985 ( .C1(n559), .C2(n4194), .A(n4614), .B(n4615), .ZN(n4610) );
  AOI22_X1 U1984 ( .A1(net644821), .A2(n6389), .B1(n6388), .B2(n4124), .ZN(
        n4612) );
  OAI21_X1 U1983 ( .B1(n621), .B2(n4189), .A(n4612), .ZN(n4611) );
  AOI211_X1 U1982 ( .C1(net644726), .C2(n6390), .A(n4610), .B(n4611), .ZN(
        n4609) );
  NAND4_X1 U1981 ( .A1(n4606), .A2(n4607), .A3(n4608), .A4(n4609), .ZN(n2764)
         );
  AOI22_X1 U1977 ( .A1(n6376), .A2(n4017), .B1(n6375), .B2(n3937), .ZN(n4576)
         );
  AOI22_X1 U1976 ( .A1(net644888), .A2(n6378), .B1(net644854), .B2(n6377), 
        .ZN(n4577) );
  AOI22_X1 U1975 ( .A1(net644470), .A2(n6380), .B1(DATAIN[19]), .B2(n6379), 
        .ZN(n4602) );
  OAI21_X1 U1974 ( .B1(n4235), .B2(net644406), .A(n4602), .ZN(n4600) );
  OAI22_X1 U1973 ( .A1(n652), .A2(n4233), .B1(n527), .B2(n4234), .ZN(n4601) );
  AOI211_X1 U1972 ( .C1(net644662), .C2(n6381), .A(n4600), .B(n4601), .ZN(
        n4578) );
  AOI22_X1 U1971 ( .A1(net644566), .A2(n6382), .B1(net644534), .B2(n3880), 
        .ZN(n4584) );
  AOI22_X1 U1970 ( .A1(n423), .A2(n4225), .B1(n3896), .B2(n4125), .ZN(n4594)
         );
  AOI22_X1 U1969 ( .A1(net644631), .A2(n3895), .B1(net644502), .B2(n3894), 
        .ZN(n4595) );
  AOI22_X1 U1968 ( .A1(n6384), .A2(n365), .B1(n3891), .B2(n4018), .ZN(n4596)
         );
  AOI22_X1 U1967 ( .A1(net644599), .A2(n3890), .B1(net644695), .B2(n3897), 
        .ZN(n4597) );
  NAND4_X1 U1966 ( .A1(n4594), .A2(n4595), .A3(n4596), .A4(n4597), .ZN(n4586)
         );
  AOI22_X1 U1965 ( .A1(n425), .A2(n3904), .B1(n3903), .B2(n4126), .ZN(n4588)
         );
  AOI22_X1 U1964 ( .A1(net644791), .A2(n3902), .B1(net644759), .B2(n3901), 
        .ZN(n4589) );
  AOI22_X1 U1963 ( .A1(net644921), .A2(n3900), .B1(net644438), .B2(n3899), 
        .ZN(n4590) );
  AOI22_X1 U1962 ( .A1(n6385), .A2(n424), .B1(n3898), .B2(n4019), .ZN(n4591)
         );
  NAND4_X1 U1961 ( .A1(n4588), .A2(n4589), .A3(n4590), .A4(n4591), .ZN(n4587)
         );
  OAI21_X1 U1960 ( .B1(n4586), .B2(n4587), .A(n6386), .ZN(n4585) );
  OAI211_X1 U1959 ( .C1(n558), .C2(n4194), .A(n4584), .B(n4585), .ZN(n4580) );
  AOI22_X1 U1958 ( .A1(net644822), .A2(n6389), .B1(n6388), .B2(n4127), .ZN(
        n4582) );
  OAI21_X1 U1957 ( .B1(n620), .B2(n4189), .A(n4582), .ZN(n4581) );
  AOI211_X1 U1956 ( .C1(net644727), .C2(n6390), .A(n4580), .B(n4581), .ZN(
        n4579) );
  NAND4_X1 U1955 ( .A1(n4576), .A2(n4577), .A3(n4578), .A4(n4579), .ZN(n2766)
         );
  AOI22_X1 U1951 ( .A1(n6376), .A2(n4020), .B1(n6375), .B2(n3938), .ZN(n4546)
         );
  AOI22_X1 U1950 ( .A1(net644889), .A2(n4239), .B1(net644855), .B2(n4240), 
        .ZN(n4547) );
  AOI22_X1 U1949 ( .A1(net644471), .A2(n6380), .B1(DATAIN[20]), .B2(n6379), 
        .ZN(n4572) );
  OAI21_X1 U1948 ( .B1(n4235), .B2(net644407), .A(n4572), .ZN(n4570) );
  OAI22_X1 U1947 ( .A1(n651), .A2(n4233), .B1(n526), .B2(n4234), .ZN(n4571) );
  AOI211_X1 U1946 ( .C1(net644663), .C2(n6381), .A(n4570), .B(n4571), .ZN(
        n4548) );
  AOI22_X1 U1945 ( .A1(net644567), .A2(n6382), .B1(net644535), .B2(n4229), 
        .ZN(n4554) );
  AOI22_X1 U1944 ( .A1(n420), .A2(n6383), .B1(n3896), .B2(n4128), .ZN(n4564)
         );
  AOI22_X1 U1943 ( .A1(net644632), .A2(n3895), .B1(net644503), .B2(n4224), 
        .ZN(n4565) );
  AOI22_X1 U1942 ( .A1(n4220), .A2(n364), .B1(n3891), .B2(n4021), .ZN(n4566)
         );
  AOI22_X1 U1941 ( .A1(net644600), .A2(n3890), .B1(net644696), .B2(n3897), 
        .ZN(n4567) );
  NAND4_X1 U1940 ( .A1(n4564), .A2(n4565), .A3(n4566), .A4(n4567), .ZN(n4556)
         );
  AOI22_X1 U1939 ( .A1(n422), .A2(n3904), .B1(n3903), .B2(n4129), .ZN(n4558)
         );
  AOI22_X1 U1938 ( .A1(net644792), .A2(n3902), .B1(net644760), .B2(n4210), 
        .ZN(n4559) );
  AOI22_X1 U1937 ( .A1(net644922), .A2(n3900), .B1(net644439), .B2(n4208), 
        .ZN(n4560) );
  AOI22_X1 U1936 ( .A1(n4204), .A2(n421), .B1(n3898), .B2(n4022), .ZN(n4561)
         );
  NAND4_X1 U1935 ( .A1(n4558), .A2(n4559), .A3(n4560), .A4(n4561), .ZN(n4557)
         );
  OAI21_X1 U1934 ( .B1(n4556), .B2(n4557), .A(n6386), .ZN(n4555) );
  OAI211_X1 U1933 ( .C1(n557), .C2(n4194), .A(n4554), .B(n4555), .ZN(n4550) );
  AOI22_X1 U1932 ( .A1(net644823), .A2(n6389), .B1(n6388), .B2(n4130), .ZN(
        n4552) );
  OAI21_X1 U1931 ( .B1(n619), .B2(n4189), .A(n4552), .ZN(n4551) );
  AOI211_X1 U1930 ( .C1(net644728), .C2(n6390), .A(n4550), .B(n4551), .ZN(
        n4549) );
  NAND4_X1 U1929 ( .A1(n4546), .A2(n4547), .A3(n4548), .A4(n4549), .ZN(n2768)
         );
  AOI22_X1 U1769 ( .A1(n4241), .A2(n4044), .B1(n4243), .B2(n3945), .ZN(n4336)
         );
  AOI22_X1 U1768 ( .A1(net644896), .A2(n4239), .B1(net644862), .B2(n6377), 
        .ZN(n4337) );
  AOI22_X1 U1767 ( .A1(net644478), .A2(n6380), .B1(DATAIN[27]), .B2(n6379), 
        .ZN(n4362) );
  OAI21_X1 U1766 ( .B1(n4235), .B2(net644414), .A(n4362), .ZN(n4360) );
  OAI22_X1 U1765 ( .A1(n644), .A2(n4233), .B1(n519), .B2(n4234), .ZN(n4361) );
  AOI211_X1 U1764 ( .C1(net644670), .C2(n6381), .A(n4360), .B(n4361), .ZN(
        n4338) );
  AOI22_X1 U1763 ( .A1(net644574), .A2(n6382), .B1(net644542), .B2(n3880), 
        .ZN(n4344) );
  AOI22_X1 U1762 ( .A1(n399), .A2(n6383), .B1(n3896), .B2(n4152), .ZN(n4354)
         );
  AOI22_X1 U1761 ( .A1(net644639), .A2(n3895), .B1(net644510), .B2(n3894), 
        .ZN(n4355) );
  AOI22_X1 U1760 ( .A1(n4220), .A2(n357), .B1(n4221), .B2(n4045), .ZN(n4356)
         );
  AOI22_X1 U1759 ( .A1(net644607), .A2(n3890), .B1(net644703), .B2(n3897), 
        .ZN(n4357) );
  NAND4_X1 U1758 ( .A1(n4354), .A2(n4355), .A3(n4356), .A4(n4357), .ZN(n4346)
         );
  AOI22_X1 U1757 ( .A1(n401), .A2(n4211), .B1(n4212), .B2(n4153), .ZN(n4348)
         );
  AOI22_X1 U1756 ( .A1(net644799), .A2(n3902), .B1(net644767), .B2(n3901), 
        .ZN(n4349) );
  AOI22_X1 U1755 ( .A1(net644929), .A2(n3900), .B1(net644446), .B2(n3899), 
        .ZN(n4350) );
  AOI22_X1 U1754 ( .A1(n4204), .A2(n400), .B1(n4205), .B2(n4046), .ZN(n4351)
         );
  NAND4_X1 U1753 ( .A1(n4348), .A2(n4349), .A3(n4350), .A4(n4351), .ZN(n4347)
         );
  OAI21_X1 U1752 ( .B1(n4346), .B2(n4347), .A(n6386), .ZN(n4345) );
  OAI211_X1 U1751 ( .C1(n550), .C2(n4194), .A(n4344), .B(n4345), .ZN(n4340) );
  AOI22_X1 U1750 ( .A1(net644830), .A2(n6389), .B1(n4192), .B2(n4154), .ZN(
        n4342) );
  OAI21_X1 U1749 ( .B1(n612), .B2(n4189), .A(n4342), .ZN(n4341) );
  AOI211_X1 U1748 ( .C1(net644735), .C2(n6390), .A(n4340), .B(n4341), .ZN(
        n4339) );
  NAND4_X1 U1747 ( .A1(n4336), .A2(n4337), .A3(n4338), .A4(n4339), .ZN(n2782)
         );
  AOI22_X1 U1899 ( .A1(n6376), .A2(n4026), .B1(n4243), .B2(n3940), .ZN(n4486)
         );
  AOI22_X1 U1898 ( .A1(net644891), .A2(n6378), .B1(net644857), .B2(n4240), 
        .ZN(n4487) );
  AOI22_X1 U1897 ( .A1(net644473), .A2(n4237), .B1(DATAIN[22]), .B2(n6379), 
        .ZN(n4512) );
  OAI21_X1 U1896 ( .B1(n4235), .B2(net644409), .A(n4512), .ZN(n4510) );
  OAI22_X1 U1895 ( .A1(n649), .A2(n4233), .B1(n524), .B2(n4234), .ZN(n4511) );
  AOI211_X1 U1894 ( .C1(net644665), .C2(n6381), .A(n4510), .B(n4511), .ZN(
        n4488) );
  AOI22_X1 U1893 ( .A1(net644569), .A2(n6382), .B1(net644537), .B2(n4229), 
        .ZN(n4494) );
  AOI22_X1 U1892 ( .A1(n414), .A2(n6383), .B1(n3896), .B2(n4134), .ZN(n4504)
         );
  AOI22_X1 U1891 ( .A1(net644634), .A2(n3895), .B1(net644505), .B2(n4224), 
        .ZN(n4505) );
  AOI22_X1 U1890 ( .A1(n4220), .A2(n362), .B1(n3891), .B2(n4027), .ZN(n4506)
         );
  AOI22_X1 U1889 ( .A1(net644602), .A2(n4218), .B1(net644698), .B2(n3897), 
        .ZN(n4507) );
  NAND4_X1 U1888 ( .A1(n4504), .A2(n4505), .A3(n4506), .A4(n4507), .ZN(n4496)
         );
  AOI22_X1 U1887 ( .A1(n416), .A2(n4211), .B1(n3903), .B2(n4135), .ZN(n4498)
         );
  AOI22_X1 U1886 ( .A1(net644794), .A2(n3902), .B1(net644762), .B2(n4210), 
        .ZN(n4499) );
  AOI22_X1 U1885 ( .A1(net644924), .A2(n3900), .B1(net644441), .B2(n4208), 
        .ZN(n4500) );
  AOI22_X1 U1884 ( .A1(n4204), .A2(n415), .B1(n3898), .B2(n4028), .ZN(n4501)
         );
  NAND4_X1 U1883 ( .A1(n4498), .A2(n4499), .A3(n4500), .A4(n4501), .ZN(n4497)
         );
  OAI21_X1 U1882 ( .B1(n4496), .B2(n4497), .A(n6386), .ZN(n4495) );
  OAI211_X1 U1881 ( .C1(n555), .C2(n4194), .A(n4494), .B(n4495), .ZN(n4490) );
  AOI22_X1 U1880 ( .A1(net644825), .A2(n6389), .B1(n6388), .B2(n4136), .ZN(
        n4492) );
  OAI21_X1 U1879 ( .B1(n617), .B2(n4189), .A(n4492), .ZN(n4491) );
  AOI211_X1 U1878 ( .C1(net644730), .C2(n4186), .A(n4490), .B(n4491), .ZN(
        n4489) );
  NAND4_X1 U1877 ( .A1(n4486), .A2(n4487), .A3(n4488), .A4(n4489), .ZN(n2772)
         );
  AOI22_X1 U1795 ( .A1(n4241), .A2(n4041), .B1(n6375), .B2(n3944), .ZN(n4366)
         );
  AOI22_X1 U1794 ( .A1(net644895), .A2(n6378), .B1(net644861), .B2(n6377), 
        .ZN(n4367) );
  AOI22_X1 U1793 ( .A1(net644477), .A2(n6380), .B1(DATAIN[26]), .B2(n6379), 
        .ZN(n4392) );
  OAI21_X1 U1792 ( .B1(n4235), .B2(net644413), .A(n4392), .ZN(n4390) );
  OAI22_X1 U1791 ( .A1(n645), .A2(n4233), .B1(n520), .B2(n4234), .ZN(n4391) );
  AOI211_X1 U1790 ( .C1(net644669), .C2(n6381), .A(n4390), .B(n4391), .ZN(
        n4368) );
  AOI22_X1 U1789 ( .A1(net644573), .A2(n6382), .B1(net644541), .B2(n3880), 
        .ZN(n4374) );
  AOI22_X1 U1788 ( .A1(n402), .A2(n6383), .B1(n3896), .B2(n4149), .ZN(n4384)
         );
  AOI22_X1 U1787 ( .A1(net644638), .A2(n3895), .B1(net644509), .B2(n3894), 
        .ZN(n4385) );
  AOI22_X1 U1786 ( .A1(n4220), .A2(n358), .B1(n4221), .B2(n4042), .ZN(n4386)
         );
  AOI22_X1 U1785 ( .A1(net644606), .A2(n3890), .B1(net644702), .B2(n3897), 
        .ZN(n4387) );
  NAND4_X1 U1784 ( .A1(n4384), .A2(n4385), .A3(n4386), .A4(n4387), .ZN(n4376)
         );
  AOI22_X1 U1783 ( .A1(n404), .A2(n4211), .B1(n4212), .B2(n4150), .ZN(n4378)
         );
  AOI22_X1 U1782 ( .A1(net644798), .A2(n3902), .B1(net644766), .B2(n3901), 
        .ZN(n4379) );
  AOI22_X1 U1781 ( .A1(net644928), .A2(n3900), .B1(net644445), .B2(n3899), 
        .ZN(n4380) );
  AOI22_X1 U1780 ( .A1(n4204), .A2(n403), .B1(n3898), .B2(n4043), .ZN(n4381)
         );
  NAND4_X1 U1779 ( .A1(n4378), .A2(n4379), .A3(n4380), .A4(n4381), .ZN(n4377)
         );
  OAI21_X1 U1778 ( .B1(n4376), .B2(n4377), .A(n6386), .ZN(n4375) );
  OAI211_X1 U1777 ( .C1(n551), .C2(n4194), .A(n4374), .B(n4375), .ZN(n4370) );
  AOI22_X1 U1776 ( .A1(net644829), .A2(n6389), .B1(n4192), .B2(n4151), .ZN(
        n4372) );
  OAI21_X1 U1775 ( .B1(n613), .B2(n4189), .A(n4372), .ZN(n4371) );
  AOI211_X1 U1774 ( .C1(net644734), .C2(n6390), .A(n4370), .B(n4371), .ZN(
        n4369) );
  NAND4_X1 U1773 ( .A1(n4366), .A2(n4367), .A3(n4368), .A4(n4369), .ZN(n2780)
         );
  AOI22_X1 U3467 ( .A1(n6356), .A2(n3916), .B1(n6355), .B2(n3954), .ZN(n5903)
         );
  AOI22_X1 U3466 ( .A1(n6358), .A2(net644870), .B1(n5262), .B2(net644836), 
        .ZN(n5904) );
  AOI22_X1 U3465 ( .A1(n6360), .A2(net644452), .B1(n6359), .B2(DATAIN[1]), 
        .ZN(n5926) );
  OAI21_X1 U3464 ( .B1(n5257), .B2(net644357), .A(n5926), .ZN(n5923) );
  OAI22_X1 U3462 ( .A1(n545), .A2(n5255), .B1(n670), .B2(n5256), .ZN(n5924) );
  AOI211_X1 U3461 ( .C1(n6361), .C2(net644644), .A(n5923), .B(n5924), .ZN(
        n5905) );
  AOI22_X1 U3460 ( .A1(n6363), .A2(net644516), .B1(n6362), .B2(net644548), 
        .ZN(n5911) );
  AOI22_X1 U3459 ( .A1(n5248), .A2(n477), .B1(n6364), .B2(n222), .ZN(n5919) );
  AOI22_X1 U3458 ( .A1(n3911), .A2(net644613), .B1(n3912), .B2(net644484), 
        .ZN(n5920) );
  AOI22_X1 U3456 ( .A1(n5244), .A2(n3955), .B1(n6366), .B2(n383), .ZN(n5921)
         );
  AOI22_X1 U3455 ( .A1(n3913), .A2(net644581), .B1(n3914), .B2(net644677), 
        .ZN(n5922) );
  NAND4_X1 U3454 ( .A1(n5919), .A2(n5920), .A3(n5921), .A4(n5922), .ZN(n5913)
         );
  AOI22_X1 U3452 ( .A1(n5236), .A2(n479), .B1(n6368), .B2(n4063), .ZN(n5915)
         );
  AOI22_X1 U3451 ( .A1(n3910), .A2(net644773), .B1(n3909), .B2(net644741), 
        .ZN(n5916) );
  AOI22_X1 U3450 ( .A1(n3908), .A2(net644903), .B1(n3907), .B2(net644420), 
        .ZN(n5917) );
  AOI22_X1 U3448 ( .A1(n3906), .A2(n3956), .B1(n3905), .B2(n478), .ZN(n5918)
         );
  NAND4_X1 U3447 ( .A1(n5915), .A2(n5916), .A3(n5917), .A4(n5918), .ZN(n5914)
         );
  OAI21_X1 U3446 ( .B1(n5913), .B2(n5914), .A(n6370), .ZN(n5912) );
  OAI211_X1 U3445 ( .C1(n576), .C2(n5220), .A(n5911), .B(n5912), .ZN(n5907) );
  AOI22_X1 U3442 ( .A1(n6373), .A2(net644804), .B1(n5219), .B2(n4064), .ZN(
        n5909) );
  OAI21_X1 U3441 ( .B1(n638), .B2(n5216), .A(n5909), .ZN(n5908) );
  AOI211_X1 U3440 ( .C1(n6374), .C2(net644709), .A(n5907), .B(n5908), .ZN(
        n5906) );
  NAND4_X1 U3439 ( .A1(n5903), .A2(n5904), .A3(n5905), .A4(n5906), .ZN(n2697)
         );
  AOI22_X1 U3286 ( .A1(n6356), .A2(n3922), .B1(n6355), .B2(n3975), .ZN(n5771)
         );
  AOI22_X1 U3285 ( .A1(n6358), .A2(net644876), .B1(n6357), .B2(net644842), 
        .ZN(n5772) );
  AOI22_X1 U3284 ( .A1(n6360), .A2(net644458), .B1(n6359), .B2(DATAIN[7]), 
        .ZN(n5792) );
  OAI21_X1 U3283 ( .B1(n5257), .B2(net644363), .A(n5792), .ZN(n5790) );
  OAI22_X1 U3282 ( .A1(n539), .A2(n5255), .B1(n664), .B2(n5256), .ZN(n5791) );
  AOI211_X1 U3281 ( .C1(n6361), .C2(net644650), .A(n5790), .B(n5791), .ZN(
        n5773) );
  AOI22_X1 U3280 ( .A1(n6363), .A2(net644522), .B1(n6362), .B2(net644554), 
        .ZN(n5778) );
  AOI22_X1 U3278 ( .A1(n5248), .A2(n459), .B1(n6364), .B2(n4084), .ZN(n5786)
         );
  AOI22_X1 U3277 ( .A1(n3911), .A2(net644619), .B1(n3912), .B2(net644490), 
        .ZN(n5787) );
  AOI22_X1 U3275 ( .A1(n5244), .A2(n3976), .B1(n6366), .B2(n377), .ZN(n5788)
         );
  AOI22_X1 U3274 ( .A1(n3913), .A2(net644587), .B1(n3914), .B2(net644683), 
        .ZN(n5789) );
  NAND4_X1 U3273 ( .A1(n5786), .A2(n5787), .A3(n5788), .A4(n5789), .ZN(n5780)
         );
  AOI22_X1 U3271 ( .A1(n5236), .A2(n461), .B1(n6368), .B2(n4085), .ZN(n5782)
         );
  AOI22_X1 U3270 ( .A1(n3910), .A2(net644779), .B1(n3909), .B2(net644747), 
        .ZN(n5783) );
  AOI22_X1 U3269 ( .A1(n3908), .A2(net644909), .B1(n3907), .B2(net644426), 
        .ZN(n5784) );
  AOI22_X1 U3267 ( .A1(n3906), .A2(n3977), .B1(n3905), .B2(n460), .ZN(n5785)
         );
  NAND4_X1 U3266 ( .A1(n5782), .A2(n5783), .A3(n5784), .A4(n5785), .ZN(n5781)
         );
  OAI21_X1 U3265 ( .B1(n5780), .B2(n5781), .A(n6370), .ZN(n5779) );
  OAI211_X1 U3264 ( .C1(n570), .C2(n5220), .A(n5778), .B(n5779), .ZN(n5775) );
  AOI22_X1 U3262 ( .A1(n6373), .A2(net644810), .B1(n5219), .B2(n4086), .ZN(
        n5777) );
  OAI21_X1 U3261 ( .B1(n632), .B2(n5216), .A(n5777), .ZN(n5776) );
  AOI211_X1 U3260 ( .C1(n6374), .C2(net644715), .A(n5775), .B(n5776), .ZN(
        n5774) );
  NAND4_X1 U3259 ( .A1(n5771), .A2(n5772), .A3(n5773), .A4(n5774), .ZN(n2703)
         );
  AOI22_X1 U3346 ( .A1(n6356), .A2(n3920), .B1(n6355), .B2(n3969), .ZN(n5815)
         );
  AOI22_X1 U3345 ( .A1(n6358), .A2(net644874), .B1(n5262), .B2(net644840), 
        .ZN(n5816) );
  AOI22_X1 U3344 ( .A1(n6360), .A2(net644456), .B1(n6359), .B2(DATAIN[5]), 
        .ZN(n5836) );
  OAI21_X1 U3343 ( .B1(n5257), .B2(net644361), .A(n5836), .ZN(n5834) );
  OAI22_X1 U3342 ( .A1(n541), .A2(n5255), .B1(n666), .B2(n5256), .ZN(n5835) );
  AOI211_X1 U3341 ( .C1(n6361), .C2(net644648), .A(n5834), .B(n5835), .ZN(
        n5817) );
  AOI22_X1 U3340 ( .A1(n6363), .A2(net644520), .B1(n6362), .B2(net644552), 
        .ZN(n5822) );
  AOI22_X1 U3338 ( .A1(n5248), .A2(n465), .B1(n6364), .B2(n4078), .ZN(n5830)
         );
  AOI22_X1 U3337 ( .A1(n3911), .A2(net644617), .B1(n3912), .B2(net644488), 
        .ZN(n5831) );
  AOI22_X1 U3335 ( .A1(n5244), .A2(n3970), .B1(n6366), .B2(n379), .ZN(n5832)
         );
  AOI22_X1 U3334 ( .A1(n3913), .A2(net644585), .B1(n3914), .B2(net644681), 
        .ZN(n5833) );
  NAND4_X1 U3333 ( .A1(n5830), .A2(n5831), .A3(n5832), .A4(n5833), .ZN(n5824)
         );
  AOI22_X1 U3331 ( .A1(n5236), .A2(n467), .B1(n6368), .B2(n4079), .ZN(n5826)
         );
  AOI22_X1 U3330 ( .A1(n3910), .A2(net644777), .B1(n3909), .B2(net644745), 
        .ZN(n5827) );
  AOI22_X1 U3329 ( .A1(n3908), .A2(net644907), .B1(n3907), .B2(net644424), 
        .ZN(n5828) );
  AOI22_X1 U3327 ( .A1(n3906), .A2(n3971), .B1(n3905), .B2(n466), .ZN(n5829)
         );
  NAND4_X1 U3326 ( .A1(n5826), .A2(n5827), .A3(n5828), .A4(n5829), .ZN(n5825)
         );
  OAI21_X1 U3325 ( .B1(n5824), .B2(n5825), .A(n6370), .ZN(n5823) );
  OAI211_X1 U3324 ( .C1(n572), .C2(n5220), .A(n5822), .B(n5823), .ZN(n5819) );
  AOI22_X1 U3322 ( .A1(n6373), .A2(net644808), .B1(n5219), .B2(n4080), .ZN(
        n5821) );
  OAI21_X1 U3321 ( .B1(n634), .B2(n5216), .A(n5821), .ZN(n5820) );
  AOI211_X1 U3320 ( .C1(n6374), .C2(net644713), .A(n5819), .B(n5820), .ZN(
        n5818) );
  NAND4_X1 U3319 ( .A1(n5815), .A2(n5816), .A3(n5817), .A4(n5818), .ZN(n2701)
         );
  AOI22_X1 U3376 ( .A1(n6356), .A2(n3919), .B1(n6355), .B2(n3966), .ZN(n5837)
         );
  AOI22_X1 U3375 ( .A1(n6358), .A2(net644873), .B1(n5262), .B2(net644839), 
        .ZN(n5838) );
  AOI22_X1 U3374 ( .A1(n6360), .A2(net644455), .B1(n6359), .B2(DATAIN[4]), 
        .ZN(n5858) );
  OAI21_X1 U3373 ( .B1(n5257), .B2(net644360), .A(n5858), .ZN(n5856) );
  OAI22_X1 U3372 ( .A1(n542), .A2(n5255), .B1(n667), .B2(n5256), .ZN(n5857) );
  AOI211_X1 U3371 ( .C1(n6361), .C2(net644647), .A(n5856), .B(n5857), .ZN(
        n5839) );
  AOI22_X1 U3370 ( .A1(n6363), .A2(net644519), .B1(n6362), .B2(net644551), 
        .ZN(n5844) );
  AOI22_X1 U3368 ( .A1(n5248), .A2(n468), .B1(n6364), .B2(n4075), .ZN(n5852)
         );
  AOI22_X1 U3367 ( .A1(n3911), .A2(net644616), .B1(n3912), .B2(net644487), 
        .ZN(n5853) );
  AOI22_X1 U3365 ( .A1(n5244), .A2(n3967), .B1(n6366), .B2(n380), .ZN(n5854)
         );
  AOI22_X1 U3364 ( .A1(n3913), .A2(net644584), .B1(n3914), .B2(net644680), 
        .ZN(n5855) );
  NAND4_X1 U3363 ( .A1(n5852), .A2(n5853), .A3(n5854), .A4(n5855), .ZN(n5846)
         );
  AOI22_X1 U3361 ( .A1(n5236), .A2(n470), .B1(n6368), .B2(n4076), .ZN(n5848)
         );
  AOI22_X1 U3360 ( .A1(n3910), .A2(net644776), .B1(n3909), .B2(net644744), 
        .ZN(n5849) );
  AOI22_X1 U3359 ( .A1(n3908), .A2(net644906), .B1(n3907), .B2(net644423), 
        .ZN(n5850) );
  AOI22_X1 U3357 ( .A1(n3906), .A2(n3968), .B1(n3905), .B2(n469), .ZN(n5851)
         );
  NAND4_X1 U3356 ( .A1(n5848), .A2(n5849), .A3(n5850), .A4(n5851), .ZN(n5847)
         );
  OAI21_X1 U3355 ( .B1(n5846), .B2(n5847), .A(n6370), .ZN(n5845) );
  OAI211_X1 U3354 ( .C1(n573), .C2(n5220), .A(n5844), .B(n5845), .ZN(n5841) );
  AOI22_X1 U3352 ( .A1(n6373), .A2(net644807), .B1(n5219), .B2(n4077), .ZN(
        n5843) );
  OAI21_X1 U3351 ( .B1(n635), .B2(n5216), .A(n5843), .ZN(n5842) );
  AOI211_X1 U3350 ( .C1(n6374), .C2(net644712), .A(n5841), .B(n5842), .ZN(
        n5840) );
  NAND4_X1 U3349 ( .A1(n5837), .A2(n5838), .A3(n5839), .A4(n5840), .ZN(n2700)
         );
  AOI22_X1 U2716 ( .A1(n6356), .A2(n3944), .B1(n5264), .B2(n4041), .ZN(n5353)
         );
  AOI22_X1 U2715 ( .A1(n6358), .A2(net644895), .B1(n5262), .B2(net644861), 
        .ZN(n5354) );
  AOI22_X1 U2714 ( .A1(n5259), .A2(net644477), .B1(n5260), .B2(DATAIN[26]), 
        .ZN(n5374) );
  OAI21_X1 U2713 ( .B1(n5257), .B2(net644382), .A(n5374), .ZN(n5372) );
  OAI22_X1 U2712 ( .A1(n520), .A2(n5255), .B1(n645), .B2(n5256), .ZN(n5373) );
  AOI211_X1 U2711 ( .C1(n6361), .C2(net644669), .A(n5372), .B(n5373), .ZN(
        n5355) );
  AOI22_X1 U2710 ( .A1(n5250), .A2(net644541), .B1(n5251), .B2(net644573), 
        .ZN(n5360) );
  AOI22_X1 U2708 ( .A1(n5248), .A2(n402), .B1(n5249), .B2(n4149), .ZN(n5368)
         );
  AOI22_X1 U2707 ( .A1(n5246), .A2(net644638), .B1(n5247), .B2(net644509), 
        .ZN(n5369) );
  AOI22_X1 U2705 ( .A1(n5244), .A2(n4042), .B1(n5245), .B2(n358), .ZN(n5370)
         );
  AOI22_X1 U2704 ( .A1(n5242), .A2(net644606), .B1(n5243), .B2(net644702), 
        .ZN(n5371) );
  NAND4_X1 U2703 ( .A1(n5368), .A2(n5369), .A3(n5370), .A4(n5371), .ZN(n5362)
         );
  AOI22_X1 U2701 ( .A1(n5236), .A2(n404), .B1(n5237), .B2(n4150), .ZN(n5364)
         );
  AOI22_X1 U2700 ( .A1(n5234), .A2(net644798), .B1(n5235), .B2(net644766), 
        .ZN(n5365) );
  AOI22_X1 U2699 ( .A1(n5232), .A2(net644928), .B1(n5233), .B2(net644445), 
        .ZN(n5366) );
  AOI22_X1 U2697 ( .A1(n5230), .A2(n4043), .B1(n5231), .B2(n403), .ZN(n5367)
         );
  NAND4_X1 U2696 ( .A1(n5364), .A2(n5365), .A3(n5366), .A4(n5367), .ZN(n5363)
         );
  OAI21_X1 U2695 ( .B1(n5362), .B2(n5363), .A(n6370), .ZN(n5361) );
  OAI211_X1 U2694 ( .C1(n551), .C2(n5220), .A(n5360), .B(n5361), .ZN(n5357) );
  AOI22_X1 U2692 ( .A1(n6373), .A2(net644829), .B1(n5219), .B2(n4151), .ZN(
        n5359) );
  OAI21_X1 U2691 ( .B1(n613), .B2(n5216), .A(n5359), .ZN(n5358) );
  AOI211_X1 U2690 ( .C1(n5213), .C2(net644734), .A(n5357), .B(n5358), .ZN(
        n5356) );
  NAND4_X1 U2689 ( .A1(n5353), .A2(n5354), .A3(n5355), .A4(n5356), .ZN(n2722)
         );
  OAI22_X1 U496 ( .A1(n5063), .A2(n6431), .B1(n1688), .B2(n6430), .ZN(n3451)
         );
  OAI22_X1 U484 ( .A1(n5084), .A2(n1885), .B1(n1676), .B2(n6430), .ZN(n3457)
         );
  OAI22_X1 U431 ( .A1(n5252), .A2(n6433), .B1(n1688), .B2(n6432), .ZN(n3483)
         );
  OAI22_X1 U518 ( .A1(n5023), .A2(n6431), .B1(n1710), .B2(n6430), .ZN(n3440)
         );
  OAI22_X1 U478 ( .A1(n5102), .A2(n1885), .B1(n1670), .B2(n6430), .ZN(n3460)
         );
  OAI22_X1 U453 ( .A1(n5144), .A2(n6433), .B1(n1710), .B2(n6432), .ZN(n3472)
         );
  OAI22_X1 U498 ( .A1(n5055), .A2(n6431), .B1(n1690), .B2(n6430), .ZN(n3450)
         );
  OAI22_X1 U502 ( .A1(n5053), .A2(n6431), .B1(n1694), .B2(n6430), .ZN(n3448)
         );
  OAI22_X1 U486 ( .A1(n5083), .A2(n1885), .B1(n1678), .B2(n6430), .ZN(n3456)
         );
  OAI22_X1 U506 ( .A1(n5048), .A2(n6431), .B1(n1698), .B2(n6430), .ZN(n3446)
         );
  OAI22_X1 U445 ( .A1(n5180), .A2(n6433), .B1(n1702), .B2(n6432), .ZN(n3476)
         );
  OAI22_X1 U516 ( .A1(n5024), .A2(n6431), .B1(n1708), .B2(n6430), .ZN(n3441)
         );
  OAI22_X1 U441 ( .A1(n5188), .A2(n6433), .B1(n1698), .B2(n6432), .ZN(n3478)
         );
  OAI22_X1 U451 ( .A1(n5145), .A2(n6433), .B1(n1708), .B2(n6432), .ZN(n3473)
         );
  OAI22_X1 U439 ( .A1(n5193), .A2(n6433), .B1(n1696), .B2(n6432), .ZN(n3479)
         );
  OAI22_X1 U500 ( .A1(n5054), .A2(n6431), .B1(n1692), .B2(n6430), .ZN(n3449)
         );
  OAI22_X1 U512 ( .A1(n5033), .A2(n6431), .B1(n1704), .B2(n6430), .ZN(n3443)
         );
  OAI22_X1 U474 ( .A1(n5108), .A2(n6431), .B1(n1666), .B2(n6430), .ZN(n3462)
         );
  OAI22_X1 U443 ( .A1(n5183), .A2(n6433), .B1(n1700), .B2(n6432), .ZN(n3477)
         );
  OAI22_X1 U476 ( .A1(n5103), .A2(n1885), .B1(n1668), .B2(n6430), .ZN(n3461)
         );
  OAI22_X1 U504 ( .A1(n5049), .A2(n6431), .B1(n1696), .B2(n6430), .ZN(n3447)
         );
  OAI22_X1 U435 ( .A1(n5204), .A2(n6433), .B1(n1692), .B2(n6432), .ZN(n3481)
         );
  OAI22_X1 U514 ( .A1(n5025), .A2(n6431), .B1(n1706), .B2(n6430), .ZN(n3442)
         );
  OAI22_X1 U411 ( .A1(n5991), .A2(n1852), .B1(n1668), .B2(n6432), .ZN(n3493)
         );
  OAI22_X1 U510 ( .A1(n5042), .A2(n6431), .B1(n1702), .B2(n6430), .ZN(n3444)
         );
  OAI22_X1 U508 ( .A1(n5043), .A2(n6431), .B1(n1700), .B2(n6430), .ZN(n3445)
         );
  OAI22_X1 U413 ( .A1(n5990), .A2(n1852), .B1(n1670), .B2(n6432), .ZN(n3492)
         );
  OAI22_X1 U421 ( .A1(n5986), .A2(n1852), .B1(n1678), .B2(n6432), .ZN(n3488)
         );
  OAI22_X1 U449 ( .A1(n5153), .A2(n6433), .B1(n1706), .B2(n6432), .ZN(n3474)
         );
  OAI22_X1 U447 ( .A1(n5174), .A2(n6433), .B1(n1704), .B2(n6432), .ZN(n3475)
         );
  OAI22_X1 U437 ( .A1(n5203), .A2(n6433), .B1(n1694), .B2(n6432), .ZN(n3480)
         );
  OAI22_X1 U433 ( .A1(n5218), .A2(n6433), .B1(n1690), .B2(n6432), .ZN(n3482)
         );
  OAI22_X1 U409 ( .A1(n5992), .A2(n6433), .B1(n1666), .B2(n6432), .ZN(n3494)
         );
  OAI22_X1 U419 ( .A1(n5987), .A2(n1852), .B1(n1676), .B2(n6432), .ZN(n3489)
         );
  OAI22_X1 U469 ( .A1(n2601), .A2(n6433), .B1(n6432), .B2(n1726), .ZN(n3464)
         );
  OAI22_X1 U534 ( .A1(n481), .A2(n6431), .B1(n6430), .B2(n1726), .ZN(n3432) );
  OAI22_X1 U1444 ( .A1(n6223), .A2(n6400), .B1(n1702), .B2(n6399), .ZN(n2900)
         );
  OAI22_X1 U1436 ( .A1(n6227), .A2(n6400), .B1(n1694), .B2(n6399), .ZN(n2904)
         );
  OAI22_X1 U1456 ( .A1(n6217), .A2(n6400), .B1(n1714), .B2(n6399), .ZN(n2894)
         );
  OAI22_X1 U1438 ( .A1(n6226), .A2(n6400), .B1(n1696), .B2(n6399), .ZN(n2903)
         );
  OAI22_X1 U1440 ( .A1(n6225), .A2(n6400), .B1(n1698), .B2(n6399), .ZN(n2902)
         );
  OAI22_X1 U1466 ( .A1(n6212), .A2(n6400), .B1(n1724), .B2(n6399), .ZN(n2889)
         );
  OAI22_X1 U1452 ( .A1(n6219), .A2(n6400), .B1(n1710), .B2(n6399), .ZN(n2896)
         );
  OAI22_X1 U1442 ( .A1(n6224), .A2(n6400), .B1(n1700), .B2(n6399), .ZN(n2901)
         );
  OAI22_X1 U1364 ( .A1(n6150), .A2(n6403), .B1(n1724), .B2(n6402), .ZN(n2953)
         );
  OAI22_X1 U1362 ( .A1(n6151), .A2(n6403), .B1(n1722), .B2(n6402), .ZN(n2954)
         );
  OAI22_X1 U1360 ( .A1(n6152), .A2(n6403), .B1(n1720), .B2(n6402), .ZN(n2955)
         );
  OAI22_X1 U1354 ( .A1(n6155), .A2(n6403), .B1(n1714), .B2(n6402), .ZN(n2958)
         );
  OAI22_X1 U1352 ( .A1(n6156), .A2(n6403), .B1(n1712), .B2(n6402), .ZN(n2959)
         );
  OAI22_X1 U1350 ( .A1(n6157), .A2(n6403), .B1(n1710), .B2(n6402), .ZN(n2960)
         );
  OAI22_X1 U1430 ( .A1(n6230), .A2(n6400), .B1(n1688), .B2(n6399), .ZN(n2907)
         );
  OAI22_X1 U1454 ( .A1(n6218), .A2(n6400), .B1(n1712), .B2(n6399), .ZN(n2895)
         );
  OAI22_X1 U1434 ( .A1(n6228), .A2(n6400), .B1(n1692), .B2(n6399), .ZN(n2905)
         );
  OAI22_X1 U1432 ( .A1(n6229), .A2(n6400), .B1(n1690), .B2(n6399), .ZN(n2906)
         );
  OAI22_X1 U1462 ( .A1(n6214), .A2(n6400), .B1(n1720), .B2(n6399), .ZN(n2891)
         );
  OAI22_X1 U1428 ( .A1(n6231), .A2(n6400), .B1(n1686), .B2(n6399), .ZN(n2908)
         );
  OAI22_X1 U1426 ( .A1(n6232), .A2(n6400), .B1(n1684), .B2(n6399), .ZN(n2909)
         );
  OAI22_X1 U1424 ( .A1(n6233), .A2(n6400), .B1(n1682), .B2(n6399), .ZN(n2910)
         );
  OAI22_X1 U1422 ( .A1(n6234), .A2(n4073), .B1(n1680), .B2(n6399), .ZN(n2911)
         );
  OAI22_X1 U1342 ( .A1(n6161), .A2(n6403), .B1(n1702), .B2(n6402), .ZN(n2964)
         );
  OAI22_X1 U1464 ( .A1(n6213), .A2(n6400), .B1(n1722), .B2(n6399), .ZN(n2890)
         );
  OAI22_X1 U1320 ( .A1(n6172), .A2(n4035), .B1(n1680), .B2(n6402), .ZN(n2975)
         );
  OAI22_X1 U1340 ( .A1(n6162), .A2(n6403), .B1(n1700), .B2(n6402), .ZN(n2965)
         );
  OAI22_X1 U1322 ( .A1(n6171), .A2(n6403), .B1(n1682), .B2(n6402), .ZN(n2974)
         );
  OAI22_X1 U1338 ( .A1(n6163), .A2(n6403), .B1(n1698), .B2(n6402), .ZN(n2966)
         );
  OAI22_X1 U1324 ( .A1(n6170), .A2(n6403), .B1(n1684), .B2(n6402), .ZN(n2973)
         );
  OAI22_X1 U1326 ( .A1(n6169), .A2(n6403), .B1(n1686), .B2(n6402), .ZN(n2972)
         );
  OAI22_X1 U1328 ( .A1(n6168), .A2(n6403), .B1(n1688), .B2(n6402), .ZN(n2971)
         );
  OAI22_X1 U1330 ( .A1(n6167), .A2(n6403), .B1(n1690), .B2(n6402), .ZN(n2970)
         );
  OAI22_X1 U1332 ( .A1(n6166), .A2(n6403), .B1(n1692), .B2(n6402), .ZN(n2969)
         );
  OAI22_X1 U1334 ( .A1(n6165), .A2(n6403), .B1(n1694), .B2(n6402), .ZN(n2968)
         );
  OAI22_X1 U1336 ( .A1(n6164), .A2(n6403), .B1(n1696), .B2(n6402), .ZN(n2967)
         );
  OAI22_X1 U1256 ( .A1(n6140), .A2(n6405), .B1(n1682), .B2(n6404), .ZN(n3006)
         );
  OAI22_X1 U1274 ( .A1(n6131), .A2(n6405), .B1(n1700), .B2(n6404), .ZN(n2997)
         );
  OAI22_X1 U1272 ( .A1(n6132), .A2(n6405), .B1(n1698), .B2(n6404), .ZN(n2998)
         );
  OAI22_X1 U1270 ( .A1(n6133), .A2(n6405), .B1(n1696), .B2(n6404), .ZN(n2999)
         );
  OAI22_X1 U1268 ( .A1(n6134), .A2(n6405), .B1(n1694), .B2(n6404), .ZN(n3000)
         );
  OAI22_X1 U1300 ( .A1(n6349), .A2(n6405), .B1(n1726), .B2(n6404), .ZN(n2984)
         );
  OAI22_X1 U1266 ( .A1(n6135), .A2(n6405), .B1(n1692), .B2(n6404), .ZN(n3001)
         );
  OAI22_X1 U1296 ( .A1(n6120), .A2(n6405), .B1(n1722), .B2(n6404), .ZN(n2986)
         );
  OAI22_X1 U1262 ( .A1(n6137), .A2(n6405), .B1(n1688), .B2(n6404), .ZN(n3003)
         );
  OAI22_X1 U1294 ( .A1(n6121), .A2(n6405), .B1(n1720), .B2(n6404), .ZN(n2987)
         );
  OAI22_X1 U1258 ( .A1(n6139), .A2(n6405), .B1(n1684), .B2(n6404), .ZN(n3005)
         );
  OAI22_X1 U1254 ( .A1(n6141), .A2(n4000), .B1(n1680), .B2(n6404), .ZN(n3007)
         );
  OAI22_X1 U1260 ( .A1(n6138), .A2(n6405), .B1(n1686), .B2(n6404), .ZN(n3004)
         );
  OAI22_X1 U1288 ( .A1(n6124), .A2(n6405), .B1(n1714), .B2(n6404), .ZN(n2990)
         );
  OAI22_X1 U1284 ( .A1(n6126), .A2(n6405), .B1(n1710), .B2(n6404), .ZN(n2992)
         );
  OAI22_X1 U1286 ( .A1(n6125), .A2(n6405), .B1(n1712), .B2(n6404), .ZN(n2991)
         );
  OAI22_X1 U1276 ( .A1(n6130), .A2(n6405), .B1(n1702), .B2(n6404), .ZN(n2996)
         );
  OAI22_X1 U1264 ( .A1(n6136), .A2(n6405), .B1(n1690), .B2(n6404), .ZN(n3002)
         );
  OAI22_X1 U308 ( .A1(n6318), .A2(n6437), .B1(n1700), .B2(n6436), .ZN(n3573)
         );
  OAI22_X1 U304 ( .A1(n6320), .A2(n6437), .B1(n1696), .B2(n6436), .ZN(n3575)
         );
  OAI22_X1 U274 ( .A1(n6335), .A2(n6437), .B1(n1666), .B2(n6436), .ZN(n3590)
         );
  OAI22_X1 U318 ( .A1(n6313), .A2(n6437), .B1(n1710), .B2(n6436), .ZN(n3568)
         );
  OAI22_X1 U316 ( .A1(n6314), .A2(n6437), .B1(n1708), .B2(n6436), .ZN(n3569)
         );
  OAI22_X1 U314 ( .A1(n6315), .A2(n6437), .B1(n1706), .B2(n6436), .ZN(n3570)
         );
  OAI22_X1 U300 ( .A1(n6322), .A2(n6437), .B1(n1692), .B2(n6436), .ZN(n3577)
         );
  OAI22_X1 U312 ( .A1(n6316), .A2(n6437), .B1(n1704), .B2(n6436), .ZN(n3571)
         );
  OAI22_X1 U306 ( .A1(n6319), .A2(n6437), .B1(n1698), .B2(n6436), .ZN(n3574)
         );
  OAI22_X1 U278 ( .A1(n6333), .A2(n1811), .B1(n1670), .B2(n6436), .ZN(n3588)
         );
  OAI22_X1 U302 ( .A1(n6321), .A2(n6437), .B1(n1694), .B2(n6436), .ZN(n3576)
         );
  OAI22_X1 U286 ( .A1(n6329), .A2(n1811), .B1(n1678), .B2(n6436), .ZN(n3584)
         );
  OAI22_X1 U310 ( .A1(n6317), .A2(n6437), .B1(n1702), .B2(n6436), .ZN(n3572)
         );
  OAI22_X1 U296 ( .A1(n6324), .A2(n6437), .B1(n1688), .B2(n6436), .ZN(n3579)
         );
  OAI22_X1 U284 ( .A1(n6330), .A2(n1811), .B1(n1676), .B2(n6436), .ZN(n3585)
         );
  OAI22_X1 U298 ( .A1(n6323), .A2(n6437), .B1(n1690), .B2(n6436), .ZN(n3578)
         );
  OAI22_X1 U276 ( .A1(n6334), .A2(n1811), .B1(n1668), .B2(n6436), .ZN(n3589)
         );
  OAI22_X1 U334 ( .A1(n480), .A2(n6437), .B1(n6436), .B2(n1726), .ZN(n3560) );
  NAND2_X1 U169 ( .A1(n1769), .A2(n1770), .ZN(n1729) );
  OAI22_X1 U31 ( .A1(n6041), .A2(n6445), .B1(n1692), .B2(n6444), .ZN(n3737) );
  OAI22_X1 U37 ( .A1(n6038), .A2(n6445), .B1(n1698), .B2(n6444), .ZN(n3734) );
  OAI22_X1 U33 ( .A1(n6040), .A2(n6445), .B1(n1694), .B2(n6444), .ZN(n3736) );
  OAI22_X1 U63 ( .A1(n6025), .A2(n6445), .B1(n1724), .B2(n6444), .ZN(n3721) );
  OAI22_X1 U25 ( .A1(n6044), .A2(n6445), .B1(n1686), .B2(n6444), .ZN(n3740) );
  OAI22_X1 U61 ( .A1(n6026), .A2(n6445), .B1(n1722), .B2(n6444), .ZN(n3722) );
  OAI22_X1 U21 ( .A1(n6046), .A2(n6445), .B1(n1682), .B2(n6444), .ZN(n3742) );
  OAI22_X1 U35 ( .A1(n6039), .A2(n6445), .B1(n1696), .B2(n6444), .ZN(n3735) );
  OAI22_X1 U23 ( .A1(n6045), .A2(n6445), .B1(n1684), .B2(n6444), .ZN(n3741) );
  OAI22_X1 U27 ( .A1(n6043), .A2(n6445), .B1(n1688), .B2(n6444), .ZN(n3739) );
  OAI22_X1 U49 ( .A1(n6032), .A2(n6445), .B1(n1710), .B2(n6444), .ZN(n3728) );
  OAI22_X1 U41 ( .A1(n6036), .A2(n6445), .B1(n1702), .B2(n6444), .ZN(n3732) );
  OAI22_X1 U29 ( .A1(n6042), .A2(n6445), .B1(n1690), .B2(n6444), .ZN(n3738) );
  OAI22_X1 U39 ( .A1(n6037), .A2(n6445), .B1(n1700), .B2(n6444), .ZN(n3733) );
  OAI22_X1 U53 ( .A1(n6030), .A2(n6445), .B1(n1714), .B2(n6444), .ZN(n3726) );
  OAI22_X1 U59 ( .A1(n6027), .A2(n6445), .B1(n1720), .B2(n6444), .ZN(n3723) );
  OAI22_X1 U19 ( .A1(n6047), .A2(n1662), .B1(n1680), .B2(n6444), .ZN(n3743) );
  OAI22_X1 U51 ( .A1(n6031), .A2(n6445), .B1(n1712), .B2(n6444), .ZN(n3727) );
  OAI22_X1 U565 ( .A1(n510), .A2(n6429), .B1(n6428), .B2(n1720), .ZN(n3403) );
  OAI22_X1 U552 ( .A1(n497), .A2(n6429), .B1(n6428), .B2(n1694), .ZN(n3416) );
  OAI22_X1 U557 ( .A1(n502), .A2(n6429), .B1(n6428), .B2(n1704), .ZN(n3411) );
  OAI22_X1 U547 ( .A1(n492), .A2(n6429), .B1(n6428), .B2(n1684), .ZN(n3421) );
  OAI22_X1 U549 ( .A1(n494), .A2(n6429), .B1(n6428), .B2(n1688), .ZN(n3419) );
  OAI22_X1 U562 ( .A1(n507), .A2(n6429), .B1(n6428), .B2(n1714), .ZN(n3406) );
  OAI22_X1 U554 ( .A1(n499), .A2(n6429), .B1(n6428), .B2(n1698), .ZN(n3414) );
  OAI22_X1 U550 ( .A1(n495), .A2(n6429), .B1(n6428), .B2(n1690), .ZN(n3418) );
  OAI22_X1 U553 ( .A1(n498), .A2(n6429), .B1(n6428), .B2(n1696), .ZN(n3415) );
  OAI22_X1 U548 ( .A1(n493), .A2(n6429), .B1(n6428), .B2(n1686), .ZN(n3420) );
  OAI22_X1 U545 ( .A1(n490), .A2(n1917), .B1(n6428), .B2(n1680), .ZN(n3423) );
  OAI22_X1 U560 ( .A1(n505), .A2(n6429), .B1(n6428), .B2(n1710), .ZN(n3408) );
  OAI22_X1 U561 ( .A1(n506), .A2(n6429), .B1(n6428), .B2(n1712), .ZN(n3407) );
  OAI22_X1 U546 ( .A1(n491), .A2(n6429), .B1(n6428), .B2(n1682), .ZN(n3422) );
  OAI22_X1 U555 ( .A1(n500), .A2(n6429), .B1(n6428), .B2(n1700), .ZN(n3413) );
  OAI22_X1 U556 ( .A1(n501), .A2(n6429), .B1(n6428), .B2(n1702), .ZN(n3412) );
  OAI22_X1 U566 ( .A1(n511), .A2(n6429), .B1(n6428), .B2(n1722), .ZN(n3402) );
  OAI22_X1 U551 ( .A1(n496), .A2(n6429), .B1(n6428), .B2(n1692), .ZN(n3417) );
  OAI22_X1 U195 ( .A1(n4364), .A2(n6440), .B1(n1688), .B2(n6439), .ZN(n3643)
         );
  OAI22_X1 U199 ( .A1(n4359), .A2(n6440), .B1(n1692), .B2(n6439), .ZN(n3641)
         );
  OAI22_X1 U227 ( .A1(n4304), .A2(n6440), .B1(n1720), .B2(n6439), .ZN(n3627)
         );
  OAI22_X1 U191 ( .A1(n4373), .A2(n6440), .B1(n1684), .B2(n6439), .ZN(n3645)
         );
  OAI22_X1 U193 ( .A1(n4365), .A2(n6440), .B1(n1686), .B2(n6439), .ZN(n3644)
         );
  OAI22_X1 U201 ( .A1(n4358), .A2(n6440), .B1(n1694), .B2(n6439), .ZN(n3640)
         );
  OAI22_X1 U221 ( .A1(n4322), .A2(n6440), .B1(n1714), .B2(n6439), .ZN(n3630)
         );
  OAI22_X1 U203 ( .A1(n4353), .A2(n6440), .B1(n1696), .B2(n6439), .ZN(n3639)
         );
  OAI22_X1 U197 ( .A1(n4363), .A2(n6440), .B1(n1690), .B2(n6439), .ZN(n3642)
         );
  OAI22_X1 U205 ( .A1(n4352), .A2(n6440), .B1(n1698), .B2(n6439), .ZN(n3638)
         );
  OAI22_X1 U219 ( .A1(n4323), .A2(n6440), .B1(n1712), .B2(n6439), .ZN(n3631)
         );
  OAI22_X1 U217 ( .A1(n4328), .A2(n6440), .B1(n1710), .B2(n6439), .ZN(n3632)
         );
  OAI22_X1 U189 ( .A1(n4382), .A2(n6440), .B1(n1682), .B2(n6439), .ZN(n3646)
         );
  OAI22_X1 U233 ( .A1(n6353), .A2(n6440), .B1(n1726), .B2(n6439), .ZN(n3624)
         );
  OAI22_X1 U209 ( .A1(n4335), .A2(n6440), .B1(n1702), .B2(n6439), .ZN(n3636)
         );
  OAI22_X1 U187 ( .A1(n4383), .A2(n1772), .B1(n1680), .B2(n6439), .ZN(n3647)
         );
  OAI22_X1 U207 ( .A1(n4343), .A2(n6440), .B1(n1700), .B2(n6439), .ZN(n3637)
         );
  OAI22_X1 U229 ( .A1(n4303), .A2(n6440), .B1(n1722), .B2(n6439), .ZN(n3626)
         );
  OAI22_X1 U1536 ( .A1(n4592), .A2(n6396), .B1(n1694), .B2(n6395), .ZN(n2840)
         );
  OAI22_X1 U1542 ( .A1(n4574), .A2(n6396), .B1(n1700), .B2(n6395), .ZN(n2837)
         );
  OAI22_X1 U1534 ( .A1(n4593), .A2(n6396), .B1(n1692), .B2(n6395), .ZN(n2841)
         );
  OAI22_X1 U1532 ( .A1(n4598), .A2(n6396), .B1(n1690), .B2(n6395), .ZN(n2842)
         );
  OAI22_X1 U1544 ( .A1(n4573), .A2(n6396), .B1(n1702), .B2(n6395), .ZN(n2836)
         );
  OAI22_X1 U1528 ( .A1(n4603), .A2(n6396), .B1(n1686), .B2(n6395), .ZN(n2844)
         );
  OAI22_X1 U1530 ( .A1(n4599), .A2(n6396), .B1(n1688), .B2(n6395), .ZN(n2843)
         );
  OAI22_X1 U1562 ( .A1(n4539), .A2(n6396), .B1(n1720), .B2(n6395), .ZN(n2827)
         );
  OAI22_X1 U1538 ( .A1(n4583), .A2(n6396), .B1(n1696), .B2(n6395), .ZN(n2839)
         );
  OAI22_X1 U1526 ( .A1(n4604), .A2(n6396), .B1(n1684), .B2(n6395), .ZN(n2845)
         );
  OAI22_X1 U1546 ( .A1(n4569), .A2(n6396), .B1(n1704), .B2(n6395), .ZN(n2835)
         );
  OAI22_X1 U1540 ( .A1(n4575), .A2(n6396), .B1(n1698), .B2(n6395), .ZN(n2838)
         );
  OAI22_X1 U1556 ( .A1(n4545), .A2(n6396), .B1(n1714), .B2(n6395), .ZN(n2830)
         );
  OAI22_X1 U1522 ( .A1(n4613), .A2(n4110), .B1(n1680), .B2(n6395), .ZN(n2847)
         );
  OAI22_X1 U1554 ( .A1(n4553), .A2(n6396), .B1(n1712), .B2(n6395), .ZN(n2831)
         );
  OAI22_X1 U1552 ( .A1(n4562), .A2(n6396), .B1(n1710), .B2(n6395), .ZN(n2832)
         );
  OAI22_X1 U1524 ( .A1(n4605), .A2(n6396), .B1(n1682), .B2(n6395), .ZN(n2846)
         );
  OAI22_X1 U1564 ( .A1(n4538), .A2(n6396), .B1(n1722), .B2(n6395), .ZN(n2826)
         );
  OAI22_X1 U1075 ( .A1(n4808), .A2(n6412), .B1(n1702), .B2(n6411), .ZN(n3124)
         );
  OAI22_X1 U1071 ( .A1(n4813), .A2(n6412), .B1(n1698), .B2(n6411), .ZN(n3126)
         );
  OAI22_X1 U1073 ( .A1(n4809), .A2(n6412), .B1(n1700), .B2(n6411), .ZN(n3125)
         );
  OAI22_X1 U1069 ( .A1(n4814), .A2(n6412), .B1(n1696), .B2(n6411), .ZN(n3127)
         );
  OAI22_X1 U1067 ( .A1(n4815), .A2(n6412), .B1(n1694), .B2(n6411), .ZN(n3128)
         );
  OAI22_X1 U1065 ( .A1(n4823), .A2(n6412), .B1(n1692), .B2(n6411), .ZN(n3129)
         );
  OAI22_X1 U1055 ( .A1(n4843), .A2(n6412), .B1(n1682), .B2(n6411), .ZN(n3134)
         );
  OAI22_X1 U1063 ( .A1(n4832), .A2(n6412), .B1(n1690), .B2(n6411), .ZN(n3130)
         );
  OAI22_X1 U1061 ( .A1(n4833), .A2(n6412), .B1(n1688), .B2(n6411), .ZN(n3131)
         );
  OAI22_X1 U1059 ( .A1(n4838), .A2(n6412), .B1(n1686), .B2(n6411), .ZN(n3132)
         );
  OAI22_X1 U1095 ( .A1(n4772), .A2(n6412), .B1(n1722), .B2(n6411), .ZN(n3114)
         );
  OAI22_X1 U1057 ( .A1(n4839), .A2(n6412), .B1(n1684), .B2(n6411), .ZN(n3133)
         );
  OAI22_X1 U1087 ( .A1(n4783), .A2(n6412), .B1(n1714), .B2(n6411), .ZN(n3118)
         );
  OAI22_X1 U1053 ( .A1(n4844), .A2(n3926), .B1(n1680), .B2(n6411), .ZN(n3135)
         );
  OAI22_X1 U1083 ( .A1(n4785), .A2(n6412), .B1(n1710), .B2(n6411), .ZN(n3120)
         );
  OAI22_X1 U1085 ( .A1(n4784), .A2(n6412), .B1(n1712), .B2(n6411), .ZN(n3119)
         );
  OAI22_X1 U1097 ( .A1(n4763), .A2(n6412), .B1(n1724), .B2(n6411), .ZN(n3113)
         );
  OAI22_X1 U1093 ( .A1(n4773), .A2(n6412), .B1(n1720), .B2(n6411), .ZN(n3115)
         );
  OAI22_X1 U667 ( .A1(n6290), .A2(n6425), .B1(n1694), .B2(n6424), .ZN(n3352)
         );
  OAI22_X1 U653 ( .A1(n6297), .A2(n1956), .B1(n1680), .B2(n6424), .ZN(n3359)
         );
  OAI22_X1 U657 ( .A1(n6295), .A2(n6425), .B1(n1684), .B2(n6424), .ZN(n3357)
         );
  OAI22_X1 U655 ( .A1(n6296), .A2(n6425), .B1(n1682), .B2(n6424), .ZN(n3358)
         );
  OAI22_X1 U659 ( .A1(n6294), .A2(n6425), .B1(n1686), .B2(n6424), .ZN(n3356)
         );
  OAI22_X1 U753 ( .A1(n6093), .A2(n6423), .B1(n1714), .B2(n6422), .ZN(n3310)
         );
  OAI22_X1 U661 ( .A1(n6293), .A2(n6425), .B1(n1688), .B2(n6424), .ZN(n3355)
         );
  OAI22_X1 U669 ( .A1(n6289), .A2(n6425), .B1(n1696), .B2(n6424), .ZN(n3351)
         );
  OAI22_X1 U671 ( .A1(n6288), .A2(n6425), .B1(n1698), .B2(n6424), .ZN(n3350)
         );
  OAI22_X1 U739 ( .A1(n6100), .A2(n6423), .B1(n1700), .B2(n6422), .ZN(n3317)
         );
  OAI22_X1 U663 ( .A1(n6292), .A2(n6425), .B1(n1690), .B2(n6424), .ZN(n3354)
         );
  OAI22_X1 U763 ( .A1(n6088), .A2(n6423), .B1(n1724), .B2(n6422), .ZN(n3305)
         );
  OAI22_X1 U761 ( .A1(n6089), .A2(n6423), .B1(n1722), .B2(n6422), .ZN(n3306)
         );
  OAI22_X1 U759 ( .A1(n6090), .A2(n6423), .B1(n1720), .B2(n6422), .ZN(n3307)
         );
  OAI22_X1 U721 ( .A1(n6109), .A2(n6423), .B1(n1682), .B2(n6422), .ZN(n3326)
         );
  OAI22_X1 U719 ( .A1(n6110), .A2(n1990), .B1(n1680), .B2(n6422), .ZN(n3327)
         );
  OAI22_X1 U675 ( .A1(n6286), .A2(n6425), .B1(n1702), .B2(n6424), .ZN(n3348)
         );
  OAI22_X1 U697 ( .A1(n6275), .A2(n6425), .B1(n1724), .B2(n6424), .ZN(n3337)
         );
  OAI22_X1 U665 ( .A1(n6291), .A2(n6425), .B1(n1692), .B2(n6424), .ZN(n3353)
         );
  OAI22_X1 U693 ( .A1(n6277), .A2(n6425), .B1(n1720), .B2(n6424), .ZN(n3339)
         );
  OAI22_X1 U687 ( .A1(n6280), .A2(n6425), .B1(n1714), .B2(n6424), .ZN(n3342)
         );
  OAI22_X1 U685 ( .A1(n6281), .A2(n6425), .B1(n1712), .B2(n6424), .ZN(n3343)
         );
  OAI22_X1 U683 ( .A1(n6282), .A2(n6425), .B1(n1710), .B2(n6424), .ZN(n3344)
         );
  OAI22_X1 U737 ( .A1(n6101), .A2(n6423), .B1(n1698), .B2(n6422), .ZN(n3318)
         );
  OAI22_X1 U735 ( .A1(n6102), .A2(n6423), .B1(n1696), .B2(n6422), .ZN(n3319)
         );
  OAI22_X1 U733 ( .A1(n6103), .A2(n6423), .B1(n1694), .B2(n6422), .ZN(n3320)
         );
  OAI22_X1 U731 ( .A1(n6104), .A2(n6423), .B1(n1692), .B2(n6422), .ZN(n3321)
         );
  OAI22_X1 U727 ( .A1(n6106), .A2(n6423), .B1(n1688), .B2(n6422), .ZN(n3323)
         );
  OAI22_X1 U729 ( .A1(n6105), .A2(n6423), .B1(n1690), .B2(n6422), .ZN(n3322)
         );
  OAI22_X1 U673 ( .A1(n6287), .A2(n6425), .B1(n1700), .B2(n6424), .ZN(n3349)
         );
  OAI22_X1 U725 ( .A1(n6107), .A2(n6423), .B1(n1686), .B2(n6422), .ZN(n3324)
         );
  OAI22_X1 U749 ( .A1(n6095), .A2(n6423), .B1(n1710), .B2(n6422), .ZN(n3312)
         );
  OAI22_X1 U723 ( .A1(n6108), .A2(n6423), .B1(n1684), .B2(n6422), .ZN(n3325)
         );
  OAI22_X1 U695 ( .A1(n6276), .A2(n6425), .B1(n1722), .B2(n6424), .ZN(n3338)
         );
  OAI22_X1 U751 ( .A1(n6094), .A2(n6423), .B1(n1712), .B2(n6422), .ZN(n3311)
         );
  OAI22_X1 U741 ( .A1(n6099), .A2(n6423), .B1(n1702), .B2(n6422), .ZN(n3316)
         );
  OAI22_X1 U617 ( .A1(n4904), .A2(n6427), .B1(n1710), .B2(n6426), .ZN(n3376)
         );
  OAI22_X1 U605 ( .A1(n4929), .A2(n6427), .B1(n1698), .B2(n6426), .ZN(n3382)
         );
  OAI22_X1 U603 ( .A1(n4933), .A2(n6427), .B1(n1696), .B2(n6426), .ZN(n3383)
         );
  OAI22_X1 U627 ( .A1(n4892), .A2(n6427), .B1(n1720), .B2(n6426), .ZN(n3371)
         );
  OAI22_X1 U607 ( .A1(n4928), .A2(n6427), .B1(n1700), .B2(n6426), .ZN(n3381)
         );
  OAI22_X1 U609 ( .A1(n4923), .A2(n6427), .B1(n1702), .B2(n6426), .ZN(n3380)
         );
  OAI22_X1 U591 ( .A1(n4958), .A2(n6427), .B1(n1684), .B2(n6426), .ZN(n3389)
         );
  OAI22_X1 U619 ( .A1(n4903), .A2(n6427), .B1(n1712), .B2(n6426), .ZN(n3375)
         );
  OAI22_X1 U621 ( .A1(n4899), .A2(n6427), .B1(n1714), .B2(n6426), .ZN(n3374)
         );
  OAI22_X1 U587 ( .A1(n4963), .A2(n1921), .B1(n1680), .B2(n6426), .ZN(n3391)
         );
  OAI22_X1 U629 ( .A1(n4883), .A2(n6427), .B1(n1722), .B2(n6426), .ZN(n3370)
         );
  OAI22_X1 U631 ( .A1(n4875), .A2(n6427), .B1(n1724), .B2(n6426), .ZN(n3369)
         );
  OAI22_X1 U597 ( .A1(n4943), .A2(n6427), .B1(n1690), .B2(n6426), .ZN(n3386)
         );
  OAI22_X1 U589 ( .A1(n4959), .A2(n6427), .B1(n1682), .B2(n6426), .ZN(n3390)
         );
  OAI22_X1 U593 ( .A1(n4953), .A2(n6427), .B1(n1686), .B2(n6426), .ZN(n3388)
         );
  OAI22_X1 U595 ( .A1(n4952), .A2(n6427), .B1(n1688), .B2(n6426), .ZN(n3387)
         );
  OAI22_X1 U601 ( .A1(n4934), .A2(n6427), .B1(n1694), .B2(n6426), .ZN(n3384)
         );
  OAI22_X1 U599 ( .A1(n4935), .A2(n6427), .B1(n1692), .B2(n6426), .ZN(n3385)
         );
  OAI22_X1 U1692 ( .A1(n4515), .A2(n6392), .B1(n1668), .B2(n6391), .ZN(n2787)
         );
  OAI22_X1 U1666 ( .A1(n4523), .A2(n4180), .B1(n1666), .B2(n6391), .ZN(n2789)
         );
  OAI22_X1 U1718 ( .A1(n4514), .A2(n6392), .B1(n1670), .B2(n6391), .ZN(n2785)
         );
  OAI22_X1 U2160 ( .A1(n4453), .A2(n6392), .B1(n1704), .B2(n6391), .ZN(n2751)
         );
  OAI22_X1 U1796 ( .A1(n4508), .A2(n6392), .B1(n1676), .B2(n6391), .ZN(n2779)
         );
  OAI22_X1 U1822 ( .A1(n4503), .A2(n4180), .B1(n1678), .B2(n6391), .ZN(n2777)
         );
  OAI22_X1 U1848 ( .A1(n4502), .A2(n4180), .B1(n1680), .B2(n6391), .ZN(n2775)
         );
  OAI22_X1 U1952 ( .A1(n4483), .A2(n6392), .B1(n1688), .B2(n6391), .ZN(n2767)
         );
  OAI22_X1 U1978 ( .A1(n4479), .A2(n6392), .B1(n1690), .B2(n6391), .ZN(n2765)
         );
  OAI22_X1 U2004 ( .A1(n4478), .A2(n6392), .B1(n1692), .B2(n6391), .ZN(n2763)
         );
  OAI22_X1 U2030 ( .A1(n4473), .A2(n6392), .B1(n1694), .B2(n6391), .ZN(n2761)
         );
  OAI22_X1 U2056 ( .A1(n4472), .A2(n6392), .B1(n1696), .B2(n6391), .ZN(n2759)
         );
  OAI22_X1 U2082 ( .A1(n4463), .A2(n6392), .B1(n1698), .B2(n6391), .ZN(n2757)
         );
  OAI22_X1 U2186 ( .A1(n4449), .A2(n6392), .B1(n1706), .B2(n6391), .ZN(n2749)
         );
  OAI22_X1 U2238 ( .A1(n4443), .A2(n6392), .B1(n1710), .B2(n6391), .ZN(n2745)
         );
  OAI22_X1 U2108 ( .A1(n4455), .A2(n6392), .B1(n1700), .B2(n6391), .ZN(n2755)
         );
  OAI22_X1 U2212 ( .A1(n4448), .A2(n6392), .B1(n1708), .B2(n6391), .ZN(n2747)
         );
  OAI22_X1 U2134 ( .A1(n4454), .A2(n6392), .B1(n1702), .B2(n6391), .ZN(n2753)
         );
  OAI22_X1 U1179 ( .A1(n525), .A2(n6408), .B1(n6407), .B2(n1684), .ZN(n3069)
         );
  OAI22_X1 U1181 ( .A1(n527), .A2(n6408), .B1(n6407), .B2(n1688), .ZN(n3067)
         );
  OAI22_X1 U1178 ( .A1(n524), .A2(n6408), .B1(n6407), .B2(n1682), .ZN(n3070)
         );
  OAI22_X1 U1183 ( .A1(n529), .A2(n6408), .B1(n6407), .B2(n1692), .ZN(n3065)
         );
  OAI22_X1 U1184 ( .A1(n530), .A2(n6408), .B1(n6407), .B2(n1694), .ZN(n3064)
         );
  OAI22_X1 U1198 ( .A1(n544), .A2(n6408), .B1(n6407), .B2(n1722), .ZN(n3050)
         );
  OAI22_X1 U1185 ( .A1(n531), .A2(n6408), .B1(n6407), .B2(n1696), .ZN(n3063)
         );
  OAI22_X1 U1186 ( .A1(n532), .A2(n6408), .B1(n6407), .B2(n1698), .ZN(n3062)
         );
  OAI22_X1 U1187 ( .A1(n533), .A2(n6408), .B1(n6407), .B2(n1700), .ZN(n3061)
         );
  OAI22_X1 U1177 ( .A1(n523), .A2(n3994), .B1(n6407), .B2(n1680), .ZN(n3071)
         );
  OAI22_X1 U1188 ( .A1(n534), .A2(n6408), .B1(n6407), .B2(n1702), .ZN(n3060)
         );
  OAI22_X1 U1192 ( .A1(n538), .A2(n6408), .B1(n6407), .B2(n1710), .ZN(n3056)
         );
  OAI22_X1 U1193 ( .A1(n539), .A2(n6408), .B1(n6407), .B2(n1712), .ZN(n3055)
         );
  OAI22_X1 U1180 ( .A1(n526), .A2(n6408), .B1(n6407), .B2(n1686), .ZN(n3068)
         );
  OAI22_X1 U1194 ( .A1(n540), .A2(n6408), .B1(n6407), .B2(n1714), .ZN(n3054)
         );
  OAI22_X1 U1197 ( .A1(n543), .A2(n6408), .B1(n6407), .B2(n1720), .ZN(n3051)
         );
  OAI22_X1 U1182 ( .A1(n528), .A2(n6408), .B1(n6407), .B2(n1690), .ZN(n3066)
         );
  OAI22_X1 U1189 ( .A1(n535), .A2(n6408), .B1(n6407), .B2(n1704), .ZN(n3059)
         );
  OAI22_X1 U783 ( .A1(n718), .A2(n6421), .B1(n6420), .B2(n1692), .ZN(n3289) );
  OAI22_X1 U786 ( .A1(n721), .A2(n6421), .B1(n6420), .B2(n1698), .ZN(n3286) );
  OAI22_X1 U782 ( .A1(n717), .A2(n6421), .B1(n6420), .B2(n1690), .ZN(n3290) );
  OAI22_X1 U781 ( .A1(n716), .A2(n6421), .B1(n6420), .B2(n1688), .ZN(n3291) );
  OAI22_X1 U780 ( .A1(n715), .A2(n6421), .B1(n6420), .B2(n1686), .ZN(n3292) );
  OAI22_X1 U779 ( .A1(n714), .A2(n6421), .B1(n6420), .B2(n1684), .ZN(n3293) );
  OAI22_X1 U778 ( .A1(n713), .A2(n6421), .B1(n6420), .B2(n1682), .ZN(n3294) );
  OAI22_X1 U777 ( .A1(n712), .A2(n2023), .B1(n6420), .B2(n1680), .ZN(n3295) );
  OAI22_X1 U788 ( .A1(n723), .A2(n6421), .B1(n6420), .B2(n1702), .ZN(n3284) );
  OAI22_X1 U798 ( .A1(n733), .A2(n6421), .B1(n6420), .B2(n1722), .ZN(n3274) );
  OAI22_X1 U797 ( .A1(n732), .A2(n6421), .B1(n6420), .B2(n1720), .ZN(n3275) );
  OAI22_X1 U794 ( .A1(n729), .A2(n6421), .B1(n6420), .B2(n1714), .ZN(n3278) );
  OAI22_X1 U793 ( .A1(n728), .A2(n6421), .B1(n6420), .B2(n1712), .ZN(n3279) );
  OAI22_X1 U792 ( .A1(n727), .A2(n6421), .B1(n6420), .B2(n1710), .ZN(n3280) );
  OAI22_X1 U789 ( .A1(n724), .A2(n6421), .B1(n6420), .B2(n1704), .ZN(n3283) );
  OAI22_X1 U785 ( .A1(n720), .A2(n6421), .B1(n6420), .B2(n1696), .ZN(n3287) );
  OAI22_X1 U787 ( .A1(n722), .A2(n6421), .B1(n6420), .B2(n1700), .ZN(n3285) );
  OAI22_X1 U784 ( .A1(n719), .A2(n6421), .B1(n6420), .B2(n1694), .ZN(n3288) );
  OAI22_X1 U1609 ( .A1(n6193), .A2(n6394), .B1(n1700), .B2(n6393), .ZN(n2805)
         );
  OAI22_X1 U1629 ( .A1(n6183), .A2(n6394), .B1(n1720), .B2(n6393), .ZN(n2795)
         );
  OAI22_X1 U1619 ( .A1(n6188), .A2(n6394), .B1(n1710), .B2(n6393), .ZN(n2800)
         );
  OAI22_X1 U1605 ( .A1(n6195), .A2(n6394), .B1(n1696), .B2(n6393), .ZN(n2807)
         );
  OAI22_X1 U1603 ( .A1(n6196), .A2(n6394), .B1(n1694), .B2(n6393), .ZN(n2808)
         );
  OAI22_X1 U1601 ( .A1(n6197), .A2(n6394), .B1(n1692), .B2(n6393), .ZN(n2809)
         );
  OAI22_X1 U1595 ( .A1(n6200), .A2(n6394), .B1(n1686), .B2(n6393), .ZN(n2812)
         );
  OAI22_X1 U1631 ( .A1(n6182), .A2(n6394), .B1(n1722), .B2(n6393), .ZN(n2794)
         );
  OAI22_X1 U1621 ( .A1(n6187), .A2(n6394), .B1(n1712), .B2(n6393), .ZN(n2799)
         );
  OAI22_X1 U1607 ( .A1(n6194), .A2(n6394), .B1(n1698), .B2(n6393), .ZN(n2806)
         );
  OAI22_X1 U1613 ( .A1(n6191), .A2(n6394), .B1(n1704), .B2(n6393), .ZN(n2803)
         );
  OAI22_X1 U1599 ( .A1(n6198), .A2(n6394), .B1(n1690), .B2(n6393), .ZN(n2810)
         );
  OAI22_X1 U1597 ( .A1(n6199), .A2(n6394), .B1(n1688), .B2(n6393), .ZN(n2811)
         );
  OAI22_X1 U1593 ( .A1(n6201), .A2(n6394), .B1(n1684), .B2(n6393), .ZN(n2813)
         );
  OAI22_X1 U1611 ( .A1(n6192), .A2(n6394), .B1(n1702), .B2(n6393), .ZN(n2804)
         );
  OAI22_X1 U1591 ( .A1(n6202), .A2(n6394), .B1(n1682), .B2(n6393), .ZN(n2814)
         );
  OAI22_X1 U1623 ( .A1(n6186), .A2(n6394), .B1(n1714), .B2(n6393), .ZN(n2798)
         );
  OAI22_X1 U1589 ( .A1(n6203), .A2(n4145), .B1(n1680), .B2(n6393), .ZN(n2815)
         );
  OAI22_X1 U1163 ( .A1(n4652), .A2(n6410), .B1(n1724), .B2(n6409), .ZN(n3081)
         );
  OAI22_X1 U1109 ( .A1(n4749), .A2(n6410), .B1(n1670), .B2(n6409), .ZN(n3108)
         );
  OAI22_X1 U1165 ( .A1(n6340), .A2(n6410), .B1(n1726), .B2(n6409), .ZN(n3080)
         );
  OAI22_X1 U1113 ( .A1(n4743), .A2(n6410), .B1(n1674), .B2(n6409), .ZN(n3106)
         );
  OAI22_X1 U1151 ( .A1(n4665), .A2(n6410), .B1(n1712), .B2(n6409), .ZN(n3087)
         );
  OAI22_X1 U1137 ( .A1(n4694), .A2(n6410), .B1(n1698), .B2(n6409), .ZN(n3094)
         );
  OAI22_X1 U1135 ( .A1(n4695), .A2(n6410), .B1(n1696), .B2(n6409), .ZN(n3095)
         );
  OAI22_X1 U1155 ( .A1(n4663), .A2(n6410), .B1(n1716), .B2(n6409), .ZN(n3085)
         );
  OAI22_X1 U1139 ( .A1(n4693), .A2(n6410), .B1(n1700), .B2(n6409), .ZN(n3093)
         );
  OAI22_X1 U1157 ( .A1(n4659), .A2(n6410), .B1(n1718), .B2(n6409), .ZN(n3084)
         );
  OAI22_X1 U1159 ( .A1(n4658), .A2(n6410), .B1(n1720), .B2(n6409), .ZN(n3083)
         );
  OAI22_X1 U1161 ( .A1(n4653), .A2(n6410), .B1(n1722), .B2(n6409), .ZN(n3082)
         );
  OAI22_X1 U1125 ( .A1(n4719), .A2(n6410), .B1(n1686), .B2(n6409), .ZN(n3100)
         );
  OAI22_X1 U1149 ( .A1(n4673), .A2(n6410), .B1(n1710), .B2(n6409), .ZN(n3088)
         );
  OAI22_X1 U1153 ( .A1(n4664), .A2(n6410), .B1(n1714), .B2(n6409), .ZN(n3086)
         );
  OAI22_X1 U1145 ( .A1(n4683), .A2(n6410), .B1(n1706), .B2(n6409), .ZN(n3090)
         );
  OAI22_X1 U1143 ( .A1(n4688), .A2(n6410), .B1(n1704), .B2(n6409), .ZN(n3091)
         );
  OAI22_X1 U1127 ( .A1(n4718), .A2(n6410), .B1(n1688), .B2(n6409), .ZN(n3099)
         );
  OAI22_X1 U1147 ( .A1(n4682), .A2(n6410), .B1(n1708), .B2(n6409), .ZN(n3089)
         );
  OAI22_X1 U1490 ( .A1(n564), .A2(n6398), .B1(n6397), .B2(n1700), .ZN(n2869)
         );
  OAI22_X1 U1489 ( .A1(n563), .A2(n6398), .B1(n6397), .B2(n1698), .ZN(n2870)
         );
  OAI22_X1 U1487 ( .A1(n561), .A2(n6398), .B1(n6397), .B2(n1694), .ZN(n2872)
         );
  OAI22_X1 U1486 ( .A1(n560), .A2(n6398), .B1(n6397), .B2(n1692), .ZN(n2873)
         );
  OAI22_X1 U1500 ( .A1(n574), .A2(n6398), .B1(n6397), .B2(n1720), .ZN(n2859)
         );
  OAI22_X1 U1488 ( .A1(n562), .A2(n6398), .B1(n6397), .B2(n1696), .ZN(n2871)
         );
  OAI22_X1 U1483 ( .A1(n557), .A2(n6398), .B1(n6397), .B2(n1686), .ZN(n2876)
         );
  OAI22_X1 U1482 ( .A1(n556), .A2(n6398), .B1(n6397), .B2(n1684), .ZN(n2877)
         );
  OAI22_X1 U1481 ( .A1(n555), .A2(n6398), .B1(n6397), .B2(n1682), .ZN(n2878)
         );
  OAI22_X1 U1480 ( .A1(n554), .A2(n4106), .B1(n6397), .B2(n1680), .ZN(n2879)
         );
  OAI22_X1 U1491 ( .A1(n565), .A2(n6398), .B1(n6397), .B2(n1702), .ZN(n2868)
         );
  OAI22_X1 U1485 ( .A1(n559), .A2(n6398), .B1(n6397), .B2(n1690), .ZN(n2874)
         );
  OAI22_X1 U1502 ( .A1(n576), .A2(n6398), .B1(n6397), .B2(n1724), .ZN(n2857)
         );
  OAI22_X1 U1501 ( .A1(n575), .A2(n6398), .B1(n6397), .B2(n1722), .ZN(n2858)
         );
  OAI22_X1 U1495 ( .A1(n569), .A2(n6398), .B1(n6397), .B2(n1710), .ZN(n2864)
         );
  OAI22_X1 U1499 ( .A1(n573), .A2(n6398), .B1(n6397), .B2(n1718), .ZN(n2860)
         );
  OAI22_X1 U1496 ( .A1(n570), .A2(n6398), .B1(n6397), .B2(n1712), .ZN(n2863)
         );
  OAI22_X1 U1484 ( .A1(n558), .A2(n6398), .B1(n6397), .B2(n1688), .ZN(n2875)
         );
  OAI22_X1 U1373 ( .A1(n2245), .A2(n6401), .B1(n3886), .B2(n1670), .ZN(n2948)
         );
  OAI22_X1 U1389 ( .A1(n2229), .A2(n6401), .B1(n3886), .B2(n1702), .ZN(n2932)
         );
  OAI22_X1 U1383 ( .A1(n2235), .A2(n6401), .B1(n3886), .B2(n1690), .ZN(n2938)
         );
  OAI22_X1 U1380 ( .A1(n2238), .A2(n6401), .B1(n3886), .B2(n1684), .ZN(n2941)
         );
  OAI22_X1 U1377 ( .A1(n2241), .A2(n4068), .B1(n3886), .B2(n1678), .ZN(n2944)
         );
  OAI22_X1 U1378 ( .A1(n2240), .A2(n4068), .B1(n3886), .B2(n1680), .ZN(n2943)
         );
  OAI22_X1 U1384 ( .A1(n2234), .A2(n6401), .B1(n3886), .B2(n1692), .ZN(n2937)
         );
  OAI22_X1 U1385 ( .A1(n2233), .A2(n6401), .B1(n3886), .B2(n1694), .ZN(n2936)
         );
  OAI22_X1 U1379 ( .A1(n2239), .A2(n6401), .B1(n3886), .B2(n1682), .ZN(n2942)
         );
  OAI22_X1 U1387 ( .A1(n2231), .A2(n6401), .B1(n3886), .B2(n1698), .ZN(n2934)
         );
  OAI22_X1 U1375 ( .A1(n2243), .A2(n4068), .B1(n3886), .B2(n1674), .ZN(n2946)
         );
  OAI22_X1 U1386 ( .A1(n2232), .A2(n6401), .B1(n3886), .B2(n1696), .ZN(n2935)
         );
  OAI22_X1 U1381 ( .A1(n2237), .A2(n6401), .B1(n3886), .B2(n1686), .ZN(n2940)
         );
  OAI22_X1 U1382 ( .A1(n2236), .A2(n6401), .B1(n3886), .B2(n1688), .ZN(n2939)
         );
  OAI22_X1 U1388 ( .A1(n2230), .A2(n6401), .B1(n3886), .B2(n1700), .ZN(n2933)
         );
  OAI22_X1 U383 ( .A1(n2653), .A2(n6434), .B1(n3881), .B2(n1686), .ZN(n3516)
         );
  OAI22_X1 U379 ( .A1(n2657), .A2(n1847), .B1(n3881), .B2(n1678), .ZN(n3520)
         );
  OAI22_X1 U382 ( .A1(n2654), .A2(n6434), .B1(n3881), .B2(n1684), .ZN(n3517)
         );
  OAI22_X1 U380 ( .A1(n2656), .A2(n1847), .B1(n3881), .B2(n1680), .ZN(n3519)
         );
  OAI22_X1 U384 ( .A1(n2652), .A2(n6434), .B1(n3881), .B2(n1688), .ZN(n3515)
         );
  OAI22_X1 U385 ( .A1(n2651), .A2(n6434), .B1(n3881), .B2(n1690), .ZN(n3514)
         );
  OAI22_X1 U377 ( .A1(n2659), .A2(n1847), .B1(n3881), .B2(n1674), .ZN(n3522)
         );
  OAI22_X1 U388 ( .A1(n2648), .A2(n6434), .B1(n3881), .B2(n1696), .ZN(n3511)
         );
  OAI22_X1 U389 ( .A1(n2647), .A2(n6434), .B1(n3881), .B2(n1698), .ZN(n3510)
         );
  OAI22_X1 U386 ( .A1(n2650), .A2(n6434), .B1(n3881), .B2(n1692), .ZN(n3513)
         );
  OAI22_X1 U381 ( .A1(n2655), .A2(n6434), .B1(n3881), .B2(n1682), .ZN(n3518)
         );
  OAI22_X1 U375 ( .A1(n2661), .A2(n6434), .B1(n3881), .B2(n1670), .ZN(n3524)
         );
  OAI22_X1 U387 ( .A1(n2649), .A2(n6434), .B1(n3881), .B2(n1694), .ZN(n3512)
         );
  OAI22_X1 U390 ( .A1(n2646), .A2(n6434), .B1(n3881), .B2(n1700), .ZN(n3509)
         );
  OAI22_X1 U391 ( .A1(n2645), .A2(n6434), .B1(n3881), .B2(n1702), .ZN(n3508)
         );
  OAI22_X1 U1400 ( .A1(n6243), .A2(n6401), .B1(n1724), .B2(n3886), .ZN(n2921)
         );
  OAI22_X1 U1402 ( .A1(n4167), .A2(n6401), .B1(n1726), .B2(n3886), .ZN(n2920)
         );
  OAI22_X1 U403 ( .A1(n4169), .A2(n6434), .B1(n1726), .B2(n3881), .ZN(n3496)
         );
  OAI22_X1 U1348 ( .A1(n6158), .A2(n6403), .B1(n1708), .B2(n4036), .ZN(n2961)
         );
  OAI22_X1 U1304 ( .A1(n6180), .A2(n4035), .B1(n1663), .B2(n4036), .ZN(n2983)
         );
  OAI22_X1 U1306 ( .A1(n6179), .A2(n4035), .B1(n1666), .B2(n4036), .ZN(n2982)
         );
  OAI22_X1 U1312 ( .A1(n6176), .A2(n6403), .B1(n1672), .B2(n4036), .ZN(n2979)
         );
  OAI22_X1 U1356 ( .A1(n6154), .A2(n6403), .B1(n1716), .B2(n4036), .ZN(n2957)
         );
  OAI22_X1 U1406 ( .A1(n6242), .A2(n4073), .B1(n1663), .B2(n4074), .ZN(n2919)
         );
  OAI22_X1 U1346 ( .A1(n6159), .A2(n6403), .B1(n1706), .B2(n4036), .ZN(n2962)
         );
  OAI22_X1 U1344 ( .A1(n6160), .A2(n6403), .B1(n1704), .B2(n4036), .ZN(n2963)
         );
  OAI22_X1 U1318 ( .A1(n6173), .A2(n4035), .B1(n1678), .B2(n4036), .ZN(n2976)
         );
  OAI22_X1 U1316 ( .A1(n6174), .A2(n4035), .B1(n1676), .B2(n4036), .ZN(n2977)
         );
  OAI22_X1 U1314 ( .A1(n6175), .A2(n6403), .B1(n1674), .B2(n4036), .ZN(n2978)
         );
  OAI22_X1 U1366 ( .A1(n6339), .A2(n6403), .B1(n1726), .B2(n4036), .ZN(n2952)
         );
  OAI22_X1 U1358 ( .A1(n6153), .A2(n6403), .B1(n1718), .B2(n4036), .ZN(n2956)
         );
  OAI22_X1 U1418 ( .A1(n6236), .A2(n4073), .B1(n1676), .B2(n4074), .ZN(n2913)
         );
  OAI22_X1 U1420 ( .A1(n6235), .A2(n4073), .B1(n1678), .B2(n4074), .ZN(n2912)
         );
  OAI22_X1 U1446 ( .A1(n6222), .A2(n6400), .B1(n1704), .B2(n4074), .ZN(n2899)
         );
  OAI22_X1 U1448 ( .A1(n6221), .A2(n6400), .B1(n1706), .B2(n4074), .ZN(n2898)
         );
  OAI22_X1 U1450 ( .A1(n6220), .A2(n6400), .B1(n1708), .B2(n4074), .ZN(n2897)
         );
  OAI22_X1 U1458 ( .A1(n6216), .A2(n6400), .B1(n1716), .B2(n4074), .ZN(n2893)
         );
  OAI22_X1 U1460 ( .A1(n6215), .A2(n6400), .B1(n1718), .B2(n4074), .ZN(n2892)
         );
  OAI22_X1 U1468 ( .A1(n6348), .A2(n6400), .B1(n1726), .B2(n4074), .ZN(n2888)
         );
  OAI22_X1 U1310 ( .A1(n6177), .A2(n6403), .B1(n1670), .B2(n4036), .ZN(n2980)
         );
  OAI22_X1 U1308 ( .A1(n6178), .A2(n6403), .B1(n1668), .B2(n4036), .ZN(n2981)
         );
  OAI22_X1 U1408 ( .A1(n6241), .A2(n4073), .B1(n1666), .B2(n4074), .ZN(n2918)
         );
  OAI22_X1 U1410 ( .A1(n6240), .A2(n6400), .B1(n1668), .B2(n4074), .ZN(n2917)
         );
  OAI22_X1 U1412 ( .A1(n6239), .A2(n6400), .B1(n1670), .B2(n4074), .ZN(n2916)
         );
  OAI22_X1 U1414 ( .A1(n6238), .A2(n6400), .B1(n1672), .B2(n4074), .ZN(n2915)
         );
  OAI22_X1 U1416 ( .A1(n6237), .A2(n6400), .B1(n1674), .B2(n4074), .ZN(n2914)
         );
  OAI22_X1 U1250 ( .A1(n6143), .A2(n4000), .B1(n1676), .B2(n4001), .ZN(n3009)
         );
  OAI22_X1 U1252 ( .A1(n6142), .A2(n4000), .B1(n1678), .B2(n4001), .ZN(n3008)
         );
  OAI22_X1 U1278 ( .A1(n6129), .A2(n6405), .B1(n1704), .B2(n4001), .ZN(n2995)
         );
  OAI22_X1 U1238 ( .A1(n6149), .A2(n4000), .B1(n1663), .B2(n4001), .ZN(n3015)
         );
  OAI22_X1 U1240 ( .A1(n6148), .A2(n4000), .B1(n1666), .B2(n4001), .ZN(n3014)
         );
  OAI22_X1 U1242 ( .A1(n6147), .A2(n6405), .B1(n1668), .B2(n4001), .ZN(n3013)
         );
  OAI22_X1 U1244 ( .A1(n6146), .A2(n6405), .B1(n1670), .B2(n4001), .ZN(n3012)
         );
  OAI22_X1 U1246 ( .A1(n6145), .A2(n6405), .B1(n1672), .B2(n4001), .ZN(n3011)
         );
  OAI22_X1 U1248 ( .A1(n6144), .A2(n6405), .B1(n1674), .B2(n4001), .ZN(n3010)
         );
  OAI22_X1 U1282 ( .A1(n6127), .A2(n6405), .B1(n1708), .B2(n4001), .ZN(n2993)
         );
  OAI22_X1 U1290 ( .A1(n6123), .A2(n6405), .B1(n1716), .B2(n4001), .ZN(n2989)
         );
  OAI22_X1 U1280 ( .A1(n6128), .A2(n6405), .B1(n1706), .B2(n4001), .ZN(n2994)
         );
  OAI22_X1 U1292 ( .A1(n6122), .A2(n6405), .B1(n1718), .B2(n4001), .ZN(n2988)
         );
  OAI22_X1 U1298 ( .A1(n6119), .A2(n6405), .B1(n1724), .B2(n4001), .ZN(n2985)
         );
  OAI22_X1 U1391 ( .A1(n2227), .A2(n6401), .B1(n3886), .B2(n1706), .ZN(n2930)
         );
  OAI22_X1 U1374 ( .A1(n2244), .A2(n6401), .B1(n3886), .B2(n1672), .ZN(n2947)
         );
  OAI22_X1 U1390 ( .A1(n2228), .A2(n6401), .B1(n3886), .B2(n1704), .ZN(n2931)
         );
  OAI22_X1 U1394 ( .A1(n2224), .A2(n6401), .B1(n3886), .B2(n1712), .ZN(n2927)
         );
  OAI22_X1 U1372 ( .A1(n2246), .A2(n6401), .B1(n3886), .B2(n1668), .ZN(n2949)
         );
  OAI22_X1 U1396 ( .A1(n2222), .A2(n6401), .B1(n3886), .B2(n1716), .ZN(n2925)
         );
  OAI22_X1 U1397 ( .A1(n2221), .A2(n6401), .B1(n3886), .B2(n1718), .ZN(n2924)
         );
  OAI22_X1 U1398 ( .A1(n2220), .A2(n6401), .B1(n3886), .B2(n1720), .ZN(n2923)
         );
  OAI22_X1 U1399 ( .A1(n2219), .A2(n6401), .B1(n3886), .B2(n1722), .ZN(n2922)
         );
  OAI22_X1 U1392 ( .A1(n2226), .A2(n6401), .B1(n3886), .B2(n1708), .ZN(n2929)
         );
  OAI22_X1 U1393 ( .A1(n2225), .A2(n6401), .B1(n3886), .B2(n1710), .ZN(n2928)
         );
  OAI22_X1 U1395 ( .A1(n2223), .A2(n6401), .B1(n3886), .B2(n1714), .ZN(n2926)
         );
  OAI22_X1 U374 ( .A1(n2662), .A2(n6434), .B1(n3881), .B2(n1668), .ZN(n3525)
         );
  OAI22_X1 U376 ( .A1(n2660), .A2(n6434), .B1(n3881), .B2(n1672), .ZN(n3523)
         );
  OAI22_X1 U401 ( .A1(n2635), .A2(n6434), .B1(n3881), .B2(n1722), .ZN(n3498)
         );
  OAI22_X1 U402 ( .A1(n2634), .A2(n6434), .B1(n3881), .B2(n1724), .ZN(n3497)
         );
  OAI22_X1 U395 ( .A1(n2641), .A2(n6434), .B1(n3881), .B2(n1710), .ZN(n3504)
         );
  OAI22_X1 U396 ( .A1(n2640), .A2(n6434), .B1(n3881), .B2(n1712), .ZN(n3503)
         );
  OAI22_X1 U397 ( .A1(n2639), .A2(n6434), .B1(n3881), .B2(n1714), .ZN(n3502)
         );
  OAI22_X1 U398 ( .A1(n2638), .A2(n6434), .B1(n3881), .B2(n1716), .ZN(n3501)
         );
  OAI22_X1 U399 ( .A1(n2637), .A2(n6434), .B1(n3881), .B2(n1718), .ZN(n3500)
         );
  OAI22_X1 U392 ( .A1(n2644), .A2(n6434), .B1(n3881), .B2(n1704), .ZN(n3507)
         );
  OAI22_X1 U393 ( .A1(n2643), .A2(n6434), .B1(n3881), .B2(n1706), .ZN(n3506)
         );
  OAI22_X1 U394 ( .A1(n2642), .A2(n6434), .B1(n3881), .B2(n1708), .ZN(n3505)
         );
  OAI22_X1 U400 ( .A1(n2636), .A2(n6434), .B1(n3881), .B2(n1720), .ZN(n3499)
         );
  OAI22_X1 U429 ( .A1(n5933), .A2(n6433), .B1(n1686), .B2(n1853), .ZN(n3484)
         );
  OAI22_X1 U490 ( .A1(n5078), .A2(n1885), .B1(n1682), .B2(n1886), .ZN(n3454)
         );
  OAI22_X1 U528 ( .A1(n5003), .A2(n6431), .B1(n1720), .B2(n1886), .ZN(n3435)
         );
  OAI22_X1 U427 ( .A1(n5965), .A2(n6433), .B1(n1684), .B2(n1853), .ZN(n3485)
         );
  OAI22_X1 U488 ( .A1(n5079), .A2(n6431), .B1(n1680), .B2(n1886), .ZN(n3455)
         );
  OAI22_X1 U520 ( .A1(n5019), .A2(n6431), .B1(n1712), .B2(n1886), .ZN(n3439)
         );
  OAI22_X1 U522 ( .A1(n5018), .A2(n6431), .B1(n1714), .B2(n1886), .ZN(n3438)
         );
  OAI22_X1 U524 ( .A1(n5013), .A2(n6431), .B1(n1716), .B2(n1886), .ZN(n3437)
         );
  OAI22_X1 U526 ( .A1(n5012), .A2(n6431), .B1(n1718), .B2(n1886), .ZN(n3436)
         );
  OAI22_X1 U494 ( .A1(n5072), .A2(n6431), .B1(n1686), .B2(n1886), .ZN(n3452)
         );
  OAI22_X1 U492 ( .A1(n5073), .A2(n6431), .B1(n1684), .B2(n1886), .ZN(n3453)
         );
  OAI22_X1 U457 ( .A1(n5134), .A2(n6433), .B1(n1714), .B2(n1853), .ZN(n3470)
         );
  OAI22_X1 U425 ( .A1(n5970), .A2(n1852), .B1(n1682), .B2(n1853), .ZN(n3486)
         );
  OAI22_X1 U407 ( .A1(n5993), .A2(n6433), .B1(n1663), .B2(n1853), .ZN(n3495)
         );
  OAI22_X1 U530 ( .A1(n4995), .A2(n6431), .B1(n1722), .B2(n1886), .ZN(n3434)
         );
  OAI22_X1 U482 ( .A1(n5085), .A2(n6431), .B1(n1674), .B2(n1886), .ZN(n3458)
         );
  OAI22_X1 U480 ( .A1(n5093), .A2(n6431), .B1(n1672), .B2(n1886), .ZN(n3459)
         );
  OAI22_X1 U532 ( .A1(n4994), .A2(n6431), .B1(n1724), .B2(n1886), .ZN(n3433)
         );
  OAI22_X1 U417 ( .A1(n5988), .A2(n6433), .B1(n1674), .B2(n1853), .ZN(n3490)
         );
  OAI22_X1 U467 ( .A1(n5113), .A2(n6433), .B1(n1724), .B2(n1853), .ZN(n3465)
         );
  OAI22_X1 U472 ( .A1(n5109), .A2(n6431), .B1(n1663), .B2(n1886), .ZN(n3463)
         );
  OAI22_X1 U463 ( .A1(n5115), .A2(n6433), .B1(n1720), .B2(n1853), .ZN(n3467)
         );
  OAI22_X1 U461 ( .A1(n5123), .A2(n6433), .B1(n1718), .B2(n1853), .ZN(n3468)
         );
  OAI22_X1 U465 ( .A1(n5114), .A2(n6433), .B1(n1722), .B2(n1853), .ZN(n3466)
         );
  OAI22_X1 U423 ( .A1(n5985), .A2(n6433), .B1(n1680), .B2(n1853), .ZN(n3487)
         );
  OAI22_X1 U455 ( .A1(n5139), .A2(n6433), .B1(n1712), .B2(n1853), .ZN(n3471)
         );
  OAI22_X1 U459 ( .A1(n5133), .A2(n6433), .B1(n1716), .B2(n1853), .ZN(n3469)
         );
  OAI22_X1 U415 ( .A1(n5989), .A2(n6433), .B1(n1672), .B2(n1853), .ZN(n3491)
         );
  OAI22_X1 U563 ( .A1(n508), .A2(n6429), .B1(n1918), .B2(n1716), .ZN(n3405) );
  OAI22_X1 U540 ( .A1(n485), .A2(n6429), .B1(n1918), .B2(n1670), .ZN(n3428) );
  OAI22_X1 U539 ( .A1(n484), .A2(n6429), .B1(n1918), .B2(n1668), .ZN(n3429) );
  OAI22_X1 U558 ( .A1(n503), .A2(n6429), .B1(n1918), .B2(n1706), .ZN(n3410) );
  OAI22_X1 U537 ( .A1(n482), .A2(n1917), .B1(n1918), .B2(n1663), .ZN(n3431) );
  OAI22_X1 U538 ( .A1(n483), .A2(n1917), .B1(n1918), .B2(n1666), .ZN(n3430) );
  OAI22_X1 U544 ( .A1(n489), .A2(n1917), .B1(n1918), .B2(n1678), .ZN(n3424) );
  OAI22_X1 U568 ( .A1(n639), .A2(n6429), .B1(n1918), .B2(n1726), .ZN(n3400) );
  OAI22_X1 U541 ( .A1(n486), .A2(n6429), .B1(n1918), .B2(n1672), .ZN(n3427) );
  OAI22_X1 U559 ( .A1(n504), .A2(n6429), .B1(n1918), .B2(n1708), .ZN(n3409) );
  OAI22_X1 U564 ( .A1(n509), .A2(n6429), .B1(n1918), .B2(n1718), .ZN(n3404) );
  OAI22_X1 U543 ( .A1(n488), .A2(n1917), .B1(n1918), .B2(n1676), .ZN(n3425) );
  OAI22_X1 U542 ( .A1(n487), .A2(n6429), .B1(n1918), .B2(n1674), .ZN(n3426) );
  OAI22_X1 U567 ( .A1(n512), .A2(n6429), .B1(n1918), .B2(n1724), .ZN(n3401) );
  OAI22_X1 U345 ( .A1(n616), .A2(n1843), .B1(n3883), .B2(n1680), .ZN(n3551) );
  OAI22_X1 U348 ( .A1(n619), .A2(n6435), .B1(n3883), .B2(n1686), .ZN(n3548) );
  OAI22_X1 U347 ( .A1(n618), .A2(n6435), .B1(n3883), .B2(n1684), .ZN(n3549) );
  OAI22_X1 U351 ( .A1(n622), .A2(n6435), .B1(n3883), .B2(n1692), .ZN(n3545) );
  OAI22_X1 U353 ( .A1(n624), .A2(n6435), .B1(n3883), .B2(n1696), .ZN(n3543) );
  OAI22_X1 U346 ( .A1(n617), .A2(n6435), .B1(n3883), .B2(n1682), .ZN(n3550) );
  OAI22_X1 U355 ( .A1(n626), .A2(n6435), .B1(n3883), .B2(n1700), .ZN(n3541) );
  OAI22_X1 U356 ( .A1(n627), .A2(n6435), .B1(n3883), .B2(n1702), .ZN(n3540) );
  OAI22_X1 U349 ( .A1(n620), .A2(n6435), .B1(n3883), .B2(n1688), .ZN(n3547) );
  OAI22_X1 U350 ( .A1(n621), .A2(n6435), .B1(n3883), .B2(n1690), .ZN(n3546) );
  OAI22_X1 U340 ( .A1(n611), .A2(n6435), .B1(n3883), .B2(n1670), .ZN(n3556) );
  OAI22_X1 U352 ( .A1(n623), .A2(n6435), .B1(n3883), .B2(n1694), .ZN(n3544) );
  OAI22_X1 U342 ( .A1(n613), .A2(n1843), .B1(n3883), .B2(n1674), .ZN(n3554) );
  OAI22_X1 U354 ( .A1(n625), .A2(n6435), .B1(n3883), .B2(n1698), .ZN(n3542) );
  OAI22_X1 U344 ( .A1(n615), .A2(n1843), .B1(n3883), .B2(n1678), .ZN(n3552) );
  OAI22_X1 U250 ( .A1(n3771), .A2(n6438), .B1(n3882), .B2(n1690), .ZN(n3610)
         );
  OAI22_X1 U245 ( .A1(n3776), .A2(n1807), .B1(n3882), .B2(n1680), .ZN(n3615)
         );
  OAI22_X1 U246 ( .A1(n3775), .A2(n6438), .B1(n3882), .B2(n1682), .ZN(n3614)
         );
  OAI22_X1 U247 ( .A1(n3774), .A2(n6438), .B1(n3882), .B2(n1684), .ZN(n3613)
         );
  OAI22_X1 U248 ( .A1(n3773), .A2(n6438), .B1(n3882), .B2(n1686), .ZN(n3612)
         );
  OAI22_X1 U249 ( .A1(n3772), .A2(n6438), .B1(n3882), .B2(n1688), .ZN(n3611)
         );
  OAI22_X1 U253 ( .A1(n3768), .A2(n6438), .B1(n3882), .B2(n1696), .ZN(n3607)
         );
  OAI22_X1 U251 ( .A1(n3770), .A2(n6438), .B1(n3882), .B2(n1692), .ZN(n3609)
         );
  OAI22_X1 U252 ( .A1(n3769), .A2(n6438), .B1(n3882), .B2(n1694), .ZN(n3608)
         );
  OAI22_X1 U256 ( .A1(n3765), .A2(n6438), .B1(n3882), .B2(n1702), .ZN(n3604)
         );
  OAI22_X1 U254 ( .A1(n3767), .A2(n6438), .B1(n3882), .B2(n1698), .ZN(n3606)
         );
  OAI22_X1 U255 ( .A1(n3766), .A2(n6438), .B1(n3882), .B2(n1700), .ZN(n3605)
         );
  OAI22_X1 U240 ( .A1(n3781), .A2(n6438), .B1(n3882), .B2(n1670), .ZN(n3620)
         );
  OAI22_X1 U244 ( .A1(n3777), .A2(n1807), .B1(n3882), .B2(n1678), .ZN(n3616)
         );
  OAI22_X1 U242 ( .A1(n3779), .A2(n1807), .B1(n3882), .B2(n1674), .ZN(n3618)
         );
  OAI22_X1 U368 ( .A1(n6343), .A2(n6435), .B1(n1726), .B2(n3883), .ZN(n3528)
         );
  OAI22_X1 U55 ( .A1(n6029), .A2(n6445), .B1(n1716), .B2(n1664), .ZN(n3725) );
  OAI22_X1 U3 ( .A1(n6055), .A2(n1662), .B1(n1663), .B2(n1664), .ZN(n3751) );
  OAI22_X1 U17 ( .A1(n6048), .A2(n1662), .B1(n1678), .B2(n1664), .ZN(n3744) );
  OAI22_X1 U47 ( .A1(n6033), .A2(n6445), .B1(n1708), .B2(n1664), .ZN(n3729) );
  OAI22_X1 U43 ( .A1(n6035), .A2(n6445), .B1(n1704), .B2(n1664), .ZN(n3731) );
  OAI22_X1 U7 ( .A1(n6053), .A2(n6445), .B1(n1668), .B2(n1664), .ZN(n3749) );
  OAI22_X1 U9 ( .A1(n6052), .A2(n6445), .B1(n1670), .B2(n1664), .ZN(n3748) );
  OAI22_X1 U45 ( .A1(n6034), .A2(n6445), .B1(n1706), .B2(n1664), .ZN(n3730) );
  OAI22_X1 U65 ( .A1(n6346), .A2(n6445), .B1(n1726), .B2(n1664), .ZN(n3720) );
  OAI22_X1 U5 ( .A1(n6054), .A2(n1662), .B1(n1666), .B2(n1664), .ZN(n3750) );
  OAI22_X1 U57 ( .A1(n6028), .A2(n6445), .B1(n1718), .B2(n1664), .ZN(n3724) );
  OAI22_X1 U11 ( .A1(n6051), .A2(n6445), .B1(n1672), .B2(n1664), .ZN(n3747) );
  OAI22_X1 U15 ( .A1(n6049), .A2(n1662), .B1(n1676), .B2(n1664), .ZN(n3745) );
  OAI22_X1 U13 ( .A1(n6050), .A2(n6445), .B1(n1674), .B2(n1664), .ZN(n3746) );
  OAI22_X1 U1220 ( .A1(n689), .A2(n6406), .B1(n3887), .B2(n1698), .ZN(n3030)
         );
  OAI22_X1 U1221 ( .A1(n690), .A2(n6406), .B1(n3887), .B2(n1700), .ZN(n3029)
         );
  OAI22_X1 U1222 ( .A1(n691), .A2(n6406), .B1(n3887), .B2(n1702), .ZN(n3028)
         );
  OAI22_X1 U1217 ( .A1(n686), .A2(n6406), .B1(n3887), .B2(n1692), .ZN(n3033)
         );
  OAI22_X1 U1206 ( .A1(n675), .A2(n6406), .B1(n3887), .B2(n1670), .ZN(n3044)
         );
  OAI22_X1 U1218 ( .A1(n687), .A2(n6406), .B1(n3887), .B2(n1694), .ZN(n3032)
         );
  OAI22_X1 U1214 ( .A1(n683), .A2(n6406), .B1(n3887), .B2(n1686), .ZN(n3036)
         );
  OAI22_X1 U1213 ( .A1(n682), .A2(n6406), .B1(n3887), .B2(n1684), .ZN(n3037)
         );
  OAI22_X1 U1212 ( .A1(n681), .A2(n6406), .B1(n3887), .B2(n1682), .ZN(n3038)
         );
  OAI22_X1 U1211 ( .A1(n680), .A2(n3996), .B1(n3887), .B2(n1680), .ZN(n3039)
         );
  OAI22_X1 U1210 ( .A1(n679), .A2(n3996), .B1(n3887), .B2(n1678), .ZN(n3040)
         );
  OAI22_X1 U1208 ( .A1(n677), .A2(n3996), .B1(n3887), .B2(n1674), .ZN(n3042)
         );
  OAI22_X1 U1216 ( .A1(n685), .A2(n6406), .B1(n3887), .B2(n1690), .ZN(n3034)
         );
  OAI22_X1 U1215 ( .A1(n684), .A2(n6406), .B1(n3887), .B2(n1688), .ZN(n3035)
         );
  OAI22_X1 U1219 ( .A1(n688), .A2(n6406), .B1(n3887), .B2(n1696), .ZN(n3031)
         );
  OAI22_X1 U268 ( .A1(n6344), .A2(n6438), .B1(n1726), .B2(n3882), .ZN(n3592)
         );
  OAI22_X1 U920 ( .A1(n4175), .A2(n6417), .B1(n1714), .B2(n6416), .ZN(n3214)
         );
  OAI22_X1 U926 ( .A1(n4172), .A2(n6417), .B1(n1720), .B2(n6416), .ZN(n3211)
         );
  OAI22_X1 U928 ( .A1(n4171), .A2(n6417), .B1(n1722), .B2(n6416), .ZN(n3210)
         );
  OAI22_X1 U930 ( .A1(n4170), .A2(n6417), .B1(n1724), .B2(n6416), .ZN(n3209)
         );
  OAI22_X1 U898 ( .A1(n4242), .A2(n6417), .B1(n1692), .B2(n6416), .ZN(n3225)
         );
  OAI22_X1 U900 ( .A1(n4230), .A2(n6417), .B1(n1694), .B2(n6416), .ZN(n3224)
         );
  OAI22_X1 U892 ( .A1(n4253), .A2(n6417), .B1(n1686), .B2(n6416), .ZN(n3228)
         );
  OAI22_X1 U894 ( .A1(n4245), .A2(n6417), .B1(n1688), .B2(n6416), .ZN(n3227)
         );
  OAI22_X1 U906 ( .A1(n4213), .A2(n6417), .B1(n1700), .B2(n6416), .ZN(n3221)
         );
  OAI22_X1 U904 ( .A1(n4222), .A2(n2062), .B1(n1698), .B2(n6416), .ZN(n3222)
         );
  OAI22_X1 U918 ( .A1(n4176), .A2(n6417), .B1(n1712), .B2(n6416), .ZN(n3215)
         );
  OAI22_X1 U886 ( .A1(n4268), .A2(n2062), .B1(n1680), .B2(n6416), .ZN(n3231)
         );
  OAI22_X1 U888 ( .A1(n4263), .A2(n6417), .B1(n1682), .B2(n6416), .ZN(n3230)
         );
  OAI22_X1 U890 ( .A1(n4262), .A2(n6417), .B1(n1684), .B2(n6416), .ZN(n3229)
         );
  OAI22_X1 U908 ( .A1(n4206), .A2(n6417), .B1(n1702), .B2(n6416), .ZN(n3220)
         );
  OAI22_X1 U902 ( .A1(n4227), .A2(n6417), .B1(n1696), .B2(n6416), .ZN(n3223)
         );
  OAI22_X1 U884 ( .A1(n4269), .A2(n2062), .B1(n1678), .B2(n6416), .ZN(n3232)
         );
  OAI22_X1 U896 ( .A1(n4244), .A2(n2062), .B1(n1690), .B2(n6416), .ZN(n3226)
         );
  OAI22_X1 U838 ( .A1(n6257), .A2(n6419), .B1(n1698), .B2(n6418), .ZN(n3254)
         );
  OAI22_X1 U824 ( .A1(n6264), .A2(n6419), .B1(n1684), .B2(n6418), .ZN(n3261)
         );
  OAI22_X1 U822 ( .A1(n6265), .A2(n6419), .B1(n1682), .B2(n6418), .ZN(n3262)
         );
  OAI22_X1 U836 ( .A1(n6258), .A2(n6419), .B1(n1696), .B2(n6418), .ZN(n3255)
         );
  OAI22_X1 U860 ( .A1(n6246), .A2(n6419), .B1(n1720), .B2(n6418), .ZN(n3243)
         );
  OAI22_X1 U826 ( .A1(n6263), .A2(n6419), .B1(n1686), .B2(n6418), .ZN(n3260)
         );
  OAI22_X1 U818 ( .A1(n6267), .A2(n2027), .B1(n1678), .B2(n6418), .ZN(n3264)
         );
  OAI22_X1 U864 ( .A1(n6244), .A2(n6419), .B1(n1724), .B2(n6418), .ZN(n3241)
         );
  OAI22_X1 U840 ( .A1(n6256), .A2(n2027), .B1(n1700), .B2(n6418), .ZN(n3253)
         );
  OAI22_X1 U820 ( .A1(n6266), .A2(n6419), .B1(n1680), .B2(n6418), .ZN(n3263)
         );
  OAI22_X1 U862 ( .A1(n6245), .A2(n6419), .B1(n1722), .B2(n6418), .ZN(n3242)
         );
  OAI22_X1 U834 ( .A1(n6259), .A2(n6419), .B1(n1694), .B2(n6418), .ZN(n3256)
         );
  OAI22_X1 U832 ( .A1(n6260), .A2(n6419), .B1(n1692), .B2(n6418), .ZN(n3257)
         );
  OAI22_X1 U854 ( .A1(n6249), .A2(n6419), .B1(n1714), .B2(n6418), .ZN(n3246)
         );
  OAI22_X1 U828 ( .A1(n6262), .A2(n6419), .B1(n1688), .B2(n6418), .ZN(n3259)
         );
  OAI22_X1 U830 ( .A1(n6261), .A2(n2027), .B1(n1690), .B2(n6418), .ZN(n3258)
         );
  OAI22_X1 U842 ( .A1(n6255), .A2(n2027), .B1(n1702), .B2(n6418), .ZN(n3252)
         );
  OAI22_X1 U852 ( .A1(n6250), .A2(n6419), .B1(n1712), .B2(n6418), .ZN(n3247)
         );
  OAI22_X1 U223 ( .A1(n4313), .A2(n6440), .B1(n1716), .B2(n1773), .ZN(n3629)
         );
  OAI22_X1 U173 ( .A1(n4412), .A2(n1772), .B1(n1666), .B2(n1773), .ZN(n3654)
         );
  OAI22_X1 U179 ( .A1(n4394), .A2(n6440), .B1(n1672), .B2(n1773), .ZN(n3651)
         );
  OAI22_X1 U231 ( .A1(n4299), .A2(n6440), .B1(n1724), .B2(n1773), .ZN(n3625)
         );
  OAI22_X1 U183 ( .A1(n4389), .A2(n6440), .B1(n1676), .B2(n1773), .ZN(n3649)
         );
  OAI22_X1 U181 ( .A1(n4393), .A2(n1772), .B1(n1674), .B2(n1773), .ZN(n3650)
         );
  OAI22_X1 U171 ( .A1(n4413), .A2(n1772), .B1(n1663), .B2(n1773), .ZN(n3655)
         );
  OAI22_X1 U177 ( .A1(n4395), .A2(n6440), .B1(n1670), .B2(n1773), .ZN(n3652)
         );
  OAI22_X1 U211 ( .A1(n4334), .A2(n6440), .B1(n1704), .B2(n1773), .ZN(n3635)
         );
  OAI22_X1 U175 ( .A1(n4403), .A2(n6440), .B1(n1668), .B2(n1773), .ZN(n3653)
         );
  OAI22_X1 U225 ( .A1(n4305), .A2(n6440), .B1(n1718), .B2(n1773), .ZN(n3628)
         );
  OAI22_X1 U215 ( .A1(n4329), .A2(n6440), .B1(n1708), .B2(n1773), .ZN(n3633)
         );
  OAI22_X1 U213 ( .A1(n4333), .A2(n6440), .B1(n1706), .B2(n1773), .ZN(n3634)
         );
  OAI22_X1 U185 ( .A1(n4388), .A2(n1772), .B1(n1678), .B2(n1773), .ZN(n3648)
         );
  OAI22_X1 U358 ( .A1(n629), .A2(n6435), .B1(n3883), .B2(n1706), .ZN(n3538) );
  OAI22_X1 U362 ( .A1(n633), .A2(n6435), .B1(n3883), .B2(n1714), .ZN(n3534) );
  OAI22_X1 U363 ( .A1(n634), .A2(n6435), .B1(n3883), .B2(n1716), .ZN(n3533) );
  OAI22_X1 U360 ( .A1(n631), .A2(n6435), .B1(n3883), .B2(n1710), .ZN(n3536) );
  OAI22_X1 U359 ( .A1(n630), .A2(n6435), .B1(n3883), .B2(n1708), .ZN(n3537) );
  OAI22_X1 U357 ( .A1(n628), .A2(n6435), .B1(n3883), .B2(n1704), .ZN(n3539) );
  OAI22_X1 U361 ( .A1(n632), .A2(n6435), .B1(n3883), .B2(n1712), .ZN(n3535) );
  OAI22_X1 U339 ( .A1(n610), .A2(n6435), .B1(n3883), .B2(n1668), .ZN(n3557) );
  OAI22_X1 U341 ( .A1(n612), .A2(n6435), .B1(n3883), .B2(n1672), .ZN(n3555) );
  OAI22_X1 U366 ( .A1(n637), .A2(n6435), .B1(n3883), .B2(n1722), .ZN(n3530) );
  OAI22_X1 U365 ( .A1(n636), .A2(n6435), .B1(n3883), .B2(n1720), .ZN(n3531) );
  OAI22_X1 U367 ( .A1(n638), .A2(n6435), .B1(n3883), .B2(n1724), .ZN(n3529) );
  OAI22_X1 U364 ( .A1(n635), .A2(n6435), .B1(n3883), .B2(n1718), .ZN(n3532) );
  OAI22_X1 U257 ( .A1(n3764), .A2(n6438), .B1(n3882), .B2(n1704), .ZN(n3603)
         );
  OAI22_X1 U259 ( .A1(n3762), .A2(n6438), .B1(n3882), .B2(n1708), .ZN(n3601)
         );
  OAI22_X1 U258 ( .A1(n3763), .A2(n6438), .B1(n3882), .B2(n1706), .ZN(n3602)
         );
  OAI22_X1 U267 ( .A1(n3754), .A2(n6438), .B1(n3882), .B2(n1724), .ZN(n3593)
         );
  OAI22_X1 U263 ( .A1(n3758), .A2(n6438), .B1(n3882), .B2(n1716), .ZN(n3597)
         );
  OAI22_X1 U265 ( .A1(n3756), .A2(n6438), .B1(n3882), .B2(n1720), .ZN(n3595)
         );
  OAI22_X1 U264 ( .A1(n3757), .A2(n6438), .B1(n3882), .B2(n1718), .ZN(n3596)
         );
  OAI22_X1 U260 ( .A1(n3761), .A2(n6438), .B1(n3882), .B2(n1710), .ZN(n3600)
         );
  OAI22_X1 U239 ( .A1(n3782), .A2(n6438), .B1(n3882), .B2(n1668), .ZN(n3621)
         );
  OAI22_X1 U262 ( .A1(n3759), .A2(n6438), .B1(n3882), .B2(n1714), .ZN(n3598)
         );
  OAI22_X1 U261 ( .A1(n3760), .A2(n6438), .B1(n3882), .B2(n1712), .ZN(n3599)
         );
  OAI22_X1 U241 ( .A1(n3780), .A2(n6438), .B1(n3882), .B2(n1672), .ZN(n3619)
         );
  OAI22_X1 U266 ( .A1(n3755), .A2(n6438), .B1(n3882), .B2(n1722), .ZN(n3594)
         );
  OAI22_X1 U1558 ( .A1(n4544), .A2(n6396), .B1(n1716), .B2(n4111), .ZN(n2829)
         );
  OAI22_X1 U1510 ( .A1(n4634), .A2(n6396), .B1(n1668), .B2(n4111), .ZN(n2853)
         );
  OAI22_X1 U1508 ( .A1(n4635), .A2(n4110), .B1(n1666), .B2(n4111), .ZN(n2854)
         );
  OAI22_X1 U1568 ( .A1(n6338), .A2(n6396), .B1(n1726), .B2(n4111), .ZN(n2824)
         );
  OAI22_X1 U1566 ( .A1(n4533), .A2(n6396), .B1(n1724), .B2(n4111), .ZN(n2825)
         );
  OAI22_X1 U1520 ( .A1(n4622), .A2(n4110), .B1(n1678), .B2(n4111), .ZN(n2848)
         );
  OAI22_X1 U1518 ( .A1(n4623), .A2(n4110), .B1(n1676), .B2(n4111), .ZN(n2849)
         );
  OAI22_X1 U1516 ( .A1(n4628), .A2(n6396), .B1(n1674), .B2(n4111), .ZN(n2850)
         );
  OAI22_X1 U1514 ( .A1(n4629), .A2(n6396), .B1(n1672), .B2(n4111), .ZN(n2851)
         );
  OAI22_X1 U1506 ( .A1(n4643), .A2(n4110), .B1(n1663), .B2(n4111), .ZN(n2855)
         );
  OAI22_X1 U1550 ( .A1(n4563), .A2(n6396), .B1(n1708), .B2(n4111), .ZN(n2833)
         );
  OAI22_X1 U1548 ( .A1(n4568), .A2(n6396), .B1(n1706), .B2(n4111), .ZN(n2834)
         );
  OAI22_X1 U1560 ( .A1(n4543), .A2(n6396), .B1(n1718), .B2(n4111), .ZN(n2828)
         );
  OAI22_X1 U1512 ( .A1(n4633), .A2(n6396), .B1(n1670), .B2(n4111), .ZN(n2852)
         );
  OAI22_X1 U1234 ( .A1(n6350), .A2(n6406), .B1(n1726), .B2(n3887), .ZN(n3016)
         );
  OAI22_X1 U332 ( .A1(n6306), .A2(n6437), .B1(n1724), .B2(n1812), .ZN(n3561)
         );
  OAI22_X1 U330 ( .A1(n6307), .A2(n6437), .B1(n1722), .B2(n1812), .ZN(n3562)
         );
  OAI22_X1 U328 ( .A1(n6308), .A2(n6437), .B1(n1720), .B2(n1812), .ZN(n3563)
         );
  OAI22_X1 U326 ( .A1(n6309), .A2(n6437), .B1(n1718), .B2(n1812), .ZN(n3564)
         );
  OAI22_X1 U324 ( .A1(n6310), .A2(n6437), .B1(n1716), .B2(n1812), .ZN(n3565)
         );
  OAI22_X1 U322 ( .A1(n6311), .A2(n6437), .B1(n1714), .B2(n1812), .ZN(n3566)
         );
  OAI22_X1 U320 ( .A1(n6312), .A2(n6437), .B1(n1712), .B2(n1812), .ZN(n3567)
         );
  OAI22_X1 U280 ( .A1(n6332), .A2(n6437), .B1(n1672), .B2(n1812), .ZN(n3587)
         );
  OAI22_X1 U282 ( .A1(n6331), .A2(n6437), .B1(n1674), .B2(n1812), .ZN(n3586)
         );
  OAI22_X1 U288 ( .A1(n6328), .A2(n6437), .B1(n1680), .B2(n1812), .ZN(n3583)
         );
  OAI22_X1 U290 ( .A1(n6327), .A2(n1811), .B1(n1682), .B2(n1812), .ZN(n3582)
         );
  OAI22_X1 U1079 ( .A1(n4802), .A2(n6412), .B1(n1706), .B2(n3927), .ZN(n3122)
         );
  OAI22_X1 U1081 ( .A1(n4793), .A2(n6412), .B1(n1708), .B2(n3927), .ZN(n3121)
         );
  OAI22_X1 U1089 ( .A1(n4779), .A2(n6412), .B1(n1716), .B2(n3927), .ZN(n3117)
         );
  OAI22_X1 U1091 ( .A1(n4778), .A2(n6412), .B1(n1718), .B2(n3927), .ZN(n3116)
         );
  OAI22_X1 U1099 ( .A1(n6341), .A2(n6412), .B1(n1726), .B2(n3927), .ZN(n3112)
         );
  OAI22_X1 U1039 ( .A1(n4873), .A2(n3926), .B1(n1666), .B2(n3927), .ZN(n3142)
         );
  OAI22_X1 U1077 ( .A1(n4803), .A2(n6412), .B1(n1704), .B2(n3927), .ZN(n3123)
         );
  OAI22_X1 U1041 ( .A1(n4869), .A2(n6412), .B1(n1668), .B2(n3927), .ZN(n3141)
         );
  OAI22_X1 U1043 ( .A1(n4868), .A2(n6412), .B1(n1670), .B2(n3927), .ZN(n3140)
         );
  OAI22_X1 U1047 ( .A1(n4862), .A2(n6412), .B1(n1674), .B2(n3927), .ZN(n3138)
         );
  OAI22_X1 U1049 ( .A1(n4853), .A2(n3926), .B1(n1676), .B2(n3927), .ZN(n3137)
         );
  OAI22_X1 U294 ( .A1(n6325), .A2(n6437), .B1(n1686), .B2(n1812), .ZN(n3580)
         );
  OAI22_X1 U272 ( .A1(n6336), .A2(n6437), .B1(n1663), .B2(n1812), .ZN(n3591)
         );
  OAI22_X1 U1045 ( .A1(n4863), .A2(n6412), .B1(n1672), .B2(n3927), .ZN(n3139)
         );
  OAI22_X1 U1051 ( .A1(n4845), .A2(n3926), .B1(n1678), .B2(n3927), .ZN(n3136)
         );
  OAI22_X1 U292 ( .A1(n6326), .A2(n6437), .B1(n1684), .B2(n1812), .ZN(n3581)
         );
  OAI22_X1 U1037 ( .A1(n4874), .A2(n3926), .B1(n1663), .B2(n3927), .ZN(n3143)
         );
  OAI22_X1 U128 ( .A1(n6012), .A2(n6442), .B1(n1688), .B2(n6441), .ZN(n3675)
         );
  OAI22_X1 U122 ( .A1(n6015), .A2(n6442), .B1(n1682), .B2(n6441), .ZN(n3678)
         );
  OAI22_X1 U124 ( .A1(n6014), .A2(n6442), .B1(n1684), .B2(n6441), .ZN(n3677)
         );
  OAI22_X1 U120 ( .A1(n6016), .A2(n6442), .B1(n1680), .B2(n6441), .ZN(n3679)
         );
  OAI22_X1 U152 ( .A1(n6000), .A2(n6442), .B1(n1712), .B2(n6441), .ZN(n3663)
         );
  OAI22_X1 U134 ( .A1(n6009), .A2(n6442), .B1(n1694), .B2(n6441), .ZN(n3672)
         );
  OAI22_X1 U126 ( .A1(n6013), .A2(n1735), .B1(n1686), .B2(n6441), .ZN(n3676)
         );
  OAI22_X1 U160 ( .A1(n5996), .A2(n6442), .B1(n1720), .B2(n6441), .ZN(n3659)
         );
  OAI22_X1 U136 ( .A1(n6008), .A2(n1735), .B1(n1696), .B2(n6441), .ZN(n3671)
         );
  OAI22_X1 U162 ( .A1(n5995), .A2(n6442), .B1(n1722), .B2(n6441), .ZN(n3658)
         );
  OAI22_X1 U154 ( .A1(n5999), .A2(n6442), .B1(n1714), .B2(n6441), .ZN(n3662)
         );
  OAI22_X1 U138 ( .A1(n6007), .A2(n6442), .B1(n1698), .B2(n6441), .ZN(n3670)
         );
  OAI22_X1 U118 ( .A1(n6017), .A2(n6442), .B1(n1678), .B2(n6441), .ZN(n3680)
         );
  OAI22_X1 U130 ( .A1(n6011), .A2(n6442), .B1(n1690), .B2(n6441), .ZN(n3674)
         );
  OAI22_X1 U132 ( .A1(n6010), .A2(n6442), .B1(n1692), .B2(n6441), .ZN(n3673)
         );
  OAI22_X1 U140 ( .A1(n6006), .A2(n1735), .B1(n1700), .B2(n6441), .ZN(n3669)
         );
  OAI22_X1 U164 ( .A1(n5994), .A2(n6442), .B1(n1724), .B2(n6441), .ZN(n3657)
         );
  OAI22_X1 U142 ( .A1(n6005), .A2(n1735), .B1(n1702), .B2(n6441), .ZN(n3668)
         );
  OAI22_X1 U715 ( .A1(n6112), .A2(n1990), .B1(n1676), .B2(n1991), .ZN(n3329)
         );
  OAI22_X1 U699 ( .A1(n6352), .A2(n6425), .B1(n1726), .B2(n1957), .ZN(n3336)
         );
  OAI22_X1 U677 ( .A1(n6285), .A2(n6425), .B1(n1704), .B2(n1957), .ZN(n3347)
         );
  OAI22_X1 U717 ( .A1(n6111), .A2(n1990), .B1(n1678), .B2(n1991), .ZN(n3328)
         );
  OAI22_X1 U641 ( .A1(n6303), .A2(n6425), .B1(n1668), .B2(n1957), .ZN(n3365)
         );
  OAI22_X1 U639 ( .A1(n6304), .A2(n1956), .B1(n1666), .B2(n1957), .ZN(n3366)
         );
  OAI22_X1 U681 ( .A1(n6283), .A2(n6425), .B1(n1708), .B2(n1957), .ZN(n3345)
         );
  OAI22_X1 U689 ( .A1(n6279), .A2(n6425), .B1(n1716), .B2(n1957), .ZN(n3341)
         );
  OAI22_X1 U691 ( .A1(n6278), .A2(n6425), .B1(n1718), .B2(n1957), .ZN(n3340)
         );
  OAI22_X1 U679 ( .A1(n6284), .A2(n6425), .B1(n1706), .B2(n1957), .ZN(n3346)
         );
  OAI22_X1 U705 ( .A1(n6117), .A2(n1990), .B1(n1666), .B2(n1991), .ZN(n3334)
         );
  OAI22_X1 U713 ( .A1(n6113), .A2(n6423), .B1(n1674), .B2(n1991), .ZN(n3330)
         );
  OAI22_X1 U709 ( .A1(n6115), .A2(n6423), .B1(n1670), .B2(n1991), .ZN(n3332)
         );
  OAI22_X1 U711 ( .A1(n6114), .A2(n6423), .B1(n1672), .B2(n1991), .ZN(n3331)
         );
  OAI22_X1 U743 ( .A1(n6098), .A2(n6423), .B1(n1704), .B2(n1991), .ZN(n3315)
         );
  OAI22_X1 U745 ( .A1(n6097), .A2(n6423), .B1(n1706), .B2(n1991), .ZN(n3314)
         );
  OAI22_X1 U747 ( .A1(n6096), .A2(n6423), .B1(n1708), .B2(n1991), .ZN(n3313)
         );
  OAI22_X1 U765 ( .A1(n6087), .A2(n6423), .B1(n1726), .B2(n1991), .ZN(n3304)
         );
  OAI22_X1 U643 ( .A1(n6302), .A2(n6425), .B1(n1670), .B2(n1957), .ZN(n3364)
         );
  OAI22_X1 U651 ( .A1(n6298), .A2(n1956), .B1(n1678), .B2(n1957), .ZN(n3360)
         );
  OAI22_X1 U755 ( .A1(n6092), .A2(n6423), .B1(n1716), .B2(n1991), .ZN(n3309)
         );
  OAI22_X1 U757 ( .A1(n6091), .A2(n6423), .B1(n1718), .B2(n1991), .ZN(n3308)
         );
  OAI22_X1 U649 ( .A1(n6299), .A2(n1956), .B1(n1676), .B2(n1957), .ZN(n3361)
         );
  OAI22_X1 U647 ( .A1(n6300), .A2(n6425), .B1(n1674), .B2(n1957), .ZN(n3362)
         );
  OAI22_X1 U645 ( .A1(n6301), .A2(n6425), .B1(n1672), .B2(n1957), .ZN(n3363)
         );
  OAI22_X1 U637 ( .A1(n6305), .A2(n1956), .B1(n1663), .B2(n1957), .ZN(n3367)
         );
  OAI22_X1 U707 ( .A1(n6116), .A2(n6423), .B1(n1668), .B2(n1991), .ZN(n3333)
         );
  OAI22_X1 U703 ( .A1(n6118), .A2(n1990), .B1(n1663), .B2(n1991), .ZN(n3335)
         );
  OAI22_X1 U613 ( .A1(n4913), .A2(n6427), .B1(n1706), .B2(n1922), .ZN(n3378)
         );
  OAI22_X1 U573 ( .A1(n4989), .A2(n1921), .B1(n1666), .B2(n1922), .ZN(n3398)
         );
  OAI22_X1 U575 ( .A1(n4988), .A2(n6427), .B1(n1668), .B2(n1922), .ZN(n3397)
         );
  OAI22_X1 U623 ( .A1(n4898), .A2(n6427), .B1(n1716), .B2(n1922), .ZN(n3373)
         );
  OAI22_X1 U611 ( .A1(n4922), .A2(n6427), .B1(n1704), .B2(n1922), .ZN(n3379)
         );
  OAI22_X1 U585 ( .A1(n4964), .A2(n1921), .B1(n1678), .B2(n1922), .ZN(n3392)
         );
  OAI22_X1 U625 ( .A1(n4893), .A2(n6427), .B1(n1718), .B2(n1922), .ZN(n3372)
         );
  OAI22_X1 U615 ( .A1(n4905), .A2(n6427), .B1(n1708), .B2(n1922), .ZN(n3377)
         );
  OAI22_X1 U579 ( .A1(n4982), .A2(n6427), .B1(n1672), .B2(n1922), .ZN(n3395)
         );
  OAI22_X1 U577 ( .A1(n4983), .A2(n6427), .B1(n1670), .B2(n1922), .ZN(n3396)
         );
  OAI22_X1 U633 ( .A1(n6342), .A2(n6427), .B1(n1726), .B2(n1922), .ZN(n3368)
         );
  OAI22_X1 U583 ( .A1(n4965), .A2(n1921), .B1(n1676), .B2(n1922), .ZN(n3393)
         );
  OAI22_X1 U571 ( .A1(n4993), .A2(n1921), .B1(n1663), .B2(n1922), .ZN(n3399)
         );
  OAI22_X1 U581 ( .A1(n4973), .A2(n6427), .B1(n1674), .B2(n1922), .ZN(n3394)
         );
  OAI22_X1 U1225 ( .A1(n694), .A2(n6406), .B1(n3887), .B2(n1708), .ZN(n3025)
         );
  OAI22_X1 U1224 ( .A1(n693), .A2(n6406), .B1(n3887), .B2(n1706), .ZN(n3026)
         );
  OAI22_X1 U1233 ( .A1(n702), .A2(n6406), .B1(n3887), .B2(n1724), .ZN(n3017)
         );
  OAI22_X1 U1232 ( .A1(n701), .A2(n6406), .B1(n3887), .B2(n1722), .ZN(n3018)
         );
  OAI22_X1 U1207 ( .A1(n676), .A2(n6406), .B1(n3887), .B2(n1672), .ZN(n3043)
         );
  OAI22_X1 U1205 ( .A1(n674), .A2(n6406), .B1(n3887), .B2(n1668), .ZN(n3045)
         );
  OAI22_X1 U1223 ( .A1(n692), .A2(n6406), .B1(n3887), .B2(n1704), .ZN(n3027)
         );
  OAI22_X1 U1227 ( .A1(n696), .A2(n6406), .B1(n3887), .B2(n1712), .ZN(n3023)
         );
  OAI22_X1 U1231 ( .A1(n700), .A2(n6406), .B1(n3887), .B2(n1720), .ZN(n3019)
         );
  OAI22_X1 U1230 ( .A1(n699), .A2(n6406), .B1(n3887), .B2(n1718), .ZN(n3020)
         );
  OAI22_X1 U1229 ( .A1(n698), .A2(n6406), .B1(n3887), .B2(n1716), .ZN(n3021)
         );
  OAI22_X1 U1226 ( .A1(n695), .A2(n6406), .B1(n3887), .B2(n1710), .ZN(n3024)
         );
  OAI22_X1 U1228 ( .A1(n697), .A2(n6406), .B1(n3887), .B2(n1714), .ZN(n3022)
         );
  OAI22_X1 U2448 ( .A1(n2087), .A2(n6392), .B1(n4181), .B2(n1726), .ZN(n2729)
         );
  OAI22_X1 U1770 ( .A1(n4509), .A2(n4180), .B1(n1674), .B2(n4181), .ZN(n2781)
         );
  OAI22_X1 U2420 ( .A1(n4418), .A2(n6392), .B1(n1724), .B2(n4181), .ZN(n2731)
         );
  OAI22_X1 U1874 ( .A1(n4493), .A2(n6392), .B1(n1682), .B2(n4181), .ZN(n2773)
         );
  OAI22_X1 U1744 ( .A1(n4513), .A2(n6392), .B1(n1672), .B2(n4181), .ZN(n2783)
         );
  OAI22_X1 U1640 ( .A1(n4532), .A2(n4180), .B1(n1663), .B2(n4181), .ZN(n2791)
         );
  OAI22_X1 U2264 ( .A1(n4442), .A2(n6392), .B1(n1712), .B2(n4181), .ZN(n2743)
         );
  OAI22_X1 U1900 ( .A1(n4485), .A2(n6392), .B1(n1684), .B2(n4181), .ZN(n2771)
         );
  OAI22_X1 U1926 ( .A1(n4484), .A2(n6392), .B1(n1686), .B2(n4181), .ZN(n2769)
         );
  OAI22_X1 U2316 ( .A1(n4425), .A2(n6392), .B1(n1716), .B2(n4181), .ZN(n2739)
         );
  OAI22_X1 U2394 ( .A1(n4419), .A2(n6392), .B1(n1722), .B2(n4181), .ZN(n2733)
         );
  OAI22_X1 U2290 ( .A1(n4433), .A2(n6392), .B1(n1714), .B2(n4181), .ZN(n2741)
         );
  OAI22_X1 U2368 ( .A1(n4423), .A2(n6392), .B1(n1720), .B2(n4181), .ZN(n2735)
         );
  OAI22_X1 U2342 ( .A1(n4424), .A2(n6392), .B1(n1718), .B2(n4181), .ZN(n2737)
         );
  OAI22_X1 U1627 ( .A1(n6184), .A2(n6394), .B1(n1718), .B2(n4146), .ZN(n2796)
         );
  OAI22_X1 U1583 ( .A1(n6206), .A2(n4145), .B1(n1674), .B2(n4146), .ZN(n2818)
         );
  OAI22_X1 U1587 ( .A1(n6204), .A2(n4145), .B1(n1678), .B2(n4146), .ZN(n2816)
         );
  OAI22_X1 U1617 ( .A1(n6189), .A2(n6394), .B1(n1708), .B2(n4146), .ZN(n2801)
         );
  OAI22_X1 U1615 ( .A1(n6190), .A2(n6394), .B1(n1706), .B2(n4146), .ZN(n2802)
         );
  OAI22_X1 U1573 ( .A1(n6211), .A2(n4145), .B1(n1663), .B2(n4146), .ZN(n2823)
         );
  OAI22_X1 U1625 ( .A1(n6185), .A2(n6394), .B1(n1716), .B2(n4146), .ZN(n2797)
         );
  OAI22_X1 U1577 ( .A1(n6209), .A2(n6394), .B1(n1668), .B2(n4146), .ZN(n2821)
         );
  OAI22_X1 U1581 ( .A1(n6207), .A2(n6394), .B1(n1672), .B2(n4146), .ZN(n2819)
         );
  OAI22_X1 U1635 ( .A1(n6347), .A2(n6394), .B1(n1726), .B2(n4146), .ZN(n2792)
         );
  OAI22_X1 U1579 ( .A1(n6208), .A2(n6394), .B1(n1670), .B2(n4146), .ZN(n2820)
         );
  OAI22_X1 U1633 ( .A1(n6181), .A2(n6394), .B1(n1724), .B2(n4146), .ZN(n2793)
         );
  OAI22_X1 U1585 ( .A1(n6205), .A2(n6394), .B1(n1676), .B2(n4146), .ZN(n2817)
         );
  OAI22_X1 U1575 ( .A1(n6210), .A2(n4145), .B1(n1666), .B2(n4146), .ZN(n2822)
         );
  OAI22_X1 U1195 ( .A1(n541), .A2(n6408), .B1(n3995), .B2(n1716), .ZN(n3053)
         );
  OAI22_X1 U1190 ( .A1(n536), .A2(n6408), .B1(n3995), .B2(n1706), .ZN(n3058)
         );
  OAI22_X1 U1170 ( .A1(n516), .A2(n3994), .B1(n3995), .B2(n1666), .ZN(n3078)
         );
  OAI22_X1 U1200 ( .A1(n671), .A2(n6408), .B1(n3995), .B2(n1726), .ZN(n3048)
         );
  OAI22_X1 U1173 ( .A1(n519), .A2(n6408), .B1(n3995), .B2(n1672), .ZN(n3075)
         );
  OAI22_X1 U1174 ( .A1(n520), .A2(n6408), .B1(n3995), .B2(n1674), .ZN(n3074)
         );
  OAI22_X1 U1199 ( .A1(n545), .A2(n6408), .B1(n3995), .B2(n1724), .ZN(n3049)
         );
  OAI22_X1 U1171 ( .A1(n517), .A2(n6408), .B1(n3995), .B2(n1668), .ZN(n3077)
         );
  OAI22_X1 U1172 ( .A1(n518), .A2(n6408), .B1(n3995), .B2(n1670), .ZN(n3076)
         );
  OAI22_X1 U1196 ( .A1(n542), .A2(n6408), .B1(n3995), .B2(n1718), .ZN(n3052)
         );
  OAI22_X1 U1191 ( .A1(n537), .A2(n6408), .B1(n3995), .B2(n1708), .ZN(n3057)
         );
  OAI22_X1 U1176 ( .A1(n522), .A2(n3994), .B1(n3995), .B2(n1678), .ZN(n3072)
         );
  OAI22_X1 U1169 ( .A1(n515), .A2(n3994), .B1(n3995), .B2(n1663), .ZN(n3079)
         );
  OAI22_X1 U1175 ( .A1(n521), .A2(n3994), .B1(n3995), .B2(n1676), .ZN(n3073)
         );
  OAI22_X1 U773 ( .A1(n708), .A2(n6421), .B1(n2024), .B2(n1672), .ZN(n3299) );
  OAI22_X1 U791 ( .A1(n726), .A2(n6421), .B1(n2024), .B2(n1708), .ZN(n3281) );
  OAI22_X1 U790 ( .A1(n725), .A2(n6421), .B1(n2024), .B2(n1706), .ZN(n3282) );
  OAI22_X1 U770 ( .A1(n705), .A2(n2023), .B1(n2024), .B2(n1666), .ZN(n3302) );
  OAI22_X1 U776 ( .A1(n711), .A2(n2023), .B1(n2024), .B2(n1678), .ZN(n3296) );
  OAI22_X1 U795 ( .A1(n730), .A2(n6421), .B1(n2024), .B2(n1716), .ZN(n3277) );
  OAI22_X1 U774 ( .A1(n709), .A2(n6421), .B1(n2024), .B2(n1674), .ZN(n3298) );
  OAI22_X1 U772 ( .A1(n707), .A2(n6421), .B1(n2024), .B2(n1670), .ZN(n3300) );
  OAI22_X1 U771 ( .A1(n706), .A2(n6421), .B1(n2024), .B2(n1668), .ZN(n3301) );
  OAI22_X1 U796 ( .A1(n731), .A2(n6421), .B1(n2024), .B2(n1718), .ZN(n3276) );
  OAI22_X1 U769 ( .A1(n704), .A2(n2023), .B1(n2024), .B2(n1663), .ZN(n3303) );
  OAI22_X1 U799 ( .A1(n734), .A2(n6421), .B1(n2024), .B2(n1724), .ZN(n3273) );
  OAI22_X1 U800 ( .A1(n513), .A2(n6421), .B1(n2024), .B2(n1726), .ZN(n3272) );
  OAI22_X1 U775 ( .A1(n710), .A2(n2023), .B1(n2024), .B2(n1676), .ZN(n3297) );
  OAI22_X1 U1129 ( .A1(n4713), .A2(n6410), .B1(n1690), .B2(n3962), .ZN(n3098)
         );
  OAI22_X1 U1121 ( .A1(n4724), .A2(n6410), .B1(n1682), .B2(n3962), .ZN(n3102)
         );
  OAI22_X1 U1103 ( .A1(n4755), .A2(n3961), .B1(n1663), .B2(n3962), .ZN(n3111)
         );
  OAI22_X1 U1107 ( .A1(n4753), .A2(n6410), .B1(n1668), .B2(n3962), .ZN(n3109)
         );
  OAI22_X1 U1117 ( .A1(n4733), .A2(n3961), .B1(n1678), .B2(n3962), .ZN(n3104)
         );
  OAI22_X1 U1133 ( .A1(n4703), .A2(n6410), .B1(n1694), .B2(n3962), .ZN(n3096)
         );
  OAI22_X1 U1141 ( .A1(n4689), .A2(n6410), .B1(n1702), .B2(n3962), .ZN(n3092)
         );
  OAI22_X1 U1123 ( .A1(n4723), .A2(n6410), .B1(n1684), .B2(n3962), .ZN(n3101)
         );
  OAI22_X1 U1105 ( .A1(n4754), .A2(n3961), .B1(n1666), .B2(n3962), .ZN(n3110)
         );
  OAI22_X1 U1115 ( .A1(n4742), .A2(n3961), .B1(n1676), .B2(n3962), .ZN(n3105)
         );
  OAI22_X1 U1131 ( .A1(n4712), .A2(n6410), .B1(n1692), .B2(n3962), .ZN(n3097)
         );
  OAI22_X1 U1119 ( .A1(n4725), .A2(n3961), .B1(n1680), .B2(n3962), .ZN(n3103)
         );
  OAI22_X1 U1111 ( .A1(n4748), .A2(n6410), .B1(n1672), .B2(n3962), .ZN(n3107)
         );
  OAI22_X1 U1474 ( .A1(n548), .A2(n6398), .B1(n4107), .B2(n1668), .ZN(n2885)
         );
  OAI22_X1 U1473 ( .A1(n547), .A2(n6398), .B1(n4107), .B2(n1666), .ZN(n2886)
         );
  OAI22_X1 U1475 ( .A1(n549), .A2(n6398), .B1(n4107), .B2(n1670), .ZN(n2884)
         );
  OAI22_X1 U1498 ( .A1(n572), .A2(n6398), .B1(n4107), .B2(n1716), .ZN(n2861)
         );
  OAI22_X1 U1477 ( .A1(n551), .A2(n6398), .B1(n4107), .B2(n1674), .ZN(n2882)
         );
  OAI22_X1 U1497 ( .A1(n571), .A2(n6398), .B1(n4107), .B2(n1714), .ZN(n2862)
         );
  OAI22_X1 U1503 ( .A1(n703), .A2(n6398), .B1(n4107), .B2(n1726), .ZN(n2856)
         );
  OAI22_X1 U1479 ( .A1(n553), .A2(n4106), .B1(n4107), .B2(n1678), .ZN(n2880)
         );
  OAI22_X1 U1492 ( .A1(n566), .A2(n4106), .B1(n4107), .B2(n1704), .ZN(n2867)
         );
  OAI22_X1 U1472 ( .A1(n546), .A2(n4106), .B1(n4107), .B2(n1663), .ZN(n2887)
         );
  OAI22_X1 U1476 ( .A1(n550), .A2(n6398), .B1(n4107), .B2(n1672), .ZN(n2883)
         );
  OAI22_X1 U1494 ( .A1(n568), .A2(n6398), .B1(n4107), .B2(n1708), .ZN(n2865)
         );
  OAI22_X1 U1493 ( .A1(n567), .A2(n6398), .B1(n4107), .B2(n1706), .ZN(n2866)
         );
  OAI22_X1 U1478 ( .A1(n552), .A2(n4106), .B1(n4107), .B2(n1676), .ZN(n2881)
         );
  OAI22_X1 U1017 ( .A1(n6063), .A2(n3892), .B1(n1710), .B2(n6413), .ZN(n3152)
         );
  OAI22_X1 U1009 ( .A1(n6067), .A2(n6414), .B1(n1702), .B2(n6413), .ZN(n3156)
         );
  OAI22_X1 U1007 ( .A1(n6068), .A2(n6414), .B1(n1700), .B2(n6413), .ZN(n3157)
         );
  OAI22_X1 U973 ( .A1(n6085), .A2(n6414), .B1(n1666), .B2(n6413), .ZN(n3174)
         );
  OAI22_X1 U1015 ( .A1(n6064), .A2(n3892), .B1(n1708), .B2(n6413), .ZN(n3153)
         );
  OAI22_X1 U1013 ( .A1(n6065), .A2(n3892), .B1(n1706), .B2(n6413), .ZN(n3154)
         );
  OAI22_X1 U1005 ( .A1(n6069), .A2(n6414), .B1(n1698), .B2(n6413), .ZN(n3158)
         );
  OAI22_X1 U999 ( .A1(n6072), .A2(n6414), .B1(n1692), .B2(n6413), .ZN(n3161)
         );
  OAI22_X1 U997 ( .A1(n6073), .A2(n6414), .B1(n1690), .B2(n6413), .ZN(n3162)
         );
  OAI22_X1 U995 ( .A1(n6074), .A2(n6414), .B1(n1688), .B2(n6413), .ZN(n3163)
         );
  OAI22_X1 U1003 ( .A1(n6070), .A2(n6414), .B1(n1696), .B2(n6413), .ZN(n3159)
         );
  OAI22_X1 U1001 ( .A1(n6071), .A2(n6414), .B1(n1694), .B2(n6413), .ZN(n3160)
         );
  OAI22_X1 U985 ( .A1(n6079), .A2(n6414), .B1(n1678), .B2(n6413), .ZN(n3168)
         );
  OAI22_X1 U983 ( .A1(n6080), .A2(n6414), .B1(n1676), .B2(n6413), .ZN(n3169)
         );
  OAI22_X1 U977 ( .A1(n6083), .A2(n6414), .B1(n1670), .B2(n6413), .ZN(n3172)
         );
  OAI22_X1 U1011 ( .A1(n6066), .A2(n6414), .B1(n1704), .B2(n6413), .ZN(n3155)
         );
  OAI22_X1 U975 ( .A1(n6084), .A2(n6414), .B1(n1668), .B2(n6413), .ZN(n3173)
         );
  OAI22_X1 U1033 ( .A1(n514), .A2(n6414), .B1(n6413), .B2(n1726), .ZN(n3144)
         );
  OAI22_X1 U943 ( .A1(n647), .A2(n3888), .B1(n3884), .B2(n1678), .ZN(n3200) );
  OAI22_X1 U953 ( .A1(n657), .A2(n3888), .B1(n3884), .B2(n1698), .ZN(n3190) );
  OAI22_X1 U950 ( .A1(n654), .A2(n3888), .B1(n3884), .B2(n1692), .ZN(n3193) );
  OAI22_X1 U941 ( .A1(n645), .A2(n3888), .B1(n3884), .B2(n1674), .ZN(n3202) );
  OAI22_X1 U954 ( .A1(n658), .A2(n3888), .B1(n3884), .B2(n1700), .ZN(n3189) );
  OAI22_X1 U949 ( .A1(n653), .A2(n3888), .B1(n3884), .B2(n1690), .ZN(n3194) );
  OAI22_X1 U955 ( .A1(n659), .A2(n3888), .B1(n3884), .B2(n1702), .ZN(n3188) );
  OAI22_X1 U951 ( .A1(n655), .A2(n6415), .B1(n3884), .B2(n1694), .ZN(n3192) );
  OAI22_X1 U946 ( .A1(n650), .A2(n6415), .B1(n3884), .B2(n1684), .ZN(n3197) );
  OAI22_X1 U947 ( .A1(n651), .A2(n3888), .B1(n3884), .B2(n1686), .ZN(n3196) );
  OAI22_X1 U944 ( .A1(n648), .A2(n3888), .B1(n3884), .B2(n1680), .ZN(n3199) );
  OAI22_X1 U945 ( .A1(n649), .A2(n3888), .B1(n3884), .B2(n1682), .ZN(n3198) );
  OAI22_X1 U948 ( .A1(n652), .A2(n3888), .B1(n3884), .B2(n1688), .ZN(n3195) );
  OAI22_X1 U952 ( .A1(n656), .A2(n6415), .B1(n3884), .B2(n1696), .ZN(n3191) );
  OAI22_X1 U967 ( .A1(n6337), .A2(n6415), .B1(n1726), .B2(n3884), .ZN(n3176)
         );
  OAI22_X1 U81 ( .A1(n589), .A2(n1730), .B1(n3885), .B2(n1688), .ZN(n3707) );
  OAI22_X1 U84 ( .A1(n592), .A2(n1730), .B1(n3885), .B2(n1694), .ZN(n3704) );
  OAI22_X1 U85 ( .A1(n593), .A2(n1730), .B1(n3885), .B2(n1696), .ZN(n3703) );
  OAI22_X1 U78 ( .A1(n586), .A2(n1730), .B1(n3885), .B2(n1682), .ZN(n3710) );
  OAI22_X1 U83 ( .A1(n591), .A2(n1730), .B1(n3885), .B2(n1692), .ZN(n3705) );
  OAI22_X1 U80 ( .A1(n588), .A2(n1730), .B1(n3885), .B2(n1686), .ZN(n3708) );
  OAI22_X1 U74 ( .A1(n582), .A2(n1730), .B1(n3885), .B2(n1674), .ZN(n3714) );
  OAI22_X1 U88 ( .A1(n596), .A2(n6443), .B1(n3885), .B2(n1702), .ZN(n3700) );
  OAI22_X1 U87 ( .A1(n595), .A2(n6443), .B1(n3885), .B2(n1700), .ZN(n3701) );
  OAI22_X1 U77 ( .A1(n585), .A2(n1730), .B1(n3885), .B2(n1680), .ZN(n3711) );
  OAI22_X1 U82 ( .A1(n590), .A2(n1730), .B1(n3885), .B2(n1690), .ZN(n3706) );
  OAI22_X1 U79 ( .A1(n587), .A2(n1730), .B1(n3885), .B2(n1684), .ZN(n3709) );
  OAI22_X1 U86 ( .A1(n594), .A2(n1730), .B1(n3885), .B2(n1698), .ZN(n3702) );
  OAI22_X1 U76 ( .A1(n584), .A2(n6443), .B1(n3885), .B2(n1678), .ZN(n3712) );
  OAI22_X1 U963 ( .A1(n667), .A2(n6415), .B1(n3884), .B2(n1718), .ZN(n3180) );
  OAI22_X1 U958 ( .A1(n662), .A2(n6415), .B1(n3884), .B2(n1708), .ZN(n3185) );
  OAI22_X1 U961 ( .A1(n665), .A2(n6415), .B1(n3884), .B2(n1714), .ZN(n3182) );
  OAI22_X1 U962 ( .A1(n666), .A2(n6415), .B1(n3884), .B2(n1716), .ZN(n3181) );
  OAI22_X1 U956 ( .A1(n660), .A2(n6415), .B1(n3884), .B2(n1704), .ZN(n3187) );
  OAI22_X1 U966 ( .A1(n670), .A2(n6415), .B1(n3884), .B2(n1724), .ZN(n3177) );
  OAI22_X1 U957 ( .A1(n661), .A2(n6415), .B1(n3884), .B2(n1706), .ZN(n3186) );
  OAI22_X1 U964 ( .A1(n668), .A2(n6415), .B1(n3884), .B2(n1720), .ZN(n3179) );
  OAI22_X1 U959 ( .A1(n663), .A2(n6415), .B1(n3884), .B2(n1710), .ZN(n3184) );
  OAI22_X1 U940 ( .A1(n644), .A2(n6415), .B1(n3884), .B2(n1672), .ZN(n3203) );
  OAI22_X1 U960 ( .A1(n664), .A2(n6415), .B1(n3884), .B2(n1712), .ZN(n3183) );
  OAI22_X1 U965 ( .A1(n669), .A2(n6415), .B1(n3884), .B2(n1722), .ZN(n3178) );
  OAI22_X1 U100 ( .A1(n6345), .A2(n6443), .B1(n1726), .B2(n3885), .ZN(n3688)
         );
  OAI22_X1 U73 ( .A1(n581), .A2(n6443), .B1(n3885), .B2(n1672), .ZN(n3715) );
  OAI22_X1 U98 ( .A1(n606), .A2(n6443), .B1(n3885), .B2(n1722), .ZN(n3690) );
  OAI22_X1 U90 ( .A1(n598), .A2(n6443), .B1(n3885), .B2(n1706), .ZN(n3698) );
  OAI22_X1 U95 ( .A1(n603), .A2(n6443), .B1(n3885), .B2(n1716), .ZN(n3693) );
  OAI22_X1 U96 ( .A1(n604), .A2(n6443), .B1(n3885), .B2(n1718), .ZN(n3692) );
  OAI22_X1 U89 ( .A1(n597), .A2(n6443), .B1(n3885), .B2(n1704), .ZN(n3699) );
  OAI22_X1 U94 ( .A1(n602), .A2(n6443), .B1(n3885), .B2(n1714), .ZN(n3694) );
  OAI22_X1 U97 ( .A1(n605), .A2(n6443), .B1(n3885), .B2(n1720), .ZN(n3691) );
  OAI22_X1 U99 ( .A1(n607), .A2(n6443), .B1(n3885), .B2(n1724), .ZN(n3689) );
  OAI22_X1 U92 ( .A1(n600), .A2(n6443), .B1(n3885), .B2(n1710), .ZN(n3696) );
  OAI22_X1 U91 ( .A1(n599), .A2(n6443), .B1(n3885), .B2(n1708), .ZN(n3697) );
  OAI22_X1 U93 ( .A1(n601), .A2(n6443), .B1(n3885), .B2(n1712), .ZN(n3695) );
  OAI22_X1 U870 ( .A1(n4298), .A2(n2062), .B1(n1663), .B2(n2063), .ZN(n3239)
         );
  OAI22_X1 U912 ( .A1(n4191), .A2(n6417), .B1(n1706), .B2(n2063), .ZN(n3218)
         );
  OAI22_X1 U910 ( .A1(n4193), .A2(n6417), .B1(n1704), .B2(n2063), .ZN(n3219)
         );
  OAI22_X1 U922 ( .A1(n4174), .A2(n6417), .B1(n1716), .B2(n2063), .ZN(n3213)
         );
  OAI22_X1 U872 ( .A1(n4293), .A2(n2062), .B1(n1666), .B2(n2063), .ZN(n3238)
         );
  OAI22_X1 U874 ( .A1(n4292), .A2(n2062), .B1(n1668), .B2(n2063), .ZN(n3237)
         );
  OAI22_X1 U932 ( .A1(n4168), .A2(n6417), .B1(n1726), .B2(n2063), .ZN(n3208)
         );
  OAI22_X1 U882 ( .A1(n4273), .A2(n2062), .B1(n1676), .B2(n2063), .ZN(n3233)
         );
  OAI22_X1 U916 ( .A1(n4177), .A2(n6417), .B1(n1710), .B2(n2063), .ZN(n3216)
         );
  OAI22_X1 U914 ( .A1(n4179), .A2(n6417), .B1(n1708), .B2(n2063), .ZN(n3217)
         );
  OAI22_X1 U876 ( .A1(n4283), .A2(n2062), .B1(n1670), .B2(n2063), .ZN(n3236)
         );
  OAI22_X1 U924 ( .A1(n4173), .A2(n6417), .B1(n1718), .B2(n2063), .ZN(n3212)
         );
  OAI22_X1 U880 ( .A1(n4274), .A2(n2062), .B1(n1674), .B2(n2063), .ZN(n3234)
         );
  OAI22_X1 U878 ( .A1(n4275), .A2(n2062), .B1(n1672), .B2(n2063), .ZN(n3235)
         );
  OAI22_X1 U844 ( .A1(n6254), .A2(n2027), .B1(n1704), .B2(n2028), .ZN(n3251)
         );
  OAI22_X1 U850 ( .A1(n6251), .A2(n6419), .B1(n1710), .B2(n2028), .ZN(n3248)
         );
  OAI22_X1 U848 ( .A1(n6252), .A2(n6419), .B1(n1708), .B2(n2028), .ZN(n3249)
         );
  OAI22_X1 U846 ( .A1(n6253), .A2(n6419), .B1(n1706), .B2(n2028), .ZN(n3250)
         );
  OAI22_X1 U816 ( .A1(n6268), .A2(n6419), .B1(n1676), .B2(n2028), .ZN(n3265)
         );
  OAI22_X1 U814 ( .A1(n6269), .A2(n2027), .B1(n1674), .B2(n2028), .ZN(n3266)
         );
  OAI22_X1 U812 ( .A1(n6270), .A2(n2027), .B1(n1672), .B2(n2028), .ZN(n3267)
         );
  OAI22_X1 U866 ( .A1(n6351), .A2(n6419), .B1(n1726), .B2(n2028), .ZN(n3240)
         );
  OAI22_X1 U808 ( .A1(n6272), .A2(n2027), .B1(n1668), .B2(n2028), .ZN(n3269)
         );
  OAI22_X1 U806 ( .A1(n6273), .A2(n2027), .B1(n1666), .B2(n2028), .ZN(n3270)
         );
  OAI22_X1 U804 ( .A1(n6274), .A2(n2027), .B1(n1663), .B2(n2028), .ZN(n3271)
         );
  OAI22_X1 U856 ( .A1(n6248), .A2(n6419), .B1(n1716), .B2(n2028), .ZN(n3245)
         );
  OAI22_X1 U858 ( .A1(n6247), .A2(n6419), .B1(n1718), .B2(n2028), .ZN(n3244)
         );
  OAI22_X1 U810 ( .A1(n6271), .A2(n2027), .B1(n1670), .B2(n2028), .ZN(n3268)
         );
  OAI22_X1 U110 ( .A1(n6021), .A2(n1735), .B1(n1670), .B2(n1736), .ZN(n3684)
         );
  OAI22_X1 U144 ( .A1(n6004), .A2(n6442), .B1(n1704), .B2(n1736), .ZN(n3667)
         );
  OAI22_X1 U158 ( .A1(n5997), .A2(n6442), .B1(n1718), .B2(n1736), .ZN(n3660)
         );
  OAI22_X1 U156 ( .A1(n5998), .A2(n6442), .B1(n1716), .B2(n1736), .ZN(n3661)
         );
  OAI22_X1 U146 ( .A1(n6003), .A2(n6442), .B1(n1706), .B2(n1736), .ZN(n3666)
         );
  OAI22_X1 U116 ( .A1(n6018), .A2(n1735), .B1(n1676), .B2(n1736), .ZN(n3681)
         );
  OAI22_X1 U166 ( .A1(n6354), .A2(n6442), .B1(n1726), .B2(n1736), .ZN(n3656)
         );
  OAI22_X1 U150 ( .A1(n6001), .A2(n6442), .B1(n1710), .B2(n1736), .ZN(n3664)
         );
  OAI22_X1 U148 ( .A1(n6002), .A2(n6442), .B1(n1708), .B2(n1736), .ZN(n3665)
         );
  OAI22_X1 U108 ( .A1(n6022), .A2(n1735), .B1(n1668), .B2(n1736), .ZN(n3685)
         );
  OAI22_X1 U106 ( .A1(n6023), .A2(n1735), .B1(n1666), .B2(n1736), .ZN(n3686)
         );
  OAI22_X1 U114 ( .A1(n6019), .A2(n1735), .B1(n1674), .B2(n1736), .ZN(n3682)
         );
  OAI22_X1 U112 ( .A1(n6020), .A2(n1735), .B1(n1672), .B2(n1736), .ZN(n3683)
         );
  OAI22_X1 U104 ( .A1(n6024), .A2(n1735), .B1(n1663), .B2(n1736), .ZN(n3687)
         );
  OAI22_X1 U1376 ( .A1(n2242), .A2(n6401), .B1(n4069), .B2(n1676), .ZN(n2945)
         );
  OAI22_X1 U1370 ( .A1(n2248), .A2(n4068), .B1(n4069), .B2(n1663), .ZN(n2951)
         );
  OAI22_X1 U1371 ( .A1(n2247), .A2(n4068), .B1(n4069), .B2(n1666), .ZN(n2950)
         );
  OAI22_X1 U372 ( .A1(n2664), .A2(n1847), .B1(n1848), .B2(n1663), .ZN(n3527)
         );
  OAI22_X1 U373 ( .A1(n2663), .A2(n1847), .B1(n1848), .B2(n1666), .ZN(n3526)
         );
  OAI22_X1 U378 ( .A1(n2658), .A2(n6434), .B1(n1848), .B2(n1676), .ZN(n3521)
         );
  OAI22_X1 U338 ( .A1(n609), .A2(n1843), .B1(n1844), .B2(n1666), .ZN(n3558) );
  OAI22_X1 U337 ( .A1(n608), .A2(n1843), .B1(n1844), .B2(n1663), .ZN(n3559) );
  OAI22_X1 U343 ( .A1(n614), .A2(n6435), .B1(n1844), .B2(n1676), .ZN(n3553) );
  OAI22_X1 U237 ( .A1(n3784), .A2(n1807), .B1(n1808), .B2(n1663), .ZN(n3623)
         );
  OAI22_X1 U243 ( .A1(n3778), .A2(n6438), .B1(n1808), .B2(n1676), .ZN(n3617)
         );
  OAI22_X1 U238 ( .A1(n3783), .A2(n1807), .B1(n1808), .B2(n1666), .ZN(n3622)
         );
  OAI22_X1 U1204 ( .A1(n673), .A2(n3996), .B1(n3997), .B2(n1666), .ZN(n3046)
         );
  OAI22_X1 U1209 ( .A1(n678), .A2(n6406), .B1(n3997), .B2(n1676), .ZN(n3041)
         );
  OAI22_X1 U1203 ( .A1(n672), .A2(n3996), .B1(n3997), .B2(n1663), .ZN(n3047)
         );
  OAI22_X1 U979 ( .A1(n6082), .A2(n6414), .B1(n1672), .B2(n3893), .ZN(n3171)
         );
  OAI22_X1 U1021 ( .A1(n6061), .A2(n6414), .B1(n1714), .B2(n3893), .ZN(n3150)
         );
  OAI22_X1 U1031 ( .A1(n6056), .A2(n6414), .B1(n1724), .B2(n3893), .ZN(n3145)
         );
  OAI22_X1 U991 ( .A1(n6076), .A2(n6414), .B1(n1684), .B2(n3893), .ZN(n3165)
         );
  OAI22_X1 U1025 ( .A1(n6059), .A2(n6414), .B1(n1718), .B2(n3893), .ZN(n3148)
         );
  OAI22_X1 U971 ( .A1(n6086), .A2(n6414), .B1(n1663), .B2(n3893), .ZN(n3175)
         );
  OAI22_X1 U1019 ( .A1(n6062), .A2(n6414), .B1(n1712), .B2(n3893), .ZN(n3151)
         );
  OAI22_X1 U987 ( .A1(n6078), .A2(n6414), .B1(n1680), .B2(n3893), .ZN(n3167)
         );
  OAI22_X1 U1027 ( .A1(n6058), .A2(n6414), .B1(n1720), .B2(n3893), .ZN(n3147)
         );
  OAI22_X1 U1029 ( .A1(n6057), .A2(n6414), .B1(n1722), .B2(n3893), .ZN(n3146)
         );
  OAI22_X1 U989 ( .A1(n6077), .A2(n6414), .B1(n1682), .B2(n3893), .ZN(n3166)
         );
  OAI22_X1 U1023 ( .A1(n6060), .A2(n6414), .B1(n1716), .B2(n3893), .ZN(n3149)
         );
  OAI22_X1 U981 ( .A1(n6081), .A2(n6414), .B1(n1674), .B2(n3893), .ZN(n3170)
         );
  OAI22_X1 U993 ( .A1(n6075), .A2(n6414), .B1(n1686), .B2(n3893), .ZN(n3164)
         );
  OAI22_X1 U937 ( .A1(n641), .A2(n6415), .B1(n3889), .B2(n1666), .ZN(n3206) );
  OAI22_X1 U939 ( .A1(n643), .A2(n6415), .B1(n3889), .B2(n1670), .ZN(n3204) );
  OAI22_X1 U942 ( .A1(n646), .A2(n6415), .B1(n3889), .B2(n1676), .ZN(n3201) );
  OAI22_X1 U936 ( .A1(n640), .A2(n6415), .B1(n3889), .B2(n1663), .ZN(n3207) );
  OAI22_X1 U938 ( .A1(n642), .A2(n6415), .B1(n3889), .B2(n1668), .ZN(n3205) );
  OAI22_X1 U72 ( .A1(n580), .A2(n6443), .B1(n1731), .B2(n1670), .ZN(n3716) );
  OAI22_X1 U75 ( .A1(n583), .A2(n6443), .B1(n1731), .B2(n1676), .ZN(n3713) );
  OAI22_X1 U70 ( .A1(n578), .A2(n6443), .B1(n1731), .B2(n1666), .ZN(n3718) );
  OAI22_X1 U71 ( .A1(n579), .A2(n6443), .B1(n1731), .B2(n1668), .ZN(n3717) );
  OAI22_X1 U69 ( .A1(n577), .A2(n6443), .B1(n1731), .B2(n1663), .ZN(n3719) );
  NOR2_X2 U3540 ( .A1(n5953), .A2(n5939), .ZN(n5264) );
  NOR2_X2 U3536 ( .A1(n5949), .A2(n5936), .ZN(n5262) );
  NOR2_X2 U3515 ( .A1(n5938), .A2(n5936), .ZN(n5213) );
  NOR2_X2 U3508 ( .A1(n5950), .A2(n5960), .ZN(n5249) );
  NOR2_X2 U3507 ( .A1(n5959), .A2(n5951), .ZN(n5248) );
  NOR2_X2 U3501 ( .A1(n5952), .A2(n5935), .ZN(n5245) );
  NOR2_X2 U3500 ( .A1(n5953), .A2(n5951), .ZN(n5244) );
  NOR2_X2 U3493 ( .A1(n5952), .A2(n5938), .ZN(n5237) );
  NOR2_X2 U3492 ( .A1(n5952), .A2(n5953), .ZN(n5236) );
  NOR2_X2 U2522 ( .A1(n5173), .A2(n5159), .ZN(n4241) );
  NOR2_X2 U2518 ( .A1(n5169), .A2(n5156), .ZN(n4240) );
  NOR2_X2 U2509 ( .A1(n5168), .A2(n5185), .ZN(n4237) );
  NOR2_X2 U2498 ( .A1(n5158), .A2(n5156), .ZN(n4186) );
  NOR2_X2 U2485 ( .A1(n5172), .A2(n5155), .ZN(n4220) );
  NAND2_X1 U3542 ( .A1(n5964), .A2(ADD_RD1[1]), .ZN(n5960) );
  NAND2_X1 U3538 ( .A1(ADD_RD1[1]), .A2(ADD_RD1[2]), .ZN(n5951) );
  NAND2_X1 U3528 ( .A1(ADD_RD1[2]), .A2(n5963), .ZN(n5948) );
  NAND2_X1 U2524 ( .A1(n5186), .A2(ADD_RD2[1]), .ZN(n5182) );
  NAND2_X1 U2520 ( .A1(ADD_RD2[2]), .A2(ADD_RD2[1]), .ZN(n5171) );
  NAND2_X1 U2511 ( .A1(ADD_RD2[2]), .A2(n5187), .ZN(n5168) );
  NOR2_X1 U3547 ( .A1(n5206), .A2(n5981), .ZN(n5977) );
  NAND3_X1 U3570 ( .A1(ADD_WR[3]), .A2(ADD_WR[2]), .A3(n1770), .ZN(n1954) );
  INV_X1 U2454 ( .A(WR), .ZN(n2025) );
  NAND3_X1 U3569 ( .A1(ADD_WR[3]), .A2(n1770), .A3(n1919), .ZN(n1850) );
  NAND3_X1 U3568 ( .A1(ADD_WR[2]), .A2(n1770), .A3(n1846), .ZN(n1806) );
  NAND3_X1 U3573 ( .A1(ADD_WR[3]), .A2(ADD_WR[2]), .A3(n3924), .ZN(n4108) );
  NAND2_X1 U1036 ( .A1(n1769), .A2(n3924), .ZN(n2060) );
  OAI21_X1 U536 ( .B1(n1733), .B2(n1850), .A(n6446), .ZN(n1885) );
  OAI21_X1 U471 ( .B1(n1728), .B2(n1850), .A(n6446), .ZN(n1852) );
  NAND3_X1 U3572 ( .A1(ADD_WR[3]), .A2(n3924), .A3(n1919), .ZN(n4033) );
  OAI21_X1 U570 ( .B1(n1768), .B2(n1850), .A(n6446), .ZN(n1917) );
  NAND3_X1 U3571 ( .A1(ADD_WR[2]), .A2(n3924), .A3(n1846), .ZN(n3959) );
  OAI21_X1 U701 ( .B1(n1728), .B2(n1954), .A(n6446), .ZN(n1956) );
  OAI21_X1 U635 ( .B1(n1805), .B2(n1954), .A(n6446), .ZN(n1921) );
  OAI21_X1 U802 ( .B1(n1768), .B2(n1954), .A(n6446), .ZN(n2023) );
  NOR2_X1 U2453 ( .A1(n2025), .A2(n5146), .ZN(n3924) );
  INV_X1 U3560 ( .A(ADD_RD1[0]), .ZN(n5966) );
  INV_X1 U3563 ( .A(ADD_RD1[3]), .ZN(n5971) );
  INV_X1 U3566 ( .A(ADD_RD1[1]), .ZN(n5963) );
  INV_X1 U3567 ( .A(ADD_RD1[4]), .ZN(n5967) );
  INV_X1 U3543 ( .A(ADD_RD1[2]), .ZN(n5964) );
  INV_X1 U2535 ( .A(ADD_RD2[2]), .ZN(n5186) );
  INV_X1 U2521 ( .A(ADD_RD2[3]), .ZN(n5194) );
  INV_X1 U2533 ( .A(ADD_RD2[1]), .ZN(n5187) );
  INV_X1 U2538 ( .A(ADD_RD2[4]), .ZN(n5190) );
  INV_X1 U2537 ( .A(ADD_RD2[0]), .ZN(n5189) );
  INV_X1 U3551 ( .A(ADD_WR[2]), .ZN(n1919) );
  OAI21_X1 U2451 ( .B1(n1768), .B2(n4108), .A(n6446), .ZN(n4180) );
  OAI21_X1 U1637 ( .B1(n4108), .B2(n1733), .A(n6446), .ZN(n4145) );
  OAI21_X1 U336 ( .B1(n1733), .B2(n1806), .A(n6446), .ZN(n1811) );
  OAI21_X1 U1202 ( .B1(n1733), .B2(n3959), .A(n6446), .ZN(n3994) );
  OAI21_X1 U370 ( .B1(n1768), .B2(n1806), .A(n6446), .ZN(n1843) );
  OAI21_X1 U1236 ( .B1(n1768), .B2(n3959), .A(n6446), .ZN(n3996) );
  OAI21_X1 U1470 ( .B1(n1768), .B2(n4033), .A(n6446), .ZN(n4073) );
  OAI21_X1 U767 ( .B1(n1733), .B2(n1954), .A(n6446), .ZN(n1990) );
  OAI21_X1 U1404 ( .B1(n1733), .B2(n4033), .A(n6446), .ZN(n4068) );
  OAI21_X1 U1035 ( .B1(n1768), .B2(n2060), .A(n6446), .ZN(n3892) );
  NAND2_X1 U3556 ( .A1(n4143), .A2(n4178), .ZN(n1805) );
  OAI21_X1 U1167 ( .B1(n1728), .B2(n3959), .A(n6446), .ZN(n3961) );
  OAI21_X1 U235 ( .B1(n1805), .B2(n1806), .A(n6446), .ZN(n1772) );
  OAI21_X1 U1101 ( .B1(n1805), .B2(n3959), .A(n6446), .ZN(n3926) );
  OAI21_X1 U405 ( .B1(n1805), .B2(n1850), .A(n6446), .ZN(n1847) );
  OAI21_X1 U1505 ( .B1(n1805), .B2(n4108), .A(n6446), .ZN(n4106) );
  INV_X1 U3555 ( .A(n1805), .ZN(n5984) );
  OAI21_X1 U1570 ( .B1(n4108), .B2(n1728), .A(n6446), .ZN(n4110) );
  OAI21_X1 U270 ( .B1(n1728), .B2(n1806), .A(n6446), .ZN(n1807) );
  OAI21_X1 U1368 ( .B1(n1728), .B2(n4033), .A(n6446), .ZN(n4035) );
  OAI21_X1 U67 ( .B1(n1728), .B2(n1729), .A(n6446), .ZN(n1662) );
  OAI21_X1 U1302 ( .B1(n1805), .B2(n4033), .A(n6446), .ZN(n4000) );
  AOI211_X1 U2526 ( .C1(n5205), .C2(n5200), .A(N4487), .B(n5197), .ZN(n4199)
         );
  AOI211_X1 U3545 ( .C1(n5980), .C2(n5977), .A(N4487), .B(n5974), .ZN(n5225)
         );
  INV_X2 U2512 ( .A(n5197), .ZN(n4235) );
  OR2_X1 U2523 ( .A1(n6387), .A2(n5182), .ZN(n5159) );
  OR2_X1 U2497 ( .A1(n6387), .A2(n5170), .ZN(n5184) );
  OR2_X1 U2519 ( .A1(n6387), .A2(n5171), .ZN(n5156) );
  OR2_X1 U2510 ( .A1(n6387), .A2(n5181), .ZN(n5185) );
  OR2_X1 U3514 ( .A1(n6371), .A2(n5950), .ZN(n5961) );
  OR2_X1 U3541 ( .A1(n6371), .A2(n5960), .ZN(n5939) );
  OR2_X1 U3527 ( .A1(n6371), .A2(n5959), .ZN(n5962) );
  OR2_X1 U3537 ( .A1(n6371), .A2(n5951), .ZN(n5936) );
  NOR2_X1 U3474 ( .A1(n5935), .A2(n5936), .ZN(n5219) );
  NOR2_X1 U2460 ( .A1(n5155), .A2(n5156), .ZN(n4192) );
  NOR2_X1 U3510 ( .A1(n5961), .A2(n5952), .ZN(n5251) );
  NOR2_X1 U3511 ( .A1(n5952), .A2(n5962), .ZN(n5250) );
  NOR2_X1 U2515 ( .A1(n5157), .A2(n5159), .ZN(n4239) );
  NOR2_X1 U3533 ( .A1(n5949), .A2(n5939), .ZN(n5263) );
  NOR2_X1 U2516 ( .A1(n5169), .A2(n5159), .ZN(n4243) );
  NOR2_X1 U3532 ( .A1(n5937), .A2(n5939), .ZN(n5261) );
  NOR2_X1 U3526 ( .A1(n5948), .A2(n5962), .ZN(n5259) );
  NOR2_X1 U2493 ( .A1(n5184), .A2(n5172), .ZN(n4228) );
  NOR2_X1 U2494 ( .A1(n5172), .A2(n5185), .ZN(n4229) );
  INV_X4 U4 ( .A(n5142), .ZN(n4233) );
  INV_X4 U6 ( .A(n5124), .ZN(n4189) );
  INV_X4 U8 ( .A(n5910), .ZN(n5216) );
  INV_X4 U10 ( .A(n5925), .ZN(n5256) );
  INV_X4 U12 ( .A(N4487), .ZN(n6446) );
  BUF_X1 U14 ( .A(n4243), .Z(n6375) );
  BUF_X2 U16 ( .A(n4229), .Z(n3880) );
  BUF_X1 U18 ( .A(n1664), .Z(n6444) );
  BUF_X1 U20 ( .A(n1773), .Z(n6439) );
  BUF_X1 U22 ( .A(n4111), .Z(n6395) );
  BUF_X1 U24 ( .A(n4181), .Z(n6391) );
  BUF_X2 U26 ( .A(n1848), .Z(n3881) );
  BUF_X1 U28 ( .A(n1991), .Z(n6422) );
  BUF_X2 U30 ( .A(n1808), .Z(n3882) );
  BUF_X1 U32 ( .A(n4146), .Z(n6393) );
  BUF_X2 U34 ( .A(n1844), .Z(n3883) );
  BUF_X2 U36 ( .A(n3889), .Z(n3884) );
  BUF_X2 U38 ( .A(n1731), .Z(n3885) );
  BUF_X2 U40 ( .A(n4069), .Z(n3886) );
  BUF_X2 U42 ( .A(n3997), .Z(n3887) );
  INV_X2 U44 ( .A(DATAIN[6]), .ZN(n1714) );
  INV_X2 U46 ( .A(DATAIN[5]), .ZN(n1716) );
  INV_X2 U48 ( .A(DATAIN[26]), .ZN(n1674) );
  INV_X2 U50 ( .A(DATAIN[4]), .ZN(n1718) );
  INV_X2 U52 ( .A(DATAIN[3]), .ZN(n1720) );
  INV_X2 U54 ( .A(DATAIN[2]), .ZN(n1722) );
  INV_X2 U56 ( .A(DATAIN[1]), .ZN(n1724) );
  INV_X2 U58 ( .A(DATAIN[0]), .ZN(n1726) );
  INV_X2 U60 ( .A(DATAIN[27]), .ZN(n1672) );
  INV_X2 U62 ( .A(DATAIN[28]), .ZN(n1670) );
  INV_X2 U64 ( .A(DATAIN[29]), .ZN(n1668) );
  INV_X2 U66 ( .A(DATAIN[21]), .ZN(n1684) );
  INV_X2 U68 ( .A(DATAIN[20]), .ZN(n1686) );
  INV_X2 U101 ( .A(DATAIN[19]), .ZN(n1688) );
  INV_X2 U102 ( .A(DATAIN[18]), .ZN(n1690) );
  INV_X2 U103 ( .A(DATAIN[22]), .ZN(n1682) );
  INV_X2 U105 ( .A(DATAIN[17]), .ZN(n1692) );
  INV_X2 U107 ( .A(DATAIN[16]), .ZN(n1694) );
  INV_X2 U109 ( .A(DATAIN[15]), .ZN(n1696) );
  INV_X2 U111 ( .A(DATAIN[23]), .ZN(n1680) );
  INV_X2 U113 ( .A(DATAIN[14]), .ZN(n1698) );
  INV_X2 U115 ( .A(DATAIN[13]), .ZN(n1700) );
  INV_X2 U117 ( .A(DATAIN[24]), .ZN(n1678) );
  INV_X2 U119 ( .A(DATAIN[12]), .ZN(n1702) );
  INV_X2 U121 ( .A(DATAIN[11]), .ZN(n1704) );
  INV_X2 U123 ( .A(DATAIN[10]), .ZN(n1706) );
  INV_X2 U125 ( .A(DATAIN[9]), .ZN(n1708) );
  INV_X2 U127 ( .A(DATAIN[8]), .ZN(n1710) );
  INV_X2 U129 ( .A(DATAIN[7]), .ZN(n1712) );
  INV_X2 U131 ( .A(DATAIN[25]), .ZN(n1676) );
  INV_X2 U133 ( .A(DATAIN[31]), .ZN(n1663) );
  INV_X2 U135 ( .A(DATAIN[30]), .ZN(n1666) );
  BUF_X1 U137 ( .A(n4221), .Z(n3891) );
  BUF_X1 U139 ( .A(n4212), .Z(n3903) );
  BUF_X2 U141 ( .A(n5259), .Z(n6360) );
  BUF_X2 U143 ( .A(n5250), .Z(n6363) );
  BUF_X2 U145 ( .A(n5261), .Z(n6358) );
  BUF_X2 U147 ( .A(n5263), .Z(n6356) );
  BUF_X2 U149 ( .A(n4239), .Z(n6378) );
  OR2_X1 U151 ( .A1(n5155), .A2(n5159), .ZN(n3950) );
  OR2_X1 U153 ( .A1(n5935), .A2(n5939), .ZN(n3952) );
  OR2_X1 U155 ( .A1(n5938), .A2(n5939), .ZN(n3953) );
  OR2_X1 U157 ( .A1(n5158), .A2(n5159), .ZN(n3951) );
  INV_X1 U159 ( .A(n4199), .ZN(n6387) );
  INV_X1 U161 ( .A(n5225), .ZN(n6371) );
  NOR2_X1 U163 ( .A1(ENABLE), .A2(N4487), .ZN(n5197) );
  NOR2_X1 U165 ( .A1(ENABLE), .A2(N4487), .ZN(n5974) );
  BUF_X1 U167 ( .A(n4036), .Z(n6402) );
  BUF_X1 U168 ( .A(n4001), .Z(n6404) );
  BUF_X1 U170 ( .A(n2063), .Z(n6416) );
  BUF_X1 U172 ( .A(n4107), .Z(n6397) );
  BUF_X1 U174 ( .A(n3962), .Z(n6409) );
  BUF_X1 U176 ( .A(n3927), .Z(n6411) );
  BUF_X1 U178 ( .A(n4074), .Z(n6399) );
  NAND2_X1 U180 ( .A1(n6446), .A2(n6410), .ZN(n3962) );
  BUF_X1 U182 ( .A(n1736), .Z(n6441) );
  NAND2_X1 U184 ( .A1(n6446), .A2(n6438), .ZN(n1808) );
  NAND2_X1 U186 ( .A1(n6446), .A2(n6434), .ZN(n1848) );
  NAND2_X1 U188 ( .A1(n6446), .A2(n6405), .ZN(n4001) );
  NAND2_X1 U190 ( .A1(n6446), .A2(n6412), .ZN(n3927) );
  NAND2_X1 U192 ( .A1(n6446), .A2(n6396), .ZN(n4111) );
  BUF_X1 U194 ( .A(n1812), .Z(n6436) );
  NAND2_X1 U196 ( .A1(n6446), .A2(n6440), .ZN(n1773) );
  NAND2_X1 U198 ( .A1(n6446), .A2(n6398), .ZN(n4107) );
  NAND2_X1 U200 ( .A1(n6446), .A2(n6417), .ZN(n2063) );
  NAND2_X1 U202 ( .A1(n6446), .A2(n6403), .ZN(n4036) );
  BUF_X1 U204 ( .A(n3995), .Z(n6407) );
  NAND2_X1 U206 ( .A1(n6446), .A2(n6445), .ZN(n1664) );
  NAND2_X1 U208 ( .A1(n6446), .A2(n6419), .ZN(n2028) );
  BUF_X2 U210 ( .A(n1772), .Z(n6440) );
  BUF_X2 U212 ( .A(n4110), .Z(n6396) );
  BUF_X2 U214 ( .A(n1662), .Z(n6445) );
  BUF_X2 U216 ( .A(n1956), .Z(n6425) );
  NAND2_X1 U218 ( .A1(n6446), .A2(n6401), .ZN(n4069) );
  BUF_X2 U220 ( .A(n4106), .Z(n6398) );
  BUF_X2 U222 ( .A(n4035), .Z(n6403) );
  BUF_X2 U224 ( .A(n3926), .Z(n6412) );
  NAND2_X1 U226 ( .A1(n6446), .A2(n6392), .ZN(n4181) );
  NAND2_X1 U228 ( .A1(n6446), .A2(n6437), .ZN(n1812) );
  NAND2_X1 U230 ( .A1(n6446), .A2(n6408), .ZN(n3995) );
  BUF_X2 U232 ( .A(n1852), .Z(n6433) );
  BUF_X2 U234 ( .A(n4000), .Z(n6405) );
  BUF_X2 U236 ( .A(n1807), .Z(n6438) );
  NAND2_X1 U269 ( .A1(n6446), .A2(n6423), .ZN(n1991) );
  BUF_X1 U271 ( .A(n2062), .Z(n6417) );
  BUF_X2 U273 ( .A(n1921), .Z(n6427) );
  BUF_X2 U275 ( .A(n3961), .Z(n6410) );
  NAND2_X1 U277 ( .A1(n6446), .A2(n6415), .ZN(n3889) );
  NAND2_X1 U279 ( .A1(n6446), .A2(n6400), .ZN(n4074) );
  NAND2_X1 U281 ( .A1(n6446), .A2(n6435), .ZN(n1844) );
  BUF_X2 U283 ( .A(n1847), .Z(n6434) );
  NAND2_X1 U285 ( .A1(n6446), .A2(n6442), .ZN(n1736) );
  NAND2_X1 U287 ( .A1(n6446), .A2(n6443), .ZN(n1731) );
  NAND2_X1 U289 ( .A1(n6446), .A2(n6394), .ZN(n4146) );
  NAND2_X1 U291 ( .A1(n6446), .A2(n6406), .ZN(n3997) );
  BUF_X2 U293 ( .A(n3892), .Z(n6414) );
  NAND2_X1 U295 ( .A1(n6446), .A2(n3892), .ZN(n3893) );
  BUF_X2 U297 ( .A(n1885), .Z(n6431) );
  BUF_X2 U299 ( .A(n1990), .Z(n6423) );
  BUF_X2 U301 ( .A(n3994), .Z(n6408) );
  BUF_X2 U303 ( .A(n1917), .Z(n6429) );
  BUF_X2 U305 ( .A(n3996), .Z(n6406) );
  BUF_X2 U307 ( .A(n2023), .Z(n6421) );
  BUF_X2 U309 ( .A(n1843), .Z(n6435) );
  BUF_X1 U311 ( .A(n1735), .Z(n6442) );
  BUF_X2 U313 ( .A(n4180), .Z(n6392) );
  BUF_X2 U315 ( .A(n4145), .Z(n6394) );
  BUF_X2 U317 ( .A(n4073), .Z(n6400) );
  BUF_X2 U319 ( .A(n4068), .Z(n6401) );
  BUF_X2 U321 ( .A(n1811), .Z(n6437) );
  INV_X1 U323 ( .A(ADD_WR[1]), .ZN(n4143) );
  BUF_X2 U325 ( .A(n4204), .Z(n6385) );
  INV_X1 U327 ( .A(ADD_WR[0]), .ZN(n4178) );
  INV_X1 U329 ( .A(ADD_WR[3]), .ZN(n1846) );
  BUF_X2 U331 ( .A(n4218), .Z(n3890) );
  BUF_X2 U333 ( .A(n4224), .Z(n3894) );
  BUF_X2 U335 ( .A(n4223), .Z(n3895) );
  BUF_X2 U369 ( .A(n4226), .Z(n3896) );
  BUF_X2 U371 ( .A(n4219), .Z(n3897) );
  BUF_X2 U404 ( .A(n4205), .Z(n3898) );
  BUF_X2 U406 ( .A(n4208), .Z(n3899) );
  BUF_X2 U408 ( .A(n4207), .Z(n3900) );
  BUF_X2 U410 ( .A(n4210), .Z(n3901) );
  BUF_X2 U412 ( .A(n4209), .Z(n3902) );
  BUF_X2 U414 ( .A(n4211), .Z(n3904) );
  BUF_X2 U416 ( .A(n5231), .Z(n3905) );
  BUF_X2 U418 ( .A(n5230), .Z(n3906) );
  BUF_X2 U420 ( .A(n5233), .Z(n3907) );
  BUF_X2 U422 ( .A(n5232), .Z(n3908) );
  BUF_X2 U424 ( .A(n5235), .Z(n3909) );
  BUF_X2 U426 ( .A(n5234), .Z(n3910) );
  BUF_X2 U428 ( .A(n5246), .Z(n3911) );
  BUF_X2 U430 ( .A(n5247), .Z(n3912) );
  BUF_X2 U432 ( .A(n5242), .Z(n3913) );
  BUF_X2 U434 ( .A(n5243), .Z(n3914) );
  NOR2_X2 U436 ( .A1(n5181), .A2(n5171), .ZN(n4225) );
  BUF_X2 U438 ( .A(n5260), .Z(n6359) );
  BUF_X2 U440 ( .A(n4238), .Z(n6379) );
  NAND2_X1 U442 ( .A1(n6446), .A2(n6433), .ZN(n1853) );
  NAND2_X1 U444 ( .A1(n6446), .A2(n6431), .ZN(n1886) );
  NAND2_X1 U446 ( .A1(n6446), .A2(n6429), .ZN(n1918) );
  NAND2_X1 U448 ( .A1(n6446), .A2(n6427), .ZN(n1922) );
  NAND2_X1 U450 ( .A1(n6446), .A2(n6425), .ZN(n1957) );
  NAND2_X1 U452 ( .A1(n6446), .A2(n6421), .ZN(n2024) );
  BUF_X2 U454 ( .A(n4228), .Z(n6382) );
  BUF_X1 U456 ( .A(n1730), .Z(n6443) );
  BUF_X1 U458 ( .A(n3888), .Z(n6415) );
  BUF_X1 U460 ( .A(n3893), .Z(n6413) );
  BUF_X1 U462 ( .A(n2028), .Z(n6418) );
  BUF_X1 U464 ( .A(n2024), .Z(n6420) );
  BUF_X1 U466 ( .A(n1922), .Z(n6426) );
  BUF_X1 U468 ( .A(n1957), .Z(n6424) );
  BUF_X1 U470 ( .A(n1918), .Z(n6428) );
  BUF_X1 U473 ( .A(n1853), .Z(n6432) );
  BUF_X1 U475 ( .A(n1886), .Z(n6430) );
  BUF_X1 U477 ( .A(n4240), .Z(n6377) );
  OAI21_X1 U479 ( .B1(n1768), .B2(n1729), .A(n6446), .ZN(n1735) );
  OAI21_X1 U481 ( .B1(n1728), .B2(n2060), .A(n6446), .ZN(n2062) );
  NAND2_X1 U483 ( .A1(ADD_WR[0]), .A2(n4143), .ZN(n1728) );
  BUF_X1 U485 ( .A(n4241), .Z(n6376) );
  BUF_X1 U487 ( .A(n4192), .Z(n6388) );
  OAI21_X1 U489 ( .B1(n1733), .B2(n1729), .A(n6446), .ZN(n1730) );
  OAI21_X1 U491 ( .B1(n1733), .B2(n2060), .A(n6446), .ZN(n3888) );
  NAND2_X1 U493 ( .A1(ADD_WR[1]), .A2(ADD_WR[0]), .ZN(n1768) );
  NAND2_X1 U495 ( .A1(ADD_WR[1]), .A2(n4178), .ZN(n1733) );
  BUF_X1 U497 ( .A(n5219), .Z(n6372) );
  BUF_X1 U499 ( .A(n5262), .Z(n6357) );
  BUF_X1 U501 ( .A(n5264), .Z(n6355) );
  BUF_X1 U503 ( .A(n4186), .Z(n6390) );
  BUF_X1 U505 ( .A(n2027), .Z(n6419) );
  NOR2_X1 U507 ( .A1(ADD_WR[4]), .A2(n2025), .ZN(n1770) );
  INV_X2 U509 ( .A(n3950), .ZN(n6381) );
  BUF_X1 U511 ( .A(n5213), .Z(n6374) );
  INV_X1 U513 ( .A(ADD_WR[4]), .ZN(n5146) );
  NOR2_X1 U515 ( .A1(ADD_WR[3]), .A2(ADD_WR[2]), .ZN(n1769) );
  INV_X2 U517 ( .A(n3952), .ZN(n6361) );
  OAI21_X1 U519 ( .B1(n1805), .B2(n2060), .A(n6446), .ZN(n2027) );
  INV_X2 U521 ( .A(n3951), .ZN(n6389) );
  BUF_X1 U523 ( .A(n4225), .Z(n6383) );
  BUF_X1 U525 ( .A(n4237), .Z(n6380) );
  BUF_X1 U527 ( .A(n5236), .Z(n6369) );
  BUF_X1 U529 ( .A(n5244), .Z(n6367) );
  BUF_X1 U531 ( .A(n5248), .Z(n6365) );
  INV_X2 U533 ( .A(n3953), .ZN(n6373) );
  INV_X2 U535 ( .A(n6387), .ZN(n6386) );
  BUF_X1 U569 ( .A(n4220), .Z(n6384) );
  OR2_X2 U572 ( .A1(n5168), .A2(n5184), .ZN(n4194) );
  OR2_X2 U574 ( .A1(n5179), .A2(n5156), .ZN(n4234) );
  INV_X2 U576 ( .A(n6371), .ZN(n6370) );
  BUF_X1 U578 ( .A(n5237), .Z(n6368) );
  BUF_X1 U580 ( .A(n5245), .Z(n6366) );
  BUF_X1 U582 ( .A(n5249), .Z(n6364) );
  BUF_X1 U584 ( .A(n5251), .Z(n6362) );
  OR2_X2 U586 ( .A1(n5948), .A2(n5961), .ZN(n5220) );
  OR2_X2 U588 ( .A1(n5958), .A2(n5936), .ZN(n5255) );
  INV_X2 U590 ( .A(n5974), .ZN(n5257) );
  NOR2_X1 U592 ( .A1(n5172), .A2(n5173), .ZN(n4211) );
  NOR2_X1 U594 ( .A1(n5948), .A2(n5937), .ZN(n5230) );
  NOR2_X1 U596 ( .A1(n5172), .A2(n5157), .ZN(n4207) );
  NOR2_X1 U598 ( .A1(n5168), .A2(n5158), .ZN(n4209) );
  NOR2_X1 U600 ( .A1(n5172), .A2(n5179), .ZN(n4219) );
  NOR2_X1 U602 ( .A1(n5168), .A2(n5179), .ZN(n4223) );
  NOR2_X1 U604 ( .A1(n5173), .A2(n5171), .ZN(n4221) );
  NOR2_X1 U606 ( .A1(n5172), .A2(n5158), .ZN(n4212) );
  NOR2_X1 U608 ( .A1(n5952), .A2(n5937), .ZN(n5232) );
  NOR2_X1 U610 ( .A1(n5948), .A2(n5938), .ZN(n5234) );
  NOR2_X1 U612 ( .A1(n5948), .A2(n5958), .ZN(n5246) );
  NOR2_X1 U614 ( .A1(n5948), .A2(n5935), .ZN(n5242) );
  NOR2_X1 U616 ( .A1(n5948), .A2(n5949), .ZN(n5231) );
  NOR2_X1 U618 ( .A1(n5170), .A2(n5182), .ZN(n4226) );
  NOR2_X1 U620 ( .A1(n5168), .A2(n5157), .ZN(n4205) );
  NOR2_X1 U622 ( .A1(n5168), .A2(n5173), .ZN(n4210) );
  NOR2_X1 U624 ( .A1(n5168), .A2(n5155), .ZN(n4218) );
  NOR2_X1 U626 ( .A1(n5181), .A2(n5182), .ZN(n4224) );
  NOR2_X1 U628 ( .A1(n5170), .A2(n5171), .ZN(n4208) );
  NOR2_X1 U630 ( .A1(n5948), .A2(n5953), .ZN(n5235) );
  NOR2_X1 U632 ( .A1(n5959), .A2(n5960), .ZN(n5247) );
  NOR2_X1 U634 ( .A1(n5952), .A2(n5958), .ZN(n5243) );
  NOR2_X1 U636 ( .A1(n5950), .A2(n5951), .ZN(n5233) );
  OAI21_X1 U638 ( .B1(ADD_WR[4]), .B2(n5983), .A(WR), .ZN(n5206) );
  AOI22_X1 U640 ( .A1(ADD_WR[1]), .A2(ADD_RD1[1]), .B1(n5963), .B2(n4143), 
        .ZN(n5979) );
  AOI22_X1 U642 ( .A1(ADD_WR[1]), .A2(ADD_RD2[1]), .B1(n5187), .B2(n4143), 
        .ZN(n5201) );
  AOI22_X1 U644 ( .A1(ADD_WR[0]), .A2(ADD_RD1[0]), .B1(n5966), .B2(n4178), 
        .ZN(n5978) );
  AOI22_X1 U646 ( .A1(ADD_WR[0]), .A2(ADD_RD2[0]), .B1(n5189), .B2(n4178), 
        .ZN(n5202) );
  AOI22_X1 U648 ( .A1(ADD_WR[3]), .A2(ADD_RD1[3]), .B1(n5971), .B2(n1846), 
        .ZN(n5973) );
endmodule



    module dlx_cu_MICROCODE_MEM_SIZE64_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE13 ( 
        Clk, Rst, IR_IN, stall_exe_i, mispredict_i, D1_i, D2_i, S1_LATCH_EN, 
        S2_LATCH_EN, S3_LATCH_EN, S_MUX_PC_BUS, S_EXT, S_EXT_SIGN, S_EQ_NEQ, 
        S_MUX_DEST, S_MUX_LINK, S_MEM_W_R, S_MEM_EN, S_RF_W_wb, S_RF_W_mem, 
        S_RF_W_exe, S_MUX_ALUIN, stall_exe_o, stall_dec_o, stall_fetch_o, 
        stall_btb_o, was_branch_o, was_jmp_o, ALU_WORD_o, .ALU_OPCODE({
        \ALU_OPCODE[4] , \ALU_OPCODE[3] , \ALU_OPCODE[2] , \ALU_OPCODE[1] , 
        \ALU_OPCODE[0] }), S_MUX_MEM_BAR );
  input [31:0] IR_IN;
  input [4:0] D1_i;
  input [4:0] D2_i;
  output [1:0] S_MUX_PC_BUS;
  output [1:0] S_MUX_DEST;
  output [12:0] ALU_WORD_o;
  input Clk, Rst, stall_exe_i, mispredict_i;
  output S1_LATCH_EN, S2_LATCH_EN, S3_LATCH_EN, S_EXT, S_EXT_SIGN, S_EQ_NEQ,
         S_MUX_LINK, S_MEM_W_R, S_MEM_EN, S_RF_W_wb, S_RF_W_mem, S_RF_W_exe,
         S_MUX_ALUIN, stall_exe_o, stall_dec_o, stall_fetch_o, stall_btb_o,
         was_branch_o, was_jmp_o, \ALU_OPCODE[4] , \ALU_OPCODE[3] ,
         \ALU_OPCODE[2] , \ALU_OPCODE[1] , \ALU_OPCODE[0] , S_MUX_MEM_BAR;
  wire   IR_IN_10, IR_IN_9, IR_IN_8, IR_IN_7, IR_IN_6, IR_IN_5, IR_IN_4,
         IR_IN_3, IR_IN_2, IR_IN_1, IR_IN_0, stall_exe_i, S_MEM_LOAD,
         S_EXE_LOAD, next_bubble_dec, stall_fetch_o_TEMP, N29, N30, N31, N32,
         n138, n139, n140, n143, n150, n151, n152, n153, n154, n155, n156,
         n157, n159, n2, n119, n123, net644355, net644356, n35, n36, n37, n38,
         n39, n40, n41, n42, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n141,
         n149, n158, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n142, n147, stall_btb_o, n173, n174, n175;
  wire   [12:0] cw_from_mem;
  wire   [4:0] aluOpcode_d;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign IR_IN_10 = IR_IN[10];
  assign IR_IN_9 = IR_IN[9];
  assign IR_IN_8 = IR_IN[8];
  assign IR_IN_7 = IR_IN[7];
  assign IR_IN_6 = IR_IN[6];
  assign IR_IN_5 = IR_IN[5];
  assign IR_IN_4 = IR_IN[4];
  assign IR_IN_3 = IR_IN[3];
  assign IR_IN_2 = IR_IN[2];
  assign IR_IN_1 = IR_IN[1];
  assign IR_IN_0 = IR_IN[0];
  assign stall_exe_o = stall_exe_i;
  assign stall_dec_o = stall_btb_o;
  assign stall_fetch_o = stall_btb_o;

  DFF_X1 bubble_dec_reg ( .D(n157), .CK(Clk), .Q(n119), .QN(n173) );
  DFFR_X1 \cw_e_reg[0]  ( .D(n156), .CK(Clk), .RN(n175), .QN(n123) );
  DFFR_X1 \cw_e_reg[5]  ( .D(n154), .CK(Clk), .RN(n175), .Q(S_MUX_DEST[1]), 
        .QN(n139) );
  DFFR_X1 \cw_e_reg[4]  ( .D(n153), .CK(Clk), .RN(n175), .Q(S_MUX_DEST[0]), 
        .QN(n138) );
  DFFR_X1 \cw_e_reg[3]  ( .D(n152), .CK(Clk), .RN(n175), .QN(n2) );
  DFFR_X1 \cw_e_reg[2]  ( .D(n151), .CK(Clk), .RN(n175), .Q(net644356) );
  DFFR_X1 \cw_e_reg[1]  ( .D(n150), .CK(Clk), .RN(n175), .Q(net644355) );
  DFFR_X1 \cw_m_reg[2]  ( .D(N31), .CK(Clk), .RN(n175), .Q(S_MEM_W_R) );
  DFFR_X1 \cw_m_reg[3]  ( .D(N32), .CK(Clk), .RN(n175), .Q(S_MEM_EN), .QN(n159) );
  DFFR_X1 \cw_m_reg[0]  ( .D(N29), .CK(Clk), .RN(n175), .Q(S_RF_W_mem), .QN(
        n143) );
  XOR2_X1 U145 ( .A(S_MUX_PC_BUS[1]), .B(S_MUX_PC_BUS[0]), .Z(was_jmp_o) );
  MUX2_X1 U146 ( .A(next_bubble_dec), .B(n119), .S(Rst), .Z(n157) );
  NAND3_X1 U147 ( .A1(n174), .A2(n67), .A3(n68), .ZN(n66) );
  NAND3_X1 U148 ( .A1(IR_IN_5), .A2(IR_IN_0), .A3(IR_IN_4), .ZN(n80) );
  NAND3_X1 U149 ( .A1(n137), .A2(n77), .A3(n100), .ZN(n72) );
  NAND3_X1 U150 ( .A1(IR_IN[30]), .A2(n174), .A3(n93), .ZN(n164) );
  NAND3_X1 U151 ( .A1(n116), .A2(n117), .A3(n141), .ZN(n167) );
  NAND3_X1 U152 ( .A1(IR_IN_1), .A2(IR_IN_3), .A3(n75), .ZN(n62) );
  NAND3_X1 U153 ( .A1(IR_IN_5), .A2(IR_IN_4), .A3(n100), .ZN(n61) );
  stall_logic_FUNC_SIZE11_OP_CODE_SIZE6 STALL_L ( .OPCODE_i({IR_IN[31:29], 
        n174, n147, IR_IN[26]}), .FUNC_i({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .rA_i(IR_IN[25:21]), .rB_i(
        IR_IN[20:16]), .D1_i(D1_i), .D2_i(D2_i), .S_mem_LOAD_i(S_MEM_LOAD), 
        .S_exe_LOAD_i(S_EXE_LOAD), .S_MUX_PC_BUS_i({1'b0, 1'b0}), 
        .mispredict_i(mispredict_i), .bubble_dec_o(next_bubble_dec), 
        .stall_fetch_o(stall_fetch_o_TEMP), .S_exe_WRITE_i_BAR(n123) );
  cw_mem_MICROCODE_MEM_SIZE64_OP_CODE_SIZE6_CW_SIZE13 CWM ( .OPCODE_IN(
        IR_IN[31:26]), .CW_OUT({cw_from_mem[12:6], SYNOPSYS_UNCONNECTED__0, 
        cw_from_mem[4:0]}) );
  alu_ctrl ALU_C ( .OP(aluOpcode_d), .ALU_WORD(ALU_WORD_o) );
  DFFR_X1 \cw_m_reg[1]  ( .D(N30), .CK(Clk), .RN(n175), .QN(S_MUX_MEM_BAR) );
  AND2_X1 U137 ( .A1(cw_from_mem[8]), .A2(n173), .ZN(S_EQ_NEQ) );
  NOR4_X1 U116 ( .A1(IR_IN_7), .A2(IR_IN_9), .A3(IR_IN_8), .A4(IR_IN_6), .ZN(
        n169) );
  NAND4_X1 U112 ( .A1(n169), .A2(n170), .A3(n106), .A4(n165), .ZN(n168) );
  NAND2_X1 U37 ( .A1(IR_IN_5), .A2(IR_IN_4), .ZN(n50) );
  NAND2_X1 U70 ( .A1(IR_IN_5), .A2(IR_IN_0), .ZN(n54) );
  NAND4_X1 U77 ( .A1(IR_IN_2), .A2(n59), .A3(IR_IN_3), .A4(n99), .ZN(n55) );
  NOR2_X1 U36 ( .A1(n61), .A2(n62), .ZN(n60) );
  NAND2_X1 U52 ( .A1(IR_IN[26]), .A2(n82), .ZN(n57) );
  OAI211_X1 U34 ( .C1(n54), .C2(n55), .A(n56), .B(n57), .ZN(n52) );
  NOR2_X1 U106 ( .A1(IR_IN_0), .A2(n99), .ZN(n116) );
  NOR3_X1 U102 ( .A1(n124), .A2(n168), .A3(n75), .ZN(n117) );
  NOR3_X1 U101 ( .A1(IR_IN_5), .A2(n166), .A3(n167), .ZN(n83) );
  NAND2_X1 U64 ( .A1(n59), .A2(n76), .ZN(n114) );
  NOR2_X1 U128 ( .A1(IR_IN_5), .A2(IR_IN_4), .ZN(n115) );
  NAND4_X1 U63 ( .A1(IR_IN_3), .A2(n115), .A3(n116), .A4(n117), .ZN(n94) );
  OAI21_X1 U62 ( .B1(n62), .B2(n114), .A(n94), .ZN(n84) );
  OAI221_X1 U45 ( .B1(n55), .B2(n61), .C1(n55), .C2(n80), .A(n81), .ZN(n53) );
  NOR2_X1 U33 ( .A1(n52), .A2(n53), .ZN(n51) );
  NAND2_X1 U59 ( .A1(n106), .A2(n107), .ZN(n86) );
  NAND2_X1 U79 ( .A1(n82), .A2(n124), .ZN(n64) );
  NAND2_X1 U127 ( .A1(IR_IN_0), .A2(IR_IN_1), .ZN(n78) );
  AOI22_X1 U43 ( .A1(IR_IN_1), .A2(n76), .B1(n77), .B2(n78), .ZN(n74) );
  NOR3_X1 U42 ( .A1(IR_IN_3), .A2(n74), .A3(n75), .ZN(n69) );
  NAND2_X1 U108 ( .A1(n77), .A2(n75), .ZN(n96) );
  NOR2_X1 U107 ( .A1(n141), .A2(n96), .ZN(n73) );
  NOR3_X1 U85 ( .A1(IR_IN_1), .A2(n75), .A3(n141), .ZN(n137) );
  OAI211_X1 U40 ( .C1(n61), .C2(n62), .A(n71), .B(n72), .ZN(n70) );
  OAI21_X1 U39 ( .B1(n69), .B2(n70), .A(n59), .ZN(n65) );
  NAND4_X1 U38 ( .A1(n63), .A2(n64), .A3(n65), .A4(n66), .ZN(aluOpcode_d[3])
         );
  NAND2_X1 U124 ( .A1(n100), .A2(n99), .ZN(n133) );
  NAND2_X1 U84 ( .A1(n59), .A2(n73), .ZN(n128) );
  OAI21_X1 U81 ( .B1(n105), .B2(n87), .A(n107), .ZN(n134) );
  OAI211_X1 U78 ( .C1(n133), .C2(n128), .A(n134), .B(n64), .ZN(n131) );
  AOI221_X1 U76 ( .B1(n99), .B2(n55), .C1(n49), .C2(n55), .A(n61), .ZN(n132)
         );
  AOI211_X1 U75 ( .C1(n59), .C2(n104), .A(n131), .B(n132), .ZN(n108) );
  NOR2_X1 U73 ( .A1(n128), .A2(n78), .ZN(n127) );
  OAI21_X1 U69 ( .B1(IR_IN_5), .B2(IR_IN_2), .A(n54), .ZN(n118) );
  NOR3_X1 U68 ( .A1(n118), .A2(IR_IN_4), .A3(n99), .ZN(n112) );
  NOR2_X1 U66 ( .A1(IR_IN_1), .A2(n80), .ZN(n103) );
  AOI221_X1 U61 ( .B1(n112), .B2(n113), .C1(n103), .C2(n113), .A(n84), .ZN(
        n111) );
  NAND4_X1 U60 ( .A1(n108), .A2(n109), .A3(n110), .A4(n111), .ZN(
        aluOpcode_d[1]) );
  AOI21_X1 U122 ( .B1(n78), .B2(n133), .A(n75), .ZN(n171) );
  NOR2_X1 U121 ( .A1(IR_IN_1), .A2(n100), .ZN(n172) );
  AOI221_X1 U117 ( .B1(n115), .B2(n171), .C1(n172), .C2(n77), .A(n97), .ZN(
        n129) );
  NAND2_X1 U105 ( .A1(n73), .A2(n116), .ZN(n102) );
  OAI21_X1 U104 ( .B1(n62), .B2(n61), .A(n102), .ZN(n149) );
  NAND2_X1 U96 ( .A1(n67), .A2(n165), .ZN(n160) );
  AOI21_X1 U88 ( .B1(n162), .B2(n126), .A(n163), .ZN(n161) );
  OAI221_X1 U87 ( .B1(n124), .B2(n160), .C1(IR_IN[26]), .C2(n85), .A(n161), 
        .ZN(n158) );
  AOI211_X1 U86 ( .C1(n59), .C2(n149), .A(n83), .B(n158), .ZN(n130) );
  OAI211_X1 U74 ( .C1(n129), .C2(n49), .A(n130), .B(n108), .ZN(aluOpcode_d[0])
         );
  AOI21_X1 U57 ( .B1(IR_IN_2), .B2(n103), .A(n104), .ZN(n101) );
  OAI211_X1 U56 ( .C1(n96), .C2(n100), .A(n101), .B(n102), .ZN(n90) );
  NOR2_X1 U55 ( .A1(n99), .A2(n80), .ZN(n98) );
  AOI22_X1 U54 ( .A1(IR_IN_2), .A2(n97), .B1(n98), .B2(n75), .ZN(n95) );
  AOI21_X1 U53 ( .B1(n95), .B2(n96), .A(n49), .ZN(n91) );
  AOI211_X1 U50 ( .C1(n59), .C2(n90), .A(n91), .B(n92), .ZN(n89) );
  NOR2_X1 U19 ( .A1(n119), .A2(stall_btb_o), .ZN(n37) );
  AOI22_X1 U18 ( .A1(stall_exe_i), .A2(net644355), .B1(n37), .B2(
        cw_from_mem[1]), .ZN(n42) );
  AOI22_X1 U16 ( .A1(stall_exe_i), .A2(net644356), .B1(n37), .B2(
        cw_from_mem[2]), .ZN(n41) );
  INV_X1 U143 ( .A(stall_exe_i), .ZN(n35) );
  NAND2_X1 U10 ( .A1(n37), .A2(cw_from_mem[6]), .ZN(n38) );
  OAI21_X1 U8 ( .B1(n140), .B2(n35), .A(n38), .ZN(n155) );
  OAI21_X1 U9 ( .B1(n139), .B2(n35), .A(n38), .ZN(n154) );
  NAND2_X1 U14 ( .A1(n37), .A2(cw_from_mem[3]), .ZN(n40) );
  OAI21_X1 U13 ( .B1(n35), .B2(n2), .A(n40), .ZN(n152) );
  NAND2_X1 U12 ( .A1(n37), .A2(cw_from_mem[4]), .ZN(n39) );
  OAI21_X1 U11 ( .B1(n35), .B2(n138), .A(n39), .ZN(n153) );
  NAND2_X1 U7 ( .A1(n37), .A2(cw_from_mem[0]), .ZN(n36) );
  OAI21_X1 U6 ( .B1(n35), .B2(n123), .A(n36), .ZN(n156) );
  NOR2_X1 U140 ( .A1(stall_exe_i), .A2(n2), .ZN(N32) );
  NOR2_X1 U144 ( .A1(stall_exe_i), .A2(n123), .ZN(N29) );
  AND2_X2 U131 ( .A1(cw_from_mem[7]), .A2(n173), .ZN(S_MUX_LINK) );
  NOR2_X1 U111 ( .A1(IR_IN[26]), .A2(n168), .ZN(n59) );
  NAND2_X1 U109 ( .A1(n59), .A2(n141), .ZN(n49) );
  INV_X1 U103 ( .A(IR_IN[26]), .ZN(n124) );
  OAI21_X1 U32 ( .B1(n49), .B2(n50), .A(n51), .ZN(aluOpcode_d[4]) );
  OAI211_X1 U49 ( .C1(n87), .C2(n86), .A(n88), .B(n89), .ZN(aluOpcode_d[2]) );
  NOR2_X1 U136 ( .A1(net644356), .A2(n2), .ZN(S_EXE_LOAD) );
  DFFR_X2 \cw_e_reg[6]  ( .D(n155), .CK(Clk), .RN(n175), .Q(S_MUX_ALUIN), .QN(
        n140) );
  INV_X1 U120 ( .A(IR_IN_4), .ZN(n166) );
  INV_X1 U126 ( .A(IR_IN_0), .ZN(n100) );
  INV_X1 U125 ( .A(IR_IN_1), .ZN(n99) );
  INV_X1 U123 ( .A(IR_IN_2), .ZN(n75) );
  INV_X1 U110 ( .A(IR_IN_3), .ZN(n141) );
  INV_X1 U65 ( .A(n80), .ZN(n76) );
  AND2_X1 U119 ( .A1(n166), .A2(IR_IN_5), .ZN(n77) );
  AND2_X1 U97 ( .A1(n135), .A2(n107), .ZN(n67) );
  INV_X1 U118 ( .A(n61), .ZN(n97) );
  INV_X1 U92 ( .A(n68), .ZN(n162) );
  INV_X1 U48 ( .A(n86), .ZN(n79) );
  INV_X1 U47 ( .A(n85), .ZN(n58) );
  INV_X1 U41 ( .A(n73), .ZN(n71) );
  INV_X1 U67 ( .A(n49), .ZN(n113) );
  AND2_X1 U141 ( .A1(n35), .A2(net644356), .ZN(N31) );
  AND2_X1 U5 ( .A1(S_MUX_PC_BUS[1]), .A2(S_MUX_PC_BUS[0]), .ZN(was_branch_o)
         );
  INV_X1 U17 ( .A(n42), .ZN(n150) );
  INV_X1 U15 ( .A(n41), .ZN(n151) );
  DFFS_X1 \cw_w_reg[0]  ( .D(n143), .CK(Clk), .SN(n175), .QN(S_RF_W_wb) );
  OAI21_X1 U3 ( .B1(n78), .B2(n142), .A(n72), .ZN(n104) );
  OR2_X1 U4 ( .A1(n96), .A2(IR_IN_3), .ZN(n142) );
  AND2_X1 U20 ( .A1(n173), .A2(cw_from_mem[10]), .ZN(S_EXT) );
  AND2_X1 U21 ( .A1(n173), .A2(cw_from_mem[11]), .ZN(S_MUX_PC_BUS[0]) );
  NOR2_X1 U22 ( .A1(n159), .A2(S_MEM_W_R), .ZN(S_MEM_LOAD) );
  OR2_X2 U23 ( .A1(stall_exe_i), .A2(stall_fetch_o_TEMP), .ZN(stall_btb_o) );
  INV_X1 U24 ( .A(n165), .ZN(n147) );
  INV_X1 U25 ( .A(n174), .ZN(n106) );
  INV_X1 U26 ( .A(Rst), .ZN(n175) );
  AND2_X2 U27 ( .A1(cw_from_mem[9]), .A2(n173), .ZN(S_EXT_SIGN) );
  AND2_X1 U28 ( .A1(net644355), .A2(n35), .ZN(N30) );
  INV_X1 U29 ( .A(IR_IN[27]), .ZN(n165) );
  INV_X1 U30 ( .A(IR_IN[30]), .ZN(n135) );
  AND2_X1 U31 ( .A1(cw_from_mem[12]), .A2(n173), .ZN(S_MUX_PC_BUS[1]) );
  BUF_X1 U35 ( .A(IR_IN[28]), .Z(n174) );
  NOR2_X1 U44 ( .A1(IR_IN[29]), .A2(n164), .ZN(n126) );
  INV_X1 U46 ( .A(IR_IN[29]), .ZN(n136) );
  AOI21_X1 U51 ( .B1(n105), .B2(IR_IN[31]), .A(n83), .ZN(n88) );
  AOI22_X1 U58 ( .A1(IR_IN[31]), .A2(n58), .B1(n59), .B2(n60), .ZN(n56) );
  OAI221_X1 U71 ( .B1(IR_IN[31]), .B2(n64), .C1(n93), .C2(n57), .A(n94), .ZN(
        n92) );
  NOR2_X1 U72 ( .A1(IR_IN[31]), .A2(n136), .ZN(n107) );
  AOI211_X1 U80 ( .C1(n82), .C2(IR_IN[31]), .A(n83), .B(n84), .ZN(n81) );
  INV_X1 U82 ( .A(IR_IN[31]), .ZN(n93) );
  AOI211_X1 U83 ( .C1(IR_IN[30]), .C2(n79), .A(n58), .B(n53), .ZN(n63) );
  NOR4_X1 U89 ( .A1(IR_IN_10), .A2(IR_IN[31]), .A3(IR_IN[29]), .A4(IR_IN[30]), 
        .ZN(n170) );
  NOR3_X1 U90 ( .A1(n174), .A2(n135), .A3(n136), .ZN(n125) );
  NOR3_X1 U91 ( .A1(IR_IN[30]), .A2(n174), .A3(n68), .ZN(n105) );
  AOI21_X1 U93 ( .B1(n147), .B2(n126), .A(n127), .ZN(n109) );
  OAI221_X1 U94 ( .B1(n124), .B2(n125), .C1(IR_IN[26]), .C2(n67), .A(n147), 
        .ZN(n110) );
  NOR3_X1 U95 ( .A1(n164), .A2(IR_IN[26]), .A3(n147), .ZN(n163) );
  NAND2_X1 U98 ( .A1(n147), .A2(n125), .ZN(n85) );
  NOR3_X1 U99 ( .A1(IR_IN[26]), .A2(n147), .A3(n135), .ZN(n87) );
  NAND2_X1 U100 ( .A1(IR_IN[26]), .A2(n147), .ZN(n68) );
  NOR4_X1 U113 ( .A1(n147), .A2(n135), .A3(n136), .A4(n106), .ZN(n82) );
endmodule


module jump_logic ( NPCF_i, IR_i, A_i, A_o, rA_o, rB_o, rC_o, branch_target_o, 
        sum_addr_o, extended_imm, taken_o, FW_X_i, FW_W_i, S_FW_Adec_i, 
        S_EXT_i, S_EXT_SIGN_i, S_MUX_LINK_i, S_EQ_NEQ_i );
  input [31:0] NPCF_i;
  input [31:0] IR_i;
  input [31:0] A_i;
  output [31:0] A_o;
  output [4:0] rA_o;
  output [4:0] rB_o;
  output [4:0] rC_o;
  output [31:0] branch_target_o;
  output [31:0] sum_addr_o;
  output [31:0] extended_imm;
  input [31:0] FW_X_i;
  input [31:0] FW_W_i;
  input [1:0] S_FW_Adec_i;
  input S_EXT_i, S_EXT_SIGN_i, S_MUX_LINK_i, S_EQ_NEQ_i;
  output taken_o;
  wire   \IR_i[25] , \IR_i[24] , \IR_i[23] , \IR_i[22] , \IR_i[21] ,
         \IR_i[20] , \IR_i[19] , \IR_i[18] , \IR_i[17] , \IR_i[16] ,
         \IR_i[15] , \IR_i[14] , \IR_i[13] , \IR_i[12] , \IR_i[11] ,
         branch_sel, n1, n2;
  wire   [31:0] ext_imm;
  assign rA_o[4] = \IR_i[25] ;
  assign \IR_i[25]  = IR_i[25];
  assign rA_o[3] = \IR_i[24] ;
  assign \IR_i[24]  = IR_i[24];
  assign rA_o[2] = \IR_i[23] ;
  assign \IR_i[23]  = IR_i[23];
  assign rA_o[1] = \IR_i[22] ;
  assign \IR_i[22]  = IR_i[22];
  assign rA_o[0] = \IR_i[21] ;
  assign \IR_i[21]  = IR_i[21];
  assign rB_o[4] = \IR_i[20] ;
  assign \IR_i[20]  = IR_i[20];
  assign rB_o[3] = \IR_i[19] ;
  assign \IR_i[19]  = IR_i[19];
  assign rB_o[2] = \IR_i[18] ;
  assign \IR_i[18]  = IR_i[18];
  assign rB_o[1] = \IR_i[17] ;
  assign \IR_i[17]  = IR_i[17];
  assign rB_o[0] = \IR_i[16] ;
  assign \IR_i[16]  = IR_i[16];
  assign rC_o[4] = \IR_i[15] ;
  assign \IR_i[15]  = IR_i[15];
  assign rC_o[3] = \IR_i[14] ;
  assign \IR_i[14]  = IR_i[14];
  assign rC_o[2] = \IR_i[13] ;
  assign \IR_i[13]  = IR_i[13];
  assign rC_o[1] = \IR_i[12] ;
  assign \IR_i[12]  = IR_i[12];
  assign rC_o[0] = \IR_i[11] ;
  assign \IR_i[11]  = IR_i[11];

  extender_32 EXTENDER ( .IN1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, \IR_i[25] , 
        \IR_i[24] , \IR_i[23] , \IR_i[22] , \IR_i[21] , \IR_i[20] , \IR_i[19] , 
        \IR_i[18] , \IR_i[17] , \IR_i[16] , \IR_i[15] , \IR_i[14] , \IR_i[13] , 
        \IR_i[12] , \IR_i[11] , IR_i[10:0]}), .CTRL(S_EXT_i), .SIGN(
        S_EXT_SIGN_i), .OUT1({ext_imm[31:20], n1, ext_imm[18:0]}) );
  p4add_N32_logN5_0 JUMPADDER ( .A(NPCF_i), .B({ext_imm[31:20], n1, 
        ext_imm[18:0]}), .Cin(1'b0), .sign(1'b0), .S(sum_addr_o) );
  mux21_2 BRANCHMUX ( .IN0(sum_addr_o), .IN1(NPCF_i), .CTRL(branch_sel), 
        .OUT1(branch_target_o) );
  zerocheck ZC ( .IN0(A_o), .CTRL(S_EQ_NEQ_i), .OUT1(branch_sel) );
  mux21_4 MUXLINK ( .IN0({ext_imm[31:28], ext_imm[31], ext_imm[26:20], n1, 
        ext_imm[18:0]}), .IN1(NPCF_i), .CTRL(S_MUX_LINK_i), .OUT1(extended_imm) );
  mux41_MUX_SIZE32 MUX_FWA ( .IN0(A_i), .IN1(FW_X_i), .IN2(FW_W_i), .IN3({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CTRL(S_FW_Adec_i), .OUT1(
        A_o) );
  CLKBUF_X1 U2 ( .A(branch_sel), .Z(n2) );
  INV_X1 U3 ( .A(n2), .ZN(taken_o) );
endmodule


module fetch_regs ( NPCF_i, IR_i, NPCF_o, IR_o, stall_i, clk, rst );
  input [31:0] NPCF_i;
  input [31:0] IR_i;
  output [31:0] NPCF_o;
  output [31:0] IR_o;
  input stall_i, clk, rst;
  wire   n2;

  ff32_en_1 NPCF ( .D(NPCF_i), .en(n2), .clk(clk), .rst(rst), .Q(NPCF_o) );
  ff32_en_IR IR ( .D(IR_i), .en(n2), .clk(clk), .rst(rst), .Q(IR_o) );
  INV_X4 U1 ( .A(stall_i), .ZN(n2) );
endmodule


module btb_N_LINES4_SIZE32 ( clock, reset, stall_i, TAG_i, target_PC_i, 
        was_taken_i, predicted_next_PC_o, taken_o, mispredict_o );
  input [3:0] TAG_i;
  input [31:0] target_PC_i;
  output [31:0] predicted_next_PC_o;
  input clock, reset, stall_i, was_taken_i;
  output taken_o, mispredict_o;
  wire   \predict_PC[0][31] , \predict_PC[0][30] , \predict_PC[0][29] ,
         \predict_PC[0][28] , \predict_PC[0][27] , \predict_PC[0][26] ,
         \predict_PC[0][25] , \predict_PC[0][24] , \predict_PC[0][23] ,
         \predict_PC[0][22] , \predict_PC[0][21] , \predict_PC[0][20] ,
         \predict_PC[0][19] , \predict_PC[0][18] , \predict_PC[0][17] ,
         \predict_PC[0][16] , \predict_PC[0][15] , \predict_PC[0][14] ,
         \predict_PC[0][13] , \predict_PC[0][12] , \predict_PC[0][11] ,
         \predict_PC[0][10] , \predict_PC[0][9] , \predict_PC[0][8] ,
         \predict_PC[0][7] , \predict_PC[0][6] , \predict_PC[0][5] ,
         \predict_PC[0][4] , \predict_PC[0][3] , \predict_PC[0][2] ,
         \predict_PC[0][1] , \predict_PC[0][0] , \predict_PC[1][31] ,
         \predict_PC[1][30] , \predict_PC[1][29] , \predict_PC[1][28] ,
         \predict_PC[1][27] , \predict_PC[1][26] , \predict_PC[1][25] ,
         \predict_PC[1][24] , \predict_PC[1][23] , \predict_PC[1][22] ,
         \predict_PC[1][21] , \predict_PC[1][20] , \predict_PC[1][19] ,
         \predict_PC[1][18] , \predict_PC[1][17] , \predict_PC[1][16] ,
         \predict_PC[1][15] , \predict_PC[1][14] , \predict_PC[1][13] ,
         \predict_PC[1][12] , \predict_PC[1][11] , \predict_PC[1][10] ,
         \predict_PC[1][9] , \predict_PC[1][8] , \predict_PC[1][7] ,
         \predict_PC[1][6] , \predict_PC[1][5] , \predict_PC[1][4] ,
         \predict_PC[1][3] , \predict_PC[1][2] , \predict_PC[1][1] ,
         \predict_PC[1][0] , \predict_PC[2][31] , \predict_PC[2][30] ,
         \predict_PC[2][29] , \predict_PC[2][28] , \predict_PC[2][27] ,
         \predict_PC[2][26] , \predict_PC[2][25] , \predict_PC[2][24] ,
         \predict_PC[2][23] , \predict_PC[2][22] , \predict_PC[2][21] ,
         \predict_PC[2][20] , \predict_PC[2][19] , \predict_PC[2][18] ,
         \predict_PC[2][17] , \predict_PC[2][16] , \predict_PC[2][15] ,
         \predict_PC[2][14] , \predict_PC[2][13] , \predict_PC[2][12] ,
         \predict_PC[2][11] , \predict_PC[2][10] , \predict_PC[2][9] ,
         \predict_PC[2][8] , \predict_PC[2][7] , \predict_PC[2][6] ,
         \predict_PC[2][5] , \predict_PC[2][4] , \predict_PC[2][3] ,
         \predict_PC[2][2] , \predict_PC[2][1] , \predict_PC[2][0] ,
         \predict_PC[3][31] , \predict_PC[3][30] , \predict_PC[3][29] ,
         \predict_PC[3][28] , \predict_PC[3][27] , \predict_PC[3][26] ,
         \predict_PC[3][25] , \predict_PC[3][24] , \predict_PC[3][23] ,
         \predict_PC[3][22] , \predict_PC[3][21] , \predict_PC[3][20] ,
         \predict_PC[3][19] , \predict_PC[3][18] , \predict_PC[3][17] ,
         \predict_PC[3][16] , \predict_PC[3][15] , \predict_PC[3][14] ,
         \predict_PC[3][13] , \predict_PC[3][12] , \predict_PC[3][11] ,
         \predict_PC[3][10] , \predict_PC[3][9] , \predict_PC[3][8] ,
         \predict_PC[3][7] , \predict_PC[3][6] , \predict_PC[3][5] ,
         \predict_PC[3][4] , \predict_PC[3][3] , \predict_PC[3][2] ,
         \predict_PC[3][1] , \predict_PC[3][0] , \predict_PC[4][31] ,
         \predict_PC[4][30] , \predict_PC[4][29] , \predict_PC[4][28] ,
         \predict_PC[4][27] , \predict_PC[4][26] , \predict_PC[4][25] ,
         \predict_PC[4][24] , \predict_PC[4][23] , \predict_PC[4][22] ,
         \predict_PC[4][21] , \predict_PC[4][20] , \predict_PC[4][19] ,
         \predict_PC[4][18] , \predict_PC[4][17] , \predict_PC[4][16] ,
         \predict_PC[4][15] , \predict_PC[4][14] , \predict_PC[4][13] ,
         \predict_PC[4][12] , \predict_PC[4][11] , \predict_PC[4][10] ,
         \predict_PC[4][9] , \predict_PC[4][8] , \predict_PC[4][7] ,
         \predict_PC[4][6] , \predict_PC[4][5] , \predict_PC[4][4] ,
         \predict_PC[4][3] , \predict_PC[4][2] , \predict_PC[4][1] ,
         \predict_PC[4][0] , \predict_PC[5][31] , \predict_PC[5][30] ,
         \predict_PC[5][29] , \predict_PC[5][28] , \predict_PC[5][27] ,
         \predict_PC[5][26] , \predict_PC[5][25] , \predict_PC[5][24] ,
         \predict_PC[5][23] , \predict_PC[5][22] , \predict_PC[5][21] ,
         \predict_PC[5][20] , \predict_PC[5][19] , \predict_PC[5][18] ,
         \predict_PC[5][17] , \predict_PC[5][16] , \predict_PC[5][15] ,
         \predict_PC[5][14] , \predict_PC[5][13] , \predict_PC[5][12] ,
         \predict_PC[5][11] , \predict_PC[5][10] , \predict_PC[5][9] ,
         \predict_PC[5][8] , \predict_PC[5][7] , \predict_PC[5][6] ,
         \predict_PC[5][5] , \predict_PC[5][4] , \predict_PC[5][3] ,
         \predict_PC[5][2] , \predict_PC[5][1] , \predict_PC[5][0] ,
         \predict_PC[6][31] , \predict_PC[6][30] , \predict_PC[6][29] ,
         \predict_PC[6][28] , \predict_PC[6][27] , \predict_PC[6][26] ,
         \predict_PC[6][25] , \predict_PC[6][24] , \predict_PC[6][23] ,
         \predict_PC[6][22] , \predict_PC[6][21] , \predict_PC[6][20] ,
         \predict_PC[6][19] , \predict_PC[6][18] , \predict_PC[6][17] ,
         \predict_PC[6][16] , \predict_PC[6][15] , \predict_PC[6][14] ,
         \predict_PC[6][13] , \predict_PC[6][12] , \predict_PC[6][11] ,
         \predict_PC[6][10] , \predict_PC[6][9] , \predict_PC[6][8] ,
         \predict_PC[6][7] , \predict_PC[6][6] , \predict_PC[6][5] ,
         \predict_PC[6][4] , \predict_PC[6][3] , \predict_PC[6][2] ,
         \predict_PC[6][1] , \predict_PC[6][0] , \predict_PC[7][31] ,
         \predict_PC[7][30] , \predict_PC[7][29] , \predict_PC[7][28] ,
         \predict_PC[7][27] , \predict_PC[7][26] , \predict_PC[7][25] ,
         \predict_PC[7][24] , \predict_PC[7][23] , \predict_PC[7][22] ,
         \predict_PC[7][21] , \predict_PC[7][20] , \predict_PC[7][19] ,
         \predict_PC[7][18] , \predict_PC[7][17] , \predict_PC[7][16] ,
         \predict_PC[7][15] , \predict_PC[7][14] , \predict_PC[7][13] ,
         \predict_PC[7][12] , \predict_PC[7][11] , \predict_PC[7][10] ,
         \predict_PC[7][9] , \predict_PC[7][8] , \predict_PC[7][7] ,
         \predict_PC[7][6] , \predict_PC[7][5] , \predict_PC[7][4] ,
         \predict_PC[7][3] , \predict_PC[7][2] , \predict_PC[7][1] ,
         \predict_PC[7][0] , \predict_PC[8][31] , \predict_PC[8][30] ,
         \predict_PC[8][29] , \predict_PC[8][28] , \predict_PC[8][27] ,
         \predict_PC[8][26] , \predict_PC[8][25] , \predict_PC[8][24] ,
         \predict_PC[8][23] , \predict_PC[8][22] , \predict_PC[8][21] ,
         \predict_PC[8][20] , \predict_PC[8][19] , \predict_PC[8][18] ,
         \predict_PC[8][17] , \predict_PC[8][16] , \predict_PC[8][15] ,
         \predict_PC[8][14] , \predict_PC[8][13] , \predict_PC[8][12] ,
         \predict_PC[8][11] , \predict_PC[8][10] , \predict_PC[8][9] ,
         \predict_PC[8][8] , \predict_PC[8][7] , \predict_PC[8][6] ,
         \predict_PC[8][5] , \predict_PC[8][4] , \predict_PC[8][3] ,
         \predict_PC[8][2] , \predict_PC[8][1] , \predict_PC[8][0] ,
         \predict_PC[9][31] , \predict_PC[9][30] , \predict_PC[9][29] ,
         \predict_PC[9][28] , \predict_PC[9][27] , \predict_PC[9][26] ,
         \predict_PC[9][25] , \predict_PC[9][24] , \predict_PC[9][23] ,
         \predict_PC[9][22] , \predict_PC[9][21] , \predict_PC[9][20] ,
         \predict_PC[9][19] , \predict_PC[9][18] , \predict_PC[9][17] ,
         \predict_PC[9][16] , \predict_PC[9][15] , \predict_PC[9][14] ,
         \predict_PC[9][13] , \predict_PC[9][12] , \predict_PC[9][11] ,
         \predict_PC[9][10] , \predict_PC[9][9] , \predict_PC[9][8] ,
         \predict_PC[9][7] , \predict_PC[9][6] , \predict_PC[9][5] ,
         \predict_PC[9][4] , \predict_PC[9][3] , \predict_PC[9][2] ,
         \predict_PC[9][1] , \predict_PC[9][0] , \predict_PC[10][31] ,
         \predict_PC[10][30] , \predict_PC[10][29] , \predict_PC[10][28] ,
         \predict_PC[10][27] , \predict_PC[10][26] , \predict_PC[10][25] ,
         \predict_PC[10][24] , \predict_PC[10][23] , \predict_PC[10][22] ,
         \predict_PC[10][21] , \predict_PC[10][20] , \predict_PC[10][19] ,
         \predict_PC[10][18] , \predict_PC[10][17] , \predict_PC[10][16] ,
         \predict_PC[10][15] , \predict_PC[10][14] , \predict_PC[10][13] ,
         \predict_PC[10][12] , \predict_PC[10][11] , \predict_PC[10][10] ,
         \predict_PC[10][9] , \predict_PC[10][8] , \predict_PC[10][7] ,
         \predict_PC[10][6] , \predict_PC[10][5] , \predict_PC[10][4] ,
         \predict_PC[10][3] , \predict_PC[10][2] , \predict_PC[10][1] ,
         \predict_PC[10][0] , \predict_PC[11][31] , \predict_PC[11][30] ,
         \predict_PC[11][29] , \predict_PC[11][28] , \predict_PC[11][27] ,
         \predict_PC[11][26] , \predict_PC[11][25] , \predict_PC[11][24] ,
         \predict_PC[11][23] , \predict_PC[11][22] , \predict_PC[11][21] ,
         \predict_PC[11][20] , \predict_PC[11][19] , \predict_PC[11][18] ,
         \predict_PC[11][17] , \predict_PC[11][16] , \predict_PC[11][15] ,
         \predict_PC[11][14] , \predict_PC[11][13] , \predict_PC[11][12] ,
         \predict_PC[11][11] , \predict_PC[11][10] , \predict_PC[11][9] ,
         \predict_PC[11][8] , \predict_PC[11][7] , \predict_PC[11][6] ,
         \predict_PC[11][5] , \predict_PC[11][4] , \predict_PC[11][3] ,
         \predict_PC[11][2] , \predict_PC[11][1] , \predict_PC[11][0] ,
         \predict_PC[12][31] , \predict_PC[12][30] , \predict_PC[12][29] ,
         \predict_PC[12][28] , \predict_PC[12][27] , \predict_PC[12][26] ,
         \predict_PC[12][25] , \predict_PC[12][24] , \predict_PC[12][23] ,
         \predict_PC[12][22] , \predict_PC[12][21] , \predict_PC[12][20] ,
         \predict_PC[12][19] , \predict_PC[12][18] , \predict_PC[12][17] ,
         \predict_PC[12][16] , \predict_PC[12][15] , \predict_PC[12][14] ,
         \predict_PC[12][13] , \predict_PC[12][12] , \predict_PC[12][11] ,
         \predict_PC[12][10] , \predict_PC[12][9] , \predict_PC[12][8] ,
         \predict_PC[12][7] , \predict_PC[12][6] , \predict_PC[12][5] ,
         \predict_PC[12][4] , \predict_PC[12][3] , \predict_PC[12][2] ,
         \predict_PC[12][1] , \predict_PC[12][0] , \predict_PC[13][31] ,
         \predict_PC[13][30] , \predict_PC[13][29] , \predict_PC[13][28] ,
         \predict_PC[13][27] , \predict_PC[13][26] , \predict_PC[13][25] ,
         \predict_PC[13][24] , \predict_PC[13][23] , \predict_PC[13][22] ,
         \predict_PC[13][21] , \predict_PC[13][20] , \predict_PC[13][19] ,
         \predict_PC[13][18] , \predict_PC[13][17] , \predict_PC[13][16] ,
         \predict_PC[13][15] , \predict_PC[13][14] , \predict_PC[13][13] ,
         \predict_PC[13][12] , \predict_PC[13][11] , \predict_PC[13][10] ,
         \predict_PC[13][9] , \predict_PC[13][8] , \predict_PC[13][7] ,
         \predict_PC[13][6] , \predict_PC[13][5] , \predict_PC[13][4] ,
         \predict_PC[13][3] , \predict_PC[13][2] , \predict_PC[13][1] ,
         \predict_PC[13][0] , \predict_PC[14][31] , \predict_PC[14][30] ,
         \predict_PC[14][29] , \predict_PC[14][28] , \predict_PC[14][27] ,
         \predict_PC[14][26] , \predict_PC[14][25] , \predict_PC[14][24] ,
         \predict_PC[14][23] , \predict_PC[14][22] , \predict_PC[14][21] ,
         \predict_PC[14][20] , \predict_PC[14][19] , \predict_PC[14][18] ,
         \predict_PC[14][17] , \predict_PC[14][16] , \predict_PC[14][15] ,
         \predict_PC[14][14] , \predict_PC[14][13] , \predict_PC[14][12] ,
         \predict_PC[14][11] , \predict_PC[14][10] , \predict_PC[14][9] ,
         \predict_PC[14][8] , \predict_PC[14][7] , \predict_PC[14][6] ,
         \predict_PC[14][5] , \predict_PC[14][4] , \predict_PC[14][3] ,
         \predict_PC[14][2] , \predict_PC[14][1] , \predict_PC[14][0] ,
         \predict_PC[15][31] , \predict_PC[15][30] , \predict_PC[15][29] ,
         \predict_PC[15][28] , \predict_PC[15][27] , \predict_PC[15][26] ,
         \predict_PC[15][25] , \predict_PC[15][24] , \predict_PC[15][23] ,
         \predict_PC[15][22] , \predict_PC[15][21] , \predict_PC[15][20] ,
         \predict_PC[15][19] , \predict_PC[15][18] , \predict_PC[15][17] ,
         \predict_PC[15][16] , \predict_PC[15][15] , \predict_PC[15][14] ,
         \predict_PC[15][13] , \predict_PC[15][12] , \predict_PC[15][11] ,
         \predict_PC[15][10] , \predict_PC[15][9] , \predict_PC[15][8] ,
         \predict_PC[15][7] , \predict_PC[15][6] , \predict_PC[15][5] ,
         \predict_PC[15][4] , \predict_PC[15][3] , \predict_PC[15][2] ,
         \predict_PC[15][1] , \predict_PC[15][0] , n1535, n1536, n1537, n1538,
         n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548,
         n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558,
         n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568,
         n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578,
         n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588,
         n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598,
         n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608,
         n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618,
         n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628,
         n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638,
         n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648,
         n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658,
         n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668,
         n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678,
         n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688,
         n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698,
         n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708,
         n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718,
         n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728,
         n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738,
         n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748,
         n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758,
         n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768,
         n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778,
         n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788,
         n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798,
         n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808,
         n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818,
         n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828,
         n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838,
         n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848,
         n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858,
         n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868,
         n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878,
         n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888,
         n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898,
         n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908,
         n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918,
         n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928,
         n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938,
         n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948,
         n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958,
         n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968,
         n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978,
         n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988,
         n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998,
         n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008,
         n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018,
         n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028,
         n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038,
         n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048,
         n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058,
         n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068,
         n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078,
         n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088,
         n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098,
         n2099, n2100, n6, n7, n8, n9, n588, n589, n590, n591, n592, n593,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n696, n697, n699, n701, n703, n736, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
         n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
         n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
         n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
         n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
         n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
         n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
         n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
         n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
         n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
         n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
         n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
         n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
         n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
         n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
         n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
         n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
         n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
         n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
         n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
         n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
         n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
         n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
         n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
         n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
         n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
         n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
         n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
         n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
         n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
         n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
         n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
         n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
         n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
         n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
         n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380,
         n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390,
         n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400,
         n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410,
         n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420,
         n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430,
         n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440,
         n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450,
         n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460,
         n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470,
         n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480,
         n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490,
         n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500,
         n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510,
         n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520,
         n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530,
         n1531, n1532, n1533, n1534, n2101, n2102, n2103, n2104, n2105, n2106,
         n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116,
         n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126,
         n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136,
         n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146,
         n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156,
         n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166,
         n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176,
         n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186,
         n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196,
         n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206,
         n2207, n2208, n2209, n2210, n2221, n2222, n2224, n2225, n2252, n2251,
         n2250, n2249, n2248, n2247, n2246, n2245, n2244, n2243, n2242, n2241,
         n2240, n2239, n2238, n2237, n2236, n2235, n2234, n2233, n2232, n2231,
         n2230, n2229, n2228, n2227, n2226, n2223, n2220, n2219, n2218, n2217,
         n2212, n2211, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n694, n695, n698, n700, n702, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n737, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n2213, n2214, n2215, n2216, n2253, n2254,
         n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264,
         n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274,
         n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284,
         n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294,
         n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304,
         n2305, n2306, n2307, n2308, n2309, n2310, n2311;
  wire   [15:0] taken;
  wire   [15:0] write_enable;

  DFFR_X1 \last_TAG_reg[3]  ( .D(n2100), .CK(clock), .RN(n2288), .Q(n591), 
        .QN(n664) );
  DFFR_X1 \last_TAG_reg[2]  ( .D(n2099), .CK(clock), .RN(n2303), .Q(n590), 
        .QN(n661) );
  DFFR_X1 \last_TAG_reg[1]  ( .D(n2098), .CK(clock), .RN(n2291), .Q(n589), 
        .QN(n662) );
  DFFR_X1 \last_TAG_reg[0]  ( .D(n2097), .CK(clock), .RN(n2299), .Q(n588), 
        .QN(n660) );
  DFFR_X1 \write_enable_reg[15]  ( .D(n2096), .CK(clock), .RN(n2305), .Q(
        write_enable[15]), .QN(n713) );
  DFFR_X1 \write_enable_reg[14]  ( .D(n2095), .CK(clock), .RN(n2310), .Q(
        write_enable[14]), .QN(n712) );
  DFFR_X1 \write_enable_reg[13]  ( .D(n2094), .CK(clock), .RN(n2300), .Q(
        write_enable[13]), .QN(n711) );
  DFFR_X1 \write_enable_reg[12]  ( .D(n2093), .CK(clock), .RN(n2307), .Q(
        write_enable[12]), .QN(n710) );
  DFFR_X1 \write_enable_reg[11]  ( .D(n2092), .CK(clock), .RN(n2309), .Q(
        write_enable[11]), .QN(n709) );
  DFFR_X1 \write_enable_reg[10]  ( .D(n2091), .CK(clock), .RN(n2310), .Q(
        write_enable[10]), .QN(n708) );
  DFFR_X1 \write_enable_reg[9]  ( .D(n2090), .CK(clock), .RN(n2296), .Q(
        write_enable[9]), .QN(n707) );
  DFFR_X1 \write_enable_reg[8]  ( .D(n2089), .CK(clock), .RN(n2290), .Q(
        write_enable[8]), .QN(n706) );
  DFFR_X1 \write_enable_reg[7]  ( .D(n2088), .CK(clock), .RN(n2309), .Q(
        write_enable[7]), .QN(n705) );
  DFFR_X1 \write_enable_reg[6]  ( .D(n2087), .CK(clock), .RN(n2310), .Q(
        write_enable[6]), .QN(n704) );
  DFFR_X1 \write_enable_reg[5]  ( .D(n2086), .CK(clock), .RN(n2296), .Q(
        write_enable[5]), .QN(n702) );
  DFFR_X1 \write_enable_reg[4]  ( .D(n2085), .CK(clock), .RN(n2299), .Q(
        write_enable[4]), .QN(n700) );
  DFFR_X1 \write_enable_reg[3]  ( .D(n2084), .CK(clock), .RN(n2305), .Q(
        write_enable[3]), .QN(n698) );
  DFFR_X1 \write_enable_reg[2]  ( .D(n2083), .CK(clock), .RN(n2302), .Q(
        write_enable[2]), .QN(n695) );
  DFFR_X1 \write_enable_reg[1]  ( .D(n2082), .CK(clock), .RN(n2307), .Q(
        write_enable[1]), .QN(n694) );
  DFFR_X1 \write_enable_reg[0]  ( .D(n2081), .CK(clock), .RN(n2289), .Q(
        write_enable[0]), .QN(n665) );
  DFF_X1 last_taken_reg ( .D(n2080), .CK(clock), .Q(n663) );
  DFFR_X1 \predict_PC_reg[0][31]  ( .D(n2079), .CK(clock), .RN(n2308), .Q(
        \predict_PC[0][31] ) );
  DFFR_X1 \predict_PC_reg[0][30]  ( .D(n2078), .CK(clock), .RN(n2298), .Q(
        \predict_PC[0][30] ) );
  DFFR_X1 \predict_PC_reg[0][29]  ( .D(n2077), .CK(clock), .RN(n2303), .Q(
        \predict_PC[0][29] ) );
  DFFR_X1 \predict_PC_reg[0][28]  ( .D(n2076), .CK(clock), .RN(n2308), .Q(
        \predict_PC[0][28] ) );
  DFFR_X1 \predict_PC_reg[0][27]  ( .D(n2075), .CK(clock), .RN(n2302), .Q(
        \predict_PC[0][27] ) );
  DFFR_X1 \predict_PC_reg[0][26]  ( .D(n2074), .CK(clock), .RN(n2301), .Q(
        \predict_PC[0][26] ) );
  DFFR_X1 \predict_PC_reg[0][25]  ( .D(n2073), .CK(clock), .RN(n2309), .Q(
        \predict_PC[0][25] ) );
  DFFR_X1 \predict_PC_reg[0][24]  ( .D(n2072), .CK(clock), .RN(n2308), .Q(
        \predict_PC[0][24] ) );
  DFFR_X1 \predict_PC_reg[0][23]  ( .D(n2071), .CK(clock), .RN(n2308), .Q(
        \predict_PC[0][23] ) );
  DFFR_X1 \predict_PC_reg[0][22]  ( .D(n2070), .CK(clock), .RN(n2292), .Q(
        \predict_PC[0][22] ) );
  DFFR_X1 \predict_PC_reg[0][21]  ( .D(n2069), .CK(clock), .RN(n2292), .Q(
        \predict_PC[0][21] ) );
  DFFR_X1 \predict_PC_reg[0][20]  ( .D(n2068), .CK(clock), .RN(n2292), .Q(
        \predict_PC[0][20] ) );
  DFFR_X1 \predict_PC_reg[0][19]  ( .D(n2067), .CK(clock), .RN(n2292), .Q(
        \predict_PC[0][19] ) );
  DFFR_X1 \predict_PC_reg[0][18]  ( .D(n2066), .CK(clock), .RN(n2307), .Q(
        \predict_PC[0][18] ) );
  DFFR_X1 \predict_PC_reg[0][17]  ( .D(n2065), .CK(clock), .RN(n2292), .Q(
        \predict_PC[0][17] ) );
  DFFR_X1 \predict_PC_reg[0][16]  ( .D(n2064), .CK(clock), .RN(n2292), .Q(
        \predict_PC[0][16] ) );
  DFFR_X1 \predict_PC_reg[0][15]  ( .D(n2063), .CK(clock), .RN(n2292), .Q(
        \predict_PC[0][15] ) );
  DFFR_X1 \predict_PC_reg[0][14]  ( .D(n2062), .CK(clock), .RN(n2292), .Q(
        \predict_PC[0][14] ) );
  DFFR_X1 \predict_PC_reg[0][13]  ( .D(n2061), .CK(clock), .RN(n2292), .Q(
        \predict_PC[0][13] ) );
  DFFR_X1 \predict_PC_reg[0][12]  ( .D(n2060), .CK(clock), .RN(n2292), .Q(
        \predict_PC[0][12] ) );
  DFFR_X1 \predict_PC_reg[0][11]  ( .D(n2059), .CK(clock), .RN(n2292), .Q(
        \predict_PC[0][11] ) );
  DFFR_X1 \predict_PC_reg[0][10]  ( .D(n2058), .CK(clock), .RN(n2298), .Q(
        \predict_PC[0][10] ) );
  DFFR_X1 \predict_PC_reg[0][9]  ( .D(n2057), .CK(clock), .RN(n2297), .Q(
        \predict_PC[0][9] ) );
  DFFR_X1 \predict_PC_reg[0][8]  ( .D(n2056), .CK(clock), .RN(n2301), .Q(
        \predict_PC[0][8] ) );
  DFFR_X1 \predict_PC_reg[0][7]  ( .D(n2055), .CK(clock), .RN(n2303), .Q(
        \predict_PC[0][7] ) );
  DFFR_X1 \predict_PC_reg[0][6]  ( .D(n2054), .CK(clock), .RN(n2294), .Q(
        \predict_PC[0][6] ) );
  DFFR_X1 \predict_PC_reg[0][5]  ( .D(n2053), .CK(clock), .RN(n2306), .Q(
        \predict_PC[0][5] ) );
  DFFR_X1 \predict_PC_reg[0][4]  ( .D(n2052), .CK(clock), .RN(n2300), .Q(
        \predict_PC[0][4] ) );
  DFFR_X1 \predict_PC_reg[0][3]  ( .D(n2051), .CK(clock), .RN(n2308), .Q(
        \predict_PC[0][3] ) );
  DFFR_X1 \predict_PC_reg[0][2]  ( .D(n2050), .CK(clock), .RN(n2295), .Q(
        \predict_PC[0][2] ) );
  DFFR_X1 \predict_PC_reg[0][1]  ( .D(n2049), .CK(clock), .RN(n2295), .Q(
        \predict_PC[0][1] ) );
  DFFR_X1 \predict_PC_reg[0][0]  ( .D(n2048), .CK(clock), .RN(n2306), .Q(
        \predict_PC[0][0] ) );
  DFFR_X1 \predict_PC_reg[1][31]  ( .D(n2047), .CK(clock), .RN(n2307), .Q(
        \predict_PC[1][31] ) );
  DFFR_X1 \predict_PC_reg[1][30]  ( .D(n2046), .CK(clock), .RN(n2298), .Q(
        \predict_PC[1][30] ) );
  DFFR_X1 \predict_PC_reg[1][29]  ( .D(n2045), .CK(clock), .RN(n2303), .Q(
        \predict_PC[1][29] ) );
  DFFR_X1 \predict_PC_reg[1][28]  ( .D(n2044), .CK(clock), .RN(n2307), .Q(
        \predict_PC[1][28] ) );
  DFFR_X1 \predict_PC_reg[1][27]  ( .D(n2043), .CK(clock), .RN(n2302), .Q(
        \predict_PC[1][27] ) );
  DFFR_X1 \predict_PC_reg[1][26]  ( .D(n2042), .CK(clock), .RN(n2301), .Q(
        \predict_PC[1][26] ) );
  DFFR_X1 \predict_PC_reg[1][25]  ( .D(n2041), .CK(clock), .RN(n2299), .Q(
        \predict_PC[1][25] ) );
  DFFR_X1 \predict_PC_reg[1][24]  ( .D(n2040), .CK(clock), .RN(n2310), .Q(
        \predict_PC[1][24] ) );
  DFFR_X1 \predict_PC_reg[1][23]  ( .D(n2039), .CK(clock), .RN(n2302), .Q(
        \predict_PC[1][23] ) );
  DFFR_X1 \predict_PC_reg[1][22]  ( .D(n2038), .CK(clock), .RN(n2301), .Q(
        \predict_PC[1][22] ) );
  DFFR_X1 \predict_PC_reg[1][21]  ( .D(n2037), .CK(clock), .RN(n2303), .Q(
        \predict_PC[1][21] ) );
  DFFR_X1 \predict_PC_reg[1][20]  ( .D(n2036), .CK(clock), .RN(n2294), .Q(
        \predict_PC[1][20] ) );
  DFFR_X1 \predict_PC_reg[1][19]  ( .D(n2035), .CK(clock), .RN(n2298), .Q(
        \predict_PC[1][19] ) );
  DFFR_X1 \predict_PC_reg[1][18]  ( .D(n2034), .CK(clock), .RN(n2300), .Q(
        \predict_PC[1][18] ) );
  DFFR_X1 \predict_PC_reg[1][17]  ( .D(n2033), .CK(clock), .RN(n2308), .Q(
        \predict_PC[1][17] ) );
  DFFR_X1 \predict_PC_reg[1][16]  ( .D(n2032), .CK(clock), .RN(n2294), .Q(
        \predict_PC[1][16] ) );
  DFFR_X1 \predict_PC_reg[1][15]  ( .D(n2031), .CK(clock), .RN(n2294), .Q(
        \predict_PC[1][15] ) );
  DFFR_X1 \predict_PC_reg[1][14]  ( .D(n2030), .CK(clock), .RN(n2294), .Q(
        \predict_PC[1][14] ) );
  DFFR_X1 \predict_PC_reg[1][13]  ( .D(n2029), .CK(clock), .RN(n2294), .Q(
        \predict_PC[1][13] ) );
  DFFR_X1 \predict_PC_reg[1][12]  ( .D(n2028), .CK(clock), .RN(n2294), .Q(
        \predict_PC[1][12] ) );
  DFFR_X1 \predict_PC_reg[1][11]  ( .D(n2027), .CK(clock), .RN(n2294), .Q(
        \predict_PC[1][11] ) );
  DFFR_X1 \predict_PC_reg[1][10]  ( .D(n2026), .CK(clock), .RN(n2294), .Q(
        \predict_PC[1][10] ) );
  DFFR_X1 \predict_PC_reg[1][9]  ( .D(n2025), .CK(clock), .RN(n2304), .Q(
        \predict_PC[1][9] ) );
  DFFR_X1 \predict_PC_reg[1][8]  ( .D(n2024), .CK(clock), .RN(n2294), .Q(
        \predict_PC[1][8] ) );
  DFFR_X1 \predict_PC_reg[1][7]  ( .D(n2023), .CK(clock), .RN(n2294), .Q(
        \predict_PC[1][7] ) );
  DFFR_X1 \predict_PC_reg[1][6]  ( .D(n2022), .CK(clock), .RN(n2297), .Q(
        \predict_PC[1][6] ) );
  DFFR_X1 \predict_PC_reg[1][5]  ( .D(n2021), .CK(clock), .RN(n2306), .Q(
        \predict_PC[1][5] ) );
  DFFR_X1 \predict_PC_reg[1][4]  ( .D(n2020), .CK(clock), .RN(n2306), .Q(
        \predict_PC[1][4] ) );
  DFFR_X1 \predict_PC_reg[1][3]  ( .D(n2019), .CK(clock), .RN(n2306), .Q(
        \predict_PC[1][3] ) );
  DFFR_X1 \predict_PC_reg[1][2]  ( .D(n2018), .CK(clock), .RN(n2307), .Q(
        \predict_PC[1][2] ) );
  DFFR_X1 \predict_PC_reg[1][1]  ( .D(n2017), .CK(clock), .RN(n2295), .Q(
        \predict_PC[1][1] ) );
  DFFR_X1 \predict_PC_reg[1][0]  ( .D(n2016), .CK(clock), .RN(n2307), .Q(
        \predict_PC[1][0] ) );
  DFFR_X1 \predict_PC_reg[2][31]  ( .D(n2015), .CK(clock), .RN(n2302), .Q(
        \predict_PC[2][31] ) );
  DFFR_X1 \predict_PC_reg[2][30]  ( .D(n2014), .CK(clock), .RN(n2303), .Q(
        \predict_PC[2][30] ) );
  DFFR_X1 \predict_PC_reg[2][29]  ( .D(n2013), .CK(clock), .RN(n2302), .Q(
        \predict_PC[2][29] ) );
  DFFR_X1 \predict_PC_reg[2][28]  ( .D(n2012), .CK(clock), .RN(n2302), .Q(
        \predict_PC[2][28] ) );
  DFFR_X1 \predict_PC_reg[2][27]  ( .D(n2011), .CK(clock), .RN(n2302), .Q(
        \predict_PC[2][27] ) );
  DFFR_X1 \predict_PC_reg[2][26]  ( .D(n2010), .CK(clock), .RN(n2289), .Q(
        \predict_PC[2][26] ) );
  DFFR_X1 \predict_PC_reg[2][25]  ( .D(n2009), .CK(clock), .RN(n2299), .Q(
        \predict_PC[2][25] ) );
  DFFR_X1 \predict_PC_reg[2][24]  ( .D(n2008), .CK(clock), .RN(n2289), .Q(
        \predict_PC[2][24] ) );
  DFFR_X1 \predict_PC_reg[2][23]  ( .D(n2007), .CK(clock), .RN(n2288), .Q(
        \predict_PC[2][23] ) );
  DFFR_X1 \predict_PC_reg[2][22]  ( .D(n2006), .CK(clock), .RN(n2288), .Q(
        \predict_PC[2][22] ) );
  DFFR_X1 \predict_PC_reg[2][21]  ( .D(n2005), .CK(clock), .RN(n2311), .Q(
        \predict_PC[2][21] ) );
  DFFR_X1 \predict_PC_reg[2][20]  ( .D(n2004), .CK(clock), .RN(n2288), .Q(
        \predict_PC[2][20] ) );
  DFFR_X1 \predict_PC_reg[2][19]  ( .D(n2003), .CK(clock), .RN(n2311), .Q(
        \predict_PC[2][19] ) );
  DFFR_X1 \predict_PC_reg[2][18]  ( .D(n2002), .CK(clock), .RN(n2298), .Q(
        \predict_PC[2][18] ) );
  DFFR_X1 \predict_PC_reg[2][17]  ( .D(n2001), .CK(clock), .RN(n2301), .Q(
        \predict_PC[2][17] ) );
  DFFR_X1 \predict_PC_reg[2][16]  ( .D(n2000), .CK(clock), .RN(n2288), .Q(
        \predict_PC[2][16] ) );
  DFFR_X1 \predict_PC_reg[2][15]  ( .D(n1999), .CK(clock), .RN(n2310), .Q(
        \predict_PC[2][15] ) );
  DFFR_X1 \predict_PC_reg[2][14]  ( .D(n1998), .CK(clock), .RN(n2289), .Q(
        \predict_PC[2][14] ) );
  DFFR_X1 \predict_PC_reg[2][13]  ( .D(n1997), .CK(clock), .RN(n2310), .Q(
        \predict_PC[2][13] ) );
  DFFR_X1 \predict_PC_reg[2][12]  ( .D(n1996), .CK(clock), .RN(n2311), .Q(
        \predict_PC[2][12] ) );
  DFFR_X1 \predict_PC_reg[2][11]  ( .D(n1995), .CK(clock), .RN(n2311), .Q(
        \predict_PC[2][11] ) );
  DFFR_X1 \predict_PC_reg[2][10]  ( .D(n1994), .CK(clock), .RN(n2311), .Q(
        \predict_PC[2][10] ) );
  DFFR_X1 \predict_PC_reg[2][9]  ( .D(n1993), .CK(clock), .RN(n2304), .Q(
        \predict_PC[2][9] ) );
  DFFR_X1 \predict_PC_reg[2][8]  ( .D(n1992), .CK(clock), .RN(n2311), .Q(
        \predict_PC[2][8] ) );
  DFFR_X1 \predict_PC_reg[2][7]  ( .D(n1991), .CK(clock), .RN(n2289), .Q(
        \predict_PC[2][7] ) );
  DFFR_X1 \predict_PC_reg[2][6]  ( .D(n1990), .CK(clock), .RN(n2295), .Q(
        \predict_PC[2][6] ) );
  DFFR_X1 \predict_PC_reg[2][5]  ( .D(n1989), .CK(clock), .RN(n2306), .Q(
        \predict_PC[2][5] ) );
  DFFR_X1 \predict_PC_reg[2][4]  ( .D(n1988), .CK(clock), .RN(n2311), .Q(
        \predict_PC[2][4] ) );
  DFFR_X1 \predict_PC_reg[2][3]  ( .D(n1987), .CK(clock), .RN(n2311), .Q(
        \predict_PC[2][3] ) );
  DFFR_X1 \predict_PC_reg[2][2]  ( .D(n1986), .CK(clock), .RN(n2300), .Q(
        \predict_PC[2][2] ) );
  DFFR_X1 \predict_PC_reg[2][1]  ( .D(n1985), .CK(clock), .RN(n2295), .Q(
        \predict_PC[2][1] ) );
  DFFR_X1 \predict_PC_reg[2][0]  ( .D(n1984), .CK(clock), .RN(n2311), .Q(
        \predict_PC[2][0] ) );
  DFFR_X1 \predict_PC_reg[3][31]  ( .D(n1983), .CK(clock), .RN(n2309), .Q(
        \predict_PC[3][31] ) );
  DFFR_X1 \predict_PC_reg[3][30]  ( .D(n1982), .CK(clock), .RN(n2303), .Q(
        \predict_PC[3][30] ) );
  DFFR_X1 \predict_PC_reg[3][29]  ( .D(n1981), .CK(clock), .RN(n2302), .Q(
        \predict_PC[3][29] ) );
  DFFR_X1 \predict_PC_reg[3][28]  ( .D(n1980), .CK(clock), .RN(n2297), .Q(
        \predict_PC[3][28] ) );
  DFFR_X1 \predict_PC_reg[3][27]  ( .D(n1979), .CK(clock), .RN(n2302), .Q(
        \predict_PC[3][27] ) );
  DFFR_X1 \predict_PC_reg[3][26]  ( .D(n1978), .CK(clock), .RN(n2299), .Q(
        \predict_PC[3][26] ) );
  DFFR_X1 \predict_PC_reg[3][25]  ( .D(n1977), .CK(clock), .RN(n2299), .Q(
        \predict_PC[3][25] ) );
  DFFR_X1 \predict_PC_reg[3][24]  ( .D(n1976), .CK(clock), .RN(n2299), .Q(
        \predict_PC[3][24] ) );
  DFFR_X1 \predict_PC_reg[3][23]  ( .D(n1975), .CK(clock), .RN(n2306), .Q(
        \predict_PC[3][23] ) );
  DFFR_X1 \predict_PC_reg[3][22]  ( .D(n1974), .CK(clock), .RN(n2295), .Q(
        \predict_PC[3][22] ) );
  DFFR_X1 \predict_PC_reg[3][21]  ( .D(n1973), .CK(clock), .RN(n2308), .Q(
        \predict_PC[3][21] ) );
  DFFR_X1 \predict_PC_reg[3][20]  ( .D(n1972), .CK(clock), .RN(n2295), .Q(
        \predict_PC[3][20] ) );
  DFFR_X1 \predict_PC_reg[3][19]  ( .D(n1971), .CK(clock), .RN(n2291), .Q(
        \predict_PC[3][19] ) );
  DFFR_X1 \predict_PC_reg[3][18]  ( .D(n1970), .CK(clock), .RN(n2300), .Q(
        \predict_PC[3][18] ) );
  DFFR_X1 \predict_PC_reg[3][17]  ( .D(n1969), .CK(clock), .RN(n2290), .Q(
        \predict_PC[3][17] ) );
  DFFR_X1 \predict_PC_reg[3][16]  ( .D(n1968), .CK(clock), .RN(n2290), .Q(
        \predict_PC[3][16] ) );
  DFFR_X1 \predict_PC_reg[3][15]  ( .D(n1967), .CK(clock), .RN(n2290), .Q(
        \predict_PC[3][15] ) );
  DFFR_X1 \predict_PC_reg[3][14]  ( .D(n1966), .CK(clock), .RN(n2290), .Q(
        \predict_PC[3][14] ) );
  DFFR_X1 \predict_PC_reg[3][13]  ( .D(n1965), .CK(clock), .RN(n2290), .Q(
        \predict_PC[3][13] ) );
  DFFR_X1 \predict_PC_reg[3][12]  ( .D(n1964), .CK(clock), .RN(n2290), .Q(
        \predict_PC[3][12] ) );
  DFFR_X1 \predict_PC_reg[3][11]  ( .D(n1963), .CK(clock), .RN(n2290), .Q(
        \predict_PC[3][11] ) );
  DFFR_X1 \predict_PC_reg[3][10]  ( .D(n1962), .CK(clock), .RN(n2290), .Q(
        \predict_PC[3][10] ) );
  DFFR_X1 \predict_PC_reg[3][9]  ( .D(n1961), .CK(clock), .RN(n2304), .Q(
        \predict_PC[3][9] ) );
  DFFR_X1 \predict_PC_reg[3][8]  ( .D(n1960), .CK(clock), .RN(n2290), .Q(
        \predict_PC[3][8] ) );
  DFFR_X1 \predict_PC_reg[3][7]  ( .D(n1959), .CK(clock), .RN(n2309), .Q(
        \predict_PC[3][7] ) );
  DFFR_X1 \predict_PC_reg[3][6]  ( .D(n1958), .CK(clock), .RN(n2309), .Q(
        \predict_PC[3][6] ) );
  DFFR_X1 \predict_PC_reg[3][5]  ( .D(n1957), .CK(clock), .RN(n2306), .Q(
        \predict_PC[3][5] ) );
  DFFR_X1 \predict_PC_reg[3][4]  ( .D(n1956), .CK(clock), .RN(n2309), .Q(
        \predict_PC[3][4] ) );
  DFFR_X1 \predict_PC_reg[3][3]  ( .D(n1955), .CK(clock), .RN(n2309), .Q(
        \predict_PC[3][3] ) );
  DFFR_X1 \predict_PC_reg[3][2]  ( .D(n1954), .CK(clock), .RN(n2309), .Q(
        \predict_PC[3][2] ) );
  DFFR_X1 \predict_PC_reg[3][1]  ( .D(n1953), .CK(clock), .RN(n2295), .Q(
        \predict_PC[3][1] ) );
  DFFR_X1 \predict_PC_reg[3][0]  ( .D(n1952), .CK(clock), .RN(n2309), .Q(
        \predict_PC[3][0] ) );
  DFFR_X1 \predict_PC_reg[4][31]  ( .D(n1951), .CK(clock), .RN(n2297), .Q(
        \predict_PC[4][31] ) );
  DFFR_X1 \predict_PC_reg[4][30]  ( .D(n1950), .CK(clock), .RN(n2303), .Q(
        \predict_PC[4][30] ) );
  DFFR_X1 \predict_PC_reg[4][29]  ( .D(n1949), .CK(clock), .RN(n2302), .Q(
        \predict_PC[4][29] ) );
  DFFR_X1 \predict_PC_reg[4][28]  ( .D(n1948), .CK(clock), .RN(n2309), .Q(
        \predict_PC[4][28] ) );
  DFFR_X1 \predict_PC_reg[4][27]  ( .D(n1947), .CK(clock), .RN(n2302), .Q(
        \predict_PC[4][27] ) );
  DFFR_X1 \predict_PC_reg[4][26]  ( .D(n1946), .CK(clock), .RN(n2299), .Q(
        \predict_PC[4][26] ) );
  DFFR_X1 \predict_PC_reg[4][25]  ( .D(n1945), .CK(clock), .RN(n2300), .Q(
        \predict_PC[4][25] ) );
  DFFR_X1 \predict_PC_reg[4][24]  ( .D(n1944), .CK(clock), .RN(n2302), .Q(
        \predict_PC[4][24] ) );
  DFFR_X1 \predict_PC_reg[4][23]  ( .D(n1943), .CK(clock), .RN(n2293), .Q(
        \predict_PC[4][23] ) );
  DFFR_X1 \predict_PC_reg[4][22]  ( .D(n1942), .CK(clock), .RN(n2293), .Q(
        \predict_PC[4][22] ) );
  DFFR_X1 \predict_PC_reg[4][21]  ( .D(n1941), .CK(clock), .RN(n2293), .Q(
        \predict_PC[4][21] ) );
  DFFR_X1 \predict_PC_reg[4][20]  ( .D(n1940), .CK(clock), .RN(n2293), .Q(
        \predict_PC[4][20] ) );
  DFFR_X1 \predict_PC_reg[4][19]  ( .D(n1939), .CK(clock), .RN(n2293), .Q(
        \predict_PC[4][19] ) );
  DFFR_X1 \predict_PC_reg[4][18]  ( .D(n1938), .CK(clock), .RN(n2290), .Q(
        \predict_PC[4][18] ) );
  DFFR_X1 \predict_PC_reg[4][17]  ( .D(n1937), .CK(clock), .RN(n2293), .Q(
        \predict_PC[4][17] ) );
  DFFR_X1 \predict_PC_reg[4][16]  ( .D(n1936), .CK(clock), .RN(n2293), .Q(
        \predict_PC[4][16] ) );
  DFFR_X1 \predict_PC_reg[4][15]  ( .D(n1935), .CK(clock), .RN(n2293), .Q(
        \predict_PC[4][15] ) );
  DFFR_X1 \predict_PC_reg[4][14]  ( .D(n1934), .CK(clock), .RN(n2293), .Q(
        \predict_PC[4][14] ) );
  DFFR_X1 \predict_PC_reg[4][13]  ( .D(n1933), .CK(clock), .RN(n2293), .Q(
        \predict_PC[4][13] ) );
  DFFR_X1 \predict_PC_reg[4][12]  ( .D(n1932), .CK(clock), .RN(n2293), .Q(
        \predict_PC[4][12] ) );
  DFFR_X1 \predict_PC_reg[4][11]  ( .D(n1931), .CK(clock), .RN(n2292), .Q(
        \predict_PC[4][11] ) );
  DFFR_X1 \predict_PC_reg[4][10]  ( .D(n1930), .CK(clock), .RN(n2304), .Q(
        \predict_PC[4][10] ) );
  DFFR_X1 \predict_PC_reg[4][9]  ( .D(n1929), .CK(clock), .RN(n2304), .Q(
        \predict_PC[4][9] ) );
  DFFR_X1 \predict_PC_reg[4][8]  ( .D(n1928), .CK(clock), .RN(n2307), .Q(
        \predict_PC[4][8] ) );
  DFFR_X1 \predict_PC_reg[4][7]  ( .D(n1927), .CK(clock), .RN(n2302), .Q(
        \predict_PC[4][7] ) );
  DFFR_X1 \predict_PC_reg[4][6]  ( .D(n1926), .CK(clock), .RN(n2290), .Q(
        \predict_PC[4][6] ) );
  DFFR_X1 \predict_PC_reg[4][5]  ( .D(n1925), .CK(clock), .RN(n2306), .Q(
        \predict_PC[4][5] ) );
  DFFR_X1 \predict_PC_reg[4][4]  ( .D(n1924), .CK(clock), .RN(n2293), .Q(
        \predict_PC[4][4] ) );
  DFFR_X1 \predict_PC_reg[4][3]  ( .D(n1923), .CK(clock), .RN(n2291), .Q(
        \predict_PC[4][3] ) );
  DFFR_X1 \predict_PC_reg[4][2]  ( .D(n1922), .CK(clock), .RN(n2311), .Q(
        \predict_PC[4][2] ) );
  DFFR_X1 \predict_PC_reg[4][1]  ( .D(n1921), .CK(clock), .RN(n2307), .Q(
        \predict_PC[4][1] ) );
  DFFR_X1 \predict_PC_reg[4][0]  ( .D(n1920), .CK(clock), .RN(n2292), .Q(
        \predict_PC[4][0] ) );
  DFFR_X1 \predict_PC_reg[5][31]  ( .D(n1919), .CK(clock), .RN(n2296), .Q(
        \predict_PC[5][31] ) );
  DFFR_X1 \predict_PC_reg[5][30]  ( .D(n1918), .CK(clock), .RN(n2303), .Q(
        \predict_PC[5][30] ) );
  DFFR_X1 \predict_PC_reg[5][29]  ( .D(n1917), .CK(clock), .RN(n2302), .Q(
        \predict_PC[5][29] ) );
  DFFR_X1 \predict_PC_reg[5][28]  ( .D(n1916), .CK(clock), .RN(n2296), .Q(
        \predict_PC[5][28] ) );
  DFFR_X1 \predict_PC_reg[5][27]  ( .D(n1915), .CK(clock), .RN(n2298), .Q(
        \predict_PC[5][27] ) );
  DFFR_X1 \predict_PC_reg[5][26]  ( .D(n1914), .CK(clock), .RN(n2299), .Q(
        \predict_PC[5][26] ) );
  DFFR_X1 \predict_PC_reg[5][25]  ( .D(n1913), .CK(clock), .RN(n2300), .Q(
        \predict_PC[5][25] ) );
  DFFR_X1 \predict_PC_reg[5][24]  ( .D(n1912), .CK(clock), .RN(n2296), .Q(
        \predict_PC[5][24] ) );
  DFFR_X1 \predict_PC_reg[5][23]  ( .D(n1911), .CK(clock), .RN(n2296), .Q(
        \predict_PC[5][23] ) );
  DFFR_X1 \predict_PC_reg[5][22]  ( .D(n1910), .CK(clock), .RN(n2296), .Q(
        \predict_PC[5][22] ) );
  DFFR_X1 \predict_PC_reg[5][21]  ( .D(n1909), .CK(clock), .RN(n2296), .Q(
        \predict_PC[5][21] ) );
  DFFR_X1 \predict_PC_reg[5][20]  ( .D(n1908), .CK(clock), .RN(n2295), .Q(
        \predict_PC[5][20] ) );
  DFFR_X1 \predict_PC_reg[5][19]  ( .D(n1907), .CK(clock), .RN(n2295), .Q(
        \predict_PC[5][19] ) );
  DFFR_X1 \predict_PC_reg[5][18]  ( .D(n1906), .CK(clock), .RN(n2288), .Q(
        \predict_PC[5][18] ) );
  DFFR_X1 \predict_PC_reg[5][17]  ( .D(n1905), .CK(clock), .RN(n2295), .Q(
        \predict_PC[5][17] ) );
  DFFR_X1 \predict_PC_reg[5][16]  ( .D(n1904), .CK(clock), .RN(n2295), .Q(
        \predict_PC[5][16] ) );
  DFFR_X1 \predict_PC_reg[5][15]  ( .D(n1903), .CK(clock), .RN(n2305), .Q(
        \predict_PC[5][15] ) );
  DFFR_X1 \predict_PC_reg[5][14]  ( .D(n1902), .CK(clock), .RN(n2305), .Q(
        \predict_PC[5][14] ) );
  DFFR_X1 \predict_PC_reg[5][13]  ( .D(n1901), .CK(clock), .RN(n2305), .Q(
        \predict_PC[5][13] ) );
  DFFR_X1 \predict_PC_reg[5][12]  ( .D(n1900), .CK(clock), .RN(n2306), .Q(
        \predict_PC[5][12] ) );
  DFFR_X1 \predict_PC_reg[5][11]  ( .D(n1899), .CK(clock), .RN(n2306), .Q(
        \predict_PC[5][11] ) );
  DFFR_X1 \predict_PC_reg[5][10]  ( .D(n1898), .CK(clock), .RN(n2306), .Q(
        \predict_PC[5][10] ) );
  DFFR_X1 \predict_PC_reg[5][9]  ( .D(n1897), .CK(clock), .RN(n2304), .Q(
        \predict_PC[5][9] ) );
  DFFR_X1 \predict_PC_reg[5][8]  ( .D(n1896), .CK(clock), .RN(n2306), .Q(
        \predict_PC[5][8] ) );
  DFFR_X1 \predict_PC_reg[5][7]  ( .D(n1895), .CK(clock), .RN(n2306), .Q(
        \predict_PC[5][7] ) );
  DFFR_X1 \predict_PC_reg[5][6]  ( .D(n1894), .CK(clock), .RN(n2306), .Q(
        \predict_PC[5][6] ) );
  DFFR_X1 \predict_PC_reg[5][5]  ( .D(n1893), .CK(clock), .RN(n2306), .Q(
        \predict_PC[5][5] ) );
  DFFR_X1 \predict_PC_reg[5][4]  ( .D(n1892), .CK(clock), .RN(n2306), .Q(
        \predict_PC[5][4] ) );
  DFFR_X1 \predict_PC_reg[5][3]  ( .D(n1891), .CK(clock), .RN(n2306), .Q(
        \predict_PC[5][3] ) );
  DFFR_X1 \predict_PC_reg[5][2]  ( .D(n1890), .CK(clock), .RN(n2306), .Q(
        \predict_PC[5][2] ) );
  DFFR_X1 \predict_PC_reg[5][1]  ( .D(n1889), .CK(clock), .RN(n2307), .Q(
        \predict_PC[5][1] ) );
  DFFR_X1 \predict_PC_reg[5][0]  ( .D(n1888), .CK(clock), .RN(n2296), .Q(
        \predict_PC[5][0] ) );
  DFFR_X1 \predict_PC_reg[6][31]  ( .D(n1887), .CK(clock), .RN(n2310), .Q(
        \predict_PC[6][31] ) );
  DFFR_X1 \predict_PC_reg[6][30]  ( .D(n1886), .CK(clock), .RN(n2303), .Q(
        \predict_PC[6][30] ) );
  DFFR_X1 \predict_PC_reg[6][29]  ( .D(n1885), .CK(clock), .RN(n2302), .Q(
        \predict_PC[6][29] ) );
  DFFR_X1 \predict_PC_reg[6][28]  ( .D(n1884), .CK(clock), .RN(n2310), .Q(
        \predict_PC[6][28] ) );
  DFFR_X1 \predict_PC_reg[6][27]  ( .D(n1883), .CK(clock), .RN(n2298), .Q(
        \predict_PC[6][27] ) );
  DFFR_X1 \predict_PC_reg[6][26]  ( .D(n1882), .CK(clock), .RN(n2299), .Q(
        \predict_PC[6][26] ) );
  DFFR_X1 \predict_PC_reg[6][25]  ( .D(n1881), .CK(clock), .RN(n2300), .Q(
        \predict_PC[6][25] ) );
  DFFR_X1 \predict_PC_reg[6][24]  ( .D(n1880), .CK(clock), .RN(n2311), .Q(
        \predict_PC[6][24] ) );
  DFFR_X1 \predict_PC_reg[6][23]  ( .D(n1879), .CK(clock), .RN(n2288), .Q(
        \predict_PC[6][23] ) );
  DFFR_X1 \predict_PC_reg[6][22]  ( .D(n1878), .CK(clock), .RN(n2288), .Q(
        \predict_PC[6][22] ) );
  DFFR_X1 \predict_PC_reg[6][21]  ( .D(n1877), .CK(clock), .RN(n2311), .Q(
        \predict_PC[6][21] ) );
  DFFR_X1 \predict_PC_reg[6][20]  ( .D(n1876), .CK(clock), .RN(n2308), .Q(
        \predict_PC[6][20] ) );
  DFFR_X1 \predict_PC_reg[6][19]  ( .D(n1875), .CK(clock), .RN(n2311), .Q(
        \predict_PC[6][19] ) );
  DFFR_X1 \predict_PC_reg[6][18]  ( .D(n1874), .CK(clock), .RN(n2288), .Q(
        \predict_PC[6][18] ) );
  DFFR_X1 \predict_PC_reg[6][17]  ( .D(n1873), .CK(clock), .RN(n2304), .Q(
        \predict_PC[6][17] ) );
  DFFR_X1 \predict_PC_reg[6][16]  ( .D(n1872), .CK(clock), .RN(n2289), .Q(
        \predict_PC[6][16] ) );
  DFFR_X1 \predict_PC_reg[6][15]  ( .D(n1871), .CK(clock), .RN(n2289), .Q(
        \predict_PC[6][15] ) );
  DFFR_X1 \predict_PC_reg[6][14]  ( .D(n1870), .CK(clock), .RN(n2289), .Q(
        \predict_PC[6][14] ) );
  DFFR_X1 \predict_PC_reg[6][13]  ( .D(n1869), .CK(clock), .RN(n2289), .Q(
        \predict_PC[6][13] ) );
  DFFR_X1 \predict_PC_reg[6][12]  ( .D(n1868), .CK(clock), .RN(n2289), .Q(
        \predict_PC[6][12] ) );
  DFFR_X1 \predict_PC_reg[6][11]  ( .D(n1867), .CK(clock), .RN(n2289), .Q(
        \predict_PC[6][11] ) );
  DFFR_X1 \predict_PC_reg[6][10]  ( .D(n1866), .CK(clock), .RN(n2289), .Q(
        \predict_PC[6][10] ) );
  DFFR_X1 \predict_PC_reg[6][9]  ( .D(n1865), .CK(clock), .RN(n2304), .Q(
        \predict_PC[6][9] ) );
  DFFR_X1 \predict_PC_reg[6][8]  ( .D(n1864), .CK(clock), .RN(n2289), .Q(
        \predict_PC[6][8] ) );
  DFFR_X1 \predict_PC_reg[6][7]  ( .D(n1863), .CK(clock), .RN(n2289), .Q(
        \predict_PC[6][7] ) );
  DFFR_X1 \predict_PC_reg[6][6]  ( .D(n1862), .CK(clock), .RN(n2308), .Q(
        \predict_PC[6][6] ) );
  DFFR_X1 \predict_PC_reg[6][5]  ( .D(n1861), .CK(clock), .RN(n2306), .Q(
        \predict_PC[6][5] ) );
  DFFR_X1 \predict_PC_reg[6][4]  ( .D(n1860), .CK(clock), .RN(n2289), .Q(
        \predict_PC[6][4] ) );
  DFFR_X1 \predict_PC_reg[6][3]  ( .D(n1859), .CK(clock), .RN(n2289), .Q(
        \predict_PC[6][3] ) );
  DFFR_X1 \predict_PC_reg[6][2]  ( .D(n1858), .CK(clock), .RN(n2300), .Q(
        \predict_PC[6][2] ) );
  DFFR_X1 \predict_PC_reg[6][1]  ( .D(n1857), .CK(clock), .RN(n2307), .Q(
        \predict_PC[6][1] ) );
  DFFR_X1 \predict_PC_reg[6][0]  ( .D(n1856), .CK(clock), .RN(n2310), .Q(
        \predict_PC[6][0] ) );
  DFFR_X1 \predict_PC_reg[7][31]  ( .D(n1855), .CK(clock), .RN(n2309), .Q(
        \predict_PC[7][31] ) );
  DFFR_X1 \predict_PC_reg[7][30]  ( .D(n1854), .CK(clock), .RN(n2303), .Q(
        \predict_PC[7][30] ) );
  DFFR_X1 \predict_PC_reg[7][29]  ( .D(n1853), .CK(clock), .RN(n2302), .Q(
        \predict_PC[7][29] ) );
  DFFR_X1 \predict_PC_reg[7][28]  ( .D(n1852), .CK(clock), .RN(n2309), .Q(
        \predict_PC[7][28] ) );
  DFFR_X1 \predict_PC_reg[7][27]  ( .D(n1851), .CK(clock), .RN(n2298), .Q(
        \predict_PC[7][27] ) );
  DFFR_X1 \predict_PC_reg[7][26]  ( .D(n1850), .CK(clock), .RN(n2299), .Q(
        \predict_PC[7][26] ) );
  DFFR_X1 \predict_PC_reg[7][25]  ( .D(n1849), .CK(clock), .RN(n2300), .Q(
        \predict_PC[7][25] ) );
  DFFR_X1 \predict_PC_reg[7][24]  ( .D(n1848), .CK(clock), .RN(n2309), .Q(
        \predict_PC[7][24] ) );
  DFFR_X1 \predict_PC_reg[7][23]  ( .D(n1847), .CK(clock), .RN(n2309), .Q(
        \predict_PC[7][23] ) );
  DFFR_X1 \predict_PC_reg[7][22]  ( .D(n1846), .CK(clock), .RN(n2309), .Q(
        \predict_PC[7][22] ) );
  DFFR_X1 \predict_PC_reg[7][21]  ( .D(n1845), .CK(clock), .RN(n2291), .Q(
        \predict_PC[7][21] ) );
  DFFR_X1 \predict_PC_reg[7][20]  ( .D(n1844), .CK(clock), .RN(n2291), .Q(
        \predict_PC[7][20] ) );
  DFFR_X1 \predict_PC_reg[7][19]  ( .D(n1843), .CK(clock), .RN(n2291), .Q(
        \predict_PC[7][19] ) );
  DFFR_X1 \predict_PC_reg[7][18]  ( .D(n1842), .CK(clock), .RN(n2288), .Q(
        \predict_PC[7][18] ) );
  DFFR_X1 \predict_PC_reg[7][17]  ( .D(n1841), .CK(clock), .RN(n2291), .Q(
        \predict_PC[7][17] ) );
  DFFR_X1 \predict_PC_reg[7][16]  ( .D(n1840), .CK(clock), .RN(n2291), .Q(
        \predict_PC[7][16] ) );
  DFFR_X1 \predict_PC_reg[7][15]  ( .D(n1839), .CK(clock), .RN(n2291), .Q(
        \predict_PC[7][15] ) );
  DFFR_X1 \predict_PC_reg[7][14]  ( .D(n1838), .CK(clock), .RN(n2291), .Q(
        \predict_PC[7][14] ) );
  DFFR_X1 \predict_PC_reg[7][13]  ( .D(n1837), .CK(clock), .RN(n2291), .Q(
        \predict_PC[7][13] ) );
  DFFR_X1 \predict_PC_reg[7][12]  ( .D(n1836), .CK(clock), .RN(n2291), .Q(
        \predict_PC[7][12] ) );
  DFFR_X1 \predict_PC_reg[7][11]  ( .D(n1835), .CK(clock), .RN(n2291), .Q(
        \predict_PC[7][11] ) );
  DFFR_X1 \predict_PC_reg[7][10]  ( .D(n1834), .CK(clock), .RN(n2291), .Q(
        \predict_PC[7][10] ) );
  DFFR_X1 \predict_PC_reg[7][9]  ( .D(n1833), .CK(clock), .RN(n2304), .Q(
        \predict_PC[7][9] ) );
  DFFR_X1 \predict_PC_reg[7][8]  ( .D(n1832), .CK(clock), .RN(n2291), .Q(
        \predict_PC[7][8] ) );
  DFFR_X1 \predict_PC_reg[7][7]  ( .D(n1831), .CK(clock), .RN(n2308), .Q(
        \predict_PC[7][7] ) );
  DFFR_X1 \predict_PC_reg[7][6]  ( .D(n1830), .CK(clock), .RN(n2308), .Q(
        \predict_PC[7][6] ) );
  DFFR_X1 \predict_PC_reg[7][5]  ( .D(n1829), .CK(clock), .RN(n2306), .Q(
        \predict_PC[7][5] ) );
  DFFR_X1 \predict_PC_reg[7][4]  ( .D(n1828), .CK(clock), .RN(n2308), .Q(
        \predict_PC[7][4] ) );
  DFFR_X1 \predict_PC_reg[7][3]  ( .D(n1827), .CK(clock), .RN(n2308), .Q(
        \predict_PC[7][3] ) );
  DFFR_X1 \predict_PC_reg[7][2]  ( .D(n1826), .CK(clock), .RN(n2308), .Q(
        \predict_PC[7][2] ) );
  DFFR_X1 \predict_PC_reg[7][1]  ( .D(n1825), .CK(clock), .RN(n2307), .Q(
        \predict_PC[7][1] ) );
  DFFR_X1 \predict_PC_reg[7][0]  ( .D(n1824), .CK(clock), .RN(n2308), .Q(
        \predict_PC[7][0] ) );
  DFFR_X1 \predict_PC_reg[8][31]  ( .D(n1823), .CK(clock), .RN(n2309), .Q(
        \predict_PC[8][31] ) );
  DFFR_X1 \predict_PC_reg[8][30]  ( .D(n1822), .CK(clock), .RN(n2303), .Q(
        \predict_PC[8][30] ) );
  DFFR_X1 \predict_PC_reg[8][29]  ( .D(n1821), .CK(clock), .RN(n2302), .Q(
        \predict_PC[8][29] ) );
  DFFR_X1 \predict_PC_reg[8][28]  ( .D(n1820), .CK(clock), .RN(n2309), .Q(
        \predict_PC[8][28] ) );
  DFFR_X1 \predict_PC_reg[8][27]  ( .D(n1819), .CK(clock), .RN(n2298), .Q(
        \predict_PC[8][27] ) );
  DFFR_X1 \predict_PC_reg[8][26]  ( .D(n1818), .CK(clock), .RN(n2299), .Q(
        \predict_PC[8][26] ) );
  DFFR_X1 \predict_PC_reg[8][25]  ( .D(n1817), .CK(clock), .RN(n2300), .Q(
        \predict_PC[8][25] ) );
  DFFR_X1 \predict_PC_reg[8][24]  ( .D(n1816), .CK(clock), .RN(n2309), .Q(
        \predict_PC[8][24] ) );
  DFFR_X1 \predict_PC_reg[8][23]  ( .D(n1815), .CK(clock), .RN(n2290), .Q(
        \predict_PC[8][23] ) );
  DFFR_X1 \predict_PC_reg[8][22]  ( .D(n1814), .CK(clock), .RN(n2288), .Q(
        \predict_PC[8][22] ) );
  DFFR_X1 \predict_PC_reg[8][21]  ( .D(n1813), .CK(clock), .RN(n2288), .Q(
        \predict_PC[8][21] ) );
  DFFR_X1 \predict_PC_reg[8][20]  ( .D(n1812), .CK(clock), .RN(n2309), .Q(
        \predict_PC[8][20] ) );
  DFFR_X1 \predict_PC_reg[8][19]  ( .D(n1811), .CK(clock), .RN(n2311), .Q(
        \predict_PC[8][19] ) );
  DFFR_X1 \predict_PC_reg[8][18]  ( .D(n1810), .CK(clock), .RN(n2301), .Q(
        \predict_PC[8][18] ) );
  DFFR_X1 \predict_PC_reg[8][17]  ( .D(n1809), .CK(clock), .RN(n2300), .Q(
        \predict_PC[8][17] ) );
  DFFR_X1 \predict_PC_reg[8][16]  ( .D(n1808), .CK(clock), .RN(n2292), .Q(
        \predict_PC[8][16] ) );
  DFFR_X1 \predict_PC_reg[8][15]  ( .D(n1807), .CK(clock), .RN(n2290), .Q(
        \predict_PC[8][15] ) );
  DFFR_X1 \predict_PC_reg[8][14]  ( .D(n1806), .CK(clock), .RN(n2311), .Q(
        \predict_PC[8][14] ) );
  DFFR_X1 \predict_PC_reg[8][13]  ( .D(n1805), .CK(clock), .RN(n2290), .Q(
        \predict_PC[8][13] ) );
  DFFR_X1 \predict_PC_reg[8][12]  ( .D(n1804), .CK(clock), .RN(n2290), .Q(
        \predict_PC[8][12] ) );
  DFFR_X1 \predict_PC_reg[8][11]  ( .D(n1803), .CK(clock), .RN(n2290), .Q(
        \predict_PC[8][11] ) );
  DFFR_X1 \predict_PC_reg[8][10]  ( .D(n1802), .CK(clock), .RN(n2305), .Q(
        \predict_PC[8][10] ) );
  DFFR_X1 \predict_PC_reg[8][9]  ( .D(n1801), .CK(clock), .RN(n2304), .Q(
        \predict_PC[8][9] ) );
  DFFR_X1 \predict_PC_reg[8][8]  ( .D(n1800), .CK(clock), .RN(n2290), .Q(
        \predict_PC[8][8] ) );
  DFFR_X1 \predict_PC_reg[8][7]  ( .D(n1799), .CK(clock), .RN(n2289), .Q(
        \predict_PC[8][7] ) );
  DFFR_X1 \predict_PC_reg[8][6]  ( .D(n1798), .CK(clock), .RN(n2292), .Q(
        \predict_PC[8][6] ) );
  DFFR_X1 \predict_PC_reg[8][5]  ( .D(n1797), .CK(clock), .RN(n2295), .Q(
        \predict_PC[8][5] ) );
  DFFR_X1 \predict_PC_reg[8][4]  ( .D(n1796), .CK(clock), .RN(n2290), .Q(
        \predict_PC[8][4] ) );
  DFFR_X1 \predict_PC_reg[8][3]  ( .D(n1795), .CK(clock), .RN(n2289), .Q(
        \predict_PC[8][3] ) );
  DFFR_X1 \predict_PC_reg[8][2]  ( .D(n1794), .CK(clock), .RN(n2300), .Q(
        \predict_PC[8][2] ) );
  DFFR_X1 \predict_PC_reg[8][1]  ( .D(n1793), .CK(clock), .RN(n2307), .Q(
        \predict_PC[8][1] ) );
  DFFR_X1 \predict_PC_reg[8][0]  ( .D(n1792), .CK(clock), .RN(n2306), .Q(
        \predict_PC[8][0] ) );
  DFFR_X1 \predict_PC_reg[9][31]  ( .D(n1791), .CK(clock), .RN(n2296), .Q(
        \predict_PC[9][31] ) );
  DFFR_X1 \predict_PC_reg[9][30]  ( .D(n1790), .CK(clock), .RN(n2303), .Q(
        \predict_PC[9][30] ) );
  DFFR_X1 \predict_PC_reg[9][29]  ( .D(n1789), .CK(clock), .RN(n2297), .Q(
        \predict_PC[9][29] ) );
  DFFR_X1 \predict_PC_reg[9][28]  ( .D(n1788), .CK(clock), .RN(n2296), .Q(
        \predict_PC[9][28] ) );
  DFFR_X1 \predict_PC_reg[9][27]  ( .D(n1787), .CK(clock), .RN(n2298), .Q(
        \predict_PC[9][27] ) );
  DFFR_X1 \predict_PC_reg[9][26]  ( .D(n1786), .CK(clock), .RN(n2299), .Q(
        \predict_PC[9][26] ) );
  DFFR_X1 \predict_PC_reg[9][25]  ( .D(n1785), .CK(clock), .RN(n2300), .Q(
        \predict_PC[9][25] ) );
  DFFR_X1 \predict_PC_reg[9][24]  ( .D(n1784), .CK(clock), .RN(n2296), .Q(
        \predict_PC[9][24] ) );
  DFFR_X1 \predict_PC_reg[9][23]  ( .D(n1783), .CK(clock), .RN(n2296), .Q(
        \predict_PC[9][23] ) );
  DFFR_X1 \predict_PC_reg[9][22]  ( .D(n1782), .CK(clock), .RN(n2296), .Q(
        \predict_PC[9][22] ) );
  DFFR_X1 \predict_PC_reg[9][21]  ( .D(n1781), .CK(clock), .RN(n2296), .Q(
        \predict_PC[9][21] ) );
  DFFR_X1 \predict_PC_reg[9][20]  ( .D(n1780), .CK(clock), .RN(n2296), .Q(
        \predict_PC[9][20] ) );
  DFFR_X1 \predict_PC_reg[9][19]  ( .D(n1779), .CK(clock), .RN(n2296), .Q(
        \predict_PC[9][19] ) );
  DFFR_X1 \predict_PC_reg[9][18]  ( .D(n1778), .CK(clock), .RN(n2301), .Q(
        \predict_PC[9][18] ) );
  DFFR_X1 \predict_PC_reg[9][17]  ( .D(n1777), .CK(clock), .RN(n2296), .Q(
        \predict_PC[9][17] ) );
  DFFR_X1 \predict_PC_reg[9][16]  ( .D(n1776), .CK(clock), .RN(n2296), .Q(
        \predict_PC[9][16] ) );
  DFFR_X1 \predict_PC_reg[9][15]  ( .D(n1775), .CK(clock), .RN(n2305), .Q(
        \predict_PC[9][15] ) );
  DFFR_X1 \predict_PC_reg[9][14]  ( .D(n1774), .CK(clock), .RN(n2305), .Q(
        \predict_PC[9][14] ) );
  DFFR_X1 \predict_PC_reg[9][13]  ( .D(n1773), .CK(clock), .RN(n2305), .Q(
        \predict_PC[9][13] ) );
  DFFR_X1 \predict_PC_reg[9][12]  ( .D(n1772), .CK(clock), .RN(n2305), .Q(
        \predict_PC[9][12] ) );
  DFFR_X1 \predict_PC_reg[9][11]  ( .D(n1771), .CK(clock), .RN(n2305), .Q(
        \predict_PC[9][11] ) );
  DFFR_X1 \predict_PC_reg[9][10]  ( .D(n1770), .CK(clock), .RN(n2305), .Q(
        \predict_PC[9][10] ) );
  DFFR_X1 \predict_PC_reg[9][9]  ( .D(n1769), .CK(clock), .RN(n2304), .Q(
        \predict_PC[9][9] ) );
  DFFR_X1 \predict_PC_reg[9][8]  ( .D(n1768), .CK(clock), .RN(n2305), .Q(
        \predict_PC[9][8] ) );
  DFFR_X1 \predict_PC_reg[9][7]  ( .D(n1767), .CK(clock), .RN(n2305), .Q(
        \predict_PC[9][7] ) );
  DFFR_X1 \predict_PC_reg[9][6]  ( .D(n1766), .CK(clock), .RN(n2305), .Q(
        \predict_PC[9][6] ) );
  DFFR_X1 \predict_PC_reg[9][5]  ( .D(n1765), .CK(clock), .RN(n2295), .Q(
        \predict_PC[9][5] ) );
  DFFR_X1 \predict_PC_reg[9][4]  ( .D(n1764), .CK(clock), .RN(n2305), .Q(
        \predict_PC[9][4] ) );
  DFFR_X1 \predict_PC_reg[9][3]  ( .D(n1763), .CK(clock), .RN(n2305), .Q(
        \predict_PC[9][3] ) );
  DFFR_X1 \predict_PC_reg[9][2]  ( .D(n1762), .CK(clock), .RN(n2305), .Q(
        \predict_PC[9][2] ) );
  DFFR_X1 \predict_PC_reg[9][1]  ( .D(n1761), .CK(clock), .RN(n2307), .Q(
        \predict_PC[9][1] ) );
  DFFR_X1 \predict_PC_reg[9][0]  ( .D(n1760), .CK(clock), .RN(n2290), .Q(
        \predict_PC[9][0] ) );
  DFFR_X1 \predict_PC_reg[10][31]  ( .D(n1759), .CK(clock), .RN(n2310), .Q(
        \predict_PC[10][31] ) );
  DFFR_X1 \predict_PC_reg[10][30]  ( .D(n1758), .CK(clock), .RN(n2303), .Q(
        \predict_PC[10][30] ) );
  DFFR_X1 \predict_PC_reg[10][29]  ( .D(n1757), .CK(clock), .RN(n2298), .Q(
        \predict_PC[10][29] ) );
  DFFR_X1 \predict_PC_reg[10][28]  ( .D(n1756), .CK(clock), .RN(n2310), .Q(
        \predict_PC[10][28] ) );
  DFFR_X1 \predict_PC_reg[10][27]  ( .D(n1755), .CK(clock), .RN(n2298), .Q(
        \predict_PC[10][27] ) );
  DFFR_X1 \predict_PC_reg[10][26]  ( .D(n1754), .CK(clock), .RN(n2299), .Q(
        \predict_PC[10][26] ) );
  DFFR_X1 \predict_PC_reg[10][25]  ( .D(n1753), .CK(clock), .RN(n2300), .Q(
        \predict_PC[10][25] ) );
  DFFR_X1 \predict_PC_reg[10][24]  ( .D(n1752), .CK(clock), .RN(n2310), .Q(
        \predict_PC[10][24] ) );
  DFFR_X1 \predict_PC_reg[10][23]  ( .D(n1751), .CK(clock), .RN(n2297), .Q(
        \predict_PC[10][23] ) );
  DFFR_X1 \predict_PC_reg[10][22]  ( .D(n1750), .CK(clock), .RN(n2288), .Q(
        \predict_PC[10][22] ) );
  DFFR_X1 \predict_PC_reg[10][21]  ( .D(n1749), .CK(clock), .RN(n2288), .Q(
        \predict_PC[10][21] ) );
  DFFR_X1 \predict_PC_reg[10][20]  ( .D(n1748), .CK(clock), .RN(n2310), .Q(
        \predict_PC[10][20] ) );
  DFFR_X1 \predict_PC_reg[10][19]  ( .D(n1747), .CK(clock), .RN(n2311), .Q(
        \predict_PC[10][19] ) );
  DFFR_X1 \predict_PC_reg[10][18]  ( .D(n1746), .CK(clock), .RN(n2301), .Q(
        \predict_PC[10][18] ) );
  DFFR_X1 \predict_PC_reg[10][17]  ( .D(n1745), .CK(clock), .RN(n2300), .Q(
        \predict_PC[10][17] ) );
  DFFR_X1 \predict_PC_reg[10][16]  ( .D(n1744), .CK(clock), .RN(n2310), .Q(
        \predict_PC[10][16] ) );
  DFFR_X1 \predict_PC_reg[10][15]  ( .D(n1743), .CK(clock), .RN(n2310), .Q(
        \predict_PC[10][15] ) );
  DFFR_X1 \predict_PC_reg[10][14]  ( .D(n1742), .CK(clock), .RN(n2311), .Q(
        \predict_PC[10][14] ) );
  DFFR_X1 \predict_PC_reg[10][13]  ( .D(n1741), .CK(clock), .RN(n2310), .Q(
        \predict_PC[10][13] ) );
  DFFR_X1 \predict_PC_reg[10][12]  ( .D(n1740), .CK(clock), .RN(n2310), .Q(
        \predict_PC[10][12] ) );
  DFFR_X1 \predict_PC_reg[10][11]  ( .D(n1739), .CK(clock), .RN(n2310), .Q(
        \predict_PC[10][11] ) );
  DFFR_X1 \predict_PC_reg[10][10]  ( .D(n1738), .CK(clock), .RN(n2310), .Q(
        \predict_PC[10][10] ) );
  DFFR_X1 \predict_PC_reg[10][9]  ( .D(n1737), .CK(clock), .RN(n2304), .Q(
        \predict_PC[10][9] ) );
  DFFR_X1 \predict_PC_reg[10][8]  ( .D(n1736), .CK(clock), .RN(n2292), .Q(
        \predict_PC[10][8] ) );
  DFFR_X1 \predict_PC_reg[10][7]  ( .D(n1735), .CK(clock), .RN(n2289), .Q(
        \predict_PC[10][7] ) );
  DFFR_X1 \predict_PC_reg[10][6]  ( .D(n1734), .CK(clock), .RN(n2298), .Q(
        \predict_PC[10][6] ) );
  DFFR_X1 \predict_PC_reg[10][5]  ( .D(n1733), .CK(clock), .RN(n2295), .Q(
        \predict_PC[10][5] ) );
  DFFR_X1 \predict_PC_reg[10][4]  ( .D(n1732), .CK(clock), .RN(n2311), .Q(
        \predict_PC[10][4] ) );
  DFFR_X1 \predict_PC_reg[10][3]  ( .D(n1731), .CK(clock), .RN(n2291), .Q(
        \predict_PC[10][3] ) );
  DFFR_X1 \predict_PC_reg[10][2]  ( .D(n1730), .CK(clock), .RN(n2292), .Q(
        \predict_PC[10][2] ) );
  DFFR_X1 \predict_PC_reg[10][1]  ( .D(n1729), .CK(clock), .RN(n2307), .Q(
        \predict_PC[10][1] ) );
  DFFR_X1 \predict_PC_reg[10][0]  ( .D(n1728), .CK(clock), .RN(n2293), .Q(
        \predict_PC[10][0] ) );
  DFFR_X1 \predict_PC_reg[11][31]  ( .D(n1727), .CK(clock), .RN(n2308), .Q(
        \predict_PC[11][31] ) );
  DFFR_X1 \predict_PC_reg[11][30]  ( .D(n1726), .CK(clock), .RN(n2303), .Q(
        \predict_PC[11][30] ) );
  DFFR_X1 \predict_PC_reg[11][29]  ( .D(n1725), .CK(clock), .RN(n2298), .Q(
        \predict_PC[11][29] ) );
  DFFR_X1 \predict_PC_reg[11][28]  ( .D(n1724), .CK(clock), .RN(n2309), .Q(
        \predict_PC[11][28] ) );
  DFFR_X1 \predict_PC_reg[11][27]  ( .D(n1723), .CK(clock), .RN(n2298), .Q(
        \predict_PC[11][27] ) );
  DFFR_X1 \predict_PC_reg[11][26]  ( .D(n1722), .CK(clock), .RN(n2299), .Q(
        \predict_PC[11][26] ) );
  DFFR_X1 \predict_PC_reg[11][25]  ( .D(n1721), .CK(clock), .RN(n2300), .Q(
        \predict_PC[11][25] ) );
  DFFR_X1 \predict_PC_reg[11][24]  ( .D(n1720), .CK(clock), .RN(n2309), .Q(
        \predict_PC[11][24] ) );
  DFFR_X1 \predict_PC_reg[11][23]  ( .D(n1719), .CK(clock), .RN(n2308), .Q(
        \predict_PC[11][23] ) );
  DFFR_X1 \predict_PC_reg[11][22]  ( .D(n1718), .CK(clock), .RN(n2308), .Q(
        \predict_PC[11][22] ) );
  DFFR_X1 \predict_PC_reg[11][21]  ( .D(n1717), .CK(clock), .RN(n2292), .Q(
        \predict_PC[11][21] ) );
  DFFR_X1 \predict_PC_reg[11][20]  ( .D(n1716), .CK(clock), .RN(n2291), .Q(
        \predict_PC[11][20] ) );
  DFFR_X1 \predict_PC_reg[11][19]  ( .D(n1715), .CK(clock), .RN(n2292), .Q(
        \predict_PC[11][19] ) );
  DFFR_X1 \predict_PC_reg[11][18]  ( .D(n1714), .CK(clock), .RN(n2301), .Q(
        \predict_PC[11][18] ) );
  DFFR_X1 \predict_PC_reg[11][17]  ( .D(n1713), .CK(clock), .RN(n2292), .Q(
        \predict_PC[11][17] ) );
  DFFR_X1 \predict_PC_reg[11][16]  ( .D(n1712), .CK(clock), .RN(n2291), .Q(
        \predict_PC[11][16] ) );
  DFFR_X1 \predict_PC_reg[11][15]  ( .D(n1711), .CK(clock), .RN(n2292), .Q(
        \predict_PC[11][15] ) );
  DFFR_X1 \predict_PC_reg[11][14]  ( .D(n1710), .CK(clock), .RN(n2292), .Q(
        \predict_PC[11][14] ) );
  DFFR_X1 \predict_PC_reg[11][13]  ( .D(n1709), .CK(clock), .RN(n2291), .Q(
        \predict_PC[11][13] ) );
  DFFR_X1 \predict_PC_reg[11][12]  ( .D(n1708), .CK(clock), .RN(n2291), .Q(
        \predict_PC[11][12] ) );
  DFFR_X1 \predict_PC_reg[11][11]  ( .D(n1707), .CK(clock), .RN(n2291), .Q(
        \predict_PC[11][11] ) );
  DFFR_X1 \predict_PC_reg[11][10]  ( .D(n1706), .CK(clock), .RN(n2292), .Q(
        \predict_PC[11][10] ) );
  DFFR_X1 \predict_PC_reg[11][9]  ( .D(n1705), .CK(clock), .RN(n2303), .Q(
        \predict_PC[11][9] ) );
  DFFR_X1 \predict_PC_reg[11][8]  ( .D(n1704), .CK(clock), .RN(n2291), .Q(
        \predict_PC[11][8] ) );
  DFFR_X1 \predict_PC_reg[11][7]  ( .D(n1703), .CK(clock), .RN(n2308), .Q(
        \predict_PC[11][7] ) );
  DFFR_X1 \predict_PC_reg[11][6]  ( .D(n1702), .CK(clock), .RN(n2308), .Q(
        \predict_PC[11][6] ) );
  DFFR_X1 \predict_PC_reg[11][5]  ( .D(n1701), .CK(clock), .RN(n2295), .Q(
        \predict_PC[11][5] ) );
  DFFR_X1 \predict_PC_reg[11][4]  ( .D(n1700), .CK(clock), .RN(n2308), .Q(
        \predict_PC[11][4] ) );
  DFFR_X1 \predict_PC_reg[11][3]  ( .D(n1699), .CK(clock), .RN(n2308), .Q(
        \predict_PC[11][3] ) );
  DFFR_X1 \predict_PC_reg[11][2]  ( .D(n1698), .CK(clock), .RN(n2308), .Q(
        \predict_PC[11][2] ) );
  DFFR_X1 \predict_PC_reg[11][1]  ( .D(n1697), .CK(clock), .RN(n2307), .Q(
        \predict_PC[11][1] ) );
  DFFR_X1 \predict_PC_reg[11][0]  ( .D(n1696), .CK(clock), .RN(n2308), .Q(
        \predict_PC[11][0] ) );
  DFFR_X1 \predict_PC_reg[12][31]  ( .D(n1695), .CK(clock), .RN(n2300), .Q(
        \predict_PC[12][31] ) );
  DFFR_X1 \predict_PC_reg[12][30]  ( .D(n1694), .CK(clock), .RN(n2303), .Q(
        \predict_PC[12][30] ) );
  DFFR_X1 \predict_PC_reg[12][29]  ( .D(n1693), .CK(clock), .RN(n2298), .Q(
        \predict_PC[12][29] ) );
  DFFR_X1 \predict_PC_reg[12][28]  ( .D(n1692), .CK(clock), .RN(n2305), .Q(
        \predict_PC[12][28] ) );
  DFFR_X1 \predict_PC_reg[12][27]  ( .D(n1691), .CK(clock), .RN(n2299), .Q(
        \predict_PC[12][27] ) );
  DFFR_X1 \predict_PC_reg[12][26]  ( .D(n1690), .CK(clock), .RN(n2299), .Q(
        \predict_PC[12][26] ) );
  DFFR_X1 \predict_PC_reg[12][25]  ( .D(n1689), .CK(clock), .RN(n2300), .Q(
        \predict_PC[12][25] ) );
  DFFR_X1 \predict_PC_reg[12][24]  ( .D(n1688), .CK(clock), .RN(n2289), .Q(
        \predict_PC[12][24] ) );
  DFFR_X1 \predict_PC_reg[12][23]  ( .D(n1687), .CK(clock), .RN(n2294), .Q(
        \predict_PC[12][23] ) );
  DFFR_X1 \predict_PC_reg[12][22]  ( .D(n1686), .CK(clock), .RN(n2294), .Q(
        \predict_PC[12][22] ) );
  DFFR_X1 \predict_PC_reg[12][21]  ( .D(n1685), .CK(clock), .RN(n2294), .Q(
        \predict_PC[12][21] ) );
  DFFR_X1 \predict_PC_reg[12][20]  ( .D(n1684), .CK(clock), .RN(n2294), .Q(
        \predict_PC[12][20] ) );
  DFFR_X1 \predict_PC_reg[12][19]  ( .D(n1683), .CK(clock), .RN(n2293), .Q(
        \predict_PC[12][19] ) );
  DFFR_X1 \predict_PC_reg[12][18]  ( .D(n1682), .CK(clock), .RN(n2301), .Q(
        \predict_PC[12][18] ) );
  DFFR_X1 \predict_PC_reg[12][17]  ( .D(n1681), .CK(clock), .RN(n2293), .Q(
        \predict_PC[12][17] ) );
  DFFR_X1 \predict_PC_reg[12][16]  ( .D(n1680), .CK(clock), .RN(n2293), .Q(
        \predict_PC[12][16] ) );
  DFFR_X1 \predict_PC_reg[12][15]  ( .D(n1679), .CK(clock), .RN(n2293), .Q(
        \predict_PC[12][15] ) );
  DFFR_X1 \predict_PC_reg[12][14]  ( .D(n1678), .CK(clock), .RN(n2293), .Q(
        \predict_PC[12][14] ) );
  DFFR_X1 \predict_PC_reg[12][13]  ( .D(n1677), .CK(clock), .RN(n2293), .Q(
        \predict_PC[12][13] ) );
  DFFR_X1 \predict_PC_reg[12][12]  ( .D(n1676), .CK(clock), .RN(n2293), .Q(
        \predict_PC[12][12] ) );
  DFFR_X1 \predict_PC_reg[12][11]  ( .D(n1675), .CK(clock), .RN(n2293), .Q(
        \predict_PC[12][11] ) );
  DFFR_X1 \predict_PC_reg[12][10]  ( .D(n1674), .CK(clock), .RN(n2294), .Q(
        \predict_PC[12][10] ) );
  DFFR_X1 \predict_PC_reg[12][9]  ( .D(n1673), .CK(clock), .RN(n2303), .Q(
        \predict_PC[12][9] ) );
  DFFR_X1 \predict_PC_reg[12][8]  ( .D(n1672), .CK(clock), .RN(n2294), .Q(
        \predict_PC[12][8] ) );
  DFFR_X1 \predict_PC_reg[12][7]  ( .D(n1671), .CK(clock), .RN(n2294), .Q(
        \predict_PC[12][7] ) );
  DFFR_X1 \predict_PC_reg[12][6]  ( .D(n1670), .CK(clock), .RN(n2294), .Q(
        \predict_PC[12][6] ) );
  DFFR_X1 \predict_PC_reg[12][5]  ( .D(n1669), .CK(clock), .RN(n2295), .Q(
        \predict_PC[12][5] ) );
  DFFR_X1 \predict_PC_reg[12][4]  ( .D(n1668), .CK(clock), .RN(n2294), .Q(
        \predict_PC[12][4] ) );
  DFFR_X1 \predict_PC_reg[12][3]  ( .D(n1667), .CK(clock), .RN(n2295), .Q(
        \predict_PC[12][3] ) );
  DFFR_X1 \predict_PC_reg[12][2]  ( .D(n1666), .CK(clock), .RN(n2295), .Q(
        \predict_PC[12][2] ) );
  DFFR_X1 \predict_PC_reg[12][1]  ( .D(n1665), .CK(clock), .RN(n2307), .Q(
        \predict_PC[12][1] ) );
  DFFR_X1 \predict_PC_reg[12][0]  ( .D(n1664), .CK(clock), .RN(n2306), .Q(
        \predict_PC[12][0] ) );
  DFFR_X1 \predict_PC_reg[13][31]  ( .D(n1663), .CK(clock), .RN(n2294), .Q(
        \predict_PC[13][31] ) );
  DFFR_X1 \predict_PC_reg[13][30]  ( .D(n1662), .CK(clock), .RN(n2303), .Q(
        \predict_PC[13][30] ) );
  DFFR_X1 \predict_PC_reg[13][29]  ( .D(n1661), .CK(clock), .RN(n2298), .Q(
        \predict_PC[13][29] ) );
  DFFR_X1 \predict_PC_reg[13][28]  ( .D(n1660), .CK(clock), .RN(n2303), .Q(
        \predict_PC[13][28] ) );
  DFFR_X1 \predict_PC_reg[13][27]  ( .D(n1659), .CK(clock), .RN(n2299), .Q(
        \predict_PC[13][27] ) );
  DFFR_X1 \predict_PC_reg[13][26]  ( .D(n1658), .CK(clock), .RN(n2299), .Q(
        \predict_PC[13][26] ) );
  DFFR_X1 \predict_PC_reg[13][25]  ( .D(n1657), .CK(clock), .RN(n2301), .Q(
        \predict_PC[13][25] ) );
  DFFR_X1 \predict_PC_reg[13][24]  ( .D(n1656), .CK(clock), .RN(n2301), .Q(
        \predict_PC[13][24] ) );
  DFFR_X1 \predict_PC_reg[13][23]  ( .D(n1655), .CK(clock), .RN(n2298), .Q(
        \predict_PC[13][23] ) );
  DFFR_X1 \predict_PC_reg[13][22]  ( .D(n1654), .CK(clock), .RN(n2292), .Q(
        \predict_PC[13][22] ) );
  DFFR_X1 \predict_PC_reg[13][21]  ( .D(n1653), .CK(clock), .RN(n2311), .Q(
        \predict_PC[13][21] ) );
  DFFR_X1 \predict_PC_reg[13][20]  ( .D(n1652), .CK(clock), .RN(n2291), .Q(
        \predict_PC[13][20] ) );
  DFFR_X1 \predict_PC_reg[13][19]  ( .D(n1651), .CK(clock), .RN(n2293), .Q(
        \predict_PC[13][19] ) );
  DFFR_X1 \predict_PC_reg[13][18]  ( .D(n1650), .CK(clock), .RN(n2301), .Q(
        \predict_PC[13][18] ) );
  DFFR_X1 \predict_PC_reg[13][17]  ( .D(n1649), .CK(clock), .RN(n2310), .Q(
        \predict_PC[13][17] ) );
  DFFR_X1 \predict_PC_reg[13][16]  ( .D(n1648), .CK(clock), .RN(n2296), .Q(
        \predict_PC[13][16] ) );
  DFFR_X1 \predict_PC_reg[13][15]  ( .D(n1647), .CK(clock), .RN(n2304), .Q(
        \predict_PC[13][15] ) );
  DFFR_X1 \predict_PC_reg[13][14]  ( .D(n1646), .CK(clock), .RN(n2304), .Q(
        \predict_PC[13][14] ) );
  DFFR_X1 \predict_PC_reg[13][13]  ( .D(n1645), .CK(clock), .RN(n2304), .Q(
        \predict_PC[13][13] ) );
  DFFR_X1 \predict_PC_reg[13][12]  ( .D(n1644), .CK(clock), .RN(n2304), .Q(
        \predict_PC[13][12] ) );
  DFFR_X1 \predict_PC_reg[13][11]  ( .D(n1643), .CK(clock), .RN(n2304), .Q(
        \predict_PC[13][11] ) );
  DFFR_X1 \predict_PC_reg[13][10]  ( .D(n1642), .CK(clock), .RN(n2304), .Q(
        \predict_PC[13][10] ) );
  DFFR_X1 \predict_PC_reg[13][9]  ( .D(n1641), .CK(clock), .RN(n2297), .Q(
        \predict_PC[13][9] ) );
  DFFR_X1 \predict_PC_reg[13][8]  ( .D(n1640), .CK(clock), .RN(n2304), .Q(
        \predict_PC[13][8] ) );
  DFFR_X1 \predict_PC_reg[13][7]  ( .D(n1639), .CK(clock), .RN(n2304), .Q(
        \predict_PC[13][7] ) );
  DFFR_X1 \predict_PC_reg[13][6]  ( .D(n1638), .CK(clock), .RN(n2305), .Q(
        \predict_PC[13][6] ) );
  DFFR_X1 \predict_PC_reg[13][5]  ( .D(n1637), .CK(clock), .RN(n2295), .Q(
        \predict_PC[13][5] ) );
  DFFR_X1 \predict_PC_reg[13][4]  ( .D(n1636), .CK(clock), .RN(n2305), .Q(
        \predict_PC[13][4] ) );
  DFFR_X1 \predict_PC_reg[13][3]  ( .D(n1635), .CK(clock), .RN(n2305), .Q(
        \predict_PC[13][3] ) );
  DFFR_X1 \predict_PC_reg[13][2]  ( .D(n1634), .CK(clock), .RN(n2305), .Q(
        \predict_PC[13][2] ) );
  DFFR_X1 \predict_PC_reg[13][1]  ( .D(n1633), .CK(clock), .RN(n2307), .Q(
        \predict_PC[13][1] ) );
  DFFR_X1 \predict_PC_reg[13][0]  ( .D(n1632), .CK(clock), .RN(n2297), .Q(
        \predict_PC[13][0] ) );
  DFFR_X1 \predict_PC_reg[14][31]  ( .D(n1631), .CK(clock), .RN(n2296), .Q(
        \predict_PC[14][31] ) );
  DFFR_X1 \predict_PC_reg[14][30]  ( .D(n1630), .CK(clock), .RN(n2297), .Q(
        \predict_PC[14][30] ) );
  DFFR_X1 \predict_PC_reg[14][29]  ( .D(n1629), .CK(clock), .RN(n2298), .Q(
        \predict_PC[14][29] ) );
  DFFR_X1 \predict_PC_reg[14][28]  ( .D(n1628), .CK(clock), .RN(n2290), .Q(
        \predict_PC[14][28] ) );
  DFFR_X1 \predict_PC_reg[14][27]  ( .D(n1627), .CK(clock), .RN(n2299), .Q(
        \predict_PC[14][27] ) );
  DFFR_X1 \predict_PC_reg[14][26]  ( .D(n1626), .CK(clock), .RN(n2299), .Q(
        \predict_PC[14][26] ) );
  DFFR_X1 \predict_PC_reg[14][25]  ( .D(n1625), .CK(clock), .RN(n2301), .Q(
        \predict_PC[14][25] ) );
  DFFR_X1 \predict_PC_reg[14][24]  ( .D(n1624), .CK(clock), .RN(n2302), .Q(
        \predict_PC[14][24] ) );
  DFFR_X1 \predict_PC_reg[14][23]  ( .D(n1623), .CK(clock), .RN(n2299), .Q(
        \predict_PC[14][23] ) );
  DFFR_X1 \predict_PC_reg[14][22]  ( .D(n1622), .CK(clock), .RN(n2288), .Q(
        \predict_PC[14][22] ) );
  DFFR_X1 \predict_PC_reg[14][21]  ( .D(n1621), .CK(clock), .RN(n2288), .Q(
        \predict_PC[14][21] ) );
  DFFR_X1 \predict_PC_reg[14][20]  ( .D(n1620), .CK(clock), .RN(n2307), .Q(
        \predict_PC[14][20] ) );
  DFFR_X1 \predict_PC_reg[14][19]  ( .D(n1619), .CK(clock), .RN(n2311), .Q(
        \predict_PC[14][19] ) );
  DFFR_X1 \predict_PC_reg[14][18]  ( .D(n1618), .CK(clock), .RN(n2301), .Q(
        \predict_PC[14][18] ) );
  DFFR_X1 \predict_PC_reg[14][17]  ( .D(n1617), .CK(clock), .RN(n2300), .Q(
        \predict_PC[14][17] ) );
  DFFR_X1 \predict_PC_reg[14][16]  ( .D(n1616), .CK(clock), .RN(n2304), .Q(
        \predict_PC[14][16] ) );
  DFFR_X1 \predict_PC_reg[14][15]  ( .D(n1615), .CK(clock), .RN(n2289), .Q(
        \predict_PC[14][15] ) );
  DFFR_X1 \predict_PC_reg[14][14]  ( .D(n1614), .CK(clock), .RN(n2311), .Q(
        \predict_PC[14][14] ) );
  DFFR_X1 \predict_PC_reg[14][13]  ( .D(n1613), .CK(clock), .RN(n2305), .Q(
        \predict_PC[14][13] ) );
  DFFR_X1 \predict_PC_reg[14][12]  ( .D(n1612), .CK(clock), .RN(n2304), .Q(
        \predict_PC[14][12] ) );
  DFFR_X1 \predict_PC_reg[14][11]  ( .D(n1611), .CK(clock), .RN(n2307), .Q(
        \predict_PC[14][11] ) );
  DFFR_X1 \predict_PC_reg[14][10]  ( .D(n1610), .CK(clock), .RN(n2302), .Q(
        \predict_PC[14][10] ) );
  DFFR_X1 \predict_PC_reg[14][9]  ( .D(n1609), .CK(clock), .RN(n2297), .Q(
        \predict_PC[14][9] ) );
  DFFR_X1 \predict_PC_reg[14][8]  ( .D(n1608), .CK(clock), .RN(n2290), .Q(
        \predict_PC[14][8] ) );
  DFFR_X1 \predict_PC_reg[14][7]  ( .D(n1607), .CK(clock), .RN(n2289), .Q(
        \predict_PC[14][7] ) );
  DFFR_X1 \predict_PC_reg[14][6]  ( .D(n1606), .CK(clock), .RN(n2294), .Q(
        \predict_PC[14][6] ) );
  DFFR_X1 \predict_PC_reg[14][5]  ( .D(n1605), .CK(clock), .RN(n2295), .Q(
        \predict_PC[14][5] ) );
  DFFR_X1 \predict_PC_reg[14][4]  ( .D(n1604), .CK(clock), .RN(n2296), .Q(
        \predict_PC[14][4] ) );
  DFFR_X1 \predict_PC_reg[14][3]  ( .D(n1603), .CK(clock), .RN(n2310), .Q(
        \predict_PC[14][3] ) );
  DFFR_X1 \predict_PC_reg[14][2]  ( .D(n1602), .CK(clock), .RN(n2309), .Q(
        \predict_PC[14][2] ) );
  DFFR_X1 \predict_PC_reg[14][1]  ( .D(n1601), .CK(clock), .RN(n2307), .Q(
        \predict_PC[14][1] ) );
  DFFR_X1 \predict_PC_reg[14][0]  ( .D(n1600), .CK(clock), .RN(n2293), .Q(
        \predict_PC[14][0] ) );
  DFFR_X1 \predict_PC_reg[15][31]  ( .D(n1599), .CK(clock), .RN(n2299), .Q(
        \predict_PC[15][31] ) );
  DFFR_X1 \last_PC_reg[31]  ( .D(n1598), .CK(clock), .RN(n2297), .QN(n593) );
  DFFR_X1 \predict_PC_reg[15][30]  ( .D(n1597), .CK(clock), .RN(n2297), .Q(
        \predict_PC[15][30] ) );
  DFFR_X1 \last_PC_reg[30]  ( .D(n1596), .CK(clock), .RN(n2297), .Q(n6) );
  DFFR_X1 \predict_PC_reg[15][29]  ( .D(n1595), .CK(clock), .RN(n2298), .Q(
        \predict_PC[15][29] ) );
  DFFR_X1 \last_PC_reg[29]  ( .D(n1594), .CK(clock), .RN(n2298), .Q(n7) );
  DFFR_X1 \predict_PC_reg[15][28]  ( .D(n1593), .CK(clock), .RN(n2297), .Q(
        \predict_PC[15][28] ) );
  DFFR_X1 \last_PC_reg[28]  ( .D(n1592), .CK(clock), .RN(n2297), .Q(n8) );
  DFFR_X1 \predict_PC_reg[15][27]  ( .D(n1591), .CK(clock), .RN(n2299), .Q(
        \predict_PC[15][27] ) );
  DFFR_X1 \last_PC_reg[27]  ( .D(n1590), .CK(clock), .RN(n2303), .Q(n9) );
  DFFR_X1 \predict_PC_reg[15][26]  ( .D(n1589), .CK(clock), .RN(n2302), .Q(
        \predict_PC[15][26] ) );
  DFFR_X1 \last_PC_reg[26]  ( .D(n1588), .CK(clock), .RN(n2302), .QN(n598) );
  DFFR_X1 \predict_PC_reg[15][25]  ( .D(n1587), .CK(clock), .RN(n2301), .Q(
        \predict_PC[15][25] ) );
  DFFR_X1 \last_PC_reg[25]  ( .D(n1586), .CK(clock), .RN(n2301), .QN(n599) );
  DFFR_X1 \predict_PC_reg[15][24]  ( .D(n1585), .CK(clock), .RN(n2309), .Q(
        \predict_PC[15][24] ) );
  DFFR_X1 \last_PC_reg[24]  ( .D(n1584), .CK(clock), .RN(n2297), .QN(n600) );
  DFFR_X1 \predict_PC_reg[15][23]  ( .D(n1583), .CK(clock), .RN(n2306), .Q(
        \predict_PC[15][23] ) );
  DFFR_X1 \last_PC_reg[23]  ( .D(n1582), .CK(clock), .RN(n2301), .QN(n601) );
  DFFR_X1 \predict_PC_reg[15][22]  ( .D(n1581), .CK(clock), .RN(n2288), .Q(
        \predict_PC[15][22] ) );
  DFFR_X1 \last_PC_reg[22]  ( .D(n1580), .CK(clock), .RN(n2301), .QN(n602) );
  DFFR_X1 \predict_PC_reg[15][21]  ( .D(n1579), .CK(clock), .RN(n2288), .Q(
        \predict_PC[15][21] ) );
  DFFR_X1 \last_PC_reg[21]  ( .D(n1578), .CK(clock), .RN(n2301), .QN(n603) );
  DFFR_X1 \predict_PC_reg[15][20]  ( .D(n1577), .CK(clock), .RN(n2304), .Q(
        \predict_PC[15][20] ) );
  DFFR_X1 \last_PC_reg[20]  ( .D(n1576), .CK(clock), .RN(n2297), .QN(n604) );
  DFFR_X1 \predict_PC_reg[15][19]  ( .D(n1575), .CK(clock), .RN(n2311), .Q(
        \predict_PC[15][19] ) );
  DFFR_X1 \last_PC_reg[19]  ( .D(n1574), .CK(clock), .RN(n2301), .QN(n605) );
  DFFR_X1 \predict_PC_reg[15][18]  ( .D(n1573), .CK(clock), .RN(n2300), .Q(
        \predict_PC[15][18] ) );
  DFFR_X1 \last_PC_reg[18]  ( .D(n1572), .CK(clock), .RN(n2304), .QN(n606) );
  DFFR_X1 \predict_PC_reg[15][17]  ( .D(n1571), .CK(clock), .RN(n2300), .Q(
        \predict_PC[15][17] ) );
  DFFR_X1 \last_PC_reg[17]  ( .D(n1570), .CK(clock), .RN(n2300), .QN(n607) );
  DFFR_X1 \predict_PC_reg[15][16]  ( .D(n1569), .CK(clock), .RN(n2300), .Q(
        \predict_PC[15][16] ) );
  DFFR_X1 \last_PC_reg[16]  ( .D(n1568), .CK(clock), .RN(n2297), .QN(n608) );
  DFFR_X1 \predict_PC_reg[15][15]  ( .D(n1567), .CK(clock), .RN(n2290), .Q(
        \predict_PC[15][15] ) );
  DFFR_X1 \last_PC_reg[15]  ( .D(n1566), .CK(clock), .RN(n2303), .QN(n609) );
  DFFR_X1 \predict_PC_reg[15][14]  ( .D(n1565), .CK(clock), .RN(n2311), .Q(
        \predict_PC[15][14] ) );
  DFFR_X1 \last_PC_reg[14]  ( .D(n1564), .CK(clock), .RN(n2301), .QN(n610) );
  DFFR_X1 \predict_PC_reg[15][13]  ( .D(n1563), .CK(clock), .RN(n2290), .Q(
        \predict_PC[15][13] ) );
  DFFR_X1 \last_PC_reg[13]  ( .D(n1562), .CK(clock), .RN(n2303), .QN(n611) );
  DFFR_X1 \predict_PC_reg[15][12]  ( .D(n1561), .CK(clock), .RN(n2296), .Q(
        \predict_PC[15][12] ) );
  DFFR_X1 \last_PC_reg[12]  ( .D(n1560), .CK(clock), .RN(n2297), .QN(n612) );
  DFFR_X1 \predict_PC_reg[15][11]  ( .D(n1559), .CK(clock), .RN(n2298), .Q(
        \predict_PC[15][11] ) );
  DFFR_X1 \last_PC_reg[11]  ( .D(n1558), .CK(clock), .RN(n2298), .QN(n613) );
  DFFR_X1 \predict_PC_reg[15][10]  ( .D(n1557), .CK(clock), .RN(n2310), .Q(
        \predict_PC[15][10] ) );
  DFFR_X1 \last_PC_reg[10]  ( .D(n1556), .CK(clock), .RN(n2302), .QN(n614) );
  DFFR_X1 \predict_PC_reg[15][9]  ( .D(n1555), .CK(clock), .RN(n2297), .Q(
        \predict_PC[15][9] ) );
  DFFR_X1 \last_PC_reg[9]  ( .D(n1554), .CK(clock), .RN(n2297), .QN(n615) );
  DFFR_X1 \predict_PC_reg[15][8]  ( .D(n1553), .CK(clock), .RN(n2294), .Q(
        \predict_PC[15][8] ) );
  DFFR_X1 \last_PC_reg[8]  ( .D(n1552), .CK(clock), .RN(n2298), .QN(n616) );
  DFFR_X1 \predict_PC_reg[15][7]  ( .D(n1551), .CK(clock), .RN(n2289), .Q(
        \predict_PC[15][7] ) );
  DFFR_X1 \last_PC_reg[7]  ( .D(n1550), .CK(clock), .RN(n2301), .QN(n617) );
  DFFR_X1 \predict_PC_reg[15][6]  ( .D(n1549), .CK(clock), .RN(n2303), .Q(
        \predict_PC[15][6] ) );
  DFFR_X1 \last_PC_reg[6]  ( .D(n1548), .CK(clock), .RN(n2289), .QN(n618) );
  DFFR_X1 \predict_PC_reg[15][5]  ( .D(n1547), .CK(clock), .RN(n2295), .Q(
        \predict_PC[15][5] ) );
  DFFR_X1 \last_PC_reg[5]  ( .D(n1546), .CK(clock), .RN(n2295), .QN(n619) );
  DFFR_X1 \predict_PC_reg[15][4]  ( .D(n1545), .CK(clock), .RN(n2301), .Q(
        \predict_PC[15][4] ) );
  DFFR_X1 \last_PC_reg[4]  ( .D(n1544), .CK(clock), .RN(n2297), .QN(n620) );
  DFFR_X1 \predict_PC_reg[15][3]  ( .D(n1543), .CK(clock), .RN(n2310), .Q(
        \predict_PC[15][3] ) );
  DFFR_X1 \last_PC_reg[3]  ( .D(n1542), .CK(clock), .RN(n2302), .QN(n621) );
  DFFR_X1 \predict_PC_reg[15][2]  ( .D(n1541), .CK(clock), .RN(n2297), .Q(
        \predict_PC[15][2] ) );
  DFFR_X1 \last_PC_reg[2]  ( .D(n1540), .CK(clock), .RN(n2307), .QN(n622) );
  DFFR_X1 \predict_PC_reg[15][1]  ( .D(n1539), .CK(clock), .RN(n2307), .Q(
        \predict_PC[15][1] ) );
  DFFR_X1 \last_PC_reg[1]  ( .D(n1538), .CK(clock), .RN(n2295), .QN(n623) );
  DFFR_X1 \predict_PC_reg[15][0]  ( .D(n1537), .CK(clock), .RN(n2307), .Q(
        \predict_PC[15][0] ) );
  DFFR_X1 \last_PC_reg[0]  ( .D(n1536), .CK(clock), .RN(n2297), .QN(n624) );
  DFFR_X1 last_mispredict_reg ( .D(n1535), .CK(clock), .RN(n2294), .QN(n592)
         );
  MUX2_X1 U1603 ( .A(n6), .B(predicted_next_PC_o[30]), .S(n2286), .Z(n1596) );
  MUX2_X1 U1604 ( .A(n7), .B(predicted_next_PC_o[29]), .S(n2286), .Z(n1594) );
  MUX2_X1 U1605 ( .A(n8), .B(predicted_next_PC_o[28]), .S(n2286), .Z(n1592) );
  MUX2_X1 U1606 ( .A(n9), .B(predicted_next_PC_o[27]), .S(n2286), .Z(n1590) );
  predictor_2_0 pred_x_0 ( .clock(clock), .reset(reset), .enable(
        write_enable[0]), .taken_i(was_taken_i), .prediction_o(taken[0]) );
  predictor_2_15 pred_x_1 ( .clock(clock), .reset(reset), .enable(
        write_enable[1]), .taken_i(was_taken_i), .prediction_o(taken[1]) );
  predictor_2_14 pred_x_2 ( .clock(clock), .reset(reset), .enable(
        write_enable[2]), .taken_i(was_taken_i), .prediction_o(taken[2]) );
  predictor_2_13 pred_x_3 ( .clock(clock), .reset(reset), .enable(
        write_enable[3]), .taken_i(was_taken_i), .prediction_o(taken[3]) );
  predictor_2_12 pred_x_4 ( .clock(clock), .reset(reset), .enable(
        write_enable[4]), .taken_i(was_taken_i), .prediction_o(taken[4]) );
  predictor_2_11 pred_x_5 ( .clock(clock), .reset(reset), .enable(
        write_enable[5]), .taken_i(was_taken_i), .prediction_o(taken[5]) );
  predictor_2_10 pred_x_6 ( .clock(clock), .reset(reset), .enable(
        write_enable[6]), .taken_i(was_taken_i), .prediction_o(taken[6]) );
  predictor_2_9 pred_x_7 ( .clock(clock), .reset(reset), .enable(
        write_enable[7]), .taken_i(was_taken_i), .prediction_o(taken[7]) );
  predictor_2_8 pred_x_8 ( .clock(clock), .reset(reset), .enable(
        write_enable[8]), .taken_i(was_taken_i), .prediction_o(taken[8]) );
  predictor_2_7 pred_x_9 ( .clock(clock), .reset(reset), .enable(
        write_enable[9]), .taken_i(was_taken_i), .prediction_o(taken[9]) );
  predictor_2_6 pred_x_10 ( .clock(clock), .reset(reset), .enable(
        write_enable[10]), .taken_i(was_taken_i), .prediction_o(taken[10]) );
  predictor_2_5 pred_x_11 ( .clock(clock), .reset(reset), .enable(
        write_enable[11]), .taken_i(was_taken_i), .prediction_o(taken[11]) );
  predictor_2_4 pred_x_12 ( .clock(clock), .reset(reset), .enable(
        write_enable[12]), .taken_i(was_taken_i), .prediction_o(taken[12]) );
  predictor_2_3 pred_x_13 ( .clock(clock), .reset(reset), .enable(
        write_enable[13]), .taken_i(was_taken_i), .prediction_o(taken[13]) );
  predictor_2_2 pred_x_14 ( .clock(clock), .reset(reset), .enable(
        write_enable[14]), .taken_i(was_taken_i), .prediction_o(taken[14]) );
  predictor_2_1 pred_x_15 ( .clock(clock), .reset(reset), .enable(
        write_enable[15]), .taken_i(was_taken_i), .prediction_o(taken[15]) );
  NAND2_X1 U1552 ( .A1(TAG_i[2]), .A2(TAG_i[3]), .ZN(n2209) );
  NAND2_X1 U1542 ( .A1(TAG_i[0]), .A2(n701), .ZN(n2200) );
  AOI22_X1 U80 ( .A1(n2270), .A2(taken[12]), .B1(n763), .B2(taken[13]), .ZN(
        n752) );
  NAND2_X1 U1548 ( .A1(TAG_i[1]), .A2(TAG_i[0]), .ZN(n2202) );
  AOI22_X1 U79 ( .A1(n2272), .A2(taken[14]), .B1(n761), .B2(taken[15]), .ZN(
        n753) );
  AOI22_X1 U78 ( .A1(n2274), .A2(taken[10]), .B1(n759), .B2(taken[11]), .ZN(
        n754) );
  AOI22_X1 U77 ( .A1(n2276), .A2(taken[8]), .B1(n757), .B2(taken[9]), .ZN(n755) );
  AOI22_X1 U75 ( .A1(n2278), .A2(taken[4]), .B1(n751), .B2(taken[5]), .ZN(n740) );
  AOI22_X1 U74 ( .A1(n2280), .A2(taken[6]), .B1(n749), .B2(taken[7]), .ZN(n741) );
  AOI22_X1 U73 ( .A1(n746), .A2(taken[1]), .B1(n2281), .B2(taken[0]), .ZN(n742) );
  AOI22_X1 U72 ( .A1(n744), .A2(taken[3]), .B1(n745), .B2(taken[2]), .ZN(n743)
         );
  AOI22_X1 U1367 ( .A1(n2272), .A2(\predict_PC[14][11] ), .B1(n2271), .B2(
        \predict_PC[15][11] ), .ZN(n1511) );
  AOI22_X1 U1366 ( .A1(n2270), .A2(\predict_PC[12][11] ), .B1(n2269), .B2(
        \predict_PC[13][11] ), .ZN(n1512) );
  AOI22_X1 U1365 ( .A1(n2276), .A2(\predict_PC[8][11] ), .B1(n2275), .B2(
        \predict_PC[9][11] ), .ZN(n1513) );
  AOI22_X1 U1364 ( .A1(n2274), .A2(\predict_PC[10][11] ), .B1(n2273), .B2(
        \predict_PC[11][11] ), .ZN(n1514) );
  NAND4_X1 U1363 ( .A1(n1511), .A2(n1512), .A3(n1513), .A4(n1514), .ZN(n1505)
         );
  AOI22_X1 U1362 ( .A1(n2280), .A2(\predict_PC[6][11] ), .B1(n2279), .B2(
        \predict_PC[7][11] ), .ZN(n1507) );
  AOI22_X1 U1361 ( .A1(n2278), .A2(\predict_PC[4][11] ), .B1(n2277), .B2(
        \predict_PC[5][11] ), .ZN(n1508) );
  AOI22_X1 U1360 ( .A1(n2284), .A2(\predict_PC[3][11] ), .B1(n2283), .B2(
        \predict_PC[2][11] ), .ZN(n1509) );
  AOI22_X1 U1359 ( .A1(n2282), .A2(\predict_PC[1][11] ), .B1(n2281), .B2(
        \predict_PC[0][11] ), .ZN(n1510) );
  NAND4_X1 U1358 ( .A1(n1507), .A2(n1508), .A3(n1509), .A4(n1510), .ZN(n1506)
         );
  NOR2_X1 U1357 ( .A1(n1505), .A2(n1506), .ZN(n691) );
  AOI22_X1 U1325 ( .A1(n2272), .A2(\predict_PC[14][14] ), .B1(n2271), .B2(
        \predict_PC[15][14] ), .ZN(n1478) );
  AOI22_X1 U1324 ( .A1(n2270), .A2(\predict_PC[12][14] ), .B1(n2269), .B2(
        \predict_PC[13][14] ), .ZN(n1479) );
  AOI22_X1 U1323 ( .A1(n2276), .A2(\predict_PC[8][14] ), .B1(n2275), .B2(
        \predict_PC[9][14] ), .ZN(n1480) );
  AOI22_X1 U1322 ( .A1(n2274), .A2(\predict_PC[10][14] ), .B1(n2273), .B2(
        \predict_PC[11][14] ), .ZN(n1481) );
  NAND4_X1 U1321 ( .A1(n1478), .A2(n1479), .A3(n1480), .A4(n1481), .ZN(n1472)
         );
  AOI22_X1 U1320 ( .A1(n2280), .A2(\predict_PC[6][14] ), .B1(n2279), .B2(
        \predict_PC[7][14] ), .ZN(n1474) );
  AOI22_X1 U1319 ( .A1(n2278), .A2(\predict_PC[4][14] ), .B1(n2277), .B2(
        \predict_PC[5][14] ), .ZN(n1475) );
  AOI22_X1 U1318 ( .A1(n2284), .A2(\predict_PC[3][14] ), .B1(n2283), .B2(
        \predict_PC[2][14] ), .ZN(n1476) );
  AOI22_X1 U1317 ( .A1(n2282), .A2(\predict_PC[1][14] ), .B1(n2281), .B2(
        \predict_PC[0][14] ), .ZN(n1477) );
  NAND4_X1 U1316 ( .A1(n1474), .A2(n1475), .A3(n1476), .A4(n1477), .ZN(n1473)
         );
  NOR2_X1 U1315 ( .A1(n1472), .A2(n1473), .ZN(n688) );
  AOI22_X1 U1381 ( .A1(n2272), .A2(\predict_PC[14][10] ), .B1(n2271), .B2(
        \predict_PC[15][10] ), .ZN(n1522) );
  AOI22_X1 U1380 ( .A1(n2270), .A2(\predict_PC[12][10] ), .B1(n2269), .B2(
        \predict_PC[13][10] ), .ZN(n1523) );
  AOI22_X1 U1379 ( .A1(n2276), .A2(\predict_PC[8][10] ), .B1(n2275), .B2(
        \predict_PC[9][10] ), .ZN(n1524) );
  AOI22_X1 U1378 ( .A1(n2274), .A2(\predict_PC[10][10] ), .B1(n2273), .B2(
        \predict_PC[11][10] ), .ZN(n1525) );
  NAND4_X1 U1377 ( .A1(n1522), .A2(n1523), .A3(n1524), .A4(n1525), .ZN(n1516)
         );
  AOI22_X1 U1376 ( .A1(n2280), .A2(\predict_PC[6][10] ), .B1(n2279), .B2(
        \predict_PC[7][10] ), .ZN(n1518) );
  AOI22_X1 U1375 ( .A1(n2278), .A2(\predict_PC[4][10] ), .B1(n2277), .B2(
        \predict_PC[5][10] ), .ZN(n1519) );
  AOI22_X1 U1374 ( .A1(n2284), .A2(\predict_PC[3][10] ), .B1(n2283), .B2(
        \predict_PC[2][10] ), .ZN(n1520) );
  AOI22_X1 U1373 ( .A1(n2282), .A2(\predict_PC[1][10] ), .B1(n2281), .B2(
        \predict_PC[0][10] ), .ZN(n1521) );
  NAND4_X1 U1372 ( .A1(n1518), .A2(n1519), .A3(n1520), .A4(n1521), .ZN(n1517)
         );
  NOR2_X1 U1371 ( .A1(n1516), .A2(n1517), .ZN(n692) );
  AOI22_X1 U1091 ( .A1(n2272), .A2(\predict_PC[14][31] ), .B1(n2271), .B2(
        \predict_PC[15][31] ), .ZN(n1291) );
  AOI22_X1 U1090 ( .A1(n2270), .A2(\predict_PC[12][31] ), .B1(n2269), .B2(
        \predict_PC[13][31] ), .ZN(n1292) );
  AOI22_X1 U1089 ( .A1(n2276), .A2(\predict_PC[8][31] ), .B1(n2275), .B2(
        \predict_PC[9][31] ), .ZN(n1293) );
  AOI22_X1 U1088 ( .A1(n2274), .A2(\predict_PC[10][31] ), .B1(n2273), .B2(
        \predict_PC[11][31] ), .ZN(n1294) );
  NAND4_X1 U1087 ( .A1(n1291), .A2(n1292), .A3(n1293), .A4(n1294), .ZN(n1285)
         );
  AOI22_X1 U1086 ( .A1(n2280), .A2(\predict_PC[6][31] ), .B1(n2279), .B2(
        \predict_PC[7][31] ), .ZN(n1287) );
  AOI22_X1 U1085 ( .A1(n2278), .A2(\predict_PC[4][31] ), .B1(n2277), .B2(
        \predict_PC[5][31] ), .ZN(n1288) );
  AOI22_X1 U1084 ( .A1(n2284), .A2(\predict_PC[3][31] ), .B1(n2283), .B2(
        \predict_PC[2][31] ), .ZN(n1289) );
  AOI22_X1 U1083 ( .A1(n2282), .A2(\predict_PC[1][31] ), .B1(n2281), .B2(
        \predict_PC[0][31] ), .ZN(n1290) );
  NAND4_X1 U1082 ( .A1(n1287), .A2(n1288), .A3(n1289), .A4(n1290), .ZN(n1286)
         );
  NOR2_X1 U1081 ( .A1(n1285), .A2(n1286), .ZN(n673) );
  AOI22_X1 U1297 ( .A1(n760), .A2(\predict_PC[14][16] ), .B1(n2271), .B2(
        \predict_PC[15][16] ), .ZN(n1456) );
  AOI22_X1 U1296 ( .A1(n762), .A2(\predict_PC[12][16] ), .B1(n2269), .B2(
        \predict_PC[13][16] ), .ZN(n1457) );
  AOI22_X1 U1295 ( .A1(n756), .A2(\predict_PC[8][16] ), .B1(n2275), .B2(
        \predict_PC[9][16] ), .ZN(n1458) );
  AOI22_X1 U1294 ( .A1(n758), .A2(\predict_PC[10][16] ), .B1(n2273), .B2(
        \predict_PC[11][16] ), .ZN(n1459) );
  NAND4_X1 U1293 ( .A1(n1456), .A2(n1457), .A3(n1458), .A4(n1459), .ZN(n1450)
         );
  AOI22_X1 U1292 ( .A1(n748), .A2(\predict_PC[6][16] ), .B1(n2279), .B2(
        \predict_PC[7][16] ), .ZN(n1452) );
  AOI22_X1 U1291 ( .A1(n750), .A2(\predict_PC[4][16] ), .B1(n2277), .B2(
        \predict_PC[5][16] ), .ZN(n1453) );
  AOI22_X1 U1290 ( .A1(n2284), .A2(\predict_PC[3][16] ), .B1(n2283), .B2(
        \predict_PC[2][16] ), .ZN(n1454) );
  AOI22_X1 U1289 ( .A1(n2282), .A2(\predict_PC[1][16] ), .B1(n747), .B2(
        \predict_PC[0][16] ), .ZN(n1455) );
  NAND4_X1 U1288 ( .A1(n1452), .A2(n1453), .A3(n1454), .A4(n1455), .ZN(n1451)
         );
  NOR2_X1 U1287 ( .A1(n1450), .A2(n1451), .ZN(n686) );
  AOI22_X1 U1311 ( .A1(n760), .A2(\predict_PC[14][15] ), .B1(n2271), .B2(
        \predict_PC[15][15] ), .ZN(n1467) );
  AOI22_X1 U1310 ( .A1(n2270), .A2(\predict_PC[12][15] ), .B1(n2269), .B2(
        \predict_PC[13][15] ), .ZN(n1468) );
  AOI22_X1 U1309 ( .A1(n2276), .A2(\predict_PC[8][15] ), .B1(n2275), .B2(
        \predict_PC[9][15] ), .ZN(n1469) );
  AOI22_X1 U1308 ( .A1(n2274), .A2(\predict_PC[10][15] ), .B1(n2273), .B2(
        \predict_PC[11][15] ), .ZN(n1470) );
  NAND4_X1 U1307 ( .A1(n1467), .A2(n1468), .A3(n1469), .A4(n1470), .ZN(n1461)
         );
  AOI22_X1 U1306 ( .A1(n748), .A2(\predict_PC[6][15] ), .B1(n2279), .B2(
        \predict_PC[7][15] ), .ZN(n1463) );
  AOI22_X1 U1305 ( .A1(n750), .A2(\predict_PC[4][15] ), .B1(n2277), .B2(
        \predict_PC[5][15] ), .ZN(n1464) );
  AOI22_X1 U1304 ( .A1(n2284), .A2(\predict_PC[3][15] ), .B1(n2283), .B2(
        \predict_PC[2][15] ), .ZN(n1465) );
  AOI22_X1 U1303 ( .A1(n2282), .A2(\predict_PC[1][15] ), .B1(n747), .B2(
        \predict_PC[0][15] ), .ZN(n1466) );
  NAND4_X1 U1302 ( .A1(n1463), .A2(n1464), .A3(n1465), .A4(n1466), .ZN(n1462)
         );
  NOR2_X1 U1301 ( .A1(n1461), .A2(n1462), .ZN(n687) );
  AOI22_X1 U1269 ( .A1(n2272), .A2(\predict_PC[14][18] ), .B1(n2271), .B2(
        \predict_PC[15][18] ), .ZN(n1434) );
  AOI22_X1 U1268 ( .A1(n762), .A2(\predict_PC[12][18] ), .B1(n2269), .B2(
        \predict_PC[13][18] ), .ZN(n1435) );
  AOI22_X1 U1267 ( .A1(n756), .A2(\predict_PC[8][18] ), .B1(n2275), .B2(
        \predict_PC[9][18] ), .ZN(n1436) );
  AOI22_X1 U1266 ( .A1(n758), .A2(\predict_PC[10][18] ), .B1(n2273), .B2(
        \predict_PC[11][18] ), .ZN(n1437) );
  NAND4_X1 U1265 ( .A1(n1434), .A2(n1435), .A3(n1436), .A4(n1437), .ZN(n1428)
         );
  AOI22_X1 U1264 ( .A1(n748), .A2(\predict_PC[6][18] ), .B1(n2279), .B2(
        \predict_PC[7][18] ), .ZN(n1430) );
  AOI22_X1 U1263 ( .A1(n2278), .A2(\predict_PC[4][18] ), .B1(n2277), .B2(
        \predict_PC[5][18] ), .ZN(n1431) );
  AOI22_X1 U1262 ( .A1(n2284), .A2(\predict_PC[3][18] ), .B1(n2283), .B2(
        \predict_PC[2][18] ), .ZN(n1432) );
  AOI22_X1 U1261 ( .A1(n2282), .A2(\predict_PC[1][18] ), .B1(n747), .B2(
        \predict_PC[0][18] ), .ZN(n1433) );
  NAND4_X1 U1260 ( .A1(n1430), .A2(n1431), .A3(n1432), .A4(n1433), .ZN(n1429)
         );
  NOR2_X1 U1259 ( .A1(n1428), .A2(n1429), .ZN(n684) );
  AOI22_X1 U1283 ( .A1(n760), .A2(\predict_PC[14][17] ), .B1(n2271), .B2(
        \predict_PC[15][17] ), .ZN(n1445) );
  AOI22_X1 U1282 ( .A1(n762), .A2(\predict_PC[12][17] ), .B1(n2269), .B2(
        \predict_PC[13][17] ), .ZN(n1446) );
  AOI22_X1 U1281 ( .A1(n756), .A2(\predict_PC[8][17] ), .B1(n2275), .B2(
        \predict_PC[9][17] ), .ZN(n1447) );
  AOI22_X1 U1280 ( .A1(n758), .A2(\predict_PC[10][17] ), .B1(n2273), .B2(
        \predict_PC[11][17] ), .ZN(n1448) );
  NAND4_X1 U1279 ( .A1(n1445), .A2(n1446), .A3(n1447), .A4(n1448), .ZN(n1439)
         );
  AOI22_X1 U1278 ( .A1(n2280), .A2(\predict_PC[6][17] ), .B1(n2279), .B2(
        \predict_PC[7][17] ), .ZN(n1441) );
  AOI22_X1 U1277 ( .A1(n750), .A2(\predict_PC[4][17] ), .B1(n2277), .B2(
        \predict_PC[5][17] ), .ZN(n1442) );
  AOI22_X1 U1276 ( .A1(n2284), .A2(\predict_PC[3][17] ), .B1(n2283), .B2(
        \predict_PC[2][17] ), .ZN(n1443) );
  AOI22_X1 U1275 ( .A1(n2282), .A2(\predict_PC[1][17] ), .B1(n747), .B2(
        \predict_PC[0][17] ), .ZN(n1444) );
  NAND4_X1 U1274 ( .A1(n1441), .A2(n1442), .A3(n1443), .A4(n1444), .ZN(n1440)
         );
  NOR2_X1 U1273 ( .A1(n1439), .A2(n1440), .ZN(n685) );
  AOI22_X1 U1185 ( .A1(n2272), .A2(\predict_PC[14][24] ), .B1(n2271), .B2(
        \predict_PC[15][24] ), .ZN(n1368) );
  AOI22_X1 U1184 ( .A1(n2270), .A2(\predict_PC[12][24] ), .B1(n2269), .B2(
        \predict_PC[13][24] ), .ZN(n1369) );
  AOI22_X1 U1183 ( .A1(n2276), .A2(\predict_PC[8][24] ), .B1(n2275), .B2(
        \predict_PC[9][24] ), .ZN(n1370) );
  AOI22_X1 U1182 ( .A1(n2274), .A2(\predict_PC[10][24] ), .B1(n2273), .B2(
        \predict_PC[11][24] ), .ZN(n1371) );
  NAND4_X1 U1181 ( .A1(n1368), .A2(n1369), .A3(n1370), .A4(n1371), .ZN(n1362)
         );
  AOI22_X1 U1180 ( .A1(n2280), .A2(\predict_PC[6][24] ), .B1(n2279), .B2(
        \predict_PC[7][24] ), .ZN(n1364) );
  AOI22_X1 U1179 ( .A1(n2278), .A2(\predict_PC[4][24] ), .B1(n2277), .B2(
        \predict_PC[5][24] ), .ZN(n1365) );
  AOI22_X1 U1178 ( .A1(n2284), .A2(\predict_PC[3][24] ), .B1(n2283), .B2(
        \predict_PC[2][24] ), .ZN(n1366) );
  AOI22_X1 U1177 ( .A1(n2282), .A2(\predict_PC[1][24] ), .B1(n2281), .B2(
        \predict_PC[0][24] ), .ZN(n1367) );
  NAND4_X1 U1176 ( .A1(n1364), .A2(n1365), .A3(n1366), .A4(n1367), .ZN(n1363)
         );
  NOR2_X1 U1175 ( .A1(n1362), .A2(n1363), .ZN(n677) );
  AOI22_X1 U1143 ( .A1(n2272), .A2(\predict_PC[14][27] ), .B1(n2271), .B2(
        \predict_PC[15][27] ), .ZN(n1335) );
  AOI22_X1 U1142 ( .A1(n2270), .A2(\predict_PC[12][27] ), .B1(n2269), .B2(
        \predict_PC[13][27] ), .ZN(n1336) );
  AOI22_X1 U1141 ( .A1(n2276), .A2(\predict_PC[8][27] ), .B1(n2275), .B2(
        \predict_PC[9][27] ), .ZN(n1337) );
  AOI22_X1 U1140 ( .A1(n2274), .A2(\predict_PC[10][27] ), .B1(n2273), .B2(
        \predict_PC[11][27] ), .ZN(n1338) );
  NAND4_X1 U1139 ( .A1(n1335), .A2(n1336), .A3(n1337), .A4(n1338), .ZN(n1329)
         );
  AOI22_X1 U1138 ( .A1(n2280), .A2(\predict_PC[6][27] ), .B1(n2279), .B2(
        \predict_PC[7][27] ), .ZN(n1331) );
  AOI22_X1 U1137 ( .A1(n2278), .A2(\predict_PC[4][27] ), .B1(n2277), .B2(
        \predict_PC[5][27] ), .ZN(n1332) );
  AOI22_X1 U1136 ( .A1(n2284), .A2(\predict_PC[3][27] ), .B1(n2283), .B2(
        \predict_PC[2][27] ), .ZN(n1333) );
  AOI22_X1 U1135 ( .A1(n2282), .A2(\predict_PC[1][27] ), .B1(n2281), .B2(
        \predict_PC[0][27] ), .ZN(n1334) );
  NAND4_X1 U1134 ( .A1(n1331), .A2(n1332), .A3(n1333), .A4(n1334), .ZN(n1330)
         );
  AOI22_X1 U1213 ( .A1(n2272), .A2(\predict_PC[14][22] ), .B1(n2271), .B2(
        \predict_PC[15][22] ), .ZN(n1390) );
  AOI22_X1 U1212 ( .A1(n2270), .A2(\predict_PC[12][22] ), .B1(n2269), .B2(
        \predict_PC[13][22] ), .ZN(n1391) );
  AOI22_X1 U1211 ( .A1(n2276), .A2(\predict_PC[8][22] ), .B1(n2275), .B2(
        \predict_PC[9][22] ), .ZN(n1392) );
  AOI22_X1 U1210 ( .A1(n2274), .A2(\predict_PC[10][22] ), .B1(n2273), .B2(
        \predict_PC[11][22] ), .ZN(n1393) );
  NAND4_X1 U1209 ( .A1(n1390), .A2(n1391), .A3(n1392), .A4(n1393), .ZN(n1384)
         );
  AOI22_X1 U1208 ( .A1(n2280), .A2(\predict_PC[6][22] ), .B1(n2279), .B2(
        \predict_PC[7][22] ), .ZN(n1386) );
  AOI22_X1 U1207 ( .A1(n2278), .A2(\predict_PC[4][22] ), .B1(n2277), .B2(
        \predict_PC[5][22] ), .ZN(n1387) );
  AOI22_X1 U1206 ( .A1(n2284), .A2(\predict_PC[3][22] ), .B1(n2283), .B2(
        \predict_PC[2][22] ), .ZN(n1388) );
  AOI22_X1 U1205 ( .A1(n2282), .A2(\predict_PC[1][22] ), .B1(n2281), .B2(
        \predict_PC[0][22] ), .ZN(n1389) );
  NAND4_X1 U1204 ( .A1(n1386), .A2(n1387), .A3(n1388), .A4(n1389), .ZN(n1385)
         );
  NOR2_X1 U1203 ( .A1(n1384), .A2(n1385), .ZN(n679) );
  AOI22_X1 U1255 ( .A1(n2272), .A2(\predict_PC[14][19] ), .B1(n2271), .B2(
        \predict_PC[15][19] ), .ZN(n1423) );
  AOI22_X1 U1254 ( .A1(n2270), .A2(\predict_PC[12][19] ), .B1(n2269), .B2(
        \predict_PC[13][19] ), .ZN(n1424) );
  AOI22_X1 U1253 ( .A1(n2276), .A2(\predict_PC[8][19] ), .B1(n2275), .B2(
        \predict_PC[9][19] ), .ZN(n1425) );
  AOI22_X1 U1252 ( .A1(n2274), .A2(\predict_PC[10][19] ), .B1(n2273), .B2(
        \predict_PC[11][19] ), .ZN(n1426) );
  NAND4_X1 U1251 ( .A1(n1423), .A2(n1424), .A3(n1425), .A4(n1426), .ZN(n1417)
         );
  AOI22_X1 U1250 ( .A1(n2280), .A2(\predict_PC[6][19] ), .B1(n2279), .B2(
        \predict_PC[7][19] ), .ZN(n1419) );
  AOI22_X1 U1249 ( .A1(n2278), .A2(\predict_PC[4][19] ), .B1(n2277), .B2(
        \predict_PC[5][19] ), .ZN(n1420) );
  AOI22_X1 U1248 ( .A1(n2284), .A2(\predict_PC[3][19] ), .B1(n2283), .B2(
        \predict_PC[2][19] ), .ZN(n1421) );
  AOI22_X1 U1247 ( .A1(n2282), .A2(\predict_PC[1][19] ), .B1(n2281), .B2(
        \predict_PC[0][19] ), .ZN(n1422) );
  NAND4_X1 U1246 ( .A1(n1419), .A2(n1420), .A3(n1421), .A4(n1422), .ZN(n1418)
         );
  NOR2_X1 U1245 ( .A1(n1417), .A2(n1418), .ZN(n683) );
  AOI22_X1 U1199 ( .A1(n2272), .A2(\predict_PC[14][23] ), .B1(n2271), .B2(
        \predict_PC[15][23] ), .ZN(n1379) );
  AOI22_X1 U1198 ( .A1(n2270), .A2(\predict_PC[12][23] ), .B1(n2269), .B2(
        \predict_PC[13][23] ), .ZN(n1380) );
  AOI22_X1 U1197 ( .A1(n2276), .A2(\predict_PC[8][23] ), .B1(n2275), .B2(
        \predict_PC[9][23] ), .ZN(n1381) );
  AOI22_X1 U1196 ( .A1(n2274), .A2(\predict_PC[10][23] ), .B1(n2273), .B2(
        \predict_PC[11][23] ), .ZN(n1382) );
  NAND4_X1 U1195 ( .A1(n1379), .A2(n1380), .A3(n1381), .A4(n1382), .ZN(n1373)
         );
  AOI22_X1 U1194 ( .A1(n2280), .A2(\predict_PC[6][23] ), .B1(n2279), .B2(
        \predict_PC[7][23] ), .ZN(n1375) );
  AOI22_X1 U1193 ( .A1(n2278), .A2(\predict_PC[4][23] ), .B1(n2277), .B2(
        \predict_PC[5][23] ), .ZN(n1376) );
  AOI22_X1 U1192 ( .A1(n2284), .A2(\predict_PC[3][23] ), .B1(n2283), .B2(
        \predict_PC[2][23] ), .ZN(n1377) );
  AOI22_X1 U1191 ( .A1(n2282), .A2(\predict_PC[1][23] ), .B1(n2281), .B2(
        \predict_PC[0][23] ), .ZN(n1378) );
  NAND4_X1 U1190 ( .A1(n1375), .A2(n1376), .A3(n1377), .A4(n1378), .ZN(n1374)
         );
  NOR2_X1 U1189 ( .A1(n1373), .A2(n1374), .ZN(n678) );
  AOI22_X1 U1171 ( .A1(n2272), .A2(\predict_PC[14][25] ), .B1(n2271), .B2(
        \predict_PC[15][25] ), .ZN(n1357) );
  AOI22_X1 U1170 ( .A1(n2270), .A2(\predict_PC[12][25] ), .B1(n2269), .B2(
        \predict_PC[13][25] ), .ZN(n1358) );
  AOI22_X1 U1169 ( .A1(n2276), .A2(\predict_PC[8][25] ), .B1(n2275), .B2(
        \predict_PC[9][25] ), .ZN(n1359) );
  AOI22_X1 U1168 ( .A1(n2274), .A2(\predict_PC[10][25] ), .B1(n2273), .B2(
        \predict_PC[11][25] ), .ZN(n1360) );
  NAND4_X1 U1167 ( .A1(n1357), .A2(n1358), .A3(n1359), .A4(n1360), .ZN(n1351)
         );
  AOI22_X1 U1166 ( .A1(n2280), .A2(\predict_PC[6][25] ), .B1(n2279), .B2(
        \predict_PC[7][25] ), .ZN(n1353) );
  AOI22_X1 U1165 ( .A1(n2278), .A2(\predict_PC[4][25] ), .B1(n2277), .B2(
        \predict_PC[5][25] ), .ZN(n1354) );
  AOI22_X1 U1164 ( .A1(n2284), .A2(\predict_PC[3][25] ), .B1(n2283), .B2(
        \predict_PC[2][25] ), .ZN(n1355) );
  AOI22_X1 U1163 ( .A1(n2282), .A2(\predict_PC[1][25] ), .B1(n2281), .B2(
        \predict_PC[0][25] ), .ZN(n1356) );
  NAND4_X1 U1162 ( .A1(n1353), .A2(n1354), .A3(n1355), .A4(n1356), .ZN(n1352)
         );
  NOR2_X1 U1161 ( .A1(n1351), .A2(n1352), .ZN(n676) );
  AOI22_X1 U1157 ( .A1(n2272), .A2(\predict_PC[14][26] ), .B1(n2271), .B2(
        \predict_PC[15][26] ), .ZN(n1346) );
  AOI22_X1 U1156 ( .A1(n2270), .A2(\predict_PC[12][26] ), .B1(n2269), .B2(
        \predict_PC[13][26] ), .ZN(n1347) );
  AOI22_X1 U1155 ( .A1(n2276), .A2(\predict_PC[8][26] ), .B1(n2275), .B2(
        \predict_PC[9][26] ), .ZN(n1348) );
  AOI22_X1 U1154 ( .A1(n2274), .A2(\predict_PC[10][26] ), .B1(n2273), .B2(
        \predict_PC[11][26] ), .ZN(n1349) );
  NAND4_X1 U1153 ( .A1(n1346), .A2(n1347), .A3(n1348), .A4(n1349), .ZN(n1340)
         );
  AOI22_X1 U1152 ( .A1(n2280), .A2(\predict_PC[6][26] ), .B1(n2279), .B2(
        \predict_PC[7][26] ), .ZN(n1342) );
  AOI22_X1 U1151 ( .A1(n2278), .A2(\predict_PC[4][26] ), .B1(n2277), .B2(
        \predict_PC[5][26] ), .ZN(n1343) );
  AOI22_X1 U1150 ( .A1(n2284), .A2(\predict_PC[3][26] ), .B1(n2283), .B2(
        \predict_PC[2][26] ), .ZN(n1344) );
  AOI22_X1 U1149 ( .A1(n2282), .A2(\predict_PC[1][26] ), .B1(n2281), .B2(
        \predict_PC[0][26] ), .ZN(n1345) );
  NAND4_X1 U1148 ( .A1(n1342), .A2(n1343), .A3(n1344), .A4(n1345), .ZN(n1341)
         );
  NOR2_X1 U1147 ( .A1(n1340), .A2(n1341), .ZN(n675) );
  AOI22_X1 U1423 ( .A1(n760), .A2(\predict_PC[14][7] ), .B1(n2271), .B2(
        \predict_PC[15][7] ), .ZN(n2121) );
  AOI22_X1 U1422 ( .A1(n762), .A2(\predict_PC[12][7] ), .B1(n2269), .B2(
        \predict_PC[13][7] ), .ZN(n2122) );
  AOI22_X1 U1421 ( .A1(n756), .A2(\predict_PC[8][7] ), .B1(n2275), .B2(
        \predict_PC[9][7] ), .ZN(n2123) );
  AOI22_X1 U1420 ( .A1(n758), .A2(\predict_PC[10][7] ), .B1(n2273), .B2(
        \predict_PC[11][7] ), .ZN(n2124) );
  NAND4_X1 U1419 ( .A1(n2121), .A2(n2122), .A3(n2123), .A4(n2124), .ZN(n2115)
         );
  AOI22_X1 U1418 ( .A1(n748), .A2(\predict_PC[6][7] ), .B1(n2279), .B2(
        \predict_PC[7][7] ), .ZN(n2117) );
  AOI22_X1 U1417 ( .A1(n750), .A2(\predict_PC[4][7] ), .B1(n2277), .B2(
        \predict_PC[5][7] ), .ZN(n2118) );
  AOI22_X1 U1416 ( .A1(n2284), .A2(\predict_PC[3][7] ), .B1(n2283), .B2(
        \predict_PC[2][7] ), .ZN(n2119) );
  AOI22_X1 U1415 ( .A1(n2282), .A2(\predict_PC[1][7] ), .B1(n747), .B2(
        \predict_PC[0][7] ), .ZN(n2120) );
  NAND4_X1 U1414 ( .A1(n2117), .A2(n2118), .A3(n2119), .A4(n2120), .ZN(n2116)
         );
  NOR2_X1 U1413 ( .A1(n2115), .A2(n2116), .ZN(n668) );
  AOI22_X1 U1479 ( .A1(n2272), .A2(\predict_PC[14][3] ), .B1(n2271), .B2(
        \predict_PC[15][3] ), .ZN(n2165) );
  AOI22_X1 U1478 ( .A1(n2270), .A2(\predict_PC[12][3] ), .B1(n2269), .B2(
        \predict_PC[13][3] ), .ZN(n2166) );
  AOI22_X1 U1477 ( .A1(n2276), .A2(\predict_PC[8][3] ), .B1(n2275), .B2(
        \predict_PC[9][3] ), .ZN(n2167) );
  AOI22_X1 U1476 ( .A1(n2274), .A2(\predict_PC[10][3] ), .B1(n2273), .B2(
        \predict_PC[11][3] ), .ZN(n2168) );
  NAND4_X1 U1475 ( .A1(n2165), .A2(n2166), .A3(n2167), .A4(n2168), .ZN(n2159)
         );
  AOI22_X1 U1474 ( .A1(n2280), .A2(\predict_PC[6][3] ), .B1(n2279), .B2(
        \predict_PC[7][3] ), .ZN(n2161) );
  AOI22_X1 U1473 ( .A1(n2278), .A2(\predict_PC[4][3] ), .B1(n2277), .B2(
        \predict_PC[5][3] ), .ZN(n2162) );
  AOI22_X1 U1472 ( .A1(n2284), .A2(\predict_PC[3][3] ), .B1(n2283), .B2(
        \predict_PC[2][3] ), .ZN(n2163) );
  AOI22_X1 U1471 ( .A1(n2282), .A2(\predict_PC[1][3] ), .B1(n2281), .B2(
        \predict_PC[0][3] ), .ZN(n2164) );
  NAND4_X1 U1470 ( .A1(n2161), .A2(n2162), .A3(n2163), .A4(n2164), .ZN(n2160)
         );
  NOR2_X1 U1469 ( .A1(n2159), .A2(n2160), .ZN(n672) );
  AOI22_X1 U1227 ( .A1(n2272), .A2(\predict_PC[14][21] ), .B1(n2271), .B2(
        \predict_PC[15][21] ), .ZN(n1401) );
  AOI22_X1 U1226 ( .A1(n2270), .A2(\predict_PC[12][21] ), .B1(n2269), .B2(
        \predict_PC[13][21] ), .ZN(n1402) );
  AOI22_X1 U1225 ( .A1(n2276), .A2(\predict_PC[8][21] ), .B1(n2275), .B2(
        \predict_PC[9][21] ), .ZN(n1403) );
  AOI22_X1 U1224 ( .A1(n2274), .A2(\predict_PC[10][21] ), .B1(n2273), .B2(
        \predict_PC[11][21] ), .ZN(n1404) );
  NAND4_X1 U1223 ( .A1(n1401), .A2(n1402), .A3(n1403), .A4(n1404), .ZN(n1395)
         );
  AOI22_X1 U1222 ( .A1(n2280), .A2(\predict_PC[6][21] ), .B1(n2279), .B2(
        \predict_PC[7][21] ), .ZN(n1397) );
  AOI22_X1 U1221 ( .A1(n2278), .A2(\predict_PC[4][21] ), .B1(n2277), .B2(
        \predict_PC[5][21] ), .ZN(n1398) );
  AOI22_X1 U1220 ( .A1(n2284), .A2(\predict_PC[3][21] ), .B1(n2283), .B2(
        \predict_PC[2][21] ), .ZN(n1399) );
  AOI22_X1 U1219 ( .A1(n2282), .A2(\predict_PC[1][21] ), .B1(n2281), .B2(
        \predict_PC[0][21] ), .ZN(n1400) );
  NAND4_X1 U1218 ( .A1(n1397), .A2(n1398), .A3(n1399), .A4(n1400), .ZN(n1396)
         );
  NOR2_X1 U1217 ( .A1(n1395), .A2(n1396), .ZN(n680) );
  AOI22_X1 U1241 ( .A1(n2272), .A2(\predict_PC[14][20] ), .B1(n2271), .B2(
        \predict_PC[15][20] ), .ZN(n1412) );
  AOI22_X1 U1240 ( .A1(n2270), .A2(\predict_PC[12][20] ), .B1(n2269), .B2(
        \predict_PC[13][20] ), .ZN(n1413) );
  AOI22_X1 U1239 ( .A1(n2276), .A2(\predict_PC[8][20] ), .B1(n2275), .B2(
        \predict_PC[9][20] ), .ZN(n1414) );
  AOI22_X1 U1238 ( .A1(n2274), .A2(\predict_PC[10][20] ), .B1(n2273), .B2(
        \predict_PC[11][20] ), .ZN(n1415) );
  NAND4_X1 U1237 ( .A1(n1412), .A2(n1413), .A3(n1414), .A4(n1415), .ZN(n1406)
         );
  AOI22_X1 U1236 ( .A1(n2280), .A2(\predict_PC[6][20] ), .B1(n2279), .B2(
        \predict_PC[7][20] ), .ZN(n1408) );
  AOI22_X1 U1235 ( .A1(n2278), .A2(\predict_PC[4][20] ), .B1(n2277), .B2(
        \predict_PC[5][20] ), .ZN(n1409) );
  AOI22_X1 U1234 ( .A1(n2284), .A2(\predict_PC[3][20] ), .B1(n2283), .B2(
        \predict_PC[2][20] ), .ZN(n1410) );
  AOI22_X1 U1233 ( .A1(n2282), .A2(\predict_PC[1][20] ), .B1(n2281), .B2(
        \predict_PC[0][20] ), .ZN(n1411) );
  NAND4_X1 U1232 ( .A1(n1408), .A2(n1409), .A3(n1410), .A4(n1411), .ZN(n1407)
         );
  NOR2_X1 U1231 ( .A1(n1406), .A2(n1407), .ZN(n681) );
  AOI22_X1 U1437 ( .A1(n2272), .A2(\predict_PC[14][6] ), .B1(n2271), .B2(
        \predict_PC[15][6] ), .ZN(n2132) );
  AOI22_X1 U1436 ( .A1(n2270), .A2(\predict_PC[12][6] ), .B1(n2269), .B2(
        \predict_PC[13][6] ), .ZN(n2133) );
  AOI22_X1 U1435 ( .A1(n2276), .A2(\predict_PC[8][6] ), .B1(n2275), .B2(
        \predict_PC[9][6] ), .ZN(n2134) );
  AOI22_X1 U1434 ( .A1(n2274), .A2(\predict_PC[10][6] ), .B1(n2273), .B2(
        \predict_PC[11][6] ), .ZN(n2135) );
  NAND4_X1 U1433 ( .A1(n2132), .A2(n2133), .A3(n2134), .A4(n2135), .ZN(n2126)
         );
  AOI22_X1 U1432 ( .A1(n2280), .A2(\predict_PC[6][6] ), .B1(n2279), .B2(
        \predict_PC[7][6] ), .ZN(n2128) );
  AOI22_X1 U1431 ( .A1(n2278), .A2(\predict_PC[4][6] ), .B1(n2277), .B2(
        \predict_PC[5][6] ), .ZN(n2129) );
  AOI22_X1 U1430 ( .A1(n2284), .A2(\predict_PC[3][6] ), .B1(n2283), .B2(
        \predict_PC[2][6] ), .ZN(n2130) );
  AOI22_X1 U1429 ( .A1(n2282), .A2(\predict_PC[1][6] ), .B1(n2281), .B2(
        \predict_PC[0][6] ), .ZN(n2131) );
  NAND4_X1 U1428 ( .A1(n2128), .A2(n2129), .A3(n2130), .A4(n2131), .ZN(n2127)
         );
  NOR2_X1 U1427 ( .A1(n2126), .A2(n2127), .ZN(n669) );
  AOI22_X1 U1409 ( .A1(n2272), .A2(\predict_PC[14][8] ), .B1(n2271), .B2(
        \predict_PC[15][8] ), .ZN(n2110) );
  AOI22_X1 U1408 ( .A1(n2270), .A2(\predict_PC[12][8] ), .B1(n2269), .B2(
        \predict_PC[13][8] ), .ZN(n2111) );
  AOI22_X1 U1407 ( .A1(n2276), .A2(\predict_PC[8][8] ), .B1(n2275), .B2(
        \predict_PC[9][8] ), .ZN(n2112) );
  AOI22_X1 U1406 ( .A1(n2274), .A2(\predict_PC[10][8] ), .B1(n2273), .B2(
        \predict_PC[11][8] ), .ZN(n2113) );
  NAND4_X1 U1405 ( .A1(n2110), .A2(n2111), .A3(n2112), .A4(n2113), .ZN(n2104)
         );
  AOI22_X1 U1404 ( .A1(n2280), .A2(\predict_PC[6][8] ), .B1(n2279), .B2(
        \predict_PC[7][8] ), .ZN(n2106) );
  AOI22_X1 U1403 ( .A1(n2278), .A2(\predict_PC[4][8] ), .B1(n2277), .B2(
        \predict_PC[5][8] ), .ZN(n2107) );
  AOI22_X1 U1402 ( .A1(n2284), .A2(\predict_PC[3][8] ), .B1(n2283), .B2(
        \predict_PC[2][8] ), .ZN(n2108) );
  AOI22_X1 U1401 ( .A1(n2282), .A2(\predict_PC[1][8] ), .B1(n2281), .B2(
        \predict_PC[0][8] ), .ZN(n2109) );
  NAND4_X1 U1400 ( .A1(n2106), .A2(n2107), .A3(n2108), .A4(n2109), .ZN(n2105)
         );
  NOR2_X1 U1399 ( .A1(n2104), .A2(n2105), .ZN(n667) );
  AOI22_X1 U1395 ( .A1(n760), .A2(\predict_PC[14][9] ), .B1(n2271), .B2(
        \predict_PC[15][9] ), .ZN(n1533) );
  AOI22_X1 U1394 ( .A1(n762), .A2(\predict_PC[12][9] ), .B1(n2269), .B2(
        \predict_PC[13][9] ), .ZN(n1534) );
  AOI22_X1 U1393 ( .A1(n756), .A2(\predict_PC[8][9] ), .B1(n2275), .B2(
        \predict_PC[9][9] ), .ZN(n2101) );
  AOI22_X1 U1392 ( .A1(n758), .A2(\predict_PC[10][9] ), .B1(n2273), .B2(
        \predict_PC[11][9] ), .ZN(n2102) );
  NAND4_X1 U1391 ( .A1(n1533), .A2(n1534), .A3(n2101), .A4(n2102), .ZN(n1527)
         );
  AOI22_X1 U1390 ( .A1(n748), .A2(\predict_PC[6][9] ), .B1(n2279), .B2(
        \predict_PC[7][9] ), .ZN(n1529) );
  AOI22_X1 U1389 ( .A1(n750), .A2(\predict_PC[4][9] ), .B1(n2277), .B2(
        \predict_PC[5][9] ), .ZN(n1530) );
  AOI22_X1 U1388 ( .A1(n2284), .A2(\predict_PC[3][9] ), .B1(n2283), .B2(
        \predict_PC[2][9] ), .ZN(n1531) );
  AOI22_X1 U1387 ( .A1(n2282), .A2(\predict_PC[1][9] ), .B1(n747), .B2(
        \predict_PC[0][9] ), .ZN(n1532) );
  NAND4_X1 U1386 ( .A1(n1529), .A2(n1530), .A3(n1531), .A4(n1532), .ZN(n1528)
         );
  NOR2_X1 U1385 ( .A1(n1527), .A2(n1528), .ZN(n666) );
  AOI22_X1 U1493 ( .A1(n2272), .A2(\predict_PC[14][2] ), .B1(n2271), .B2(
        \predict_PC[15][2] ), .ZN(n2176) );
  AOI22_X1 U1492 ( .A1(n2270), .A2(\predict_PC[12][2] ), .B1(n2269), .B2(
        \predict_PC[13][2] ), .ZN(n2177) );
  AOI22_X1 U1491 ( .A1(n2276), .A2(\predict_PC[8][2] ), .B1(n2275), .B2(
        \predict_PC[9][2] ), .ZN(n2178) );
  AOI22_X1 U1490 ( .A1(n2274), .A2(\predict_PC[10][2] ), .B1(n2273), .B2(
        \predict_PC[11][2] ), .ZN(n2179) );
  NAND4_X1 U1489 ( .A1(n2176), .A2(n2177), .A3(n2178), .A4(n2179), .ZN(n2170)
         );
  AOI22_X1 U1488 ( .A1(n2280), .A2(\predict_PC[6][2] ), .B1(n2279), .B2(
        \predict_PC[7][2] ), .ZN(n2172) );
  AOI22_X1 U1487 ( .A1(n2278), .A2(\predict_PC[4][2] ), .B1(n2277), .B2(
        \predict_PC[5][2] ), .ZN(n2173) );
  AOI22_X1 U1486 ( .A1(n2284), .A2(\predict_PC[3][2] ), .B1(n2283), .B2(
        \predict_PC[2][2] ), .ZN(n2174) );
  AOI22_X1 U1485 ( .A1(n2282), .A2(\predict_PC[1][2] ), .B1(n2281), .B2(
        \predict_PC[0][2] ), .ZN(n2175) );
  NAND4_X1 U1484 ( .A1(n2172), .A2(n2173), .A3(n2174), .A4(n2175), .ZN(n2171)
         );
  NOR2_X1 U1483 ( .A1(n2170), .A2(n2171), .ZN(n674) );
  AOI22_X1 U1465 ( .A1(n2272), .A2(\predict_PC[14][4] ), .B1(n2271), .B2(
        \predict_PC[15][4] ), .ZN(n2154) );
  AOI22_X1 U1464 ( .A1(n2270), .A2(\predict_PC[12][4] ), .B1(n2269), .B2(
        \predict_PC[13][4] ), .ZN(n2155) );
  AOI22_X1 U1463 ( .A1(n2276), .A2(\predict_PC[8][4] ), .B1(n2275), .B2(
        \predict_PC[9][4] ), .ZN(n2156) );
  AOI22_X1 U1462 ( .A1(n2274), .A2(\predict_PC[10][4] ), .B1(n2273), .B2(
        \predict_PC[11][4] ), .ZN(n2157) );
  NAND4_X1 U1461 ( .A1(n2154), .A2(n2155), .A3(n2156), .A4(n2157), .ZN(n2148)
         );
  AOI22_X1 U1460 ( .A1(n2280), .A2(\predict_PC[6][4] ), .B1(n2279), .B2(
        \predict_PC[7][4] ), .ZN(n2150) );
  AOI22_X1 U1459 ( .A1(n2278), .A2(\predict_PC[4][4] ), .B1(n2277), .B2(
        \predict_PC[5][4] ), .ZN(n2151) );
  AOI22_X1 U1458 ( .A1(n2284), .A2(\predict_PC[3][4] ), .B1(n2283), .B2(
        \predict_PC[2][4] ), .ZN(n2152) );
  AOI22_X1 U1457 ( .A1(n2282), .A2(\predict_PC[1][4] ), .B1(n2281), .B2(
        \predict_PC[0][4] ), .ZN(n2153) );
  NAND4_X1 U1456 ( .A1(n2150), .A2(n2151), .A3(n2152), .A4(n2153), .ZN(n2149)
         );
  NOR2_X1 U1455 ( .A1(n2148), .A2(n2149), .ZN(n671) );
  AOI22_X1 U1117 ( .A1(n2272), .A2(\predict_PC[14][29] ), .B1(n761), .B2(
        \predict_PC[15][29] ), .ZN(n1313) );
  AOI22_X1 U1116 ( .A1(n2270), .A2(\predict_PC[12][29] ), .B1(n2269), .B2(
        \predict_PC[13][29] ), .ZN(n1314) );
  AOI22_X1 U1115 ( .A1(n2276), .A2(\predict_PC[8][29] ), .B1(n2275), .B2(
        \predict_PC[9][29] ), .ZN(n1315) );
  AOI22_X1 U1114 ( .A1(n2274), .A2(\predict_PC[10][29] ), .B1(n2273), .B2(
        \predict_PC[11][29] ), .ZN(n1316) );
  NAND4_X1 U1113 ( .A1(n1313), .A2(n1314), .A3(n1315), .A4(n1316), .ZN(n1307)
         );
  AOI22_X1 U1112 ( .A1(n2280), .A2(\predict_PC[6][29] ), .B1(n2279), .B2(
        \predict_PC[7][29] ), .ZN(n1309) );
  AOI22_X1 U1111 ( .A1(n2278), .A2(\predict_PC[4][29] ), .B1(n2277), .B2(
        \predict_PC[5][29] ), .ZN(n1310) );
  AOI22_X1 U1110 ( .A1(n2284), .A2(\predict_PC[3][29] ), .B1(n2283), .B2(
        \predict_PC[2][29] ), .ZN(n1311) );
  AOI22_X1 U1109 ( .A1(n2282), .A2(\predict_PC[1][29] ), .B1(n2281), .B2(
        \predict_PC[0][29] ), .ZN(n1312) );
  NAND4_X1 U1108 ( .A1(n1309), .A2(n1310), .A3(n1311), .A4(n1312), .ZN(n1308)
         );
  AOI22_X1 U1451 ( .A1(n760), .A2(\predict_PC[14][5] ), .B1(n2271), .B2(
        \predict_PC[15][5] ), .ZN(n2143) );
  AOI22_X1 U1450 ( .A1(n762), .A2(\predict_PC[12][5] ), .B1(n2269), .B2(
        \predict_PC[13][5] ), .ZN(n2144) );
  AOI22_X1 U1449 ( .A1(n756), .A2(\predict_PC[8][5] ), .B1(n2275), .B2(
        \predict_PC[9][5] ), .ZN(n2145) );
  AOI22_X1 U1448 ( .A1(n758), .A2(\predict_PC[10][5] ), .B1(n2273), .B2(
        \predict_PC[11][5] ), .ZN(n2146) );
  NAND4_X1 U1447 ( .A1(n2143), .A2(n2144), .A3(n2145), .A4(n2146), .ZN(n2137)
         );
  AOI22_X1 U1446 ( .A1(n748), .A2(\predict_PC[6][5] ), .B1(n2279), .B2(
        \predict_PC[7][5] ), .ZN(n2139) );
  AOI22_X1 U1445 ( .A1(n750), .A2(\predict_PC[4][5] ), .B1(n2277), .B2(
        \predict_PC[5][5] ), .ZN(n2140) );
  AOI22_X1 U1444 ( .A1(n2284), .A2(\predict_PC[3][5] ), .B1(n2283), .B2(
        \predict_PC[2][5] ), .ZN(n2141) );
  AOI22_X1 U1443 ( .A1(n2282), .A2(\predict_PC[1][5] ), .B1(n747), .B2(
        \predict_PC[0][5] ), .ZN(n2142) );
  NAND4_X1 U1442 ( .A1(n2139), .A2(n2140), .A3(n2141), .A4(n2142), .ZN(n2138)
         );
  NOR2_X1 U1441 ( .A1(n2137), .A2(n2138), .ZN(n670) );
  AOI22_X1 U1130 ( .A1(n2272), .A2(\predict_PC[14][28] ), .B1(n761), .B2(
        \predict_PC[15][28] ), .ZN(n1324) );
  AOI22_X1 U1129 ( .A1(n2270), .A2(\predict_PC[12][28] ), .B1(n2269), .B2(
        \predict_PC[13][28] ), .ZN(n1325) );
  AOI22_X1 U1128 ( .A1(n2276), .A2(\predict_PC[8][28] ), .B1(n2275), .B2(
        \predict_PC[9][28] ), .ZN(n1326) );
  AOI22_X1 U1127 ( .A1(n2274), .A2(\predict_PC[10][28] ), .B1(n2273), .B2(
        \predict_PC[11][28] ), .ZN(n1327) );
  NAND4_X1 U1126 ( .A1(n1324), .A2(n1325), .A3(n1326), .A4(n1327), .ZN(n1318)
         );
  AOI22_X1 U1125 ( .A1(n2280), .A2(\predict_PC[6][28] ), .B1(n2279), .B2(
        \predict_PC[7][28] ), .ZN(n1320) );
  AOI22_X1 U1124 ( .A1(n2278), .A2(\predict_PC[4][28] ), .B1(n2277), .B2(
        \predict_PC[5][28] ), .ZN(n1321) );
  AOI22_X1 U1123 ( .A1(n2284), .A2(\predict_PC[3][28] ), .B1(n2283), .B2(
        \predict_PC[2][28] ), .ZN(n1322) );
  AOI22_X1 U1122 ( .A1(n2282), .A2(\predict_PC[1][28] ), .B1(n2281), .B2(
        \predict_PC[0][28] ), .ZN(n1323) );
  NAND4_X1 U1121 ( .A1(n1320), .A2(n1321), .A3(n1322), .A4(n1323), .ZN(n1319)
         );
  AOI22_X1 U1546 ( .A1(n2272), .A2(\predict_PC[14][0] ), .B1(n2271), .B2(
        \predict_PC[15][0] ), .ZN(n2204) );
  AOI22_X1 U1540 ( .A1(n2270), .A2(\predict_PC[12][0] ), .B1(n2269), .B2(
        \predict_PC[13][0] ), .ZN(n2205) );
  AOI22_X1 U1535 ( .A1(n2276), .A2(\predict_PC[8][0] ), .B1(n2275), .B2(
        \predict_PC[9][0] ), .ZN(n2206) );
  AOI22_X1 U1532 ( .A1(n2274), .A2(\predict_PC[10][0] ), .B1(n2273), .B2(
        \predict_PC[11][0] ), .ZN(n2207) );
  NAND4_X1 U1531 ( .A1(n2204), .A2(n2205), .A3(n2206), .A4(n2207), .ZN(n2192)
         );
  AOI22_X1 U1526 ( .A1(n2280), .A2(\predict_PC[6][0] ), .B1(n2279), .B2(
        \predict_PC[7][0] ), .ZN(n2194) );
  AOI22_X1 U1523 ( .A1(n2278), .A2(\predict_PC[4][0] ), .B1(n2277), .B2(
        \predict_PC[5][0] ), .ZN(n2195) );
  AOI22_X1 U1519 ( .A1(n2284), .A2(\predict_PC[3][0] ), .B1(n2283), .B2(
        \predict_PC[2][0] ), .ZN(n2196) );
  AOI22_X1 U1516 ( .A1(n2282), .A2(\predict_PC[1][0] ), .B1(n2281), .B2(
        \predict_PC[0][0] ), .ZN(n2197) );
  NAND4_X1 U1515 ( .A1(n2194), .A2(n2195), .A3(n2196), .A4(n2197), .ZN(n2193)
         );
  NOR2_X1 U1514 ( .A1(n2192), .A2(n2193), .ZN(n693) );
  AOI22_X1 U1507 ( .A1(n2272), .A2(\predict_PC[14][1] ), .B1(n2271), .B2(
        \predict_PC[15][1] ), .ZN(n2187) );
  AOI22_X1 U1506 ( .A1(n2270), .A2(\predict_PC[12][1] ), .B1(n2269), .B2(
        \predict_PC[13][1] ), .ZN(n2188) );
  AOI22_X1 U1505 ( .A1(n2276), .A2(\predict_PC[8][1] ), .B1(n2275), .B2(
        \predict_PC[9][1] ), .ZN(n2189) );
  AOI22_X1 U1504 ( .A1(n2274), .A2(\predict_PC[10][1] ), .B1(n2273), .B2(
        \predict_PC[11][1] ), .ZN(n2190) );
  NAND4_X1 U1503 ( .A1(n2187), .A2(n2188), .A3(n2189), .A4(n2190), .ZN(n2181)
         );
  AOI22_X1 U1502 ( .A1(n2280), .A2(\predict_PC[6][1] ), .B1(n2279), .B2(
        \predict_PC[7][1] ), .ZN(n2183) );
  AOI22_X1 U1501 ( .A1(n2278), .A2(\predict_PC[4][1] ), .B1(n2277), .B2(
        \predict_PC[5][1] ), .ZN(n2184) );
  AOI22_X1 U1500 ( .A1(n2284), .A2(\predict_PC[3][1] ), .B1(n2283), .B2(
        \predict_PC[2][1] ), .ZN(n2185) );
  AOI22_X1 U1499 ( .A1(n2282), .A2(\predict_PC[1][1] ), .B1(n2281), .B2(
        \predict_PC[0][1] ), .ZN(n2186) );
  NAND4_X1 U1498 ( .A1(n2183), .A2(n2184), .A3(n2185), .A4(n2186), .ZN(n2182)
         );
  NOR2_X1 U1497 ( .A1(n2181), .A2(n2182), .ZN(n682) );
  AOI22_X1 U1104 ( .A1(n2272), .A2(\predict_PC[14][30] ), .B1(n761), .B2(
        \predict_PC[15][30] ), .ZN(n1302) );
  AOI22_X1 U1103 ( .A1(n2270), .A2(\predict_PC[12][30] ), .B1(n2269), .B2(
        \predict_PC[13][30] ), .ZN(n1303) );
  AOI22_X1 U1102 ( .A1(n2276), .A2(\predict_PC[8][30] ), .B1(n2275), .B2(
        \predict_PC[9][30] ), .ZN(n1304) );
  AOI22_X1 U1101 ( .A1(n2274), .A2(\predict_PC[10][30] ), .B1(n2273), .B2(
        \predict_PC[11][30] ), .ZN(n1305) );
  NAND4_X1 U1100 ( .A1(n1302), .A2(n1303), .A3(n1304), .A4(n1305), .ZN(n1296)
         );
  AOI22_X1 U1099 ( .A1(n2280), .A2(\predict_PC[6][30] ), .B1(n2279), .B2(
        \predict_PC[7][30] ), .ZN(n1298) );
  AOI22_X1 U1098 ( .A1(n2278), .A2(\predict_PC[4][30] ), .B1(n2277), .B2(
        \predict_PC[5][30] ), .ZN(n1299) );
  AOI22_X1 U1097 ( .A1(n2284), .A2(\predict_PC[3][30] ), .B1(n2283), .B2(
        \predict_PC[2][30] ), .ZN(n1300) );
  AOI22_X1 U1096 ( .A1(n2282), .A2(\predict_PC[1][30] ), .B1(n2281), .B2(
        \predict_PC[0][30] ), .ZN(n1301) );
  NAND4_X1 U1095 ( .A1(n1298), .A2(n1299), .A3(n1300), .A4(n1301), .ZN(n1297)
         );
  AOI22_X1 U1339 ( .A1(n2272), .A2(\predict_PC[14][13] ), .B1(n2271), .B2(
        \predict_PC[15][13] ), .ZN(n1489) );
  AOI22_X1 U1338 ( .A1(n2270), .A2(\predict_PC[12][13] ), .B1(n2269), .B2(
        \predict_PC[13][13] ), .ZN(n1490) );
  AOI22_X1 U1337 ( .A1(n2276), .A2(\predict_PC[8][13] ), .B1(n2275), .B2(
        \predict_PC[9][13] ), .ZN(n1491) );
  AOI22_X1 U1336 ( .A1(n2274), .A2(\predict_PC[10][13] ), .B1(n2273), .B2(
        \predict_PC[11][13] ), .ZN(n1492) );
  NAND4_X1 U1335 ( .A1(n1489), .A2(n1490), .A3(n1491), .A4(n1492), .ZN(n1483)
         );
  AOI22_X1 U1334 ( .A1(n2280), .A2(\predict_PC[6][13] ), .B1(n2279), .B2(
        \predict_PC[7][13] ), .ZN(n1485) );
  AOI22_X1 U1333 ( .A1(n2278), .A2(\predict_PC[4][13] ), .B1(n2277), .B2(
        \predict_PC[5][13] ), .ZN(n1486) );
  AOI22_X1 U1332 ( .A1(n2284), .A2(\predict_PC[3][13] ), .B1(n2283), .B2(
        \predict_PC[2][13] ), .ZN(n1487) );
  AOI22_X1 U1331 ( .A1(n2282), .A2(\predict_PC[1][13] ), .B1(n2281), .B2(
        \predict_PC[0][13] ), .ZN(n1488) );
  NAND4_X1 U1330 ( .A1(n1485), .A2(n1486), .A3(n1487), .A4(n1488), .ZN(n1484)
         );
  NOR2_X1 U1329 ( .A1(n1483), .A2(n1484), .ZN(n689) );
  AOI22_X1 U1353 ( .A1(n2272), .A2(\predict_PC[14][12] ), .B1(n2271), .B2(
        \predict_PC[15][12] ), .ZN(n1500) );
  AOI22_X1 U1352 ( .A1(n2270), .A2(\predict_PC[12][12] ), .B1(n2269), .B2(
        \predict_PC[13][12] ), .ZN(n1501) );
  AOI22_X1 U1351 ( .A1(n2276), .A2(\predict_PC[8][12] ), .B1(n2275), .B2(
        \predict_PC[9][12] ), .ZN(n1502) );
  AOI22_X1 U1350 ( .A1(n2274), .A2(\predict_PC[10][12] ), .B1(n2273), .B2(
        \predict_PC[11][12] ), .ZN(n1503) );
  NAND4_X1 U1349 ( .A1(n1500), .A2(n1501), .A3(n1502), .A4(n1503), .ZN(n1494)
         );
  AOI22_X1 U1348 ( .A1(n2280), .A2(\predict_PC[6][12] ), .B1(n2279), .B2(
        \predict_PC[7][12] ), .ZN(n1496) );
  AOI22_X1 U1347 ( .A1(n2278), .A2(\predict_PC[4][12] ), .B1(n2277), .B2(
        \predict_PC[5][12] ), .ZN(n1497) );
  AOI22_X1 U1346 ( .A1(n2284), .A2(\predict_PC[3][12] ), .B1(n2283), .B2(
        \predict_PC[2][12] ), .ZN(n1498) );
  AOI22_X1 U1345 ( .A1(n2282), .A2(\predict_PC[1][12] ), .B1(n2281), .B2(
        \predict_PC[0][12] ), .ZN(n1499) );
  NAND4_X1 U1344 ( .A1(n1496), .A2(n1497), .A3(n1498), .A4(n1499), .ZN(n1495)
         );
  NOR2_X1 U1343 ( .A1(n1494), .A2(n1495), .ZN(n690) );
  AOI22_X1 U1553 ( .A1(stall_i), .A2(n592), .B1(n2210), .B2(n2285), .ZN(n1535)
         );
  OAI22_X1 U1341 ( .A1(n1284), .A2(target_PC_i[12]), .B1(\predict_PC[15][12] ), 
        .B2(n726), .ZN(n1493) );
  OAI22_X1 U1327 ( .A1(n1284), .A2(n651), .B1(\predict_PC[15][13] ), .B2(n726), 
        .ZN(n1482) );
  OAI22_X1 U1243 ( .A1(n1284), .A2(n645), .B1(\predict_PC[15][19] ), .B2(n726), 
        .ZN(n1416) );
  OAI22_X1 U1313 ( .A1(n1284), .A2(n630), .B1(\predict_PC[15][14] ), .B2(n726), 
        .ZN(n1471) );
  OAI22_X1 U1271 ( .A1(n1284), .A2(n631), .B1(\predict_PC[15][17] ), .B2(n726), 
        .ZN(n1438) );
  OAI22_X1 U1215 ( .A1(n1284), .A2(n642), .B1(\predict_PC[15][21] ), .B2(n726), 
        .ZN(n1394) );
  OAI22_X1 U1187 ( .A1(n1284), .A2(n643), .B1(\predict_PC[15][23] ), .B2(n726), 
        .ZN(n1372) );
  OAI22_X1 U1229 ( .A1(n1284), .A2(target_PC_i[20]), .B1(\predict_PC[15][20] ), 
        .B2(n726), .ZN(n1405) );
  OAI22_X1 U1285 ( .A1(n1284), .A2(target_PC_i[16]), .B1(\predict_PC[15][16] ), 
        .B2(n726), .ZN(n1449) );
  OAI22_X1 U1257 ( .A1(n1284), .A2(target_PC_i[18]), .B1(\predict_PC[15][18] ), 
        .B2(n726), .ZN(n1427) );
  OAI22_X1 U1201 ( .A1(n1284), .A2(n632), .B1(\predict_PC[15][22] ), .B2(n726), 
        .ZN(n1383) );
  OAI22_X1 U1299 ( .A1(n1284), .A2(target_PC_i[15]), .B1(\predict_PC[15][15] ), 
        .B2(n726), .ZN(n1460) );
  OAI22_X1 U914 ( .A1(n1184), .A2(n646), .B1(\predict_PC[12][12] ), .B2(n735), 
        .ZN(n1203) );
  OAI22_X1 U979 ( .A1(n1218), .A2(n651), .B1(\predict_PC[13][13] ), .B2(n732), 
        .ZN(n1236) );
  OAI22_X1 U1049 ( .A1(n1251), .A2(n646), .B1(\predict_PC[14][12] ), .B2(n729), 
        .ZN(n1270) );
  OAI22_X1 U1047 ( .A1(n1251), .A2(n651), .B1(\predict_PC[14][13] ), .B2(n729), 
        .ZN(n1269) );
  OAI22_X1 U912 ( .A1(n1184), .A2(n651), .B1(\predict_PC[12][13] ), .B2(n735), 
        .ZN(n1202) );
  OAI22_X1 U981 ( .A1(n1218), .A2(target_PC_i[12]), .B1(\predict_PC[13][12] ), 
        .B2(n732), .ZN(n1237) );
  OAI22_X1 U973 ( .A1(n1218), .A2(n637), .B1(\predict_PC[13][16] ), .B2(n732), 
        .ZN(n1233) );
  OAI22_X1 U1033 ( .A1(n1251), .A2(n638), .B1(\predict_PC[14][20] ), .B2(n729), 
        .ZN(n1262) );
  OAI22_X1 U961 ( .A1(n1218), .A2(n632), .B1(\predict_PC[13][22] ), .B2(n732), 
        .ZN(n1227) );
  OAI22_X1 U1027 ( .A1(n1251), .A2(n643), .B1(\predict_PC[14][23] ), .B2(n729), 
        .ZN(n1259) );
  OAI22_X1 U1031 ( .A1(n1251), .A2(n642), .B1(\predict_PC[14][21] ), .B2(n729), 
        .ZN(n1261) );
  OAI22_X1 U959 ( .A1(n1218), .A2(n643), .B1(\predict_PC[13][23] ), .B2(n732), 
        .ZN(n1226) );
  OAI22_X1 U1039 ( .A1(n1251), .A2(n631), .B1(\predict_PC[14][17] ), .B2(n729), 
        .ZN(n1265) );
  OAI22_X1 U908 ( .A1(n1184), .A2(target_PC_i[15]), .B1(\predict_PC[12][15] ), 
        .B2(n735), .ZN(n1200) );
  OAI22_X1 U906 ( .A1(n1184), .A2(n637), .B1(\predict_PC[12][16] ), .B2(n735), 
        .ZN(n1199) );
  OAI22_X1 U963 ( .A1(n1218), .A2(n642), .B1(\predict_PC[13][21] ), .B2(n732), 
        .ZN(n1228) );
  OAI22_X1 U965 ( .A1(n1218), .A2(n638), .B1(\predict_PC[13][20] ), .B2(n732), 
        .ZN(n1229) );
  OAI22_X1 U898 ( .A1(n1184), .A2(n638), .B1(\predict_PC[12][20] ), .B2(n735), 
        .ZN(n1195) );
  OAI22_X1 U1041 ( .A1(n1251), .A2(n637), .B1(\predict_PC[14][16] ), .B2(n729), 
        .ZN(n1266) );
  OAI22_X1 U975 ( .A1(n1218), .A2(target_PC_i[15]), .B1(\predict_PC[13][15] ), 
        .B2(n732), .ZN(n1234) );
  OAI22_X1 U910 ( .A1(n1184), .A2(n630), .B1(\predict_PC[12][14] ), .B2(n735), 
        .ZN(n1201) );
  OAI22_X1 U904 ( .A1(n1184), .A2(n631), .B1(\predict_PC[12][17] ), .B2(n735), 
        .ZN(n1198) );
  OAI22_X1 U1037 ( .A1(n1251), .A2(target_PC_i[18]), .B1(\predict_PC[14][18] ), 
        .B2(n729), .ZN(n1264) );
  OAI22_X1 U967 ( .A1(n1218), .A2(n645), .B1(\predict_PC[13][19] ), .B2(n732), 
        .ZN(n1230) );
  OAI22_X1 U892 ( .A1(n1184), .A2(n643), .B1(\predict_PC[12][23] ), .B2(n735), 
        .ZN(n1192) );
  OAI22_X1 U902 ( .A1(n1184), .A2(target_PC_i[18]), .B1(\predict_PC[12][18] ), 
        .B2(n735), .ZN(n1197) );
  OAI22_X1 U1045 ( .A1(n1251), .A2(n630), .B1(\predict_PC[14][14] ), .B2(n729), 
        .ZN(n1268) );
  OAI22_X1 U900 ( .A1(n1184), .A2(n645), .B1(\predict_PC[12][19] ), .B2(n735), 
        .ZN(n1196) );
  OAI22_X1 U1035 ( .A1(n1251), .A2(n645), .B1(\predict_PC[14][19] ), .B2(n729), 
        .ZN(n1263) );
  OAI22_X1 U969 ( .A1(n1218), .A2(target_PC_i[18]), .B1(\predict_PC[13][18] ), 
        .B2(n732), .ZN(n1231) );
  OAI22_X1 U1043 ( .A1(n1251), .A2(target_PC_i[15]), .B1(\predict_PC[14][15] ), 
        .B2(n729), .ZN(n1267) );
  OAI22_X1 U971 ( .A1(n1218), .A2(n631), .B1(\predict_PC[13][17] ), .B2(n732), 
        .ZN(n1232) );
  OAI22_X1 U977 ( .A1(n1218), .A2(n630), .B1(\predict_PC[13][14] ), .B2(n732), 
        .ZN(n1235) );
  OAI22_X1 U1029 ( .A1(n1251), .A2(n632), .B1(\predict_PC[14][22] ), .B2(n729), 
        .ZN(n1260) );
  OAI22_X1 U896 ( .A1(n1184), .A2(n642), .B1(\predict_PC[12][21] ), .B2(n735), 
        .ZN(n1194) );
  OAI22_X1 U894 ( .A1(n1184), .A2(n632), .B1(\predict_PC[12][22] ), .B2(n735), 
        .ZN(n1193) );
  OAI22_X1 U384 ( .A1(n902), .A2(n646), .B1(\predict_PC[4][12] ), .B2(n2255), 
        .ZN(n921) );
  OAI22_X1 U382 ( .A1(n902), .A2(n651), .B1(\predict_PC[4][13] ), .B2(n2255), 
        .ZN(n920) );
  OAI22_X1 U845 ( .A1(n1151), .A2(n651), .B1(\predict_PC[11][13] ), .B2(n975), 
        .ZN(n1169) );
  OAI22_X1 U847 ( .A1(n1151), .A2(n646), .B1(\predict_PC[11][12] ), .B2(n975), 
        .ZN(n1170) );
  OAI22_X1 U713 ( .A1(n1085), .A2(target_PC_i[13]), .B1(\predict_PC[9][13] ), 
        .B2(n981), .ZN(n1103) );
  OAI22_X1 U781 ( .A1(n1118), .A2(n646), .B1(\predict_PC[10][12] ), .B2(n978), 
        .ZN(n1137) );
  OAI22_X1 U649 ( .A1(n1051), .A2(n646), .B1(\predict_PC[8][12] ), .B2(n984), 
        .ZN(n1070) );
  OAI22_X1 U448 ( .A1(n936), .A2(n651), .B1(\predict_PC[5][13] ), .B2(n2216), 
        .ZN(n954) );
  OAI22_X1 U514 ( .A1(n969), .A2(n651), .B1(\predict_PC[6][13] ), .B2(n2213), 
        .ZN(n1003) );
  OAI22_X1 U779 ( .A1(n1118), .A2(n651), .B1(\predict_PC[10][13] ), .B2(n978), 
        .ZN(n1136) );
  OAI22_X1 U715 ( .A1(n1085), .A2(n646), .B1(\predict_PC[9][12] ), .B2(n981), 
        .ZN(n1104) );
  OAI22_X1 U450 ( .A1(n936), .A2(target_PC_i[12]), .B1(\predict_PC[5][12] ), 
        .B2(n2216), .ZN(n955) );
  OAI22_X1 U582 ( .A1(n1018), .A2(n646), .B1(\predict_PC[7][12] ), .B2(n987), 
        .ZN(n1037) );
  OAI22_X1 U516 ( .A1(n969), .A2(n646), .B1(\predict_PC[6][12] ), .B2(n2213), 
        .ZN(n1004) );
  OAI22_X1 U580 ( .A1(n1018), .A2(n651), .B1(\predict_PC[7][13] ), .B2(n987), 
        .ZN(n1036) );
  OAI22_X1 U647 ( .A1(n1051), .A2(n651), .B1(\predict_PC[8][13] ), .B2(n984), 
        .ZN(n1069) );
  OAI22_X1 U562 ( .A1(n1018), .A2(n632), .B1(\predict_PC[7][22] ), .B2(n987), 
        .ZN(n1027) );
  OAI22_X1 U366 ( .A1(n902), .A2(n642), .B1(\predict_PC[4][21] ), .B2(n2255), 
        .ZN(n912) );
  OAI22_X1 U370 ( .A1(n902), .A2(n645), .B1(\predict_PC[4][19] ), .B2(n2255), 
        .ZN(n914) );
  OAI22_X1 U372 ( .A1(n902), .A2(target_PC_i[18]), .B1(\predict_PC[4][18] ), 
        .B2(n2255), .ZN(n915) );
  OAI22_X1 U368 ( .A1(n902), .A2(n638), .B1(\predict_PC[4][20] ), .B2(n2255), 
        .ZN(n913) );
  OAI22_X1 U374 ( .A1(n902), .A2(n631), .B1(\predict_PC[4][17] ), .B2(n2255), 
        .ZN(n916) );
  OAI22_X1 U576 ( .A1(n1018), .A2(target_PC_i[15]), .B1(\predict_PC[7][15] ), 
        .B2(n987), .ZN(n1034) );
  OAI22_X1 U578 ( .A1(n1018), .A2(n630), .B1(\predict_PC[7][14] ), .B2(n987), 
        .ZN(n1035) );
  OAI22_X1 U572 ( .A1(n1018), .A2(n631), .B1(\predict_PC[7][17] ), .B2(n987), 
        .ZN(n1032) );
  OAI22_X1 U376 ( .A1(n902), .A2(n637), .B1(\predict_PC[4][16] ), .B2(n2255), 
        .ZN(n917) );
  OAI22_X1 U564 ( .A1(n1018), .A2(n642), .B1(\predict_PC[7][21] ), .B2(n987), 
        .ZN(n1028) );
  OAI22_X1 U627 ( .A1(n1051), .A2(n643), .B1(\predict_PC[8][23] ), .B2(n984), 
        .ZN(n1059) );
  OAI22_X1 U629 ( .A1(n1051), .A2(n632), .B1(\predict_PC[8][22] ), .B2(n984), 
        .ZN(n1060) );
  OAI22_X1 U570 ( .A1(n1018), .A2(target_PC_i[18]), .B1(\predict_PC[7][18] ), 
        .B2(n987), .ZN(n1031) );
  OAI22_X1 U631 ( .A1(n1051), .A2(n642), .B1(\predict_PC[8][21] ), .B2(n984), 
        .ZN(n1061) );
  OAI22_X1 U633 ( .A1(n1051), .A2(n638), .B1(\predict_PC[8][20] ), .B2(n984), 
        .ZN(n1062) );
  OAI22_X1 U635 ( .A1(n1051), .A2(n645), .B1(\predict_PC[8][19] ), .B2(n984), 
        .ZN(n1063) );
  OAI22_X1 U380 ( .A1(n902), .A2(n630), .B1(\predict_PC[4][14] ), .B2(n2255), 
        .ZN(n919) );
  OAI22_X1 U637 ( .A1(n1051), .A2(target_PC_i[18]), .B1(\predict_PC[8][18] ), 
        .B2(n984), .ZN(n1064) );
  OAI22_X1 U639 ( .A1(n1051), .A2(n631), .B1(\predict_PC[8][17] ), .B2(n984), 
        .ZN(n1065) );
  OAI22_X1 U641 ( .A1(n1051), .A2(n637), .B1(\predict_PC[8][16] ), .B2(n984), 
        .ZN(n1066) );
  OAI22_X1 U643 ( .A1(n1051), .A2(target_PC_i[15]), .B1(\predict_PC[8][15] ), 
        .B2(n984), .ZN(n1067) );
  OAI22_X1 U645 ( .A1(n1051), .A2(n630), .B1(\predict_PC[8][14] ), .B2(n984), 
        .ZN(n1068) );
  OAI22_X1 U378 ( .A1(n902), .A2(target_PC_i[15]), .B1(\predict_PC[4][15] ), 
        .B2(n2255), .ZN(n918) );
  OAI22_X1 U364 ( .A1(n902), .A2(n632), .B1(\predict_PC[4][22] ), .B2(n2255), 
        .ZN(n911) );
  OAI22_X1 U560 ( .A1(n1018), .A2(n643), .B1(\predict_PC[7][23] ), .B2(n987), 
        .ZN(n1026) );
  OAI22_X1 U362 ( .A1(n902), .A2(n643), .B1(\predict_PC[4][23] ), .B2(n2255), 
        .ZN(n910) );
  OAI22_X1 U512 ( .A1(n969), .A2(n630), .B1(\predict_PC[6][14] ), .B2(n2213), 
        .ZN(n1002) );
  OAI22_X1 U574 ( .A1(n1018), .A2(n637), .B1(\predict_PC[7][16] ), .B2(n987), 
        .ZN(n1033) );
  OAI22_X1 U510 ( .A1(n969), .A2(target_PC_i[15]), .B1(\predict_PC[6][15] ), 
        .B2(n2213), .ZN(n1001) );
  OAI22_X1 U693 ( .A1(n1085), .A2(n643), .B1(\predict_PC[9][23] ), .B2(n981), 
        .ZN(n1093) );
  OAI22_X1 U508 ( .A1(n969), .A2(n637), .B1(\predict_PC[6][16] ), .B2(n2213), 
        .ZN(n1000) );
  OAI22_X1 U695 ( .A1(n1085), .A2(n632), .B1(\predict_PC[9][22] ), .B2(n981), 
        .ZN(n1094) );
  OAI22_X1 U506 ( .A1(n969), .A2(n631), .B1(\predict_PC[6][17] ), .B2(n2213), 
        .ZN(n999) );
  OAI22_X1 U697 ( .A1(n1085), .A2(n642), .B1(\predict_PC[9][21] ), .B2(n981), 
        .ZN(n1095) );
  OAI22_X1 U504 ( .A1(n969), .A2(target_PC_i[18]), .B1(\predict_PC[6][18] ), 
        .B2(n2213), .ZN(n998) );
  OAI22_X1 U699 ( .A1(n1085), .A2(n638), .B1(\predict_PC[9][20] ), .B2(n981), 
        .ZN(n1096) );
  OAI22_X1 U502 ( .A1(n969), .A2(n645), .B1(\predict_PC[6][19] ), .B2(n2213), 
        .ZN(n997) );
  OAI22_X1 U701 ( .A1(n1085), .A2(n645), .B1(\predict_PC[9][19] ), .B2(n981), 
        .ZN(n1097) );
  OAI22_X1 U500 ( .A1(n969), .A2(n638), .B1(\predict_PC[6][20] ), .B2(n2213), 
        .ZN(n996) );
  OAI22_X1 U703 ( .A1(n1085), .A2(target_PC_i[18]), .B1(\predict_PC[9][18] ), 
        .B2(n981), .ZN(n1098) );
  OAI22_X1 U498 ( .A1(n969), .A2(n642), .B1(\predict_PC[6][21] ), .B2(n2213), 
        .ZN(n995) );
  OAI22_X1 U446 ( .A1(n936), .A2(n630), .B1(\predict_PC[5][14] ), .B2(n2216), 
        .ZN(n953) );
  OAI22_X1 U440 ( .A1(n936), .A2(n631), .B1(\predict_PC[5][17] ), .B2(n2216), 
        .ZN(n950) );
  OAI22_X1 U767 ( .A1(n1118), .A2(n645), .B1(\predict_PC[10][19] ), .B2(n978), 
        .ZN(n1130) );
  OAI22_X1 U442 ( .A1(n936), .A2(n637), .B1(\predict_PC[5][16] ), .B2(n2216), 
        .ZN(n951) );
  OAI22_X1 U839 ( .A1(n1151), .A2(n637), .B1(\predict_PC[11][16] ), .B2(n975), 
        .ZN(n1166) );
  OAI22_X1 U769 ( .A1(n1118), .A2(target_PC_i[18]), .B1(\predict_PC[10][18] ), 
        .B2(n978), .ZN(n1131) );
  OAI22_X1 U432 ( .A1(n936), .A2(n642), .B1(\predict_PC[5][21] ), .B2(n2216), 
        .ZN(n946) );
  OAI22_X1 U705 ( .A1(n1085), .A2(n631), .B1(\predict_PC[9][17] ), .B2(n981), 
        .ZN(n1099) );
  OAI22_X1 U833 ( .A1(n1151), .A2(n645), .B1(\predict_PC[11][19] ), .B2(n975), 
        .ZN(n1163) );
  OAI22_X1 U428 ( .A1(n936), .A2(n643), .B1(\predict_PC[5][23] ), .B2(n2216), 
        .ZN(n944) );
  OAI22_X1 U496 ( .A1(n969), .A2(n632), .B1(\predict_PC[6][22] ), .B2(n2213), 
        .ZN(n994) );
  OAI22_X1 U707 ( .A1(n1085), .A2(n637), .B1(\predict_PC[9][16] ), .B2(n981), 
        .ZN(n1100) );
  OAI22_X1 U494 ( .A1(n969), .A2(n643), .B1(\predict_PC[6][23] ), .B2(n2213), 
        .ZN(n993) );
  OAI22_X1 U430 ( .A1(n936), .A2(target_PC_i[22]), .B1(\predict_PC[5][22] ), 
        .B2(n2216), .ZN(n945) );
  OAI22_X1 U709 ( .A1(n1085), .A2(target_PC_i[15]), .B1(\predict_PC[9][15] ), 
        .B2(n981), .ZN(n1101) );
  OAI22_X1 U711 ( .A1(n1085), .A2(n630), .B1(\predict_PC[9][14] ), .B2(n981), 
        .ZN(n1102) );
  OAI22_X1 U825 ( .A1(n1151), .A2(n643), .B1(\predict_PC[11][23] ), .B2(n975), 
        .ZN(n1159) );
  OAI22_X1 U777 ( .A1(n1118), .A2(target_PC_i[14]), .B1(\predict_PC[10][14] ), 
        .B2(n978), .ZN(n1135) );
  OAI22_X1 U566 ( .A1(n1018), .A2(n638), .B1(\predict_PC[7][20] ), .B2(n987), 
        .ZN(n1029) );
  OAI22_X1 U568 ( .A1(n1018), .A2(n645), .B1(\predict_PC[7][19] ), .B2(n987), 
        .ZN(n1030) );
  OAI22_X1 U759 ( .A1(n1118), .A2(n643), .B1(\predict_PC[10][23] ), .B2(n978), 
        .ZN(n1126) );
  OAI22_X1 U761 ( .A1(n1118), .A2(n632), .B1(\predict_PC[10][22] ), .B2(n978), 
        .ZN(n1127) );
  OAI22_X1 U763 ( .A1(n1118), .A2(n642), .B1(\predict_PC[10][21] ), .B2(n978), 
        .ZN(n1128) );
  OAI22_X1 U843 ( .A1(n1151), .A2(n630), .B1(\predict_PC[11][14] ), .B2(n975), 
        .ZN(n1168) );
  OAI22_X1 U765 ( .A1(n1118), .A2(n638), .B1(\predict_PC[10][20] ), .B2(n978), 
        .ZN(n1129) );
  OAI22_X1 U841 ( .A1(n1151), .A2(target_PC_i[15]), .B1(\predict_PC[11][15] ), 
        .B2(n975), .ZN(n1167) );
  OAI22_X1 U775 ( .A1(n1118), .A2(target_PC_i[15]), .B1(\predict_PC[10][15] ), 
        .B2(n978), .ZN(n1134) );
  OAI22_X1 U438 ( .A1(n936), .A2(target_PC_i[18]), .B1(\predict_PC[5][18] ), 
        .B2(n2216), .ZN(n949) );
  OAI22_X1 U827 ( .A1(n1151), .A2(n632), .B1(\predict_PC[11][22] ), .B2(n975), 
        .ZN(n1160) );
  OAI22_X1 U444 ( .A1(n936), .A2(target_PC_i[15]), .B1(\predict_PC[5][15] ), 
        .B2(n2216), .ZN(n952) );
  OAI22_X1 U773 ( .A1(n1118), .A2(target_PC_i[16]), .B1(\predict_PC[10][16] ), 
        .B2(n978), .ZN(n1133) );
  OAI22_X1 U837 ( .A1(n1151), .A2(target_PC_i[17]), .B1(\predict_PC[11][17] ), 
        .B2(n975), .ZN(n1165) );
  OAI22_X1 U771 ( .A1(n1118), .A2(n631), .B1(\predict_PC[10][17] ), .B2(n978), 
        .ZN(n1132) );
  OAI22_X1 U835 ( .A1(n1151), .A2(target_PC_i[18]), .B1(\predict_PC[11][18] ), 
        .B2(n975), .ZN(n1164) );
  OAI22_X1 U434 ( .A1(n936), .A2(n638), .B1(\predict_PC[5][20] ), .B2(n2216), 
        .ZN(n947) );
  OAI22_X1 U829 ( .A1(n1151), .A2(n642), .B1(\predict_PC[11][21] ), .B2(n975), 
        .ZN(n1161) );
  OAI22_X1 U831 ( .A1(n1151), .A2(target_PC_i[20]), .B1(\predict_PC[11][20] ), 
        .B2(n975), .ZN(n1162) );
  OAI22_X1 U436 ( .A1(n936), .A2(n645), .B1(\predict_PC[5][19] ), .B2(n2216), 
        .ZN(n948) );
  OAI22_X1 U1355 ( .A1(n1284), .A2(n644), .B1(\predict_PC[15][11] ), .B2(n725), 
        .ZN(n1504) );
  OAI22_X1 U1439 ( .A1(n1284), .A2(target_PC_i[5]), .B1(\predict_PC[15][5] ), 
        .B2(n725), .ZN(n2136) );
  OAI22_X1 U1481 ( .A1(n1284), .A2(target_PC_i[2]), .B1(\predict_PC[15][2] ), 
        .B2(n725), .ZN(n2169) );
  OAI22_X1 U1495 ( .A1(n1284), .A2(n633), .B1(\predict_PC[15][1] ), .B2(n725), 
        .ZN(n2180) );
  OAI22_X1 U1467 ( .A1(n1284), .A2(n652), .B1(\predict_PC[15][3] ), .B2(n725), 
        .ZN(n2158) );
  OAI22_X1 U1425 ( .A1(n1284), .A2(target_PC_i[6]), .B1(\predict_PC[15][6] ), 
        .B2(n725), .ZN(n2125) );
  OAI22_X1 U1453 ( .A1(n1284), .A2(n641), .B1(\predict_PC[15][4] ), .B2(n725), 
        .ZN(n2147) );
  OAI22_X1 U1397 ( .A1(n1284), .A2(n639), .B1(\predict_PC[15][8] ), .B2(n725), 
        .ZN(n2103) );
  OAI22_X1 U1369 ( .A1(n1284), .A2(n640), .B1(\predict_PC[15][10] ), .B2(n725), 
        .ZN(n1515) );
  OAI22_X1 U118 ( .A1(n765), .A2(target_PC_i[13]), .B1(\predict_PC[0][13] ), 
        .B2(n2267), .ZN(n783) );
  OAI22_X1 U186 ( .A1(n800), .A2(n646), .B1(\predict_PC[1][12] ), .B2(n2264), 
        .ZN(n819) );
  OAI22_X1 U250 ( .A1(n834), .A2(n651), .B1(\predict_PC[2][13] ), .B2(n2261), 
        .ZN(n852) );
  OAI22_X1 U316 ( .A1(n868), .A2(n651), .B1(\predict_PC[3][13] ), .B2(n2258), 
        .ZN(n886) );
  OAI22_X1 U318 ( .A1(n868), .A2(n646), .B1(\predict_PC[3][12] ), .B2(n2258), 
        .ZN(n887) );
  OAI22_X1 U184 ( .A1(n800), .A2(target_PC_i[13]), .B1(\predict_PC[1][13] ), 
        .B2(n2264), .ZN(n818) );
  OAI22_X1 U252 ( .A1(n834), .A2(n646), .B1(\predict_PC[2][12] ), .B2(n2261), 
        .ZN(n853) );
  OAI22_X1 U120 ( .A1(n765), .A2(n646), .B1(\predict_PC[0][12] ), .B2(n2267), 
        .ZN(n784) );
  OAI22_X1 U302 ( .A1(n868), .A2(n638), .B1(\predict_PC[3][20] ), .B2(n2258), 
        .ZN(n879) );
  OAI22_X1 U238 ( .A1(n834), .A2(n645), .B1(\predict_PC[2][19] ), .B2(n2261), 
        .ZN(n846) );
  OAI22_X1 U102 ( .A1(n765), .A2(n642), .B1(\predict_PC[0][21] ), .B2(n2267), 
        .ZN(n775) );
  OAI22_X1 U240 ( .A1(n834), .A2(target_PC_i[18]), .B1(\predict_PC[2][18] ), 
        .B2(n2261), .ZN(n847) );
  OAI22_X1 U242 ( .A1(n834), .A2(n631), .B1(\predict_PC[2][17] ), .B2(n2261), 
        .ZN(n848) );
  OAI22_X1 U244 ( .A1(n834), .A2(n637), .B1(\predict_PC[2][16] ), .B2(n2261), 
        .ZN(n849) );
  OAI22_X1 U100 ( .A1(n765), .A2(n632), .B1(\predict_PC[0][22] ), .B2(n2267), 
        .ZN(n774) );
  OAI22_X1 U246 ( .A1(n834), .A2(target_PC_i[15]), .B1(\predict_PC[2][15] ), 
        .B2(n2261), .ZN(n850) );
  OAI22_X1 U104 ( .A1(n765), .A2(target_PC_i[20]), .B1(\predict_PC[0][20] ), 
        .B2(n2267), .ZN(n776) );
  OAI22_X1 U98 ( .A1(n765), .A2(n643), .B1(\predict_PC[0][23] ), .B2(n2267), 
        .ZN(n773) );
  OAI22_X1 U248 ( .A1(n834), .A2(n630), .B1(\predict_PC[2][14] ), .B2(n2261), 
        .ZN(n851) );
  OAI22_X1 U236 ( .A1(n834), .A2(n638), .B1(\predict_PC[2][20] ), .B2(n2261), 
        .ZN(n845) );
  OAI22_X1 U234 ( .A1(n834), .A2(n642), .B1(\predict_PC[2][21] ), .B2(n2261), 
        .ZN(n844) );
  OAI22_X1 U232 ( .A1(n834), .A2(n632), .B1(\predict_PC[2][22] ), .B2(n2261), 
        .ZN(n843) );
  OAI22_X1 U230 ( .A1(n834), .A2(n643), .B1(\predict_PC[2][23] ), .B2(n2261), 
        .ZN(n842) );
  OAI22_X1 U106 ( .A1(n765), .A2(n645), .B1(\predict_PC[0][19] ), .B2(n2267), 
        .ZN(n777) );
  OAI22_X1 U108 ( .A1(n765), .A2(target_PC_i[18]), .B1(\predict_PC[0][18] ), 
        .B2(n2267), .ZN(n778) );
  OAI22_X1 U110 ( .A1(n765), .A2(n631), .B1(\predict_PC[0][17] ), .B2(n2267), 
        .ZN(n779) );
  OAI22_X1 U112 ( .A1(n765), .A2(target_PC_i[16]), .B1(\predict_PC[0][16] ), 
        .B2(n2267), .ZN(n780) );
  OAI22_X1 U114 ( .A1(n765), .A2(target_PC_i[15]), .B1(\predict_PC[0][15] ), 
        .B2(n2267), .ZN(n781) );
  OAI22_X1 U170 ( .A1(n800), .A2(n638), .B1(\predict_PC[1][20] ), .B2(n2264), 
        .ZN(n811) );
  OAI22_X1 U116 ( .A1(n765), .A2(n630), .B1(\predict_PC[0][14] ), .B2(n2267), 
        .ZN(n782) );
  OAI22_X1 U182 ( .A1(n800), .A2(n630), .B1(\predict_PC[1][14] ), .B2(n2264), 
        .ZN(n817) );
  OAI22_X1 U178 ( .A1(n800), .A2(n637), .B1(\predict_PC[1][16] ), .B2(n2264), 
        .ZN(n815) );
  OAI22_X1 U180 ( .A1(n800), .A2(target_PC_i[15]), .B1(\predict_PC[1][15] ), 
        .B2(n2264), .ZN(n816) );
  OAI22_X1 U164 ( .A1(n800), .A2(n643), .B1(\predict_PC[1][23] ), .B2(n2264), 
        .ZN(n808) );
  OAI22_X1 U166 ( .A1(n800), .A2(n632), .B1(\predict_PC[1][22] ), .B2(n2264), 
        .ZN(n809) );
  OAI22_X1 U304 ( .A1(n868), .A2(n645), .B1(\predict_PC[3][19] ), .B2(n2258), 
        .ZN(n880) );
  OAI22_X1 U168 ( .A1(n800), .A2(n642), .B1(\predict_PC[1][21] ), .B2(n2264), 
        .ZN(n810) );
  OAI22_X1 U312 ( .A1(n868), .A2(target_PC_i[15]), .B1(\predict_PC[3][15] ), 
        .B2(n2258), .ZN(n884) );
  OAI22_X1 U174 ( .A1(n800), .A2(target_PC_i[18]), .B1(\predict_PC[1][18] ), 
        .B2(n2264), .ZN(n813) );
  OAI22_X1 U314 ( .A1(n868), .A2(n630), .B1(\predict_PC[3][14] ), .B2(n2258), 
        .ZN(n885) );
  OAI22_X1 U306 ( .A1(n868), .A2(target_PC_i[18]), .B1(\predict_PC[3][18] ), 
        .B2(n2258), .ZN(n881) );
  OAI22_X1 U296 ( .A1(n868), .A2(n643), .B1(\predict_PC[3][23] ), .B2(n2258), 
        .ZN(n876) );
  OAI22_X1 U310 ( .A1(n868), .A2(n637), .B1(\predict_PC[3][16] ), .B2(n2258), 
        .ZN(n883) );
  OAI22_X1 U308 ( .A1(n868), .A2(n631), .B1(\predict_PC[3][17] ), .B2(n2258), 
        .ZN(n882) );
  OAI22_X1 U298 ( .A1(n868), .A2(n632), .B1(\predict_PC[3][22] ), .B2(n2258), 
        .ZN(n877) );
  OAI22_X1 U172 ( .A1(n800), .A2(n645), .B1(\predict_PC[1][19] ), .B2(n2264), 
        .ZN(n812) );
  OAI22_X1 U176 ( .A1(n800), .A2(n631), .B1(\predict_PC[1][17] ), .B2(n2264), 
        .ZN(n814) );
  OAI22_X1 U300 ( .A1(n868), .A2(n642), .B1(\predict_PC[3][21] ), .B2(n2258), 
        .ZN(n878) );
  OAI22_X1 U1071 ( .A1(n1251), .A2(n633), .B1(\predict_PC[14][1] ), .B2(n728), 
        .ZN(n1281) );
  OAI22_X1 U995 ( .A1(n1218), .A2(target_PC_i[5]), .B1(\predict_PC[13][5] ), 
        .B2(n731), .ZN(n1244) );
  OAI22_X1 U993 ( .A1(n1218), .A2(target_PC_i[6]), .B1(\predict_PC[13][6] ), 
        .B2(n731), .ZN(n1243) );
  OAI22_X1 U989 ( .A1(n1218), .A2(n639), .B1(\predict_PC[13][8] ), .B2(n731), 
        .ZN(n1241) );
  OAI22_X1 U985 ( .A1(n1218), .A2(n640), .B1(\predict_PC[13][10] ), .B2(n731), 
        .ZN(n1239) );
  OAI22_X1 U1001 ( .A1(n1218), .A2(target_PC_i[2]), .B1(\predict_PC[13][2] ), 
        .B2(n731), .ZN(n1247) );
  OAI22_X1 U983 ( .A1(n1218), .A2(n644), .B1(\predict_PC[13][11] ), .B2(n731), 
        .ZN(n1238) );
  OAI22_X1 U999 ( .A1(n1218), .A2(n652), .B1(\predict_PC[13][3] ), .B2(n731), 
        .ZN(n1246) );
  OAI22_X1 U997 ( .A1(n1218), .A2(n641), .B1(\predict_PC[13][4] ), .B2(n731), 
        .ZN(n1245) );
  OAI22_X1 U1057 ( .A1(n1251), .A2(n639), .B1(\predict_PC[14][8] ), .B2(n728), 
        .ZN(n1274) );
  OAI22_X1 U1003 ( .A1(n1218), .A2(n633), .B1(\predict_PC[13][1] ), .B2(n731), 
        .ZN(n1248) );
  OAI22_X1 U932 ( .A1(n1184), .A2(n652), .B1(\predict_PC[12][3] ), .B2(n734), 
        .ZN(n1212) );
  OAI22_X1 U930 ( .A1(n1184), .A2(n641), .B1(\predict_PC[12][4] ), .B2(n734), 
        .ZN(n1211) );
  OAI22_X1 U1061 ( .A1(n1251), .A2(target_PC_i[6]), .B1(\predict_PC[14][6] ), 
        .B2(n728), .ZN(n1276) );
  OAI22_X1 U926 ( .A1(n1184), .A2(target_PC_i[6]), .B1(\predict_PC[12][6] ), 
        .B2(n734), .ZN(n1209) );
  OAI22_X1 U918 ( .A1(n1184), .A2(n640), .B1(\predict_PC[12][10] ), .B2(n734), 
        .ZN(n1205) );
  OAI22_X1 U1051 ( .A1(n1251), .A2(n644), .B1(\predict_PC[14][11] ), .B2(n728), 
        .ZN(n1271) );
  OAI22_X1 U922 ( .A1(n1184), .A2(n639), .B1(\predict_PC[12][8] ), .B2(n734), 
        .ZN(n1207) );
  OAI22_X1 U1069 ( .A1(n1251), .A2(n650), .B1(\predict_PC[14][2] ), .B2(n728), 
        .ZN(n1280) );
  OAI22_X1 U928 ( .A1(n1184), .A2(target_PC_i[5]), .B1(\predict_PC[12][5] ), 
        .B2(n734), .ZN(n1210) );
  OAI22_X1 U1067 ( .A1(n1251), .A2(n652), .B1(\predict_PC[14][3] ), .B2(n728), 
        .ZN(n1279) );
  OAI22_X1 U934 ( .A1(n1184), .A2(target_PC_i[2]), .B1(\predict_PC[12][2] ), 
        .B2(n734), .ZN(n1213) );
  OAI22_X1 U936 ( .A1(n1184), .A2(n633), .B1(\predict_PC[12][1] ), .B2(n734), 
        .ZN(n1214) );
  OAI22_X1 U1065 ( .A1(n1251), .A2(n641), .B1(\predict_PC[14][4] ), .B2(n728), 
        .ZN(n1278) );
  OAI22_X1 U916 ( .A1(n1184), .A2(n644), .B1(\predict_PC[12][11] ), .B2(n734), 
        .ZN(n1204) );
  OAI22_X1 U1053 ( .A1(n1251), .A2(n640), .B1(\predict_PC[14][10] ), .B2(n728), 
        .ZN(n1272) );
  OAI22_X1 U1063 ( .A1(n1251), .A2(target_PC_i[5]), .B1(\predict_PC[14][5] ), 
        .B2(n728), .ZN(n1277) );
  OAI22_X1 U663 ( .A1(n1051), .A2(target_PC_i[5]), .B1(\predict_PC[8][5] ), 
        .B2(n983), .ZN(n1077) );
  OAI22_X1 U534 ( .A1(n969), .A2(n652), .B1(\predict_PC[6][3] ), .B2(n989), 
        .ZN(n1013) );
  OAI22_X1 U520 ( .A1(n969), .A2(n640), .B1(\predict_PC[6][10] ), .B2(n989), 
        .ZN(n1006) );
  OAI22_X1 U530 ( .A1(n969), .A2(target_PC_i[5]), .B1(\predict_PC[6][5] ), 
        .B2(n989), .ZN(n1011) );
  OAI22_X1 U604 ( .A1(n1018), .A2(n633), .B1(\predict_PC[7][1] ), .B2(n986), 
        .ZN(n1048) );
  OAI22_X1 U518 ( .A1(n969), .A2(n644), .B1(\predict_PC[6][11] ), .B2(n989), 
        .ZN(n1005) );
  OAI22_X1 U532 ( .A1(n969), .A2(n641), .B1(\predict_PC[6][4] ), .B2(n989), 
        .ZN(n1012) );
  OAI22_X1 U524 ( .A1(n969), .A2(n639), .B1(\predict_PC[6][8] ), .B2(n989), 
        .ZN(n1008) );
  OAI22_X1 U653 ( .A1(n1051), .A2(n640), .B1(\predict_PC[8][10] ), .B2(n983), 
        .ZN(n1072) );
  OAI22_X1 U528 ( .A1(n969), .A2(target_PC_i[6]), .B1(\predict_PC[6][6] ), 
        .B2(n989), .ZN(n1010) );
  OAI22_X1 U651 ( .A1(n1051), .A2(n644), .B1(\predict_PC[8][11] ), .B2(n983), 
        .ZN(n1071) );
  OAI22_X1 U657 ( .A1(n1051), .A2(n639), .B1(\predict_PC[8][8] ), .B2(n983), 
        .ZN(n1074) );
  OAI22_X1 U669 ( .A1(n1051), .A2(n650), .B1(\predict_PC[8][2] ), .B2(n983), 
        .ZN(n1080) );
  OAI22_X1 U661 ( .A1(n1051), .A2(target_PC_i[6]), .B1(\predict_PC[8][6] ), 
        .B2(n983), .ZN(n1076) );
  OAI22_X1 U590 ( .A1(n1018), .A2(n639), .B1(\predict_PC[7][8] ), .B2(n986), 
        .ZN(n1041) );
  OAI22_X1 U586 ( .A1(n1018), .A2(target_PC_i[10]), .B1(\predict_PC[7][10] ), 
        .B2(n986), .ZN(n1039) );
  OAI22_X1 U602 ( .A1(n1018), .A2(target_PC_i[2]), .B1(\predict_PC[7][2] ), 
        .B2(n986), .ZN(n1047) );
  OAI22_X1 U719 ( .A1(n1085), .A2(n640), .B1(\predict_PC[9][10] ), .B2(n980), 
        .ZN(n1106) );
  OAI22_X1 U723 ( .A1(n1085), .A2(n639), .B1(\predict_PC[9][8] ), .B2(n980), 
        .ZN(n1108) );
  OAI22_X1 U584 ( .A1(n1018), .A2(n644), .B1(\predict_PC[7][11] ), .B2(n986), 
        .ZN(n1038) );
  OAI22_X1 U665 ( .A1(n1051), .A2(n641), .B1(\predict_PC[8][4] ), .B2(n983), 
        .ZN(n1078) );
  OAI22_X1 U727 ( .A1(n1085), .A2(target_PC_i[6]), .B1(\predict_PC[9][6] ), 
        .B2(n980), .ZN(n1110) );
  OAI22_X1 U594 ( .A1(n1018), .A2(target_PC_i[6]), .B1(\predict_PC[7][6] ), 
        .B2(n986), .ZN(n1043) );
  OAI22_X1 U667 ( .A1(n1051), .A2(n652), .B1(\predict_PC[8][3] ), .B2(n983), 
        .ZN(n1079) );
  OAI22_X1 U538 ( .A1(n969), .A2(n633), .B1(\predict_PC[6][1] ), .B2(n989), 
        .ZN(n1015) );
  OAI22_X1 U729 ( .A1(n1085), .A2(target_PC_i[5]), .B1(\predict_PC[9][5] ), 
        .B2(n980), .ZN(n1111) );
  OAI22_X1 U717 ( .A1(n1085), .A2(n644), .B1(\predict_PC[9][11] ), .B2(n980), 
        .ZN(n1105) );
  OAI22_X1 U731 ( .A1(n1085), .A2(target_PC_i[4]), .B1(\predict_PC[9][4] ), 
        .B2(n980), .ZN(n1112) );
  OAI22_X1 U671 ( .A1(n1051), .A2(n633), .B1(\predict_PC[8][1] ), .B2(n983), 
        .ZN(n1081) );
  OAI22_X1 U733 ( .A1(n1085), .A2(target_PC_i[3]), .B1(\predict_PC[9][3] ), 
        .B2(n980), .ZN(n1113) );
  OAI22_X1 U600 ( .A1(n1018), .A2(n652), .B1(\predict_PC[7][3] ), .B2(n986), 
        .ZN(n1046) );
  OAI22_X1 U598 ( .A1(n1018), .A2(n641), .B1(\predict_PC[7][4] ), .B2(n986), 
        .ZN(n1045) );
  OAI22_X1 U536 ( .A1(n969), .A2(n650), .B1(\predict_PC[6][2] ), .B2(n989), 
        .ZN(n1014) );
  OAI22_X1 U596 ( .A1(n1018), .A2(target_PC_i[5]), .B1(\predict_PC[7][5] ), 
        .B2(n986), .ZN(n1044) );
  OAI22_X1 U398 ( .A1(n902), .A2(target_PC_i[5]), .B1(\predict_PC[4][5] ), 
        .B2(n2254), .ZN(n928) );
  OAI22_X1 U735 ( .A1(n1085), .A2(n650), .B1(\predict_PC[9][2] ), .B2(n980), 
        .ZN(n1114) );
  OAI22_X1 U737 ( .A1(n1085), .A2(n633), .B1(\predict_PC[9][1] ), .B2(n980), 
        .ZN(n1115) );
  OAI22_X1 U472 ( .A1(n936), .A2(n633), .B1(\predict_PC[5][1] ), .B2(n2215), 
        .ZN(n966) );
  OAI22_X1 U470 ( .A1(n936), .A2(n650), .B1(\predict_PC[5][2] ), .B2(n2215), 
        .ZN(n965) );
  OAI22_X1 U468 ( .A1(n936), .A2(n652), .B1(\predict_PC[5][3] ), .B2(n2215), 
        .ZN(n964) );
  OAI22_X1 U466 ( .A1(n936), .A2(n641), .B1(\predict_PC[5][4] ), .B2(n2215), 
        .ZN(n963) );
  OAI22_X1 U464 ( .A1(n936), .A2(target_PC_i[5]), .B1(\predict_PC[5][5] ), 
        .B2(n2215), .ZN(n962) );
  OAI22_X1 U462 ( .A1(n936), .A2(target_PC_i[6]), .B1(\predict_PC[5][6] ), 
        .B2(n2215), .ZN(n961) );
  OAI22_X1 U849 ( .A1(n1151), .A2(n644), .B1(\predict_PC[11][11] ), .B2(n974), 
        .ZN(n1171) );
  OAI22_X1 U851 ( .A1(n1151), .A2(n640), .B1(\predict_PC[11][10] ), .B2(n974), 
        .ZN(n1172) );
  OAI22_X1 U855 ( .A1(n1151), .A2(n639), .B1(\predict_PC[11][8] ), .B2(n974), 
        .ZN(n1174) );
  OAI22_X1 U458 ( .A1(n936), .A2(n639), .B1(\predict_PC[5][8] ), .B2(n2215), 
        .ZN(n959) );
  OAI22_X1 U783 ( .A1(n1118), .A2(n644), .B1(\predict_PC[10][11] ), .B2(n977), 
        .ZN(n1138) );
  OAI22_X1 U785 ( .A1(n1118), .A2(n640), .B1(\predict_PC[10][10] ), .B2(n977), 
        .ZN(n1139) );
  OAI22_X1 U789 ( .A1(n1118), .A2(n639), .B1(\predict_PC[10][8] ), .B2(n977), 
        .ZN(n1141) );
  OAI22_X1 U454 ( .A1(n936), .A2(n640), .B1(\predict_PC[5][10] ), .B2(n2215), 
        .ZN(n957) );
  OAI22_X1 U793 ( .A1(n1118), .A2(target_PC_i[6]), .B1(\predict_PC[10][6] ), 
        .B2(n977), .ZN(n1143) );
  OAI22_X1 U452 ( .A1(n936), .A2(n644), .B1(\predict_PC[5][11] ), .B2(n2215), 
        .ZN(n956) );
  OAI22_X1 U795 ( .A1(n1118), .A2(target_PC_i[5]), .B1(\predict_PC[10][5] ), 
        .B2(n977), .ZN(n1144) );
  OAI22_X1 U803 ( .A1(n1118), .A2(n633), .B1(\predict_PC[10][1] ), .B2(n977), 
        .ZN(n1148) );
  OAI22_X1 U402 ( .A1(n902), .A2(n652), .B1(\predict_PC[4][3] ), .B2(n2254), 
        .ZN(n930) );
  OAI22_X1 U406 ( .A1(n902), .A2(target_PC_i[1]), .B1(\predict_PC[4][1] ), 
        .B2(n2254), .ZN(n932) );
  OAI22_X1 U400 ( .A1(n902), .A2(n641), .B1(\predict_PC[4][4] ), .B2(n2254), 
        .ZN(n929) );
  OAI22_X1 U869 ( .A1(n1151), .A2(n633), .B1(\predict_PC[11][1] ), .B2(n974), 
        .ZN(n1181) );
  OAI22_X1 U797 ( .A1(n1118), .A2(target_PC_i[4]), .B1(\predict_PC[10][4] ), 
        .B2(n977), .ZN(n1145) );
  OAI22_X1 U859 ( .A1(n1151), .A2(target_PC_i[6]), .B1(\predict_PC[11][6] ), 
        .B2(n974), .ZN(n1176) );
  OAI22_X1 U799 ( .A1(n1118), .A2(n652), .B1(\predict_PC[10][3] ), .B2(n977), 
        .ZN(n1146) );
  OAI22_X1 U801 ( .A1(n1118), .A2(target_PC_i[2]), .B1(\predict_PC[10][2] ), 
        .B2(n977), .ZN(n1147) );
  OAI22_X1 U396 ( .A1(n902), .A2(target_PC_i[6]), .B1(\predict_PC[4][6] ), 
        .B2(n2254), .ZN(n927) );
  OAI22_X1 U867 ( .A1(n1151), .A2(n650), .B1(\predict_PC[11][2] ), .B2(n974), 
        .ZN(n1180) );
  OAI22_X1 U863 ( .A1(n1151), .A2(n641), .B1(\predict_PC[11][4] ), .B2(n974), 
        .ZN(n1178) );
  OAI22_X1 U865 ( .A1(n1151), .A2(n652), .B1(\predict_PC[11][3] ), .B2(n974), 
        .ZN(n1179) );
  OAI22_X1 U404 ( .A1(n902), .A2(n650), .B1(\predict_PC[4][2] ), .B2(n2254), 
        .ZN(n931) );
  OAI22_X1 U388 ( .A1(n902), .A2(n640), .B1(\predict_PC[4][10] ), .B2(n2254), 
        .ZN(n923) );
  OAI22_X1 U392 ( .A1(n902), .A2(n639), .B1(\predict_PC[4][8] ), .B2(n2254), 
        .ZN(n925) );
  OAI22_X1 U386 ( .A1(n902), .A2(n644), .B1(\predict_PC[4][11] ), .B2(n2254), 
        .ZN(n922) );
  OAI22_X1 U861 ( .A1(n1151), .A2(target_PC_i[5]), .B1(\predict_PC[11][5] ), 
        .B2(n974), .ZN(n1177) );
  OAI22_X1 U200 ( .A1(n800), .A2(target_PC_i[5]), .B1(\predict_PC[1][5] ), 
        .B2(n2263), .ZN(n826) );
  OAI22_X1 U198 ( .A1(n800), .A2(target_PC_i[6]), .B1(\predict_PC[1][6] ), 
        .B2(n2263), .ZN(n825) );
  OAI22_X1 U194 ( .A1(n800), .A2(n639), .B1(\predict_PC[1][8] ), .B2(n2263), 
        .ZN(n823) );
  OAI22_X1 U138 ( .A1(n765), .A2(target_PC_i[3]), .B1(\predict_PC[0][3] ), 
        .B2(n2266), .ZN(n793) );
  OAI22_X1 U122 ( .A1(n765), .A2(n644), .B1(\predict_PC[0][11] ), .B2(n2266), 
        .ZN(n785) );
  OAI22_X1 U340 ( .A1(n868), .A2(n633), .B1(\predict_PC[3][1] ), .B2(n2257), 
        .ZN(n898) );
  OAI22_X1 U188 ( .A1(n800), .A2(n644), .B1(\predict_PC[1][11] ), .B2(n2263), 
        .ZN(n820) );
  OAI22_X1 U124 ( .A1(n765), .A2(n640), .B1(\predict_PC[0][10] ), .B2(n2266), 
        .ZN(n786) );
  OAI22_X1 U204 ( .A1(n800), .A2(n652), .B1(\predict_PC[1][3] ), .B2(n2263), 
        .ZN(n828) );
  OAI22_X1 U254 ( .A1(n834), .A2(n644), .B1(\predict_PC[2][11] ), .B2(n2260), 
        .ZN(n854) );
  OAI22_X1 U272 ( .A1(n834), .A2(n650), .B1(\predict_PC[2][2] ), .B2(n2260), 
        .ZN(n863) );
  OAI22_X1 U274 ( .A1(n834), .A2(n633), .B1(\predict_PC[2][1] ), .B2(n2260), 
        .ZN(n864) );
  OAI22_X1 U260 ( .A1(n834), .A2(n639), .B1(\predict_PC[2][8] ), .B2(n2260), 
        .ZN(n857) );
  OAI22_X1 U202 ( .A1(n800), .A2(target_PC_i[4]), .B1(\predict_PC[1][4] ), 
        .B2(n2263), .ZN(n827) );
  OAI22_X1 U128 ( .A1(n765), .A2(n639), .B1(\predict_PC[0][8] ), .B2(n2266), 
        .ZN(n788) );
  OAI22_X1 U140 ( .A1(n765), .A2(n650), .B1(\predict_PC[0][2] ), .B2(n2266), 
        .ZN(n794) );
  OAI22_X1 U208 ( .A1(n800), .A2(n633), .B1(\predict_PC[1][1] ), .B2(n2263), 
        .ZN(n830) );
  OAI22_X1 U256 ( .A1(n834), .A2(n640), .B1(\predict_PC[2][10] ), .B2(n2260), 
        .ZN(n855) );
  OAI22_X1 U268 ( .A1(n834), .A2(n641), .B1(\predict_PC[2][4] ), .B2(n2260), 
        .ZN(n861) );
  OAI22_X1 U270 ( .A1(n834), .A2(n652), .B1(\predict_PC[2][3] ), .B2(n2260), 
        .ZN(n862) );
  OAI22_X1 U320 ( .A1(n868), .A2(n644), .B1(\predict_PC[3][11] ), .B2(n2257), 
        .ZN(n888) );
  OAI22_X1 U206 ( .A1(n800), .A2(n650), .B1(\predict_PC[1][2] ), .B2(n2263), 
        .ZN(n829) );
  OAI22_X1 U322 ( .A1(n868), .A2(n640), .B1(\predict_PC[3][10] ), .B2(n2257), 
        .ZN(n889) );
  OAI22_X1 U136 ( .A1(n765), .A2(target_PC_i[4]), .B1(\predict_PC[0][4] ), 
        .B2(n2266), .ZN(n792) );
  OAI22_X1 U332 ( .A1(n868), .A2(target_PC_i[5]), .B1(\predict_PC[3][5] ), 
        .B2(n2257), .ZN(n894) );
  OAI22_X1 U326 ( .A1(n868), .A2(n639), .B1(\predict_PC[3][8] ), .B2(n2257), 
        .ZN(n891) );
  OAI22_X1 U132 ( .A1(n765), .A2(target_PC_i[6]), .B1(\predict_PC[0][6] ), 
        .B2(n2266), .ZN(n790) );
  OAI22_X1 U266 ( .A1(n834), .A2(target_PC_i[5]), .B1(\predict_PC[2][5] ), 
        .B2(n2260), .ZN(n860) );
  OAI22_X1 U334 ( .A1(n868), .A2(target_PC_i[4]), .B1(\predict_PC[3][4] ), 
        .B2(n2257), .ZN(n895) );
  OAI22_X1 U190 ( .A1(n800), .A2(n640), .B1(\predict_PC[1][10] ), .B2(n2263), 
        .ZN(n821) );
  OAI22_X1 U330 ( .A1(n868), .A2(target_PC_i[6]), .B1(\predict_PC[3][6] ), 
        .B2(n2257), .ZN(n893) );
  OAI22_X1 U134 ( .A1(n765), .A2(target_PC_i[5]), .B1(\predict_PC[0][5] ), 
        .B2(n2266), .ZN(n791) );
  OAI22_X1 U338 ( .A1(n868), .A2(n650), .B1(\predict_PC[3][2] ), .B2(n2257), 
        .ZN(n897) );
  OAI22_X1 U142 ( .A1(n765), .A2(n633), .B1(\predict_PC[0][1] ), .B2(n2266), 
        .ZN(n795) );
  OAI22_X1 U336 ( .A1(n868), .A2(target_PC_i[3]), .B1(\predict_PC[3][3] ), 
        .B2(n2257), .ZN(n896) );
  OAI22_X1 U264 ( .A1(n834), .A2(target_PC_i[6]), .B1(\predict_PC[2][6] ), 
        .B2(n2260), .ZN(n859) );
  OAI22_X1 U1159 ( .A1(n1284), .A2(n636), .B1(\predict_PC[15][25] ), .B2(n727), 
        .ZN(n1350) );
  OAI22_X1 U1145 ( .A1(n1284), .A2(n649), .B1(\predict_PC[15][26] ), .B2(n727), 
        .ZN(n1339) );
  OAI22_X1 U1023 ( .A1(n1251), .A2(n636), .B1(\predict_PC[14][25] ), .B2(n730), 
        .ZN(n1257) );
  OAI22_X1 U888 ( .A1(n1184), .A2(n636), .B1(\predict_PC[12][25] ), .B2(n737), 
        .ZN(n1190) );
  OAI22_X1 U1021 ( .A1(n1251), .A2(n649), .B1(\predict_PC[14][26] ), .B2(n730), 
        .ZN(n1256) );
  OAI22_X1 U955 ( .A1(n1218), .A2(n636), .B1(\predict_PC[13][25] ), .B2(n733), 
        .ZN(n1224) );
  OAI22_X1 U886 ( .A1(n1184), .A2(n649), .B1(\predict_PC[12][26] ), .B2(n737), 
        .ZN(n1189) );
  OAI22_X1 U953 ( .A1(n1218), .A2(n649), .B1(\predict_PC[13][26] ), .B2(n733), 
        .ZN(n1223) );
  OAI22_X1 U554 ( .A1(n1018), .A2(n649), .B1(\predict_PC[7][26] ), .B2(n988), 
        .ZN(n1023) );
  OAI22_X1 U422 ( .A1(n936), .A2(n649), .B1(\predict_PC[5][26] ), .B2(n2253), 
        .ZN(n941) );
  OAI22_X1 U821 ( .A1(n1151), .A2(n636), .B1(\predict_PC[11][25] ), .B2(n976), 
        .ZN(n1157) );
  OAI22_X1 U424 ( .A1(n936), .A2(n636), .B1(\predict_PC[5][25] ), .B2(n2253), 
        .ZN(n942) );
  OAI22_X1 U687 ( .A1(n1085), .A2(n649), .B1(\predict_PC[9][26] ), .B2(n982), 
        .ZN(n1090) );
  OAI22_X1 U819 ( .A1(n1151), .A2(n649), .B1(\predict_PC[11][26] ), .B2(n976), 
        .ZN(n1156) );
  OAI22_X1 U755 ( .A1(n1118), .A2(n636), .B1(\predict_PC[10][25] ), .B2(n979), 
        .ZN(n1124) );
  OAI22_X1 U556 ( .A1(n1018), .A2(n636), .B1(\predict_PC[7][25] ), .B2(n988), 
        .ZN(n1024) );
  OAI22_X1 U356 ( .A1(n902), .A2(n649), .B1(\predict_PC[4][26] ), .B2(n2256), 
        .ZN(n907) );
  OAI22_X1 U623 ( .A1(n1051), .A2(n636), .B1(\predict_PC[8][25] ), .B2(n985), 
        .ZN(n1057) );
  OAI22_X1 U753 ( .A1(n1118), .A2(n649), .B1(\predict_PC[10][26] ), .B2(n979), 
        .ZN(n1123) );
  OAI22_X1 U621 ( .A1(n1051), .A2(n649), .B1(\predict_PC[8][26] ), .B2(n985), 
        .ZN(n1056) );
  OAI22_X1 U488 ( .A1(n969), .A2(n649), .B1(\predict_PC[6][26] ), .B2(n2214), 
        .ZN(n990) );
  OAI22_X1 U490 ( .A1(n969), .A2(n636), .B1(\predict_PC[6][25] ), .B2(n2214), 
        .ZN(n991) );
  OAI22_X1 U358 ( .A1(n902), .A2(n636), .B1(\predict_PC[4][25] ), .B2(n2256), 
        .ZN(n908) );
  OAI22_X1 U689 ( .A1(n1085), .A2(n636), .B1(\predict_PC[9][25] ), .B2(n982), 
        .ZN(n1091) );
  OAI22_X1 U292 ( .A1(n868), .A2(n636), .B1(\predict_PC[3][25] ), .B2(n2259), 
        .ZN(n874) );
  OAI22_X1 U158 ( .A1(n800), .A2(n649), .B1(\predict_PC[1][26] ), .B2(n2265), 
        .ZN(n805) );
  OAI22_X1 U224 ( .A1(n834), .A2(n649), .B1(\predict_PC[2][26] ), .B2(n2262), 
        .ZN(n839) );
  OAI22_X1 U94 ( .A1(n765), .A2(n636), .B1(\predict_PC[0][25] ), .B2(n2268), 
        .ZN(n771) );
  OAI22_X1 U290 ( .A1(n868), .A2(n649), .B1(\predict_PC[3][26] ), .B2(n2259), 
        .ZN(n873) );
  OAI22_X1 U92 ( .A1(n765), .A2(n649), .B1(\predict_PC[0][26] ), .B2(n2268), 
        .ZN(n770) );
  OAI22_X1 U160 ( .A1(n800), .A2(n636), .B1(\predict_PC[1][25] ), .B2(n2265), 
        .ZN(n806) );
  OAI22_X1 U226 ( .A1(n834), .A2(n636), .B1(\predict_PC[2][25] ), .B2(n2262), 
        .ZN(n840) );
  NAND2_X1 U68 ( .A1(n2286), .A2(n2288), .ZN(n696) );
  AOI22_X1 U67 ( .A1(n2285), .A2(taken_o), .B1(n663), .B2(n696), .ZN(n736) );
  OAI21_X1 U34 ( .B1(n2285), .B2(n713), .A(n1284), .ZN(n2096) );
  OAI21_X1 U40 ( .B1(n2285), .B2(n710), .A(n1184), .ZN(n2093) );
  OAI21_X1 U38 ( .B1(n2285), .B2(n711), .A(n1218), .ZN(n2094) );
  OAI21_X1 U36 ( .B1(n2285), .B2(n712), .A(n1251), .ZN(n2095) );
  OAI21_X1 U54 ( .B1(n2285), .B2(n702), .A(n936), .ZN(n2086) );
  OAI21_X1 U44 ( .B1(n2285), .B2(n708), .A(n1118), .ZN(n2091) );
  OAI21_X1 U48 ( .B1(n2285), .B2(n706), .A(n1051), .ZN(n2089) );
  OAI21_X1 U52 ( .B1(n2285), .B2(n704), .A(n969), .ZN(n2087) );
  OAI21_X1 U46 ( .B1(n2285), .B2(n707), .A(n1085), .ZN(n2090) );
  OAI21_X1 U42 ( .B1(n2285), .B2(n709), .A(n1151), .ZN(n2092) );
  OAI21_X1 U50 ( .B1(n2285), .B2(n705), .A(n1018), .ZN(n2088) );
  OAI21_X1 U56 ( .B1(n2285), .B2(n700), .A(n902), .ZN(n2085) );
  OAI21_X1 U58 ( .B1(n2285), .B2(n698), .A(n868), .ZN(n2084) );
  OAI21_X1 U60 ( .B1(n2285), .B2(n695), .A(n834), .ZN(n2083) );
  OAI21_X1 U62 ( .B1(n2285), .B2(n694), .A(n800), .ZN(n2082) );
  OAI21_X1 U64 ( .B1(n2285), .B2(n665), .A(n765), .ZN(n2081) );
  AOI22_X1 U1188 ( .A1(n2287), .A2(n601), .B1(n678), .B2(n2285), .ZN(n1582) );
  AOI22_X1 U1244 ( .A1(n2287), .A2(n605), .B1(n683), .B2(n2285), .ZN(n1574) );
  AOI22_X1 U1216 ( .A1(n2287), .A2(n603), .B1(n680), .B2(n2285), .ZN(n1578) );
  AOI22_X1 U1272 ( .A1(n2287), .A2(n607), .B1(n685), .B2(n2285), .ZN(n1570) );
  AOI22_X1 U1356 ( .A1(n2287), .A2(n613), .B1(n691), .B2(n2285), .ZN(n1558) );
  AOI22_X1 U1412 ( .A1(n2287), .A2(n617), .B1(n668), .B2(n2285), .ZN(n1550) );
  AOI22_X1 U1230 ( .A1(n2287), .A2(n604), .B1(n681), .B2(n2285), .ZN(n1576) );
  AOI22_X1 U1258 ( .A1(n2287), .A2(n606), .B1(n684), .B2(n2285), .ZN(n1572) );
  AOI22_X1 U1342 ( .A1(n2287), .A2(n612), .B1(n690), .B2(n2285), .ZN(n1560) );
  AOI22_X1 U1314 ( .A1(n2287), .A2(n610), .B1(n688), .B2(n2285), .ZN(n1564) );
  AOI22_X1 U1300 ( .A1(n2287), .A2(n609), .B1(n687), .B2(n2285), .ZN(n1566) );
  AOI22_X1 U1202 ( .A1(n2287), .A2(n602), .B1(n679), .B2(n2285), .ZN(n1580) );
  AOI22_X1 U1286 ( .A1(n2287), .A2(n608), .B1(n686), .B2(n2285), .ZN(n1568) );
  AOI22_X1 U1328 ( .A1(n2287), .A2(n611), .B1(n689), .B2(n2285), .ZN(n1562) );
  AOI22_X1 U1454 ( .A1(n2287), .A2(n620), .B1(n671), .B2(n2285), .ZN(n1544) );
  AOI22_X1 U1146 ( .A1(n2287), .A2(n598), .B1(n675), .B2(n2285), .ZN(n1588) );
  AOI22_X1 U1426 ( .A1(stall_i), .A2(n618), .B1(n669), .B2(n2285), .ZN(n1548)
         );
  AOI22_X1 U1160 ( .A1(stall_i), .A2(n599), .B1(n676), .B2(n2285), .ZN(n1586)
         );
  AOI22_X1 U1482 ( .A1(stall_i), .A2(n622), .B1(n674), .B2(n2285), .ZN(n1540)
         );
  AOI22_X1 U1398 ( .A1(stall_i), .A2(n616), .B1(n667), .B2(n2285), .ZN(n1552)
         );
  AOI22_X1 U1384 ( .A1(stall_i), .A2(n615), .B1(n666), .B2(n2285), .ZN(n1554)
         );
  AOI22_X1 U1370 ( .A1(stall_i), .A2(n614), .B1(n692), .B2(n2285), .ZN(n1556)
         );
  AOI22_X1 U1468 ( .A1(stall_i), .A2(n621), .B1(n672), .B2(n2285), .ZN(n1542)
         );
  AOI22_X1 U1080 ( .A1(stall_i), .A2(n593), .B1(n673), .B2(n2285), .ZN(n1598)
         );
  AOI22_X1 U1174 ( .A1(stall_i), .A2(n600), .B1(n677), .B2(n2285), .ZN(n1584)
         );
  AOI22_X1 U1496 ( .A1(stall_i), .A2(n623), .B1(n682), .B2(n2285), .ZN(n1538)
         );
  AOI22_X1 U1440 ( .A1(stall_i), .A2(n619), .B1(n670), .B2(n2285), .ZN(n1546)
         );
  AOI22_X1 U1513 ( .A1(stall_i), .A2(n624), .B1(n693), .B2(n2285), .ZN(n1536)
         );
  OAI22_X1 U33 ( .A1(n2285), .A2(n660), .B1(n696), .B2(n703), .ZN(n2097) );
  OAI22_X1 U32 ( .A1(n2285), .A2(n662), .B1(n696), .B2(n701), .ZN(n2098) );
  OAI22_X1 U31 ( .A1(n2285), .A2(n661), .B1(n696), .B2(n699), .ZN(n2099) );
  OAI22_X1 U30 ( .A1(n2285), .A2(n664), .B1(n696), .B2(n697), .ZN(n2100) );
  NAND2_X1 U941 ( .A1(n662), .A2(n660), .ZN(n797) );
  NAND2_X1 U1512 ( .A1(n589), .A2(n588), .ZN(n900) );
  NAND2_X1 U1008 ( .A1(n588), .A2(n662), .ZN(n832) );
  NAND2_X1 U1076 ( .A1(n589), .A2(n660), .ZN(n866) );
  NOR2_X1 U1547 ( .A1(n2209), .A2(n2202), .ZN(n761) );
  NAND2_X1 U1538 ( .A1(TAG_i[3]), .A2(n699), .ZN(n2208) );
  NAND2_X1 U1529 ( .A1(TAG_i[2]), .A2(n697), .ZN(n2203) );
  NAND2_X1 U1550 ( .A1(TAG_i[1]), .A2(n703), .ZN(n2201) );
  NAND2_X1 U1522 ( .A1(n699), .A2(n697), .ZN(n2199) );
  NOR2_X1 U1543 ( .A1(n2198), .A2(n2209), .ZN(n762) );
  NOR2_X1 U1549 ( .A1(n2209), .A2(n2201), .ZN(n760) );
  NOR2_X1 U1534 ( .A1(n2201), .A2(n2208), .ZN(n758) );
  NOR2_X1 U1537 ( .A1(n2198), .A2(n2208), .ZN(n756) );
  NOR2_X1 U1525 ( .A1(n2198), .A2(n2203), .ZN(n750) );
  NOR2_X1 U1528 ( .A1(n2201), .A2(n2203), .ZN(n748) );
  NAND2_X1 U1544 ( .A1(n701), .A2(n703), .ZN(n2198) );
  NOR2_X1 U1517 ( .A1(n2198), .A2(n2199), .ZN(n747) );
  NAND3_X1 U1601 ( .A1(n590), .A2(n2286), .A3(n664), .ZN(n934) );
  NAND3_X1 U1602 ( .A1(n591), .A2(n2286), .A3(n661), .ZN(n1083) );
  NAND3_X1 U1600 ( .A1(n2286), .A2(n664), .A3(n661), .ZN(n798) );
  NAND3_X1 U1607 ( .A1(n591), .A2(n590), .A3(n2286), .ZN(n1216) );
  INV_X1 U1530 ( .A(TAG_i[3]), .ZN(n697) );
  INV_X1 U1539 ( .A(TAG_i[2]), .ZN(n699) );
  INV_X1 U1551 ( .A(TAG_i[0]), .ZN(n703) );
  INV_X1 U1545 ( .A(TAG_i[1]), .ZN(n701) );
  AND4_X1 U71 ( .A1(n740), .A2(n741), .A3(n742), .A4(n743), .ZN(n739) );
  AND4_X1 U76 ( .A1(n752), .A2(n753), .A3(n754), .A4(n755), .ZN(n738) );
  OR2_X1 U1107 ( .A1(n1307), .A2(n1308), .ZN(predicted_next_PC_o[29]) );
  OR2_X1 U1133 ( .A1(n1329), .A2(n1330), .ZN(predicted_next_PC_o[27]) );
  OR2_X1 U1120 ( .A1(n1318), .A2(n1319), .ZN(predicted_next_PC_o[28]) );
  OR2_X1 U1094 ( .A1(n1296), .A2(n1297), .ZN(predicted_next_PC_o[30]) );
  INV_X1 U9 ( .A(n673), .ZN(predicted_next_PC_o[31]) );
  INV_X1 U22 ( .A(n686), .ZN(predicted_next_PC_o[16]) );
  INV_X1 U6 ( .A(n670), .ZN(predicted_next_PC_o[5]) );
  INV_X1 U7 ( .A(n671), .ZN(predicted_next_PC_o[4]) );
  INV_X1 U23 ( .A(n687), .ZN(predicted_next_PC_o[15]) );
  INV_X1 U20 ( .A(n684), .ZN(predicted_next_PC_o[18]) );
  INV_X1 U21 ( .A(n685), .ZN(predicted_next_PC_o[17]) );
  INV_X1 U13 ( .A(n677), .ZN(predicted_next_PC_o[24]) );
  INV_X1 U15 ( .A(n679), .ZN(predicted_next_PC_o[22]) );
  INV_X1 U10 ( .A(n674), .ZN(predicted_next_PC_o[2]) );
  INV_X1 U2 ( .A(n666), .ZN(predicted_next_PC_o[9]) );
  INV_X1 U3 ( .A(n667), .ZN(predicted_next_PC_o[8]) );
  INV_X1 U5 ( .A(n669), .ZN(predicted_next_PC_o[6]) );
  INV_X1 U19 ( .A(n683), .ZN(predicted_next_PC_o[19]) );
  INV_X1 U17 ( .A(n681), .ZN(predicted_next_PC_o[20]) );
  INV_X1 U16 ( .A(n680), .ZN(predicted_next_PC_o[21]) );
  INV_X1 U14 ( .A(n678), .ZN(predicted_next_PC_o[23]) );
  INV_X1 U8 ( .A(n672), .ZN(predicted_next_PC_o[3]) );
  INV_X1 U4 ( .A(n668), .ZN(predicted_next_PC_o[7]) );
  INV_X1 U12 ( .A(n676), .ZN(predicted_next_PC_o[25]) );
  INV_X1 U11 ( .A(n675), .ZN(predicted_next_PC_o[26]) );
  INV_X1 U27 ( .A(n691), .ZN(predicted_next_PC_o[11]) );
  INV_X1 U25 ( .A(n689), .ZN(predicted_next_PC_o[13]) );
  INV_X1 U24 ( .A(n688), .ZN(predicted_next_PC_o[14]) );
  INV_X1 U18 ( .A(n682), .ZN(predicted_next_PC_o[1]) );
  INV_X1 U29 ( .A(n693), .ZN(predicted_next_PC_o[0]) );
  INV_X1 U28 ( .A(n692), .ZN(predicted_next_PC_o[10]) );
  INV_X1 U26 ( .A(n690), .ZN(predicted_next_PC_o[12]) );
  INV_X1 U66 ( .A(n736), .ZN(n2080) );
  OAI21_X1 U1557 ( .B1(was_taken_i), .B2(n663), .A(n592), .ZN(n2212) );
  INV_X1 U1340 ( .A(n1493), .ZN(n1561) );
  INV_X1 U800 ( .A(n1147), .ZN(n1730) );
  INV_X1 U569 ( .A(n1031), .ZN(n1842) );
  INV_X1 U429 ( .A(n945), .ZN(n1910) );
  INV_X1 U860 ( .A(n1177), .ZN(n1701) );
  INV_X1 U992 ( .A(n1243), .ZN(n1638) );
  INV_X1 U858 ( .A(n1176), .ZN(n1702) );
  INV_X1 U1062 ( .A(n1277), .ZN(n1605) );
  INV_X1 U503 ( .A(n998), .ZN(n1874) );
  INV_X1 U191 ( .A(n822), .ZN(n2025) );
  INV_X1 U804 ( .A(n1149), .ZN(n1728) );
  INV_X1 U1000 ( .A(n1247), .ZN(n1634) );
  INV_X1 U1060 ( .A(n1276), .ZN(n1606) );
  INV_X1 U636 ( .A(n1064), .ZN(n1810) );
  INV_X1 U720 ( .A(n1107), .ZN(n1769) );
  INV_X1 U197 ( .A(n825), .ZN(n2022) );
  INV_X1 U461 ( .A(n961), .ZN(n1894) );
  INV_X1 U852 ( .A(n1173), .ZN(n1705) );
  INV_X1 U463 ( .A(n962), .ZN(n1893) );
  INV_X1 U1072 ( .A(n1282), .ZN(n1600) );
  INV_X1 U305 ( .A(n881), .ZN(n1970) );
  INV_X1 U455 ( .A(n958), .ZN(n1897) );
  INV_X1 U397 ( .A(n928), .ZN(n1925) );
  INV_X1 U199 ( .A(n826), .ZN(n2021) );
  INV_X1 U449 ( .A(n955), .ZN(n1900) );
  INV_X1 U395 ( .A(n927), .ZN(n1926) );
  INV_X1 U1054 ( .A(n1273), .ZN(n1609) );
  INV_X1 U927 ( .A(n1210), .ZN(n1669) );
  INV_X1 U712 ( .A(n1103), .ZN(n1773) );
  INV_X1 U1382 ( .A(n1526), .ZN(n1555) );
  INV_X1 U994 ( .A(n1244), .ZN(n1637) );
  INV_X1 U201 ( .A(n827), .ZN(n2020) );
  INV_X1 U836 ( .A(n1165), .ZN(n1713) );
  INV_X1 U925 ( .A(n1209), .ZN(n1670) );
  INV_X1 U702 ( .A(n1098), .ZN(n1778) );
  INV_X1 U437 ( .A(n949), .ZN(n1906) );
  INV_X1 U933 ( .A(n1213), .ZN(n1666) );
  INV_X1 U323 ( .A(n890), .ZN(n1961) );
  INV_X1 U389 ( .A(n924), .ZN(n1929) );
  INV_X1 U135 ( .A(n792), .ZN(n2052) );
  INV_X1 U333 ( .A(n895), .ZN(n1956) );
  INV_X1 U137 ( .A(n793), .ZN(n2051) );
  INV_X1 U796 ( .A(n1145), .ZN(n1732) );
  INV_X1 U980 ( .A(n1237), .ZN(n1644) );
  INV_X1 U595 ( .A(n1044), .ZN(n1829) );
  INV_X1 U335 ( .A(n896), .ZN(n1955) );
  INV_X1 U660 ( .A(n1076), .ZN(n1798) );
  INV_X1 U794 ( .A(n1144), .ZN(n1733) );
  INV_X1 U792 ( .A(n1143), .ZN(n1734) );
  INV_X1 U1480 ( .A(n2169), .ZN(n1541) );
  INV_X1 U768 ( .A(n1131), .ZN(n1746) );
  INV_X1 U662 ( .A(n1077), .ZN(n1797) );
  INV_X1 U776 ( .A(n1135), .ZN(n1742) );
  INV_X1 U173 ( .A(n813), .ZN(n2034) );
  INV_X1 U521 ( .A(n1007), .ZN(n1865) );
  INV_X1 U1424 ( .A(n2125), .ZN(n1549) );
  INV_X1 U601 ( .A(n1047), .ZN(n1826) );
  INV_X1 U257 ( .A(n856), .ZN(n1993) );
  INV_X1 U529 ( .A(n1011), .ZN(n1861) );
  INV_X1 U371 ( .A(n915), .ZN(n1938) );
  INV_X1 U263 ( .A(n859), .ZN(n1990) );
  INV_X1 U265 ( .A(n860), .ZN(n1989) );
  INV_X1 U527 ( .A(n1010), .ZN(n1862) );
  INV_X1 U786 ( .A(n1140), .ZN(n1737) );
  INV_X1 U331 ( .A(n894), .ZN(n1957) );
  INV_X1 U587 ( .A(n1040), .ZN(n1833) );
  INV_X1 U732 ( .A(n1113), .ZN(n1763) );
  INV_X1 U1508 ( .A(n2191), .ZN(n1537) );
  INV_X1 U728 ( .A(n1111), .ZN(n1765) );
  INV_X1 U585 ( .A(n1039), .ZN(n1834) );
  INV_X1 U919 ( .A(n1206), .ZN(n1673) );
  INV_X1 U726 ( .A(n1110), .ZN(n1766) );
  INV_X1 U117 ( .A(n783), .ZN(n2061) );
  INV_X1 U183 ( .A(n818), .ZN(n2029) );
  INV_X1 U125 ( .A(n787), .ZN(n2057) );
  INV_X1 U1438 ( .A(n2136), .ZN(n1547) );
  INV_X1 U986 ( .A(n1240), .ZN(n1641) );
  INV_X1 U730 ( .A(n1112), .ZN(n1764) );
  INV_X1 U329 ( .A(n893), .ZN(n1958) );
  INV_X1 U654 ( .A(n1073), .ZN(n1801) );
  INV_X1 U593 ( .A(n1043), .ZN(n1830) );
  INV_X1 U1036 ( .A(n1264), .ZN(n1618) );
  INV_X1 U131 ( .A(n790), .ZN(n2054) );
  INV_X1 U133 ( .A(n791), .ZN(n2053) );
  INV_X1 U840 ( .A(n1167), .ZN(n1711) );
  INV_X1 U738 ( .A(n1116), .ZN(n1760) );
  INV_X1 U261 ( .A(n858), .ZN(n1991) );
  INV_X1 U666 ( .A(n1079), .ZN(n1795) );
  INV_X1 U788 ( .A(n1141), .ZN(n1736) );
  INV_X1 U784 ( .A(n1139), .ZN(n1738) );
  INV_X1 U982 ( .A(n1238), .ZN(n1643) );
  INV_X1 U179 ( .A(n816), .ZN(n2031) );
  INV_X1 U782 ( .A(n1138), .ZN(n1739) );
  INV_X1 U169 ( .A(n811), .ZN(n2036) );
  INV_X1 U1032 ( .A(n1262), .ZN(n1620) );
  INV_X1 U1200 ( .A(n1383), .ZN(n1581) );
  INV_X1 U605 ( .A(n1049), .ZN(n1824) );
  INV_X1 U1298 ( .A(n1460), .ZN(n1567) );
  INV_X1 U129 ( .A(n789), .ZN(n2055) );
  INV_X1 U1038 ( .A(n1265), .ZN(n1617) );
  INV_X1 U962 ( .A(n1228), .ZN(n1653) );
  INV_X1 U229 ( .A(n842), .ZN(n2007) );
  INV_X1 U1034 ( .A(n1263), .ZN(n1619) );
  INV_X1 U917 ( .A(n1205), .ZN(n1674) );
  INV_X1 U798 ( .A(n1146), .ZN(n1731) );
  INV_X1 U915 ( .A(n1204), .ZN(n1675) );
  INV_X1 U652 ( .A(n1072), .ZN(n1802) );
  INV_X1 U525 ( .A(n1009), .ZN(n1863) );
  INV_X1 U828 ( .A(n1161), .ZN(n1717) );
  INV_X1 U1270 ( .A(n1438), .ZN(n1571) );
  INV_X1 U780 ( .A(n1137), .ZN(n1740) );
  INV_X1 U167 ( .A(n810), .ZN(n2037) );
  INV_X1 U295 ( .A(n876), .ZN(n1975) );
  INV_X1 U692 ( .A(n1093), .ZN(n1783) );
  INV_X1 U231 ( .A(n843), .ZN(n2006) );
  INV_X1 U656 ( .A(n1074), .ZN(n1800) );
  INV_X1 U259 ( .A(n857), .ZN(n1992) );
  INV_X1 U341 ( .A(n899), .ZN(n1952) );
  INV_X1 U984 ( .A(n1239), .ZN(n1642) );
  INV_X1 U267 ( .A(n861), .ZN(n1988) );
  INV_X1 U523 ( .A(n1008), .ZN(n1864) );
  INV_X1 U139 ( .A(n794), .ZN(n2050) );
  INV_X1 U978 ( .A(n1236), .ZN(n1645) );
  INV_X1 U964 ( .A(n1229), .ZN(n1652) );
  INV_X1 U251 ( .A(n853), .ZN(n1996) );
  INV_X1 U513 ( .A(n1003), .ZN(n1869) );
  INV_X1 U790 ( .A(n1142), .ZN(n1735) );
  INV_X1 U511 ( .A(n1002), .ZN(n1870) );
  INV_X1 U772 ( .A(n1133), .ZN(n1744) );
  INV_X1 U958 ( .A(n1226), .ZN(n1655) );
  INV_X1 U672 ( .A(n1082), .ZN(n1792) );
  INV_X1 U175 ( .A(n814), .ZN(n2033) );
  INV_X1 U509 ( .A(n1001), .ZN(n1871) );
  INV_X1 U770 ( .A(n1132), .ZN(n1745) );
  INV_X1 U271 ( .A(n863), .ZN(n1986) );
  INV_X1 U247 ( .A(n851), .ZN(n1998) );
  INV_X1 U899 ( .A(n1196), .ZN(n1683) );
  INV_X1 U1410 ( .A(n2114), .ZN(n1551) );
  INV_X1 U515 ( .A(n1004), .ZN(n1868) );
  INV_X1 U249 ( .A(n852), .ZN(n1997) );
  INV_X1 U970 ( .A(n1232), .ZN(n1649) );
  INV_X1 U337 ( .A(n897), .ZN(n1954) );
  INV_X1 U909 ( .A(n1201), .ZN(n1678) );
  INV_X1 U517 ( .A(n1005), .ZN(n1867) );
  INV_X1 U269 ( .A(n862), .ZN(n1987) );
  INV_X1 U766 ( .A(n1130), .ZN(n1747) );
  INV_X1 U842 ( .A(n1168), .ZN(n1710) );
  INV_X1 U824 ( .A(n1159), .ZN(n1719) );
  INV_X1 U1284 ( .A(n1449), .ZN(n1569) );
  INV_X1 U764 ( .A(n1129), .ZN(n1748) );
  INV_X1 U907 ( .A(n1200), .ZN(n1679) );
  INV_X1 U762 ( .A(n1128), .ZN(n1749) );
  INV_X1 U275 ( .A(n865), .ZN(n1984) );
  INV_X1 U599 ( .A(n1046), .ZN(n1827) );
  INV_X1 U774 ( .A(n1134), .ZN(n1743) );
  INV_X1 U911 ( .A(n1202), .ZN(n1677) );
  INV_X1 U968 ( .A(n1231), .ZN(n1650) );
  INV_X1 U369 ( .A(n914), .ZN(n1939) );
  INV_X1 U531 ( .A(n1012), .ZN(n1860) );
  INV_X1 U913 ( .A(n1203), .ZN(n1676) );
  INV_X1 U373 ( .A(n916), .ZN(n1937) );
  INV_X1 U245 ( .A(n850), .ZN(n1999) );
  INV_X1 U760 ( .A(n1127), .ZN(n1750) );
  INV_X1 U972 ( .A(n1233), .ZN(n1648) );
  INV_X1 U243 ( .A(n849), .ZN(n2000) );
  INV_X1 U1026 ( .A(n1259), .ZN(n1623) );
  INV_X1 U758 ( .A(n1126), .ZN(n1751) );
  INV_X1 U1186 ( .A(n1372), .ZN(n1583) );
  INV_X1 U253 ( .A(n854), .ZN(n1995) );
  INV_X1 U960 ( .A(n1227), .ZN(n1654) );
  INV_X1 U974 ( .A(n1234), .ZN(n1647) );
  INV_X1 U519 ( .A(n1006), .ZN(n1866) );
  INV_X1 U644 ( .A(n1068), .ZN(n1806) );
  INV_X1 U241 ( .A(n848), .ZN(n2001) );
  INV_X1 U664 ( .A(n1078), .ZN(n1796) );
  INV_X1 U163 ( .A(n808), .ZN(n2039) );
  INV_X1 U597 ( .A(n1045), .ZN(n1828) );
  INV_X1 U905 ( .A(n1199), .ZN(n1680) );
  INV_X1 U255 ( .A(n855), .ZN(n1994) );
  INV_X1 U976 ( .A(n1235), .ZN(n1646) );
  INV_X1 U177 ( .A(n815), .ZN(n2032) );
  INV_X1 U239 ( .A(n847), .ZN(n2002) );
  INV_X1 U658 ( .A(n1075), .ZN(n1799) );
  INV_X1 U668 ( .A(n1080), .ZN(n1794) );
  INV_X1 U1028 ( .A(n1260), .ZN(n1622) );
  INV_X1 U143 ( .A(n796), .ZN(n2048) );
  INV_X1 U966 ( .A(n1230), .ZN(n1651) );
  INV_X1 U237 ( .A(n846), .ZN(n2003) );
  INV_X1 U778 ( .A(n1136), .ZN(n1741) );
  INV_X1 U642 ( .A(n1067), .ZN(n1807) );
  INV_X1 U235 ( .A(n845), .ZN(n2004) );
  INV_X1 U171 ( .A(n812), .ZN(n2035) );
  INV_X1 U361 ( .A(n910), .ZN(n1943) );
  INV_X1 U826 ( .A(n1160), .ZN(n1718) );
  INV_X1 U165 ( .A(n809), .ZN(n2038) );
  INV_X1 U233 ( .A(n844), .ZN(n2005) );
  INV_X1 U1030 ( .A(n1261), .ZN(n1621) );
  INV_X1 U533 ( .A(n1013), .ZN(n1859) );
  INV_X1 U433 ( .A(n947), .ZN(n1908) );
  INV_X1 U710 ( .A(n1102), .ZN(n1774) );
  INV_X1 U561 ( .A(n1027), .ZN(n1846) );
  INV_X1 U107 ( .A(n778), .ZN(n2066) );
  INV_X1 U387 ( .A(n923), .ZN(n1930) );
  INV_X1 U694 ( .A(n1094), .ZN(n1782) );
  INV_X1 U990 ( .A(n1242), .ZN(n1639) );
  INV_X1 U435 ( .A(n948), .ZN(n1907) );
  INV_X1 U209 ( .A(n831), .ZN(n2016) );
  INV_X1 U937 ( .A(n1215), .ZN(n1664) );
  INV_X1 U718 ( .A(n1106), .ZN(n1770) );
  INV_X1 U559 ( .A(n1026), .ZN(n1847) );
  INV_X1 U363 ( .A(n911), .ZN(n1942) );
  INV_X1 U309 ( .A(n883), .ZN(n1968) );
  INV_X1 U1228 ( .A(n1405), .ZN(n1577) );
  INV_X1 U921 ( .A(n1207), .ZN(n1672) );
  INV_X1 U105 ( .A(n777), .ZN(n2067) );
  INV_X1 U1050 ( .A(n1271), .ZN(n1611) );
  INV_X1 U405 ( .A(n932), .ZN(n1921) );
  INV_X1 U439 ( .A(n950), .ZN(n1905) );
  INV_X1 U317 ( .A(n887), .ZN(n1964) );
  INV_X1 U856 ( .A(n1175), .ZN(n1703) );
  INV_X1 U441 ( .A(n951), .ZN(n1904) );
  INV_X1 U205 ( .A(n829), .ZN(n2018) );
  INV_X1 U499 ( .A(n996), .ZN(n1876) );
  INV_X1 U497 ( .A(n995), .ZN(n1877) );
  INV_X1 U1396 ( .A(n2103), .ZN(n1553) );
  INV_X1 U846 ( .A(n1170), .ZN(n1708) );
  INV_X1 U903 ( .A(n1198), .ZN(n1681) );
  INV_X1 U1066 ( .A(n1279), .ZN(n1603) );
  INV_X1 U716 ( .A(n1105), .ZN(n1771) );
  INV_X1 U391 ( .A(n925), .ZN(n1928) );
  INV_X1 U495 ( .A(n994), .ZN(n1878) );
  INV_X1 U923 ( .A(n1208), .ZN(n1671) );
  INV_X1 U187 ( .A(n820), .ZN(n2027) );
  INV_X1 U193 ( .A(n823), .ZN(n2024) );
  INV_X1 U901 ( .A(n1197), .ZN(n1682) );
  INV_X1 U203 ( .A(n828), .ZN(n2019) );
  INV_X1 U696 ( .A(n1095), .ZN(n1781) );
  INV_X1 U493 ( .A(n993), .ZN(n1879) );
  INV_X1 U1052 ( .A(n1272), .ZN(n1610) );
  INV_X1 U632 ( .A(n1062), .ZN(n1812) );
  INV_X1 U403 ( .A(n931), .ZN(n1922) );
  INV_X1 U443 ( .A(n952), .ZN(n1903) );
  INV_X1 U103 ( .A(n776), .ZN(n2068) );
  INV_X1 U321 ( .A(n889), .ZN(n1962) );
  INV_X1 U393 ( .A(n926), .ZN(n1927) );
  INV_X1 U848 ( .A(n1171), .ZN(n1707) );
  INV_X1 U101 ( .A(n775), .ZN(n2069) );
  INV_X1 U996 ( .A(n1245), .ZN(n1636) );
  INV_X1 U303 ( .A(n880), .ZN(n1971) );
  INV_X1 U630 ( .A(n1061), .ZN(n1813) );
  INV_X1 U1058 ( .A(n1275), .ZN(n1607) );
  INV_X1 U1068 ( .A(n1280), .ZN(n1602) );
  INV_X1 U189 ( .A(n821), .ZN(n2026) );
  INV_X1 U99 ( .A(n774), .ZN(n2070) );
  INV_X1 U1242 ( .A(n1416), .ZN(n1575) );
  INV_X1 U473 ( .A(n967), .ZN(n1888) );
  INV_X1 U539 ( .A(n1016), .ZN(n1856) );
  INV_X1 U850 ( .A(n1172), .ZN(n1706) );
  INV_X1 U97 ( .A(n773), .ZN(n2071) );
  INV_X1 U469 ( .A(n965), .ZN(n1890) );
  INV_X1 U1452 ( .A(n2147), .ZN(n1545) );
  INV_X1 U401 ( .A(n930), .ZN(n1923) );
  INV_X1 U399 ( .A(n929), .ZN(n1924) );
  INV_X1 U445 ( .A(n953), .ZN(n1902) );
  INV_X1 U467 ( .A(n964), .ZN(n1891) );
  INV_X1 U1354 ( .A(n1504), .ZN(n1559) );
  INV_X1 U1368 ( .A(n1515), .ZN(n1557) );
  INV_X1 U1326 ( .A(n1482), .ZN(n1563) );
  INV_X1 U638 ( .A(n1065), .ZN(n1809) );
  INV_X1 U447 ( .A(n954), .ZN(n1901) );
  INV_X1 U465 ( .A(n963), .ZN(n1892) );
  INV_X1 U698 ( .A(n1096), .ZN(n1780) );
  INV_X1 U714 ( .A(n1104), .ZN(n1772) );
  INV_X1 U459 ( .A(n960), .ZN(n1895) );
  INV_X1 U998 ( .A(n1246), .ZN(n1635) );
  INV_X1 U319 ( .A(n888), .ZN(n1963) );
  INV_X1 U307 ( .A(n882), .ZN(n1969) );
  INV_X1 U457 ( .A(n959), .ZN(n1896) );
  INV_X1 U648 ( .A(n1070), .ZN(n1804) );
  INV_X1 U453 ( .A(n957), .ZN(n1898) );
  INV_X1 U854 ( .A(n1174), .ZN(n1704) );
  INV_X1 U1056 ( .A(n1274), .ZN(n1608) );
  INV_X1 U700 ( .A(n1097), .ZN(n1779) );
  INV_X1 U195 ( .A(n824), .ZN(n2023) );
  INV_X1 U451 ( .A(n956), .ZN(n1899) );
  INV_X1 U988 ( .A(n1241), .ZN(n1640) );
  INV_X1 U297 ( .A(n877), .ZN(n1974) );
  INV_X1 U591 ( .A(n1042), .ZN(n1831) );
  INV_X1 U313 ( .A(n885), .ZN(n1966) );
  INV_X1 U864 ( .A(n1179), .ZN(n1699) );
  INV_X1 U866 ( .A(n1180), .ZN(n1698) );
  INV_X1 U706 ( .A(n1100), .ZN(n1776) );
  INV_X1 U589 ( .A(n1041), .ZN(n1832) );
  INV_X1 U734 ( .A(n1114), .ZN(n1762) );
  INV_X1 U127 ( .A(n788), .ZN(n2056) );
  INV_X1 U929 ( .A(n1211), .ZN(n1668) );
  INV_X1 U646 ( .A(n1069), .ZN(n1805) );
  INV_X1 U1256 ( .A(n1427), .ZN(n1573) );
  INV_X1 U830 ( .A(n1162), .ZN(n1716) );
  INV_X1 U1312 ( .A(n1471), .ZN(n1565) );
  INV_X1 U897 ( .A(n1195), .ZN(n1684) );
  INV_X1 U535 ( .A(n1014), .ZN(n1858) );
  INV_X1 U123 ( .A(n786), .ZN(n2058) );
  INV_X1 U626 ( .A(n1059), .ZN(n1815) );
  INV_X1 U583 ( .A(n1038), .ZN(n1835) );
  INV_X1 U1040 ( .A(n1266), .ZN(n1616) );
  INV_X1 U375 ( .A(n917), .ZN(n1936) );
  INV_X1 U181 ( .A(n817), .ZN(n2030) );
  INV_X1 U895 ( .A(n1194), .ZN(n1685) );
  INV_X1 U581 ( .A(n1037), .ZN(n1836) );
  INV_X1 U708 ( .A(n1101), .ZN(n1775) );
  INV_X1 U862 ( .A(n1178), .ZN(n1700) );
  INV_X1 U1004 ( .A(n1249), .ZN(n1632) );
  INV_X1 U121 ( .A(n785), .ZN(n2059) );
  INV_X1 U579 ( .A(n1036), .ZN(n1837) );
  INV_X1 U870 ( .A(n1182), .ZN(n1696) );
  INV_X1 U1042 ( .A(n1267), .ZN(n1615) );
  INV_X1 U377 ( .A(n918), .ZN(n1935) );
  INV_X1 U931 ( .A(n1212), .ZN(n1667) );
  INV_X1 U1466 ( .A(n2158), .ZN(n1543) );
  INV_X1 U577 ( .A(n1035), .ZN(n1838) );
  INV_X1 U119 ( .A(n784), .ZN(n2060) );
  INV_X1 U379 ( .A(n919), .ZN(n1934) );
  INV_X1 U1044 ( .A(n1268), .ZN(n1614) );
  INV_X1 U315 ( .A(n886), .ZN(n1965) );
  INV_X1 U365 ( .A(n912), .ZN(n1941) );
  INV_X1 U507 ( .A(n1000), .ZN(n1872) );
  INV_X1 U381 ( .A(n920), .ZN(n1933) );
  INV_X1 U832 ( .A(n1163), .ZN(n1715) );
  INV_X1 U1064 ( .A(n1278), .ZN(n1604) );
  INV_X1 U1214 ( .A(n1394), .ZN(n1579) );
  INV_X1 U575 ( .A(n1034), .ZN(n1839) );
  INV_X1 U407 ( .A(n933), .ZN(n1920) );
  INV_X1 U650 ( .A(n1071), .ZN(n1803) );
  INV_X1 U115 ( .A(n782), .ZN(n2062) );
  INV_X1 U571 ( .A(n1032), .ZN(n1841) );
  INV_X1 U640 ( .A(n1066), .ZN(n1808) );
  INV_X1 U724 ( .A(n1109), .ZN(n1767) );
  INV_X1 U383 ( .A(n921), .ZN(n1932) );
  INV_X1 U113 ( .A(n781), .ZN(n2063) );
  INV_X1 U834 ( .A(n1164), .ZN(n1714) );
  INV_X1 U573 ( .A(n1033), .ZN(n1840) );
  INV_X1 U722 ( .A(n1108), .ZN(n1768) );
  INV_X1 U1046 ( .A(n1269), .ZN(n1613) );
  INV_X1 U427 ( .A(n944), .ZN(n1911) );
  INV_X1 U501 ( .A(n997), .ZN(n1875) );
  INV_X1 U327 ( .A(n892), .ZN(n1959) );
  INV_X1 U111 ( .A(n780), .ZN(n2064) );
  INV_X1 U844 ( .A(n1169), .ZN(n1709) );
  INV_X1 U431 ( .A(n946), .ZN(n1909) );
  INV_X1 U385 ( .A(n922), .ZN(n1931) );
  INV_X1 U628 ( .A(n1060), .ZN(n1814) );
  INV_X1 U893 ( .A(n1193), .ZN(n1686) );
  INV_X1 U185 ( .A(n819), .ZN(n2028) );
  INV_X1 U299 ( .A(n878), .ZN(n1973) );
  INV_X1 U704 ( .A(n1099), .ZN(n1777) );
  INV_X1 U311 ( .A(n884), .ZN(n1967) );
  INV_X1 U1048 ( .A(n1270), .ZN(n1612) );
  INV_X1 U563 ( .A(n1028), .ZN(n1845) );
  INV_X1 U301 ( .A(n879), .ZN(n1972) );
  INV_X1 U325 ( .A(n891), .ZN(n1960) );
  INV_X1 U838 ( .A(n1166), .ZN(n1712) );
  INV_X1 U891 ( .A(n1192), .ZN(n1687) );
  INV_X1 U367 ( .A(n913), .ZN(n1940) );
  INV_X1 U109 ( .A(n779), .ZN(n2065) );
  INV_X1 U634 ( .A(n1063), .ZN(n1811) );
  INV_X1 U505 ( .A(n999), .ZN(n1873) );
  INV_X1 U567 ( .A(n1030), .ZN(n1843) );
  INV_X1 U565 ( .A(n1029), .ZN(n1844) );
  INV_X1 U802 ( .A(n1148), .ZN(n1729) );
  INV_X1 U1494 ( .A(n2180), .ZN(n1539) );
  INV_X1 U273 ( .A(n864), .ZN(n1985) );
  INV_X1 U471 ( .A(n966), .ZN(n1889) );
  INV_X1 U221 ( .A(n838), .ZN(n2011) );
  INV_X1 U141 ( .A(n795), .ZN(n2049) );
  INV_X1 U537 ( .A(n1015), .ZN(n1857) );
  INV_X1 U736 ( .A(n1115), .ZN(n1761) );
  INV_X1 U207 ( .A(n830), .ZN(n2017) );
  INV_X1 U1002 ( .A(n1248), .ZN(n1633) );
  INV_X1 U889 ( .A(n1191), .ZN(n1688) );
  INV_X1 U935 ( .A(n1214), .ZN(n1665) );
  INV_X1 U1070 ( .A(n1281), .ZN(n1601) );
  INV_X1 U603 ( .A(n1048), .ZN(n1825) );
  INV_X1 U868 ( .A(n1181), .ZN(n1697) );
  INV_X1 U339 ( .A(n898), .ZN(n1953) );
  INV_X1 U670 ( .A(n1081), .ZN(n1793) );
  INV_X1 U950 ( .A(n1222), .ZN(n1659) );
  INV_X1 U952 ( .A(n1223), .ZN(n1658) );
  INV_X1 U1018 ( .A(n1255), .ZN(n1627) );
  INV_X1 U684 ( .A(n1089), .ZN(n1787) );
  INV_X1 U85 ( .A(n767), .ZN(n2077) );
  INV_X1 U1131 ( .A(n1328), .ZN(n1591) );
  INV_X1 U754 ( .A(n1124), .ZN(n1753) );
  INV_X1 U1020 ( .A(n1256), .ZN(n1626) );
  INV_X1 U287 ( .A(n872), .ZN(n1979) );
  INV_X1 U686 ( .A(n1090), .ZN(n1786) );
  INV_X1 U91 ( .A(n770), .ZN(n2074) );
  INV_X1 U1022 ( .A(n1257), .ZN(n1625) );
  INV_X1 U750 ( .A(n1122), .ZN(n1755) );
  INV_X1 U159 ( .A(n806), .ZN(n2041) );
  INV_X1 U1144 ( .A(n1339), .ZN(n1589) );
  INV_X1 U157 ( .A(n805), .ZN(n2042) );
  INV_X1 U155 ( .A(n804), .ZN(n2043) );
  INV_X1 U752 ( .A(n1123), .ZN(n1754) );
  INV_X1 U289 ( .A(n873), .ZN(n1978) );
  INV_X1 U225 ( .A(n840), .ZN(n2009) );
  INV_X1 U816 ( .A(n1155), .ZN(n1723) );
  INV_X1 U223 ( .A(n839), .ZN(n2010) );
  INV_X1 U291 ( .A(n874), .ZN(n1977) );
  INV_X1 U89 ( .A(n769), .ZN(n2075) );
  INV_X1 U555 ( .A(n1024), .ZN(n1849) );
  INV_X1 U885 ( .A(n1189), .ZN(n1690) );
  INV_X1 U883 ( .A(n1188), .ZN(n1691) );
  INV_X1 U553 ( .A(n1023), .ZN(n1850) );
  INV_X1 U551 ( .A(n1022), .ZN(n1851) );
  INV_X1 U419 ( .A(n940), .ZN(n1915) );
  INV_X1 U421 ( .A(n941), .ZN(n1914) );
  INV_X1 U423 ( .A(n942), .ZN(n1913) );
  INV_X1 U485 ( .A(n973), .ZN(n1883) );
  INV_X1 U487 ( .A(n990), .ZN(n1882) );
  INV_X1 U489 ( .A(n991), .ZN(n1881) );
  INV_X1 U618 ( .A(n1055), .ZN(n1819) );
  INV_X1 U353 ( .A(n906), .ZN(n1947) );
  INV_X1 U818 ( .A(n1156), .ZN(n1722) );
  INV_X1 U620 ( .A(n1056), .ZN(n1818) );
  INV_X1 U820 ( .A(n1157), .ZN(n1721) );
  INV_X1 U622 ( .A(n1057), .ZN(n1817) );
  INV_X1 U355 ( .A(n907), .ZN(n1946) );
  INV_X1 U357 ( .A(n908), .ZN(n1945) );
  INV_X1 U359 ( .A(n909), .ZN(n1944) );
  INV_X1 U491 ( .A(n992), .ZN(n1880) );
  INV_X1 U624 ( .A(n1058), .ZN(n1816) );
  INV_X1 U481 ( .A(n971), .ZN(n1885) );
  INV_X1 U1105 ( .A(n1306), .ZN(n1595) );
  INV_X1 U149 ( .A(n801), .ZN(n2046) );
  INV_X1 U217 ( .A(n836), .ZN(n2013) );
  INV_X1 U946 ( .A(n1220), .ZN(n1661) );
  INV_X1 U479 ( .A(n970), .ZN(n1886) );
  INV_X1 U1012 ( .A(n1252), .ZN(n1630) );
  INV_X1 U215 ( .A(n835), .ZN(n2014) );
  INV_X1 U293 ( .A(n875), .ZN(n1976) );
  INV_X1 U690 ( .A(n1092), .ZN(n1784) );
  INV_X1 U944 ( .A(n1219), .ZN(n1662) );
  INV_X1 U746 ( .A(n1120), .ZN(n1757) );
  INV_X1 U1024 ( .A(n1258), .ZN(n1624) );
  INV_X1 U93 ( .A(n771), .ZN(n2073) );
  INV_X1 U413 ( .A(n937), .ZN(n1918) );
  INV_X1 U756 ( .A(n1125), .ZN(n1752) );
  INV_X1 U744 ( .A(n1119), .ZN(n1758) );
  INV_X1 U283 ( .A(n870), .ZN(n1981) );
  INV_X1 U1092 ( .A(n1295), .ZN(n1597) );
  INV_X1 U415 ( .A(n938), .ZN(n1917) );
  INV_X1 U227 ( .A(n841), .ZN(n2008) );
  INV_X1 U822 ( .A(n1158), .ZN(n1720) );
  INV_X1 U425 ( .A(n943), .ZN(n1912) );
  INV_X1 U557 ( .A(n1025), .ZN(n1848) );
  INV_X1 U349 ( .A(n904), .ZN(n1949) );
  INV_X1 U151 ( .A(n802), .ZN(n2045) );
  INV_X1 U688 ( .A(n1091), .ZN(n1785) );
  INV_X1 U678 ( .A(n1086), .ZN(n1790) );
  INV_X1 U161 ( .A(n807), .ZN(n2040) );
  INV_X1 U1158 ( .A(n1350), .ZN(n1587) );
  INV_X1 U281 ( .A(n869), .ZN(n1982) );
  INV_X1 U1014 ( .A(n1253), .ZN(n1629) );
  INV_X1 U612 ( .A(n1052), .ZN(n1822) );
  INV_X1 U956 ( .A(n1225), .ZN(n1656) );
  INV_X1 U877 ( .A(n1185), .ZN(n1694) );
  INV_X1 U810 ( .A(n1152), .ZN(n1726) );
  INV_X1 U95 ( .A(n772), .ZN(n2072) );
  INV_X1 U812 ( .A(n1153), .ZN(n1725) );
  INV_X1 U610 ( .A(n1050), .ZN(n1823) );
  INV_X1 U545 ( .A(n1019), .ZN(n1854) );
  INV_X1 U1172 ( .A(n1361), .ZN(n1585) );
  INV_X1 U680 ( .A(n1087), .ZN(n1789) );
  INV_X1 U347 ( .A(n903), .ZN(n1950) );
  INV_X1 U547 ( .A(n1020), .ZN(n1853) );
  INV_X1 U887 ( .A(n1190), .ZN(n1689) );
  INV_X1 U614 ( .A(n1053), .ZN(n1821) );
  INV_X1 U954 ( .A(n1224), .ZN(n1657) );
  INV_X1 U879 ( .A(n1186), .ZN(n1693) );
  INV_X1 U83 ( .A(n766), .ZN(n2078) );
  INV_X1 U814 ( .A(n1154), .ZN(n1724) );
  INV_X1 U1016 ( .A(n1254), .ZN(n1628) );
  INV_X1 U279 ( .A(n867), .ZN(n1983) );
  INV_X1 U345 ( .A(n901), .ZN(n1951) );
  INV_X1 U1010 ( .A(n1250), .ZN(n1631) );
  INV_X1 U81 ( .A(n764), .ZN(n2079) );
  INV_X1 U616 ( .A(n1054), .ZN(n1820) );
  INV_X1 U942 ( .A(n1217), .ZN(n1663) );
  INV_X1 U682 ( .A(n1088), .ZN(n1788) );
  INV_X1 U543 ( .A(n1017), .ZN(n1855) );
  INV_X1 U1078 ( .A(n1283), .ZN(n1599) );
  INV_X1 U417 ( .A(n939), .ZN(n1916) );
  INV_X1 U881 ( .A(n1187), .ZN(n1692) );
  INV_X1 U1118 ( .A(n1317), .ZN(n1593) );
  INV_X1 U808 ( .A(n1150), .ZN(n1727) );
  INV_X1 U748 ( .A(n1121), .ZN(n1756) );
  INV_X1 U483 ( .A(n972), .ZN(n1884) );
  INV_X1 U411 ( .A(n935), .ZN(n1919) );
  INV_X1 U153 ( .A(n803), .ZN(n2044) );
  INV_X1 U213 ( .A(n833), .ZN(n2015) );
  INV_X1 U351 ( .A(n905), .ZN(n1948) );
  INV_X1 U875 ( .A(n1183), .ZN(n1695) );
  INV_X1 U742 ( .A(n1117), .ZN(n1759) );
  INV_X1 U87 ( .A(n768), .ZN(n2076) );
  INV_X1 U948 ( .A(n1221), .ZN(n1660) );
  INV_X1 U549 ( .A(n1021), .ZN(n1852) );
  INV_X1 U147 ( .A(n799), .ZN(n2047) );
  INV_X1 U676 ( .A(n1084), .ZN(n1791) );
  INV_X1 U219 ( .A(n837), .ZN(n2012) );
  INV_X1 U477 ( .A(n968), .ZN(n1887) );
  INV_X1 U285 ( .A(n871), .ZN(n1980) );
  BUF_X1 U35 ( .A(target_PC_i[23]), .Z(n643) );
  BUF_X1 U37 ( .A(target_PC_i[21]), .Z(n642) );
  CLKBUF_X1 U39 ( .A(target_PC_i[29]), .Z(n634) );
  BUF_X1 U41 ( .A(target_PC_i[25]), .Z(n636) );
  BUF_X1 U43 ( .A(target_PC_i[3]), .Z(n652) );
  BUF_X1 U45 ( .A(target_PC_i[2]), .Z(n650) );
  BUF_X1 U47 ( .A(target_PC_i[13]), .Z(n651) );
  INV_X1 U49 ( .A(stall_i), .ZN(n2286) );
  AND2_X1 U51 ( .A1(n2224), .A2(n8), .ZN(n714) );
  BUF_X1 U53 ( .A(target_PC_i[31]), .Z(n647) );
  AND2_X1 U55 ( .A1(n9), .A2(n2222), .ZN(n717) );
  BUF_X1 U57 ( .A(target_PC_i[24]), .Z(n635) );
  BUF_X1 U59 ( .A(target_PC_i[27]), .Z(n653) );
  BUF_X1 U61 ( .A(target_PC_i[1]), .Z(n633) );
  AND2_X1 U63 ( .A1(target_PC_i[6]), .A2(n618), .ZN(n720) );
  BUF_X1 U65 ( .A(target_PC_i[4]), .Z(n641) );
  BUF_X1 U69 ( .A(target_PC_i[8]), .Z(n639) );
  BUF_X1 U70 ( .A(target_PC_i[12]), .Z(n646) );
  BUF_X1 U82 ( .A(target_PC_i[0]), .Z(n648) );
  INV_X1 U84 ( .A(n765), .ZN(n2268) );
  INV_X1 U86 ( .A(n1184), .ZN(n734) );
  INV_X1 U88 ( .A(n800), .ZN(n2264) );
  INV_X1 U90 ( .A(n868), .ZN(n2259) );
  INV_X1 U96 ( .A(n1284), .ZN(n726) );
  INV_X1 U126 ( .A(n1018), .ZN(n987) );
  INV_X1 U130 ( .A(n1051), .ZN(n984) );
  INV_X1 U144 ( .A(n1085), .ZN(n982) );
  INV_X1 U145 ( .A(n902), .ZN(n2256) );
  INV_X1 U146 ( .A(n902), .ZN(n2254) );
  INV_X1 U148 ( .A(n765), .ZN(n2266) );
  INV_X1 U150 ( .A(n969), .ZN(n2214) );
  INV_X1 U152 ( .A(n834), .ZN(n2260) );
  INV_X1 U154 ( .A(n1151), .ZN(n976) );
  INV_X1 U156 ( .A(n902), .ZN(n2255) );
  INV_X1 U162 ( .A(n969), .ZN(n2213) );
  INV_X1 U192 ( .A(n1284), .ZN(n727) );
  INV_X1 U196 ( .A(n834), .ZN(n2262) );
  INV_X1 U210 ( .A(n868), .ZN(n2258) );
  INV_X1 U211 ( .A(n1184), .ZN(n735) );
  INV_X1 U212 ( .A(n1118), .ZN(n977) );
  INV_X1 U214 ( .A(n1151), .ZN(n974) );
  INV_X1 U216 ( .A(n1251), .ZN(n728) );
  INV_X1 U218 ( .A(n1218), .ZN(n732) );
  INV_X1 U220 ( .A(n1251), .ZN(n730) );
  INV_X1 U222 ( .A(n1018), .ZN(n988) );
  INV_X1 U228 ( .A(n800), .ZN(n2263) );
  INV_X1 U258 ( .A(n765), .ZN(n2267) );
  INV_X1 U262 ( .A(n1085), .ZN(n980) );
  INV_X1 U276 ( .A(n1051), .ZN(n985) );
  INV_X1 U277 ( .A(n1284), .ZN(n725) );
  INV_X1 U278 ( .A(n834), .ZN(n2261) );
  INV_X1 U280 ( .A(n1085), .ZN(n981) );
  INV_X1 U282 ( .A(n1118), .ZN(n979) );
  INV_X1 U284 ( .A(n1118), .ZN(n978) );
  INV_X1 U286 ( .A(n969), .ZN(n989) );
  INV_X1 U288 ( .A(n1184), .ZN(n737) );
  INV_X1 U294 ( .A(n936), .ZN(n2216) );
  INV_X1 U324 ( .A(n936), .ZN(n2215) );
  INV_X1 U328 ( .A(n868), .ZN(n2257) );
  INV_X1 U342 ( .A(n936), .ZN(n2253) );
  INV_X1 U343 ( .A(n1218), .ZN(n733) );
  INV_X1 U344 ( .A(n1251), .ZN(n729) );
  INV_X1 U346 ( .A(n1051), .ZN(n983) );
  INV_X1 U348 ( .A(n1151), .ZN(n975) );
  INV_X1 U350 ( .A(n1018), .ZN(n986) );
  INV_X1 U352 ( .A(n800), .ZN(n2265) );
  INV_X1 U354 ( .A(n1218), .ZN(n731) );
  OR2_X2 U360 ( .A1(n1216), .A2(n866), .ZN(n1251) );
  OR2_X2 U390 ( .A1(n900), .A2(n1083), .ZN(n1151) );
  OR2_X2 U394 ( .A1(n832), .A2(n934), .ZN(n936) );
  OR2_X2 U408 ( .A1(n866), .A2(n1083), .ZN(n1118) );
  OR2_X2 U409 ( .A1(n866), .A2(n798), .ZN(n834) );
  OR2_X2 U410 ( .A1(n900), .A2(n1216), .ZN(n1284) );
  OR2_X2 U412 ( .A1(n866), .A2(n934), .ZN(n969) );
  OR2_X2 U414 ( .A1(n832), .A2(n1083), .ZN(n1085) );
  OR2_X2 U416 ( .A1(n900), .A2(n798), .ZN(n868) );
  OR2_X2 U418 ( .A1(n1216), .A2(n797), .ZN(n1184) );
  OR2_X2 U420 ( .A1(n797), .A2(n934), .ZN(n902) );
  OR2_X2 U426 ( .A1(n797), .A2(n1083), .ZN(n1051) );
  OR2_X2 U456 ( .A1(n900), .A2(n934), .ZN(n1018) );
  OR2_X2 U460 ( .A1(n1216), .A2(n832), .ZN(n1218) );
  OR2_X2 U474 ( .A1(n832), .A2(n798), .ZN(n800) );
  OR2_X2 U475 ( .A1(n797), .A2(n798), .ZN(n765) );
  INV_X2 U476 ( .A(stall_i), .ZN(n2285) );
  BUF_X2 U478 ( .A(n762), .Z(n2270) );
  BUF_X2 U480 ( .A(n746), .Z(n2282) );
  BUF_X2 U482 ( .A(n745), .Z(n2283) );
  BUF_X2 U484 ( .A(n744), .Z(n2284) );
  BUF_X2 U486 ( .A(n751), .Z(n2277) );
  BUF_X2 U492 ( .A(n760), .Z(n2272) );
  BUF_X2 U522 ( .A(n749), .Z(n2279) );
  BUF_X2 U526 ( .A(n750), .Z(n2278) );
  BUF_X2 U540 ( .A(n748), .Z(n2280) );
  BUF_X2 U541 ( .A(n763), .Z(n2269) );
  BUF_X2 U542 ( .A(n756), .Z(n2276) );
  BUF_X2 U544 ( .A(n758), .Z(n2274) );
  BUF_X2 U546 ( .A(n757), .Z(n2275) );
  BUF_X2 U548 ( .A(n759), .Z(n2273) );
  BUF_X2 U550 ( .A(n761), .Z(n2271) );
  INV_X1 U552 ( .A(reset), .ZN(n2291) );
  INV_X1 U558 ( .A(reset), .ZN(n2293) );
  INV_X1 U588 ( .A(reset), .ZN(n2310) );
  INV_X1 U592 ( .A(reset), .ZN(n2296) );
  INV_X1 U606 ( .A(reset), .ZN(n2290) );
  INV_X1 U607 ( .A(reset), .ZN(n2302) );
  INV_X1 U608 ( .A(reset), .ZN(n2307) );
  INV_X1 U609 ( .A(reset), .ZN(n2304) );
  INV_X1 U611 ( .A(reset), .ZN(n2289) );
  INV_X1 U613 ( .A(reset), .ZN(n2288) );
  INV_X1 U615 ( .A(reset), .ZN(n2309) );
  INV_X1 U617 ( .A(reset), .ZN(n2297) );
  INV_X1 U619 ( .A(reset), .ZN(n2299) );
  INV_X1 U625 ( .A(reset), .ZN(n2306) );
  INV_X1 U655 ( .A(reset), .ZN(n2295) );
  INV_X1 U659 ( .A(reset), .ZN(n2308) );
  INV_X1 U673 ( .A(reset), .ZN(n2298) );
  INV_X1 U674 ( .A(reset), .ZN(n2294) );
  INV_X1 U675 ( .A(reset), .ZN(n2303) );
  INV_X1 U677 ( .A(reset), .ZN(n2301) );
  INV_X1 U679 ( .A(reset), .ZN(n2300) );
  INV_X1 U681 ( .A(reset), .ZN(n2292) );
  INV_X1 U683 ( .A(reset), .ZN(n2305) );
  INV_X1 U685 ( .A(reset), .ZN(n2311) );
  BUF_X1 U691 ( .A(target_PC_i[14]), .Z(n630) );
  BUF_X1 U721 ( .A(target_PC_i[19]), .Z(n645) );
  BUF_X1 U725 ( .A(target_PC_i[17]), .Z(n631) );
  BUF_X1 U739 ( .A(target_PC_i[22]), .Z(n632) );
  BUF_X1 U740 ( .A(target_PC_i[16]), .Z(n637) );
  BUF_X1 U741 ( .A(target_PC_i[20]), .Z(n638) );
  BUF_X1 U743 ( .A(target_PC_i[26]), .Z(n649) );
  BUF_X1 U745 ( .A(target_PC_i[10]), .Z(n640) );
  AND2_X1 U747 ( .A1(target_PC_i[24]), .A2(n600), .ZN(n719) );
  AND2_X1 U749 ( .A1(n7), .A2(n2225), .ZN(n715) );
  BUF_X2 U751 ( .A(target_PC_i[11]), .Z(n644) );
  AND2_X1 U757 ( .A1(n623), .A2(target_PC_i[1]), .ZN(n723) );
  AND2_X1 U787 ( .A1(target_PC_i[31]), .A2(n593), .ZN(n718) );
  AND4_X1 U791 ( .A1(n655), .A2(n654), .A3(n656), .A4(n657), .ZN(n2211) );
  AND4_X1 U805 ( .A1(n2247), .A2(n2246), .A3(n2248), .A4(n2245), .ZN(n654) );
  AND4_X1 U806 ( .A1(n2238), .A2(n2239), .A3(n2237), .A4(n2240), .ZN(n655) );
  AND4_X1 U807 ( .A1(n2232), .A2(n2229), .A3(n2231), .A4(n2230), .ZN(n656) );
  AND4_X1 U809 ( .A1(n2219), .A2(n2218), .A3(n2220), .A4(n2217), .ZN(n657) );
  INV_X1 U811 ( .A(n724), .ZN(n2210) );
  AND2_X1 U813 ( .A1(target_PC_i[0]), .A2(n624), .ZN(n722) );
  INV_X1 U815 ( .A(target_PC_i[29]), .ZN(n2225) );
  CLKBUF_X1 U817 ( .A(target_PC_i[30]), .Z(n658) );
  AND2_X1 U823 ( .A1(n2221), .A2(n6), .ZN(n716) );
  INV_X1 U853 ( .A(target_PC_i[27]), .ZN(n2222) );
  CLKBUF_X1 U857 ( .A(target_PC_i[28]), .Z(n659) );
  CLKBUF_X1 U871 ( .A(mispredict_o), .Z(n724) );
  INV_X1 U872 ( .A(target_PC_i[30]), .ZN(n2221) );
  AND2_X1 U873 ( .A1(n617), .A2(target_PC_i[7]), .ZN(n721) );
  INV_X1 U874 ( .A(target_PC_i[28]), .ZN(n2224) );
  AOI21_X1 U876 ( .B1(n2211), .B2(n663), .A(n2212), .ZN(mispredict_o) );
  AOI21_X1 U878 ( .B1(n738), .B2(n739), .A(reset), .ZN(taken_o) );
  BUF_X1 U880 ( .A(stall_i), .Z(n2287) );
  BUF_X1 U882 ( .A(n747), .Z(n2281) );
  AOI221_X1 U884 ( .B1(target_PC_i[10]), .B2(n614), .C1(n613), .C2(n644), .A(
        n2249), .ZN(n2248) );
  AOI221_X1 U890 ( .B1(target_PC_i[8]), .B2(n616), .C1(target_PC_i[9]), .C2(
        n615), .A(n2250), .ZN(n2247) );
  AOI221_X1 U920 ( .B1(target_PC_i[14]), .B2(n610), .C1(n609), .C2(
        target_PC_i[15]), .A(n2251), .ZN(n2246) );
  NOR2_X1 U924 ( .A1(n2200), .A2(n2199), .ZN(n746) );
  NOR2_X1 U938 ( .A1(n2202), .A2(n2199), .ZN(n744) );
  NOR2_X1 U939 ( .A1(n2200), .A2(n2208), .ZN(n757) );
  NOR2_X1 U940 ( .A1(n2200), .A2(n2203), .ZN(n751) );
  NOR2_X1 U943 ( .A1(n2209), .A2(n2200), .ZN(n763) );
  NOR2_X1 U945 ( .A1(n2202), .A2(n2208), .ZN(n759) );
  NOR2_X1 U947 ( .A1(n2202), .A2(n2203), .ZN(n749) );
  NOR2_X1 U949 ( .A1(n2201), .A2(n2199), .ZN(n745) );
  OAI22_X1 U951 ( .A1(target_PC_i[16]), .A2(n608), .B1(target_PC_i[17]), .B2(
        n607), .ZN(n2228) );
  OAI22_X1 U957 ( .A1(target_PC_i[18]), .A2(n606), .B1(target_PC_i[19]), .B2(
        n605), .ZN(n2227) );
  OAI22_X1 U987 ( .A1(n2224), .A2(n8), .B1(n2225), .B2(n7), .ZN(n2226) );
  OAI22_X1 U991 ( .A1(n2221), .A2(n6), .B1(n2222), .B2(n9), .ZN(n2223) );
  OAI22_X1 U1005 ( .A1(target_PC_i[22]), .A2(n602), .B1(target_PC_i[23]), .B2(
        n601), .ZN(n2233) );
  OAI22_X1 U1006 ( .A1(target_PC_i[20]), .A2(n604), .B1(target_PC_i[21]), .B2(
        n603), .ZN(n2234) );
  OAI22_X1 U1007 ( .A1(target_PC_i[25]), .A2(n599), .B1(target_PC_i[26]), .B2(
        n598), .ZN(n2235) );
  OAI22_X1 U1009 ( .A1(target_PC_i[31]), .A2(n593), .B1(target_PC_i[24]), .B2(
        n600), .ZN(n2236) );
  OAI22_X1 U1011 ( .A1(target_PC_i[2]), .A2(n622), .B1(target_PC_i[3]), .B2(
        n621), .ZN(n2241) );
  OAI22_X1 U1013 ( .A1(target_PC_i[0]), .A2(n624), .B1(target_PC_i[1]), .B2(
        n623), .ZN(n2242) );
  OAI22_X1 U1015 ( .A1(target_PC_i[6]), .A2(n618), .B1(target_PC_i[7]), .B2(
        n617), .ZN(n2243) );
  OAI22_X1 U1017 ( .A1(target_PC_i[4]), .A2(n620), .B1(target_PC_i[5]), .B2(
        n619), .ZN(n2244) );
  OAI22_X1 U1019 ( .A1(target_PC_i[10]), .A2(n614), .B1(target_PC_i[11]), .B2(
        n613), .ZN(n2249) );
  OAI22_X1 U1025 ( .A1(target_PC_i[8]), .A2(n616), .B1(target_PC_i[9]), .B2(
        n615), .ZN(n2250) );
  OAI22_X1 U1055 ( .A1(target_PC_i[14]), .A2(n610), .B1(target_PC_i[15]), .B2(
        n609), .ZN(n2251) );
  OAI22_X1 U1059 ( .A1(target_PC_i[12]), .A2(n612), .B1(target_PC_i[13]), .B2(
        n611), .ZN(n2252) );
  AOI221_X1 U1073 ( .B1(target_PC_i[16]), .B2(n608), .C1(n607), .C2(
        target_PC_i[17]), .A(n2228), .ZN(n2217) );
  AOI221_X1 U1074 ( .B1(target_PC_i[18]), .B2(n606), .C1(n605), .C2(
        target_PC_i[19]), .A(n2227), .ZN(n2218) );
  NOR3_X1 U1075 ( .A1(n2226), .A2(n715), .A3(n714), .ZN(n2219) );
  NOR3_X1 U1077 ( .A1(n2223), .A2(n717), .A3(n716), .ZN(n2220) );
  AOI221_X1 U1079 ( .B1(target_PC_i[22]), .B2(n602), .C1(target_PC_i[23]), 
        .C2(n601), .A(n2233), .ZN(n2232) );
  AOI221_X1 U1093 ( .B1(target_PC_i[20]), .B2(n604), .C1(target_PC_i[21]), 
        .C2(n603), .A(n2234), .ZN(n2231) );
  AOI221_X1 U1106 ( .B1(target_PC_i[25]), .B2(n599), .C1(n598), .C2(
        target_PC_i[26]), .A(n2235), .ZN(n2230) );
  NOR3_X1 U1119 ( .A1(n718), .A2(n719), .A3(n2236), .ZN(n2229) );
  AOI221_X1 U1132 ( .B1(target_PC_i[2]), .B2(n622), .C1(n621), .C2(
        target_PC_i[3]), .A(n2241), .ZN(n2240) );
  NOR3_X1 U1173 ( .A1(n722), .A2(n723), .A3(n2242), .ZN(n2239) );
  NOR3_X1 U1383 ( .A1(n721), .A2(n720), .A3(n2243), .ZN(n2238) );
  AOI221_X1 U1411 ( .B1(target_PC_i[4]), .B2(n620), .C1(n619), .C2(
        target_PC_i[5]), .A(n2244), .ZN(n2237) );
  AOI221_X1 U1509 ( .B1(target_PC_i[12]), .B2(n612), .C1(n611), .C2(
        target_PC_i[13]), .A(n2252), .ZN(n2245) );
  OAI22_X1 U1510 ( .A1(n1284), .A2(n647), .B1(\predict_PC[15][31] ), .B2(n727), 
        .ZN(n1283) );
  OAI22_X1 U1511 ( .A1(n1251), .A2(n647), .B1(\predict_PC[14][31] ), .B2(n730), 
        .ZN(n1250) );
  OAI22_X1 U1518 ( .A1(n969), .A2(n647), .B1(\predict_PC[6][31] ), .B2(n2214), 
        .ZN(n968) );
  OAI22_X1 U1520 ( .A1(n1118), .A2(n647), .B1(\predict_PC[10][31] ), .B2(n979), 
        .ZN(n1117) );
  OAI22_X1 U1521 ( .A1(n834), .A2(n647), .B1(\predict_PC[2][31] ), .B2(n2262), 
        .ZN(n833) );
  OAI22_X1 U1524 ( .A1(n765), .A2(n647), .B1(\predict_PC[0][31] ), .B2(n2268), 
        .ZN(n764) );
  OAI22_X1 U1527 ( .A1(n800), .A2(n647), .B1(\predict_PC[1][31] ), .B2(n2265), 
        .ZN(n799) );
  OAI22_X1 U1533 ( .A1(n868), .A2(n647), .B1(\predict_PC[3][31] ), .B2(n2259), 
        .ZN(n867) );
  OAI22_X1 U1536 ( .A1(n936), .A2(n647), .B1(\predict_PC[5][31] ), .B2(n2253), 
        .ZN(n935) );
  OAI22_X1 U1541 ( .A1(n1018), .A2(n647), .B1(\predict_PC[7][31] ), .B2(n988), 
        .ZN(n1017) );
  OAI22_X1 U1554 ( .A1(n1051), .A2(target_PC_i[31]), .B1(\predict_PC[8][31] ), 
        .B2(n985), .ZN(n1050) );
  OAI22_X1 U1555 ( .A1(n1085), .A2(n647), .B1(\predict_PC[9][31] ), .B2(n982), 
        .ZN(n1084) );
  OAI22_X1 U1556 ( .A1(n1218), .A2(n647), .B1(\predict_PC[13][31] ), .B2(n733), 
        .ZN(n1217) );
  OAI22_X1 U1558 ( .A1(n1151), .A2(n647), .B1(\predict_PC[11][31] ), .B2(n976), 
        .ZN(n1150) );
  OAI22_X1 U1559 ( .A1(n902), .A2(n647), .B1(\predict_PC[4][31] ), .B2(n2256), 
        .ZN(n901) );
  OAI22_X1 U1560 ( .A1(n1184), .A2(n647), .B1(\predict_PC[12][31] ), .B2(n737), 
        .ZN(n1183) );
  OAI22_X1 U1561 ( .A1(n765), .A2(n648), .B1(\predict_PC[0][0] ), .B2(n2266), 
        .ZN(n796) );
  OAI22_X1 U1562 ( .A1(n800), .A2(n648), .B1(\predict_PC[1][0] ), .B2(n2263), 
        .ZN(n831) );
  OAI22_X1 U1563 ( .A1(n834), .A2(n648), .B1(\predict_PC[2][0] ), .B2(n2260), 
        .ZN(n865) );
  OAI22_X1 U1564 ( .A1(n868), .A2(n648), .B1(\predict_PC[3][0] ), .B2(n2257), 
        .ZN(n899) );
  OAI22_X1 U1565 ( .A1(n902), .A2(n648), .B1(\predict_PC[4][0] ), .B2(n2254), 
        .ZN(n933) );
  OAI22_X1 U1566 ( .A1(n936), .A2(n648), .B1(\predict_PC[5][0] ), .B2(n2215), 
        .ZN(n967) );
  OAI22_X1 U1567 ( .A1(n969), .A2(n648), .B1(\predict_PC[6][0] ), .B2(n989), 
        .ZN(n1016) );
  OAI22_X1 U1568 ( .A1(n1018), .A2(n648), .B1(\predict_PC[7][0] ), .B2(n986), 
        .ZN(n1049) );
  OAI22_X1 U1569 ( .A1(n1051), .A2(n648), .B1(\predict_PC[8][0] ), .B2(n983), 
        .ZN(n1082) );
  OAI22_X1 U1570 ( .A1(n1085), .A2(n648), .B1(\predict_PC[9][0] ), .B2(n980), 
        .ZN(n1116) );
  OAI22_X1 U1571 ( .A1(n1118), .A2(target_PC_i[0]), .B1(\predict_PC[10][0] ), 
        .B2(n977), .ZN(n1149) );
  OAI22_X1 U1572 ( .A1(n1151), .A2(n648), .B1(\predict_PC[11][0] ), .B2(n974), 
        .ZN(n1182) );
  OAI22_X1 U1573 ( .A1(n1184), .A2(n648), .B1(\predict_PC[12][0] ), .B2(n734), 
        .ZN(n1215) );
  OAI22_X1 U1574 ( .A1(n1218), .A2(n648), .B1(\predict_PC[13][0] ), .B2(n731), 
        .ZN(n1249) );
  OAI22_X1 U1575 ( .A1(n1251), .A2(target_PC_i[0]), .B1(\predict_PC[14][0] ), 
        .B2(n728), .ZN(n1282) );
  OAI22_X1 U1576 ( .A1(n1284), .A2(target_PC_i[0]), .B1(\predict_PC[15][0] ), 
        .B2(n725), .ZN(n2191) );
  OAI22_X1 U1577 ( .A1(n765), .A2(target_PC_i[9]), .B1(\predict_PC[0][9] ), 
        .B2(n2266), .ZN(n787) );
  OAI22_X1 U1578 ( .A1(n1018), .A2(target_PC_i[9]), .B1(\predict_PC[7][9] ), 
        .B2(n986), .ZN(n1040) );
  OAI22_X1 U1579 ( .A1(n1251), .A2(target_PC_i[9]), .B1(\predict_PC[14][9] ), 
        .B2(n728), .ZN(n1273) );
  OAI22_X1 U1580 ( .A1(n1051), .A2(target_PC_i[9]), .B1(\predict_PC[8][9] ), 
        .B2(n983), .ZN(n1073) );
  OAI22_X1 U1581 ( .A1(n1085), .A2(target_PC_i[9]), .B1(\predict_PC[9][9] ), 
        .B2(n980), .ZN(n1107) );
  OAI22_X1 U1582 ( .A1(n1118), .A2(target_PC_i[9]), .B1(\predict_PC[10][9] ), 
        .B2(n977), .ZN(n1140) );
  OAI22_X1 U1583 ( .A1(n1151), .A2(target_PC_i[9]), .B1(\predict_PC[11][9] ), 
        .B2(n974), .ZN(n1173) );
  OAI22_X1 U1584 ( .A1(n1184), .A2(target_PC_i[9]), .B1(\predict_PC[12][9] ), 
        .B2(n734), .ZN(n1206) );
  OAI22_X1 U1585 ( .A1(n1218), .A2(target_PC_i[9]), .B1(\predict_PC[13][9] ), 
        .B2(n731), .ZN(n1240) );
  OAI22_X1 U1586 ( .A1(n1284), .A2(target_PC_i[9]), .B1(\predict_PC[15][9] ), 
        .B2(n725), .ZN(n1526) );
  OAI22_X1 U1587 ( .A1(n969), .A2(target_PC_i[9]), .B1(\predict_PC[6][9] ), 
        .B2(n989), .ZN(n1007) );
  OAI22_X1 U1588 ( .A1(n800), .A2(target_PC_i[9]), .B1(\predict_PC[1][9] ), 
        .B2(n2263), .ZN(n822) );
  OAI22_X1 U1589 ( .A1(n834), .A2(target_PC_i[9]), .B1(\predict_PC[2][9] ), 
        .B2(n2260), .ZN(n856) );
  OAI22_X1 U1590 ( .A1(n868), .A2(target_PC_i[9]), .B1(\predict_PC[3][9] ), 
        .B2(n2257), .ZN(n890) );
  OAI22_X1 U1591 ( .A1(n902), .A2(target_PC_i[9]), .B1(\predict_PC[4][9] ), 
        .B2(n2254), .ZN(n924) );
  OAI22_X1 U1592 ( .A1(n936), .A2(target_PC_i[9]), .B1(\predict_PC[5][9] ), 
        .B2(n2215), .ZN(n958) );
  OAI22_X1 U1593 ( .A1(n1284), .A2(target_PC_i[7]), .B1(\predict_PC[15][7] ), 
        .B2(n725), .ZN(n2114) );
  OAI22_X1 U1594 ( .A1(n1251), .A2(target_PC_i[7]), .B1(\predict_PC[14][7] ), 
        .B2(n728), .ZN(n1275) );
  OAI22_X1 U1595 ( .A1(n1218), .A2(target_PC_i[7]), .B1(\predict_PC[13][7] ), 
        .B2(n731), .ZN(n1242) );
  OAI22_X1 U1596 ( .A1(n1184), .A2(target_PC_i[7]), .B1(\predict_PC[12][7] ), 
        .B2(n734), .ZN(n1208) );
  OAI22_X1 U1597 ( .A1(n1151), .A2(target_PC_i[7]), .B1(\predict_PC[11][7] ), 
        .B2(n974), .ZN(n1175) );
  OAI22_X1 U1598 ( .A1(n1118), .A2(target_PC_i[7]), .B1(\predict_PC[10][7] ), 
        .B2(n977), .ZN(n1142) );
  OAI22_X1 U1599 ( .A1(n1085), .A2(target_PC_i[7]), .B1(\predict_PC[9][7] ), 
        .B2(n980), .ZN(n1109) );
  OAI22_X1 U1608 ( .A1(n1051), .A2(target_PC_i[7]), .B1(\predict_PC[8][7] ), 
        .B2(n983), .ZN(n1075) );
  OAI22_X1 U1609 ( .A1(n1018), .A2(target_PC_i[7]), .B1(\predict_PC[7][7] ), 
        .B2(n986), .ZN(n1042) );
  OAI22_X1 U1610 ( .A1(n969), .A2(target_PC_i[7]), .B1(\predict_PC[6][7] ), 
        .B2(n989), .ZN(n1009) );
  OAI22_X1 U1611 ( .A1(n936), .A2(target_PC_i[7]), .B1(\predict_PC[5][7] ), 
        .B2(n2215), .ZN(n960) );
  OAI22_X1 U1612 ( .A1(n902), .A2(target_PC_i[7]), .B1(\predict_PC[4][7] ), 
        .B2(n2254), .ZN(n926) );
  OAI22_X1 U1613 ( .A1(n868), .A2(target_PC_i[7]), .B1(\predict_PC[3][7] ), 
        .B2(n2257), .ZN(n892) );
  OAI22_X1 U1614 ( .A1(n834), .A2(target_PC_i[7]), .B1(\predict_PC[2][7] ), 
        .B2(n2260), .ZN(n858) );
  OAI22_X1 U1615 ( .A1(n800), .A2(target_PC_i[7]), .B1(\predict_PC[1][7] ), 
        .B2(n2263), .ZN(n824) );
  OAI22_X1 U1616 ( .A1(n765), .A2(target_PC_i[7]), .B1(\predict_PC[0][7] ), 
        .B2(n2266), .ZN(n789) );
  OAI22_X1 U1617 ( .A1(n1284), .A2(n635), .B1(\predict_PC[15][24] ), .B2(n727), 
        .ZN(n1361) );
  OAI22_X1 U1618 ( .A1(n1251), .A2(n635), .B1(\predict_PC[14][24] ), .B2(n730), 
        .ZN(n1258) );
  OAI22_X1 U1619 ( .A1(n1218), .A2(n635), .B1(\predict_PC[13][24] ), .B2(n733), 
        .ZN(n1225) );
  OAI22_X1 U1620 ( .A1(n1184), .A2(target_PC_i[24]), .B1(\predict_PC[12][24] ), 
        .B2(n737), .ZN(n1191) );
  OAI22_X1 U1621 ( .A1(n1151), .A2(n635), .B1(\predict_PC[11][24] ), .B2(n976), 
        .ZN(n1158) );
  OAI22_X1 U1622 ( .A1(n1118), .A2(n635), .B1(\predict_PC[10][24] ), .B2(n979), 
        .ZN(n1125) );
  OAI22_X1 U1623 ( .A1(n1085), .A2(n635), .B1(\predict_PC[9][24] ), .B2(n982), 
        .ZN(n1092) );
  OAI22_X1 U1624 ( .A1(n1051), .A2(n635), .B1(\predict_PC[8][24] ), .B2(n985), 
        .ZN(n1058) );
  OAI22_X1 U1625 ( .A1(n1018), .A2(n635), .B1(\predict_PC[7][24] ), .B2(n988), 
        .ZN(n1025) );
  OAI22_X1 U1626 ( .A1(n969), .A2(n635), .B1(\predict_PC[6][24] ), .B2(n2214), 
        .ZN(n992) );
  OAI22_X1 U1627 ( .A1(n936), .A2(n635), .B1(\predict_PC[5][24] ), .B2(n2253), 
        .ZN(n943) );
  OAI22_X1 U1628 ( .A1(n902), .A2(n635), .B1(\predict_PC[4][24] ), .B2(n2256), 
        .ZN(n909) );
  OAI22_X1 U1629 ( .A1(n868), .A2(n635), .B1(\predict_PC[3][24] ), .B2(n2259), 
        .ZN(n875) );
  OAI22_X1 U1630 ( .A1(n834), .A2(n635), .B1(\predict_PC[2][24] ), .B2(n2262), 
        .ZN(n841) );
  OAI22_X1 U1631 ( .A1(n800), .A2(n635), .B1(\predict_PC[1][24] ), .B2(n2265), 
        .ZN(n807) );
  OAI22_X1 U1632 ( .A1(n765), .A2(n635), .B1(\predict_PC[0][24] ), .B2(n2268), 
        .ZN(n772) );
  OAI22_X1 U1633 ( .A1(n1284), .A2(n653), .B1(\predict_PC[15][27] ), .B2(n727), 
        .ZN(n1328) );
  OAI22_X1 U1634 ( .A1(n765), .A2(n653), .B1(\predict_PC[0][27] ), .B2(n2268), 
        .ZN(n769) );
  OAI22_X1 U1635 ( .A1(n800), .A2(n653), .B1(\predict_PC[1][27] ), .B2(n2265), 
        .ZN(n804) );
  OAI22_X1 U1636 ( .A1(n1251), .A2(n653), .B1(\predict_PC[14][27] ), .B2(n730), 
        .ZN(n1255) );
  OAI22_X1 U1637 ( .A1(n868), .A2(n653), .B1(\predict_PC[3][27] ), .B2(n2259), 
        .ZN(n872) );
  OAI22_X1 U1638 ( .A1(n1218), .A2(n653), .B1(\predict_PC[13][27] ), .B2(n733), 
        .ZN(n1222) );
  OAI22_X1 U1639 ( .A1(n969), .A2(n653), .B1(\predict_PC[6][27] ), .B2(n2214), 
        .ZN(n973) );
  OAI22_X1 U1640 ( .A1(n936), .A2(n653), .B1(\predict_PC[5][27] ), .B2(n2253), 
        .ZN(n940) );
  OAI22_X1 U1641 ( .A1(n1018), .A2(n653), .B1(\predict_PC[7][27] ), .B2(n988), 
        .ZN(n1022) );
  OAI22_X1 U1642 ( .A1(n902), .A2(n653), .B1(\predict_PC[4][27] ), .B2(n2256), 
        .ZN(n906) );
  OAI22_X1 U1643 ( .A1(n1184), .A2(n653), .B1(\predict_PC[12][27] ), .B2(n737), 
        .ZN(n1188) );
  OAI22_X1 U1644 ( .A1(n834), .A2(target_PC_i[27]), .B1(\predict_PC[2][27] ), 
        .B2(n2262), .ZN(n838) );
  OAI22_X1 U1645 ( .A1(n1151), .A2(n653), .B1(\predict_PC[11][27] ), .B2(n976), 
        .ZN(n1155) );
  OAI22_X1 U1646 ( .A1(n1118), .A2(n653), .B1(\predict_PC[10][27] ), .B2(n979), 
        .ZN(n1122) );
  OAI22_X1 U1647 ( .A1(n1085), .A2(n653), .B1(\predict_PC[9][27] ), .B2(n982), 
        .ZN(n1089) );
  OAI22_X1 U1648 ( .A1(n1051), .A2(n653), .B1(\predict_PC[8][27] ), .B2(n985), 
        .ZN(n1055) );
  OAI22_X1 U1649 ( .A1(n1284), .A2(n658), .B1(\predict_PC[15][30] ), .B2(n727), 
        .ZN(n1295) );
  OAI22_X1 U1650 ( .A1(n1184), .A2(n658), .B1(\predict_PC[12][30] ), .B2(n737), 
        .ZN(n1185) );
  OAI22_X1 U1651 ( .A1(n1151), .A2(n658), .B1(\predict_PC[11][30] ), .B2(n976), 
        .ZN(n1152) );
  OAI22_X1 U1652 ( .A1(n800), .A2(n658), .B1(\predict_PC[1][30] ), .B2(n2265), 
        .ZN(n801) );
  OAI22_X1 U1653 ( .A1(n902), .A2(n658), .B1(\predict_PC[4][30] ), .B2(n2256), 
        .ZN(n903) );
  OAI22_X1 U1654 ( .A1(n868), .A2(n658), .B1(\predict_PC[3][30] ), .B2(n2259), 
        .ZN(n869) );
  OAI22_X1 U1655 ( .A1(n834), .A2(n658), .B1(\predict_PC[2][30] ), .B2(n2262), 
        .ZN(n835) );
  OAI22_X1 U1656 ( .A1(n936), .A2(n658), .B1(\predict_PC[5][30] ), .B2(n2253), 
        .ZN(n937) );
  OAI22_X1 U1657 ( .A1(n969), .A2(n658), .B1(\predict_PC[6][30] ), .B2(n2214), 
        .ZN(n970) );
  OAI22_X1 U1658 ( .A1(n1018), .A2(n658), .B1(\predict_PC[7][30] ), .B2(n988), 
        .ZN(n1019) );
  OAI22_X1 U1659 ( .A1(n1118), .A2(n658), .B1(\predict_PC[10][30] ), .B2(n979), 
        .ZN(n1119) );
  OAI22_X1 U1660 ( .A1(n765), .A2(n658), .B1(\predict_PC[0][30] ), .B2(n2268), 
        .ZN(n766) );
  OAI22_X1 U1661 ( .A1(n1085), .A2(n658), .B1(\predict_PC[9][30] ), .B2(n982), 
        .ZN(n1086) );
  OAI22_X1 U1662 ( .A1(n1251), .A2(n658), .B1(\predict_PC[14][30] ), .B2(n730), 
        .ZN(n1252) );
  OAI22_X1 U1663 ( .A1(n1051), .A2(n658), .B1(\predict_PC[8][30] ), .B2(n985), 
        .ZN(n1052) );
  OAI22_X1 U1664 ( .A1(n1218), .A2(n658), .B1(\predict_PC[13][30] ), .B2(n733), 
        .ZN(n1219) );
  OAI22_X1 U1665 ( .A1(n1284), .A2(n659), .B1(\predict_PC[15][28] ), .B2(n727), 
        .ZN(n1317) );
  OAI22_X1 U1666 ( .A1(n1184), .A2(n659), .B1(\predict_PC[12][28] ), .B2(n737), 
        .ZN(n1187) );
  OAI22_X1 U1667 ( .A1(n800), .A2(n659), .B1(\predict_PC[1][28] ), .B2(n2265), 
        .ZN(n803) );
  OAI22_X1 U1668 ( .A1(n1151), .A2(n659), .B1(\predict_PC[11][28] ), .B2(n976), 
        .ZN(n1154) );
  OAI22_X1 U1669 ( .A1(n902), .A2(n659), .B1(\predict_PC[4][28] ), .B2(n2256), 
        .ZN(n905) );
  OAI22_X1 U1670 ( .A1(n868), .A2(n659), .B1(\predict_PC[3][28] ), .B2(n2259), 
        .ZN(n871) );
  OAI22_X1 U1671 ( .A1(n936), .A2(n659), .B1(\predict_PC[5][28] ), .B2(n2253), 
        .ZN(n939) );
  OAI22_X1 U1672 ( .A1(n969), .A2(n659), .B1(\predict_PC[6][28] ), .B2(n2214), 
        .ZN(n972) );
  OAI22_X1 U1673 ( .A1(n1018), .A2(n659), .B1(\predict_PC[7][28] ), .B2(n988), 
        .ZN(n1021) );
  OAI22_X1 U1674 ( .A1(n834), .A2(n659), .B1(\predict_PC[2][28] ), .B2(n2262), 
        .ZN(n837) );
  OAI22_X1 U1675 ( .A1(n1085), .A2(n659), .B1(\predict_PC[9][28] ), .B2(n982), 
        .ZN(n1088) );
  OAI22_X1 U1676 ( .A1(n1118), .A2(n659), .B1(\predict_PC[10][28] ), .B2(n979), 
        .ZN(n1121) );
  OAI22_X1 U1677 ( .A1(n765), .A2(n659), .B1(\predict_PC[0][28] ), .B2(n2268), 
        .ZN(n768) );
  OAI22_X1 U1678 ( .A1(n1251), .A2(n659), .B1(\predict_PC[14][28] ), .B2(n730), 
        .ZN(n1254) );
  OAI22_X1 U1679 ( .A1(n1218), .A2(n659), .B1(\predict_PC[13][28] ), .B2(n733), 
        .ZN(n1221) );
  OAI22_X1 U1680 ( .A1(n1051), .A2(n659), .B1(\predict_PC[8][28] ), .B2(n985), 
        .ZN(n1054) );
  OAI22_X1 U1681 ( .A1(n1284), .A2(n634), .B1(\predict_PC[15][29] ), .B2(n727), 
        .ZN(n1306) );
  OAI22_X1 U1682 ( .A1(n1184), .A2(n634), .B1(\predict_PC[12][29] ), .B2(n737), 
        .ZN(n1186) );
  OAI22_X1 U1683 ( .A1(n800), .A2(n634), .B1(\predict_PC[1][29] ), .B2(n2265), 
        .ZN(n802) );
  OAI22_X1 U1684 ( .A1(n1151), .A2(n634), .B1(\predict_PC[11][29] ), .B2(n976), 
        .ZN(n1153) );
  OAI22_X1 U1685 ( .A1(n902), .A2(n634), .B1(\predict_PC[4][29] ), .B2(n2256), 
        .ZN(n904) );
  OAI22_X1 U1686 ( .A1(n868), .A2(n634), .B1(\predict_PC[3][29] ), .B2(n2259), 
        .ZN(n870) );
  OAI22_X1 U1687 ( .A1(n936), .A2(n634), .B1(\predict_PC[5][29] ), .B2(n2253), 
        .ZN(n938) );
  OAI22_X1 U1688 ( .A1(n969), .A2(n634), .B1(\predict_PC[6][29] ), .B2(n2214), 
        .ZN(n971) );
  OAI22_X1 U1689 ( .A1(n1018), .A2(n634), .B1(\predict_PC[7][29] ), .B2(n988), 
        .ZN(n1020) );
  OAI22_X1 U1690 ( .A1(n834), .A2(n634), .B1(\predict_PC[2][29] ), .B2(n2262), 
        .ZN(n836) );
  OAI22_X1 U1691 ( .A1(n1085), .A2(n634), .B1(\predict_PC[9][29] ), .B2(n982), 
        .ZN(n1087) );
  OAI22_X1 U1692 ( .A1(n1118), .A2(n634), .B1(\predict_PC[10][29] ), .B2(n979), 
        .ZN(n1120) );
  OAI22_X1 U1693 ( .A1(n765), .A2(target_PC_i[29]), .B1(\predict_PC[0][29] ), 
        .B2(n2268), .ZN(n767) );
  OAI22_X1 U1694 ( .A1(n1251), .A2(n634), .B1(\predict_PC[14][29] ), .B2(n730), 
        .ZN(n1253) );
  OAI22_X1 U1695 ( .A1(n1218), .A2(n634), .B1(\predict_PC[13][29] ), .B2(n733), 
        .ZN(n1220) );
  OAI22_X1 U1696 ( .A1(n1051), .A2(n634), .B1(\predict_PC[8][29] ), .B2(n985), 
        .ZN(n1053) );
endmodule


module fetch_block ( branch_target_i, sum_addr_i, A_i, NPC4_i, S_MUX_PC_BUS_i, 
        PC_o, PC4_o, PC_BUS_pre_BTB, stall_i, take_prediction_i, mispredict_i, 
        predicted_PC, clk, rst );
  input [31:0] branch_target_i;
  input [31:0] sum_addr_i;
  input [31:0] A_i;
  input [31:0] NPC4_i;
  input [1:0] S_MUX_PC_BUS_i;
  output [31:0] PC_o;
  output [31:0] PC4_o;
  output [31:0] PC_BUS_pre_BTB;
  input [31:0] predicted_PC;
  input stall_i, take_prediction_i, mispredict_i, clk, rst;
  wire   n5;
  wire   [31:0] PC_BUS;

  ff32_en_0 PC ( .D(PC_BUS), .en(n5), .clk(clk), .rst(rst), .Q(PC_o) );
  add4 PCADD ( .IN1(PC_o), .OUT1(PC4_o) );
  mux41_0 MUXTARGET ( .IN0(NPC4_i), .IN1(A_i), .IN2(sum_addr_i), .IN3(
        branch_target_i), .CTRL(S_MUX_PC_BUS_i), .OUT1(PC_BUS_pre_BTB) );
  mux41_1 MUXPREDICTION ( .IN0(PC4_o), .IN1(predicted_PC), .IN2(PC_BUS_pre_BTB), .IN3(PC_BUS_pre_BTB), .CTRL({mispredict_i, take_prediction_i}), .OUT1(PC_BUS) );
  INV_X1 U1 ( .A(stall_i), .ZN(n5) );
endmodule


module top_level ( clock, rst, IRAM_Addr_o, IRAM_Dout_i, DRAM_Enable_o, 
        DRAM_WR_o, DRAM_Din_o, DRAM_Addr_o, DRAM_Dout_i );
  output [31:0] IRAM_Addr_o;
  input [31:0] IRAM_Dout_i;
  output [31:0] DRAM_Din_o;
  output [31:0] DRAM_Addr_o;
  input [31:0] DRAM_Dout_i;
  input clock, rst;
  output DRAM_Enable_o, DRAM_WR_o;
  wire   was_taken_from_jl, was_branch, was_jmp, was_taken, mispredict,
         take_prediction, dummy_S_EXT, dummy_S_EXT_SIGN, dummy_S_MUX_LINK,
         dummy_S_EQ_NEQ, exe_stall_cu, dummy_S_MUX_MEM, dummy_S_RF_W_wb,
         dummy_S_RF_W_mem, dummy_S_MUX_ALUIN, stall_exe, \dummy_S_FWA2exe[1] ,
         n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22;
  wire   [31:0] dummy_branch_target;
  wire   [31:0] dummy_sum_addr;
  wire   [31:0] dummy_A;
  wire   [31:0] NPCF;
  wire   [1:0] dummy_S_MUX_PC_BUS;
  wire   [31:0] PC4;
  wire   [31:0] TARGET_PC;
  wire   [31:0] predicted_PC;
  wire   [31:0] IR;
  wire   [31:0] AtoComp;
  wire   [4:0] rA2reg;
  wire   [4:0] rB2reg;
  wire   [4:0] rC2reg;
  wire   [31:0] help_IMM;
  wire   [31:0] wb2reg;
  wire   [1:0] dummy_S_FWAdec;
  wire   [4:0] muxed_dest2exe;
  wire   [4:0] D22D3;
  wire   [1:0] dummy_S_MUX_DEST;
  wire   [12:0] ALUW_dec;
  wire   [31:0] W2wb;
  wire   [31:0] dummy_B;
  wire   [31:0] A2exe;
  wire   [31:0] B2exe;
  wire   [4:0] rA2fw;
  wire   [4:0] rB2mux;
  wire   [4:0] rC2mux;
  wire   [31:0] IMM2exe;
  wire   [12:0] ALUW;
  wire   [31:0] X2mem;
  wire   [31:0] S2mem;
  wire   [1:0] dummy_S_FWB2exe;
  wire   [4:0] D32reg;

  fetch_block UFETCH_BLOCK ( .branch_target_i(dummy_branch_target), 
        .sum_addr_i(dummy_sum_addr), .A_i(dummy_A), .NPC4_i(NPCF), 
        .S_MUX_PC_BUS_i(dummy_S_MUX_PC_BUS), .PC_o(IRAM_Addr_o), .PC4_o(PC4), 
        .PC_BUS_pre_BTB({TARGET_PC[31:21], n15, TARGET_PC[19:17], n14, 
        TARGET_PC[15:9], n16, TARGET_PC[7:0]}), .stall_i(n11), 
        .take_prediction_i(take_prediction), .mispredict_i(mispredict), 
        .predicted_PC(predicted_PC), .clk(clock), .rst(rst) );
  btb_N_LINES4_SIZE32 UBTB ( .clock(clock), .reset(rst), .stall_i(n10), 
        .TAG_i(IRAM_Addr_o[5:2]), .target_PC_i({TARGET_PC[31:21], n15, 
        TARGET_PC[19:17], n14, TARGET_PC[15:9], n16, TARGET_PC[7:0]}), 
        .was_taken_i(was_taken), .predicted_next_PC_o(predicted_PC), .taken_o(
        take_prediction), .mispredict_o(mispredict) );
  fetch_regs UFEETCH_REGS ( .NPCF_i(PC4), .IR_i(IRAM_Dout_i), .NPCF_o(NPCF), 
        .IR_o(IR), .stall_i(n12), .clk(clock), .rst(rst) );
  jump_logic UJUMP_LOGIC ( .NPCF_i(NPCF), .IR_i({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, IR[25:0]}), .A_i(AtoComp), .A_o(dummy_A), .rA_o(rA2reg), .rB_o(
        rB2reg), .rC_o(rC2reg), .branch_target_o(dummy_branch_target), 
        .sum_addr_o(dummy_sum_addr), .extended_imm(help_IMM), .taken_o(
        was_taken_from_jl), .FW_X_i(DRAM_Addr_o), .FW_W_i(wb2reg), 
        .S_FW_Adec_i(dummy_S_FWAdec), .S_EXT_i(dummy_S_EXT), .S_EXT_SIGN_i(
        dummy_S_EXT_SIGN), .S_MUX_LINK_i(dummy_S_MUX_LINK), .S_EQ_NEQ_i(
        dummy_S_EQ_NEQ) );
  dlx_cu_MICROCODE_MEM_SIZE64_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE13 UCU ( 
        .Clk(clock), .Rst(rst), .IR_IN({IR[31:16], 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, IR[10:0]}), .stall_exe_i(exe_stall_cu), .mispredict_i(n21), 
        .D1_i(muxed_dest2exe), .D2_i({D22D3[4], n19, n20, n17, n18}), 
        .S_MUX_PC_BUS(dummy_S_MUX_PC_BUS), .S_EXT(dummy_S_EXT), .S_EXT_SIGN(
        dummy_S_EXT_SIGN), .S_EQ_NEQ(dummy_S_EQ_NEQ), .S_MUX_DEST(
        dummy_S_MUX_DEST), .S_MUX_LINK(dummy_S_MUX_LINK), .S_MEM_W_R(DRAM_WR_o), .S_MEM_EN(DRAM_Enable_o), .S_RF_W_wb(dummy_S_RF_W_wb), .S_RF_W_mem(
        dummy_S_RF_W_mem), .S_MUX_ALUIN(dummy_S_MUX_ALUIN), .stall_exe_o(
        stall_exe), .stall_dec_o(n12), .stall_fetch_o(n11), .stall_btb_o(n10), 
        .was_branch_o(was_branch), .was_jmp_o(was_jmp), .ALU_WORD_o(ALUW_dec), 
        .S_MUX_MEM_BAR(dummy_S_MUX_MEM) );
  dlx_regfile RF ( .Clk(clock), .Rst(rst), .ENABLE(n22), .RD1(1'b1), .RD2(1'b1), .WR(dummy_S_RF_W_mem), .ADD_WR({D22D3[4], n19, n20, n17, n18}), .ADD_RD1(
        IRAM_Dout_i[25:21]), .ADD_RD2(IRAM_Dout_i[20:16]), .DATAIN(W2wb), 
        .OUT1(AtoComp), .OUT2(dummy_B) );
  decode_regs UDECODE_REGS ( .A_i(AtoComp), .B_i(dummy_B), .rA_i(rA2reg), 
        .rB_i(rB2reg), .rC_i(rC2reg), .IMM_i(help_IMM), .ALUW_i(ALUW_dec), 
        .A_o(A2exe), .B_o(B2exe), .rA_o(rA2fw), .rB_o(rB2mux), .rC_o(rC2mux), 
        .IMM_o(IMM2exe), .ALUW_o(ALUW), .stall_i(stall_exe), .clk(clock), 
        .rst(rst) );
  execute_regs UEXECUTE_REGS ( .X_i(X2mem), .S_i({S2mem[31:4], n9, S2mem[2:1], 
        n8}), .D2_i(muxed_dest2exe), .X_o(DRAM_Addr_o), .S_o(DRAM_Din_o), 
        .D2_o(D22D3), .stall_i(1'b0), .clk(clock), .rst(rst) );
  execute_block UEXECUTE_BLOCK ( .IMM_i(IMM2exe), .A_i(A2exe), .rB_i(rB2mux), 
        .rC_i(rC2mux), .MUXED_B_i(B2exe), .S_MUX_ALUIN_i(dummy_S_MUX_ALUIN), 
        .FW_X_i(DRAM_Addr_o), .FW_W_i(wb2reg), .S_FW_A_i({\dummy_S_FWA2exe[1] , 
        n13}), .S_FW_B_i(dummy_S_FWB2exe), .muxed_dest(muxed_dest2exe), 
        .muxed_B({S2mem[31:4], n9, S2mem[2:1], n8}), .S_MUX_DEST_i(
        dummy_S_MUX_DEST), .OP({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .ALUW_i(ALUW), 
        .DOUT(X2mem), .stall_o(exe_stall_cu), .Clock(clock), .Reset(rst) );
  mem_regs UMEM_REGS ( .W_i(W2wb), .D3_i({D22D3[4], n19, n20, n17, n18}), 
        .W_o(wb2reg), .D3_o(D32reg), .clk(clock), .rst(rst) );
  mem_block UMEM_BLOCK ( .X_i(DRAM_Addr_o), .LOAD_i(DRAM_Dout_i), .W_o(W2wb), 
        .S_MUX_MEM_i_BAR(dummy_S_MUX_MEM) );
  fw_logic UFW_LOGIC ( .D1_i({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .rAdec_i(
        IR[25:21]), .D2_i(D22D3), .D3_i(D32reg), .rA_i(rA2fw), .rB_i(rB2mux), 
        .S_mem_W(dummy_S_RF_W_mem), .S_wb_W(dummy_S_RF_W_wb), .S_exe_W(1'b0), 
        .S_FWAdec(dummy_S_FWAdec), .S_FWA({\dummy_S_FWA2exe[1] , n13}), 
        .S_FWB(dummy_S_FWB2exe), .S_mem_LOAD_BAR(dummy_S_MUX_MEM) );
  INV_X2 U9 ( .A(n7), .ZN(was_taken) );
  AOI21_X1 U10 ( .B1(was_taken_from_jl), .B2(was_branch), .A(was_jmp), .ZN(n7)
         );
  INV_X1 U11 ( .A(n12), .ZN(n22) );
  BUF_X1 U12 ( .A(D22D3[0]), .Z(n18) );
  CLKBUF_X1 U13 ( .A(mispredict), .Z(n21) );
  BUF_X1 U14 ( .A(D22D3[1]), .Z(n17) );
  BUF_X1 U15 ( .A(D22D3[3]), .Z(n19) );
  BUF_X1 U16 ( .A(D22D3[2]), .Z(n20) );
endmodule

